

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XpL1TFj1Z4ZooJGB3dSP6Pc8XBohs9jsfkhCnRPv/E0eBWI+lHNIXEa4u+PJkwlVZvWcONLhadzL
udIJCZSJZw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YotU/iVRJw4SZslAhIDvcJ/D97KMnOVr3qgyDEyjv8wq6q2fLHhj3+4ICqb6ugcylGrOPKTM6GCu
GySdwK4bI3nrS9w0oaYDzVELEOvqIm4XJLCRGucgroBYyoA8PVkBaBN/hy1UZ2eFbtpqDZTDDmUW
gnhHXGIQXAKgWs/2+Vs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FTBaXnVGlPEYCL5pjYNf/Hfv9XxLlTrcGa+WNNYupZxR3vhtfNpZc42MK/1NS/s40uJdFgxDtyJC
45US5Se8hJI4b4aDwCX364idcRnwiaGry68POf9K8M/hGFpyZ9lO5vMRxcwi4PxsPQ8qmw8HByT4
OYHJzj5VZVht/NK8xDiyoIlP036O3ULaNwMwFHKTcQi5PfIjaD1Kf2hlmMtRmABdZgxWPM2aDyjd
/VJT/RN4hCqzU/34S/Xah5tV1LyNxh8bcoQcleD/8qoNOksi1KJWJ4VINA38up8YMtfghuRTGnUb
+GbLphUSgnxkE/cYRoPFpMRVyCe+M8TQljtPag==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RVJj7ij2TGFxBIQZaIX4ashUMEnPhUxpISxR5SCF5aX5jiCNzK4ERRG6UskPCAjcM/jCqieLq27C
qmTGaTpcaUcgUesfno54IOnoTxDkZMAiDUFH/1LlefExhF1XPDvaM/vElL+mKPOPIlno9IJyNJc1
zEpJkhiPrTqkzb8KZEd0vDlGi51GzyO61dXEmY563+nDtGW0yt3UDR/7Kr4HrnSZOXgBfBllkyU/
Ltqsv1GP2HVOiHJjq73GH4jn9otgCggzWxZ2YJvkIgp/91ApwOMvBeAC4XN6dZXeU1ne9oj2vr/m
9sZH5pmnU4B5jLXGlgcB+gkSLnMODUbub08jEw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gyVZLPzK5/qGBvghd1xSzWzNxT9MZeYl7bwDM36gyqd97MSrHl5ctqmZZjV8VXmrvWlQtD5Wtf8M
Q1uYUw9jLLjLTNHK/wG1CxJ5o4twhIAQ/1VqquXRCqFkv0p3PNpB/uB9I7bTd4AWiaBbdAI7BtBw
pQG6NzdwiBg+PwPRZDs=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SLIEG44Bv4xTjB9v4fqBf1KZQbqfKca2IxfLjY4k9zESKdmwVnCmXrKEYqpYUxLJzCTdHsKD3S2n
FjbnjBB5Ipr6GLgGv0C2J70oz1d+i2v/Ude3vg89VTUFxsSxGevMvUSBnGTKAssdquUhBgmjAF7G
f249bTuKJj0kavAU86FhcUh+zwvj7mCkzuDzhzVkGMLizUdnLkDi41++Sbn49x7qC0fk9Eb9+cn5
hntm5QZ0vfbj9kz0xoreeY4r84nY12XBhaXYwSygISZfop41dAR5XcGn5qNOr/rSd8SiiAMMrDYj
bn5CvJHdPgE/d51yQsqPbl5UBX2PADtDQGjZTg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K6R6rom5y54yZsKd4jIAhbeBfM4n9MARJNMDeVGkxY2OqJ/8cW2x8wLAR43wEYFAHz2eQ8HK+Uod
wOl5zhtkBj8ASe0JmnE1aOBYUwHdGul8g2DXnoYOtrrNWJdyzb7UzcWutvF06RUuFZXUHTkTFySq
9cG/9L0pTjR1ZeNkI41RWJuoD/CLI9HUdBkfyNVMA7/98+qUdXLxPkH7NF1T17LIxenn+sQWe2Ht
xjAMgqFsM8iYLzuIO/iXG6rJy5W4SvrCeYbsRdCFERnoVKysadAJf87JmeuX7FYBbt3po4UMrumQ
UvSHKd09FRolFIgQRylhFGvGUu0A0do/Y1ezAQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ME17zFeYzdk7MyEYnQGDKeQBSCGppuWnQkdAdKigBsEhKvLNi54UcdCP533j6otidO3IOFIfZOvT
pMFZW8OTE9YcCi7t3SN3ESV4Ir5aC4TZZkHyt48WD7/CafAtx/FEQHYa2kknyjnkA9Pg5WKfZURm
dGfLQsQcFoVj/oZXtY2eqoP2S5YVXk/CrUH/dVkRBHNQEYPtWd4nn7wUI/CUNRtb+97SEHOSdvcx
q9+zdms5mWPPOj+o+NXjDwoX4ddjh04v7um6NEfjSx2nU8tdrSXSvP9FqYpHJNdEnzErIlKilsxO
5e52iv+pPKSqAPqzyQPKlRxZnf89sPbtqNrwYw==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Dl0p6TZc598ihI8QgsRd5Cxs37R2VCYY9gICl2cvqRWv2H8CrH9NUPD3aLwfUZTl+Yd8yrntWj9T
coqvorP8U4zO0oRGRPYsej4lA9y1iDlXyNcNumO9c1K3A4EiAXv5UZQEYGbDHFL1Nu2rAC+tKJEm
pe6NMC8VX4bchoEVOV1jra1Bz1ePqQ8kxNwemoTx78T1M1R5j2lBlNrk53FJuqo3P1RXoeJaZG7U
rPLzQ1j9mPvF0/mzJqfIZtE1a97g5PKv7TF/fI23MKSg3GyNJh3xu9dc97DLqEqPwYvKUgS7HKFa
oGwejJ0EI6BiVfHRcdFq6ZTSJAybKN5mf6PLjQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214096)
`protect data_block
uznzrgLas76zZ+d3UDB7OVPLENDTffoglPVhDVjWmMo5Rtgo5L9XP3ZVxj6aDq5MKSa8Uy78nOjn
UAIhbYFlCYM3AOtePj7ILrmt8k52x9eLtSgRf/fGOzI/h9osT8Dxb6gdMN7B29ZoKaKRYs8noi6n
w1aqVbOqkjPM846lCf3/1uHnHywZa3OOpawGX/rPtK6q0RU2K7TFEeD7HwOFygjVJ2FSLq6VTjyS
yyjn7X7Q82E/ubC9gH24HKO8JFqTDBdcv7hTgepQvVRLQSR5HahYKC/di/5/6DmX++T+HV4W7Q1h
22XloYdomaFCaysS0iuuSxzKs+X+jwkW3K0gGLGgGKYnQMgImvDuttstmLn196C5DYlLBd2yXMmK
vM6Mxvzl1LuVLRMJh4K0vfSeW59zqHlafPLN8rTgx9MawZL1JmCvE7MPExFfPf+/nu2aeftSoB81
S8LMKP64LYGVbUVL2QQtDhgqTXpxHln6bdf5lhtF2d6c5DJm7he/L31suiVKfswzPAl2DTuMafBZ
55J1R2RarDzj31gPJw9+tc7dAl9JGgIwPilAe/i/1q5MAuQOOjTTOO3f1l4BLGfC+KXhthtJTqAT
QBCovYBgRi8WHkDyMc9YEP2Ghn4DflGJ02aRTzllp9U7TYrA95nG/rP6o8qp21gC3sjWQEerdRJT
f751E3tzBJgIAdLYPFsOvP3ORtOL6M2vUZyAguwW9WGSjt5OigPhT2tkjopLITm2LIhZRa6IPJkX
TI+Cxa3cKwPHqKs5j/+Q5UwtUEe7txjn3MAF4PeccsZ5QlrcTE/+NzyHI6Oh/FtG9RLUrjsA3Dal
1MYRZBnsE53cTDOC1Tm0ma/ysEi++OsXZsKRvU5fsmEv/0ZdHMMWSlfGaTPPuFIS6Ol0XlR/SIxq
Fo+Utwyi0DeNLVomYXRsyZiZZeJMLOMu+VpXRt5aBj14aaSJzT/VPFJll1a76eQyKjLU+GapMOoA
uGFx2XVkITkWEVnn3sFM1H949cYkLMI+6gbM6rMqQjUcWmaAh1+uOSB5YPfbDhGK2YwttYcxBFrZ
ozb/KkT37ps4XXOK7NwVJgwXvSWCH2z//nsEgYuIdtSD2AF1/HQLKyRVBJmhVKpJ9Yjx2E2dDkbg
FE/WMEcOOZEugn5FZdMw9x6zILBwOZWArCeQqGDzAIntYqL3htvj7rQ6x5w2UVXkEMb5XxyqOsa2
liv3vHeMWLfFhPctOANWJYq10VzdaE8QfOKrw4ADiDCofo0XoR3FRs60AhOZyRqMQHoO4R1+x2OH
9gShYFWhtYmcld9gMmkzHJnmrZtKM30iJLPjTINwl0kwIqMIitseAPfDmXAkhQiQO1T4blDwX3OZ
dVpToYsCyZY8LootC87wCFkenWhg0SUqzpWBFSQnUisKuxgxyj9O0r6ZTR6iyo8io9QoixIT1LWT
4YE/LpIE6lvWztj6Gww8psxIs15Sr/1RSztzxAHz/X9ngZzpHhYTHgwLf+6oFY6JUszWSIz15Ssr
w5s5G2abvdACsEeNUUCXffodX/uizhkq2KlBUESBpG7znFr6WtChG4uotq8Qp3ayQNqXzjsgjBvF
ATuOXZqFMsJW3/7RJYx5lBJfReD42T8jdQlEkD1Xcx1nHzEwhe3p3zJzxa1BY8aQDimnCUgzMaOM
JQDS/edySVfJKNas0oWKz8qRQKoqH2lOgGJsgK6EeZ2riZqDBqzhThMl5SBSk5RAaddwV6WywL2t
1NRTGlO+n+cCDTJpaBOMHO+GH8FsQbQWG0Jadog7wM7dytti4oM1fOWWHgBTIvI7VIZ0cKB/OsVJ
de5AAUoG7QVGgP3pplNd2walP2lstfUhifxD3jOO13tUZI0geenkvAdqGh5UHwANpGxXXfpogKP8
Cre33gh5ybTFeOh/mBHwcow/FDGkjTNYR/GpaYgoq94FyVt/0L+E6OdigIL2JwE+Jmwcw+Q+6+pX
4XWYpA9sIwGv8yYh1vdXvFSr5PJsyeP/TdEkdQOPpVtJiwsNJfnnoHeW/qOo3xQ8h4KFCdutOsRN
Z1/RG4tm56Zrv4iIVEOHZkJXcx83WnfyncGyhJ1I9shOZP8IdX8QYrTF2Shvj6sNph7XNBOE3L96
VoNvVeRW4HLhuiNpObaAbxLJarssspjCofgPjmRt8q3Qgl4qKm4EGipb37ADke4oLgaqFF7jxzv/
S0a0vfB1SJKqcAreVRbgYOhEAlpEtuayq1t4WPrfEP40Ar4z/sxGdQ2hR5JeAqpvVnuieOZSPp+r
tfWaLkm/mWf2EUy0v/x7PhE7oTUzm7+dmKf3lMqxYAG8cjKM6GTP4PmonBa5EmS8oA8eCkXL1BJT
Jnrj8Z2V8zRrLp4Sztx71i1hp2pTNnoMqbXXcwJIVqB42Wj4VJdqZI0GbieQBN5NHxlrMSSmZ6Js
YuQYCWVaLc89kbmhT/8ZHxXkHtD0T+/ZpCsu7NQomdkWCaGl3vmqUYdCSUcZ4B0Z/Uql1qQBgVyZ
TfwwvXNfCGYso35/YMdiqQF24+9sKfXYOM88ijKMR0p2/hmZZ++K5KYlW8EuBpOiR+dPlVCXi/yX
hRIt7DNvVu5JKVjsMh0J6bp5aLVukXxC2wujm7FSvXEwHLxqgUbPZLwnCA+hk6bH27Kc29CDcTNU
i25yLJL/NMr2ul/sFFue8I8oF+BDmf//Areek5IclwHWkvY0nKOoCSCnSaZ8hCoi4IHLEEdNSfmu
NGVKx0TIQ54+3KuqU9lWq1Ps/wW4OsO0zH5T+g7DnceJUZSmpj50jEo2hyEVnf4Z9ZjMGrM8pLYd
NdBvUAAibXgiDq2rt+iA1DuFdVJky/hXGpgVXPapsfnPgIdmXnkI06/6h8+ffXuuMKW+M8L5+Wpu
jnwhXoNXJTs2ZExitPwv+Ag9Lr73zsQDVkR7G39XLO/6VxINEfMaVb/ckro+tX82HSPYtNKlHSdo
O1bhkpGVuUb+aIgsucx7v+pt5Wq6xoMjsSTmIPJMDT048+Z4d3UwIwLIY3TyAtRNihxfl9jcJjVX
CjYVn6C9HO6gIQrLg56VqjY1F2utIivMDpGHz84cV0EtqQTr3pUhp/EsuCSVg1Hog11a612ON+b4
g5s62TFmeRcxLYs7q31SfxAXm+SmU9R+9+Qo81MXICWv2oaoZjUr+S0kTFG5DHEfSViUw7LHvgp1
xHbyFQVtzRDht/wp3qCfp20sSw9WbH2RZt2WGxziRvFBVdS+BpimJMRZtpCLkWZGbi5jzM1I4NxD
8sBt1UeKJllGuQM4ByqilO6f9dOaCqt6a1vhOkOYFYaIKWqb+elQpX0LSzP8ECqme8pWGtmicvGO
b9KK629/AD6LN52E5akNf0DMuO2IUYNOMURfol/5jfWFm0HCLTM+yNWYBagcukoHs1gw2wrAk3CA
/Fv3ZSMJzsA3Y8TBp0fF3lUy+YUV6Sb9Hmr906eY+KijdFQLko6u84Xsal65HT+DOe2rX0/OaVlh
0FqABXjz+sfvqh5rXw3GlsGR+HxnOOyJCF85dPdbvqfP3vmkC37HL6RxakjULvXhltAUZzRDjghE
JK3cB4LbHN5GW0O18Ng6FENfLiPscQtVIlUQXeEqIB1WhNfxBmDXe288EtR+gVn2lkXz3Z1OyYqL
8kV7hXU5gAoybUc9jz7EfpfqPi5nakSGV4GTkPW+2ewewitNVr7n0Dj762KCO+wMWlnaotoxRr1i
TvAP/KR+/7C6GJlewzJifCG0tSrjFmeQY1B8R6jdNDwNoXduw6qxgeGROoDEA5r0YVg99cfzfHt8
oMpoVDPMxD9aV54nTCvW4JRXB23o8dooz7KyW0se/Nbqwdhv7fNEwAw3MtRePjyGz0+9srKjrYkB
yVVrvIMkhaiNQm077zSwma6t4mKA6d/5dSr0dFLdVgdGbxoy7vrfKvx12oQO/oTqzvaWaKG31HMb
/qT6DT3Y1/of5I/wfk9/xIewEJI6Wiu+8F2X9LoGJJDyMHy20/+dgkl15f03RJcWl11ss+IngE5w
LxMlySTxMvCBvw5xj4YF7UPQugEF8HweZRRaM63X4MpPNe+qC7EBC4lyu+z0mSiVmQoLMP0Aegl2
0D5fHzQoUgTnyNpi86PqDU+7o6j28kKyM5bTJTmi62NN2loQ0Viuvm9mxTPdH+paDO7NEIQq2hdH
GsklU3hZX9QJw7KgEAb/A1cXE3OHQ7lBmxpWwBOkH6GvY/kv9oQqCpYmqeUC9s7usB/lwqDVebZm
ZdJU2J3tDqs/Bgkjt2+FKeF8d5W87mr5xEcJ60ecS2TzFAH/HVLM1bO+VPNth2ijMNJb3rEgF/vr
Mx8GASgr/fb1XZGBrbn+Wt3fpBgrHwY1H+lLDvuAUzT+HZ5A5x039xFD4ic+mnjuD9UM4KyDOflN
vQ89cCs14pCReljkNPAzKcA/btItQxvHshmMaqFH49AqmOq8GDkoc0oQ4iVtsloADfodpD3TfYqq
MZ8iBG46GYR8ud64KlYbWyjAmc6VjNrM4HRZ/YScpwDJFetuCOArdsobegUm21gj1VPDRnPlyxkf
gy7pMiCN2Hv9/FcQ0A9ZfKuQRg3BGktC55HW+g4w/tC0o4GuGcbE1UDlVlN2pM2oi3R+kMvAqOr5
dNGF0yHzNKzolfV6O0RxGQvjExwEhIWYsiYL+DfHUHwBTgQS7JSfq/pwkYYalmswEQ2ltFSDQw0l
qAWmWoRJda168zr1Zt2Up/3meM2U5/yl+SBGdsJ1xgxX3pOjiX5lPtw7rKDjSThGhlt3w5Uf8i25
PORKiamLzaQtKeV4qw4KnoS8GM2m5x0S7NB00LukzkMpj1ujPdllyCc1ZUPP+UQ9abUV7Il+q64H
tnAwtXLnBby735BlfbPPDC9Z/uzy2Ae/iJbDaTFSc6VMdIJghz7ojPXGgfp2Ugn7F2IQb+zdX5sn
vX4vZCeJzBs10S9/AdNvQx1lvFvxtmLhtetoca8i9Czo6f48cG4hguc9yIjKMCCcWq2dvgctdmbz
a+gM/f1pZNYqLUEbv9T3qDr+G5/9htC29RFrPm7HdbS5ii08Jj7ePCbRqoqw0HCW9f2CmACss0De
H+r/mc0xLEZp8pMchU/PbDAKyrU6Ru9gPOebfnPP55AHLpPmBQAhkuYNo3YLYCz2QOwbznLaDuXD
HuZhC0/DmBuNsOIw0GwA96XrLJaoc8QSDksBwapGwmFO605XF9wcfKLPH69QREixY5HhY0aH3j38
6qGmDvlMNimRnN8JhY+EHmAL9kHrYjczJH7ksJGQB1vSOsNCEmR0RPZ9TswjIJswLnx5/mJbcHc+
HuCsoQMFBH89xwkPw17bRUWUeOwSl20pCmHAo8IZSA+8XM0TegApJktGX+JftMjwrgfxIAYe5gk/
Ya3nnF26XtT+5AGLjMXBJ04DDmOJVRiATryK00eegpscJqEIumhUUgefEYgm9JmU77FwwME/ZkJc
5DQQITM1w/NnrspOXk/AmuUU73RhG2qWWpJzBsABL9aPaXkCw24xExP+pLvKqOhX7hsYYA31GqnY
iWJq9JSgA+eRfG6ZDOuUN7cqulgJsPoXvdgElSX+iDDnjmnFnYW1tQXbkGrhb+L7ET78EduJ6sFf
J77jATmqE9JOmcIoEZwbrT/qmXCvTol7o/OHWj50PLiJS3kK4ijAX5V9n0YEIJlqGp3e3VOdGuhB
9D7VBMeLVnInJHb1rgq0fvme82WKW7hRhdZY8VJ33zIkpTevPD1zXLZQVLy171HfpoKG7m3gLr+Q
qS1mL+Nb3U6PEnKzBObRJKB7XLgF/COrUbjIUM600D5OqPD6GK1wZK0uuzhD4HZXpnXy03UVoWIY
jVCD14h+DAkygHhHRGobGK4fWmcz6ZBrg6JWGyNPCq6gzQ6BR+baEzJNMJlAsJadI+cCMxDmLU3h
5SPjVjPwzvKVNZwFjT4E3GJ61/fB57LRwXBM5/oxEMmv3yGfnZvPyLU0OltdlUQTud2iyjRbeXl8
Ede6dgxH5uGZcc9RkdP3Sm94HkbcxFyUS+CQPmcFjedxX+JVT78Kc3T4JSDhIx/jVCWNSjXnpHbd
dPjI3iDceVxl9S/YzIJBwbBvZt/yveb6cfnPOGwU9IHUbJ3TueuS4SZFRwaIxZwwOGMmB9mmHh2x
6ENQsbjBtDR6zHwQomiY8PtGZskmirATCx9WHn+Nx5RO6cm/6QCA7Ylog/HbUxVhRFqnnp6Mne+c
5U98uAE9QSr1yVz0TIH34qJXcu+S8zMuCdJiQAbtczpJeUTT+PqXP4JCBRRNTb7ZNuQvEjF2z2bN
0smmDoRLr9BQ2pATMkiOb1hnKfRXXvx9TW6S2Qs3Ai5C1cg415SLyj1SGMEfzH6lsHJPzv1lhx0F
Oj+ihuE4LSOGDa1amq9ojGKO7K2/wbXfnhr3dTsAbcTYLVW/8vT3kXjfzczZXAkaVOFLIaFaN911
cSZsEO+aO3Sw4z7tFVhpIz9kytJUWTPnMw6R/apNo26XzhWC5zMl1QsS6Iu5whMsXqo3VbM2JGdd
Tkp2mUU1K19KhSA063rO6In3awIj6n/IH7hq5p5hb8DM2iXyMgO+H+rth7Xv1nEcZRI2RKNwCQG6
w3RHO4jCY8iQapP1CxCuq+OFBKlQNBViwxPqv76xcb/0J6dn0jC6oYwX1dz9n4ClOhvwIS0+lC0p
LEe9+6GzovPGcT/JVfcrbM7PtH3/QbWoGFxI09kTZ6B8me6loB1AlIT/Pyj+4X4v1u8xEM32XzJa
HRwWuIqH7ljm66Lz0S0ECwGvDKEHafj5atP9qgrIPOMZBs5reIqrxdpST3BKdxDn7pTnDZ1uSeDt
8oEy86AZloURbhJKDLZ8Dbc5CtEzzXHEhUfM2Wzk41ZueIPsJ2NffwoTCL1ErThUMVztByTx/uiH
rB2xO17AP62cgQrIlU3kaNncr9tJ5jjt5CvYtoyoHbFy9SwPNJ83zB7FSeexnfqFm995Qg07U299
2UFairQwhmpbON8zc1Eh4FPljJYMlN28thdZbMQQe9iJrGb1nSYjpT1OzVIGy8x9oDBwJ9chFAzw
Wv9VPwEYpX3gnHOh2YP24q/RPTigg3PyE/U6rZ1zKvZ8LnRpLmY8hKtCwBbQcQt0kL9NfHJRUWbn
YfTfJrFXFUc4UuGfkcLm3tZGYBtdLDNhPKY/8NR0SoU55O/a+beAArdrvdUoMXyLCOyILsnQOBUV
iqaPOeAQHSeWn/2G0MANkI8j4OsH5te9RES3po2NsAdDL76hHJ6PnL0vSYkORKZw9/RRpTqvGJq3
5XtCBiBKIemAm/+HMTjyH9DKM25fPVrekZLZqiyNASR0j6RqnWjGKUp7bp8O9QyUpwLkih9RPTNb
u4ESL+naW6MK2Aai4mzfMOiR/uhTqFjkdgnKJPiweEZL6s6eLQxLbEDqFCyWOi0+0MrVxQUsxhg9
C5VuPDgJ/3e9471yWtS3pvsij4AyuNXH8RtEGqAqeR1V/+XmYBlVUzQNp+1S9ATs+XEIpT56kH2i
iCrvijh9z6QYFmuX2qgpRCYBKTD49uhhFzwEetBncSLSs0lcEUINpnEdGfXkz0MJIVD+Y/nO+KF6
RG60U2tZLrgBDbMwgT39fTsMAiSXfyD/hcCayfdCUeVK8L9YuxF0u24i9A96mGskAPBHG0/Ib8QX
NddQhEbMg6ht/d5NGJQcby6Jd6YU7h14yUPCkc78nDnlaeI/jMbxPMe2vC8IFZY0AkebXeXnE8IU
7mq7y4ITai3UJzVwtF4dLPkBK1WIVisqPhNWxtK26tYvzMUGQ83G1TxeclnRR0+js9JjfJeOO8LA
sgkcR3He1DLe5H7Bz+tBPVPt8zO44Ad5hjcHC18SLnFIs9yg40kNXf9gtmNjcIv+Ff6/RHryynuG
EPeZ3lbTooXuXnXUikmzfaz6kEwJl0FecuUBCoWAodiYkJ5mdiL60pcDORUCUepupDLn0xQ3tOsI
4omO41tSou94eIAhByrrgf+VS/yStJPV0bGLjFTqJYMG2+j4QtnM8i1aMxQQFwyNtLXR4m13V5Ek
ddNeccmOSOKurk1TrnE/Ds5va9wV8HUOitGw85nkou6FxGFVS7ycsw2fIOp/g+OPjRczC3AGR5nc
Mac29EsvLKe2sCvHMM6Q7kK6qESlqXjqIg4f+hT/x4Bw7b+R6XLOSRzsRMWrlMknvKyy1MjcriRW
9LNWVgUYrFOOzFW3Ct65yZWuBbzWKYinr5py5Ltgtacy4ROLhPVOH3y3wvC6z/FzKTl5DK128Ve3
Gn1Ib1S3dsLKT2azMfJ+/HRlHrPKuSF8a0k8IhU9DpdhQnu/kBRDTzTcK3umv5Uy6pPikPJp8u0z
cvwId3gN6ydeJmmd5zMD44LeZaWlQWCZRbONpSN2Gw1nxVhJDqO5E27PsGW6VT2JBWfqZOrNz2QU
cD2xQ+fAlR0hkqFhEm3wdk2LhuncH4sV1LVEkUiHOCou7hQ0VMw922Uuj1ZWSW2uxUatG5OzryQC
Qm6cKLrJnr0ZgLj9xz1gqseakeVKwlFynmgFHS3YKjifpFljoC/UDwafi0YbkTmERuhdcmGwE2YW
6NcKhh5hlziA6q/eDPB0vrd33xGsRs3VZab4gQrGtxPPRiAJOoSS+przYysL7YcDWHcTztnWvsMF
kJBDZxYjbpqllcmUTtjBYwtXx3xceCORPUgzGlxOO2QbClMYJDyyX7CjYJ5BMXP80V8qPuE3c+Vx
5L0vZ47NlI5rQLcODl1evAjOs5I64+QZE75E/VDq+l5C1I3+MzpPKLGlu4mNiVHev1XIUWeSKPPd
CS9j04gBjCYWks50/jPFJhtZcMvNXCTCkpf3S5PwLa/kGHv1Tv7dw881LNLJblLsfpbQhtci2CV4
dVOuktGgBcuXi/1C/X7pyWvm9pFFjGuVefyL8YHr/8JqGdqiJV+raozASO3tOjMtO1G/yIKZDoyC
0by11wXTELdVW0GWXmFoeqLx2s5qhWgyzzA1GZ9Ttm34AEAzQfAZrOazDgM0hAqEBdIwW3tg/wYr
I4Hogu4ESFfWG2/COaEvNY+Xoqcze4YuLQqtw9dJ8nVZmBSXt9q68KDPYgY9NdKp+u22x/wBj0Pt
AbZ2gy9+QU8rCgql71+AsAMiPVwLzxc9HO7oxsg4q0qpHCQrMPXjC6EDzV95wfcYpKqySQB4zXfe
42IOfEXFxbNuI+piFkm3jwBzyip7W565robPkdmqN8oeryyTzzUQdGY5rpNbcDDTF61OMqGDjZgQ
DAKFtZXiBaxEq5TG1Vtk7+VNe/EB8T7SnmrURjFD2+cGF6FwqS6L1GRC/wuJwpYjItHmOZITwb/i
rCaCkF5cRWtr8uwQgycERuS6TG4D79MpySCwP4Fl+6GRw/YVvD03xKv7fIbme9lV8UJOhUfO0/Cq
vftq9SXzX0lQutEO/h+jPkb1T4Z1XybNkA8ciS/8dtmB5VSeWctl6y0FKRh+O6OkaILOjDX3CTrU
fBRjwvHXirjt6Rt6H5mtkOG9ECbgEh0ViIB1czu/Ov2xx+Ht/EgwFNOPS+xF6qOXX/mGS3eYO+/a
ohcl6JRN8itMmt94awBrGqVQEBhJP89tQJ1Cj9FtyE9hy8fNP0Q9aPekNl7ZKzxkEpzQUf1HxtVe
oH/lHW0dd54ex3EWTo4T9Ospt4hjegVpdjOkR0l5W2NPx8vpl83gkNT7tMyvWbEHwy/jrrYb4pY7
FqAFfIONT7K8UCg/M3Mu/Jk53dHfb5JzEoAldtt11CuiTO1Ng05fcf+lYN5/LjX56mqETXXGmplo
3Ls/26Gk1SKtVPhBHtLrbEm9sSBFWeHU27dL+nR4sm182s6rPUBfS5nLuXdSoVYOkPxJ3waaT+18
zaUIEcYvr0t9wquCRaMQR3DYRjOWa/juRutcNg1DtGUvgrrm4Dfb1R455WnTsSZpU2K+JpIg/d/S
ZUcR7//vMrqmrAHL5RLNRgBYmpXuOAKeWmOdpb09XSNpdeJvPJI4ttTa/cMRhh7mDv2clgm9jOHV
plnqSSy7J9b1mqXpvmohYfCiFMK9sljKKShDx0urXwcrpBkp5xjiil2p7CZbsSbUl0fVxcPzw2FE
GXFVf6juBx8apq97skasyjM0I6Sd90hNaHjLP1bOKUKzFwxGbRE14XN5d4WN7CAN48ds6ojQm15D
alHCSGLd3nnFVB7Lyd2Zq2bBWL1TMUYn0An2AwH6iIFh2n9GYcvL8Xb2k+XtCC+PiOuWeL1GqfM5
pUyPS1eVwPVGlzwHvywjUJdymEIv07lqZ5pHNdsAYFTj9xc7KPEjemHmKuK9ZkVzyyjWqJWD57Mf
5B0Y7lvcVnh8qLjCWQOxT5PjMBcJzNTXGrYK+t2T7B4Bjmyo3fsvGF04hAGNsaq0D3vFt0bixIsL
+zxoOcl9rLYsEs1IXDbOmXag8Oq4kaBVA3F3Vcxls9RVHwEGxbxrsJOI0/1Ee6ypNjlZTzAHgZNg
q6c/QwlQxvOlUYVHuIygVG3fbJ2qBnj1+qMfd+mUJT4udJDEv5cRdb6qSwJt0uvyYcQVoyv647Lw
bNdS9kj3pbmtty5unMx0Ju2xknXrI46C8J7h7+1fkh3oThyjF9JB81r0UIAau91+HltjauMFzTZQ
Ki0bWOTWL8DMDYT49/0NJsvdJv6zk7JntW8PktckUxQOoXXEwQ0ws5uXmQmwjXrfHXwsRwbBfi8G
h43FroaLwsPBHFq3hADHWJUBWMa19dhbEzGoFjDju/drqt0aiusBR2AZdzP/3kZZ72PU5HxXkG58
oTc5BcVjQMH5F2vZFUciulCF2sVzbeGN4o8AXLlLf50VrU0NmhlseWYl490yMkyWbjj42t+3SHmk
T2OgSbVxeDdvONn+6mWAoEO6D3a2YAQCXHo7jqN7Jv/HfEddnz4db9CNpjFWuPV6++qjAzWebqEf
hBiTV3S/94DXssV8PKwzQYL6we6XqzLsVMGI+t4Ei1peTjpIYyPuLzaj/T13enQShcR23mbIlaze
DEj9OhcSto75R3+uqrb7fr+KJsbLKG2EgByvewxkA+HDDJjXkPJkGNd5fdK65Snld/r6BopyaYwv
D+UZS70eOMwHNITLM/6ip442gOT+91AzMchNrsIZkbP7S7oVcSk1sjUKh+cSOJFDSXspE8D1W10G
NxBjWQC7BSMjkW7SKP0qJOkJcH0vfZGGSLkzNKj2e+GthwzaUZkbJqSpM6SlwCNEcTCQRAhuSoNj
21Sd2KdnmyKbKCjxZV4cp1IhIjY+eYK/7cRTbD36bnewIczc7spHjj493cwvBmL4LQgCL5gGZBo7
bcvSXnzgVaBinslPZPnYZyQ4UxsCVnUHmHrH/V5VJIQCOhPqNiVWoby9ZwODo0AUx7OoAP7ehDny
g66VIBgjHnrRIPHhD0r00TRK2q8av333tkWaF0qe4flzFf9sEmzCZSz2HBsJd1f1eNTs5UAw4gQR
L8Bl2N0Q9vnXGG+80llJPe7y42qnZUsLVoWwOZ4IuUvG5t2lId3ekT5nVoRmcZdSz+u0BvlPB9QF
owOOd3qejiBchjmhAXDruPScsDxPoR/l7Olhu0XPxBOcCH3+u6FbHm5l/tS9UNOnHFMt3HAh6wAH
3P9gPtje2QvqC0fuaAzH56YtO0KpAk9i+Aj4P7fxXnvYx7HD594puYlQW3cb4zqxPeraMrZgctEC
7v0xTe2qR/Tk5K6bVwv405Rg9HjULtdXJsr3qhfBHvyxMfEfE3U/62CdyhI8B598jNqJM/ruiv2A
eiUz0xXx0iXUdatVwr2R0EgDp6KWyHFSCd2pkHxtHJ5QIZFxq/0hQRTYO4fBoVOGkOvkK3wMdGLq
D2GDx5oh7T9OkpDwVzcJQbzeRvxTS1nTgMOE8ba9KRIOEgHFKkmB41TsqxV6+pnxAWEfxp881kaT
DyU/jC0VOw/voQzg4JvUgGG/rgtz4uvjFjUCbzFaROTbh5u4LEewt8mSsDCY5Tzq2ctOMz09Y2oR
Lk4OtSP3VFg1prpN1A1w4/X5P/VVqBLKeuR6Qp9B643jH5omdxyMIQWi8RNDLK4B83K739P5z3+s
4gSMaPMbC9YfEt6qcB1FNN8r4q8SOr438h7ZOjV6Lajs6ajGyATtKIStYi7q1t1Xamd4eFk8Nn+y
I0CaSH7bvCUAh8e5walvvPTkmi4aiegh47rFr5hpCzie7azUcSUQPvA6+/p8cDY8n3Rxa14fNXaZ
6b6/IsCNH1QYSUcBZ1akxorTIvia9e+m0SvLegoxR/Y0RK3jTDPaBaD50cMbprxY5fCpN3gdx83N
Rd1KZBfTEREcyF0W15HRqNh42SsGDg90+5iRztAaPCdJF6xtF6jsrFmNyv3fZ3t4lbDOBZWxwlMG
JZErZO4Nvu6lCp65SFMjXvA5mt5jb5eCGaQ0W8sSBpHym+ZGnhtioTFKwzuHVFgeXiPnqGTYuA/R
n17s5ou+1HIPYkK17PCwNu3aDXJkxVDsIfzuyaO1AlWSOThRy3kDJx7eJYE4Hj/BS6QgFP+XAVMz
+jYzpMiWsrbThaCrmGjf7VmelGF1xzmAjpQMk8QNF8Tv8CbbLvhPuX8jM/m/QBgl1qFTuqVBFb1K
doAlw8mQ/nxYfPKIne5ffztM1OTAHiN/fk3c76Vn0k1nH7sSSuqYJc9DCDFhIFBwDudrnQU4Wse0
Q3uFOSPRoIctG6gOuPbRkIIqe95VS2k8K7loQTLhxHdVcgFkeN5Y/BFp3QHD6tCKVA94PJpB/MBW
fMUNYygn9cVD6HDaV0ztiyereuIzQ4307PHMsucfm7fyD5Zs1wMW8aKhQYBSTbS/nO8DUGzs7TNe
P6HgqNJ6O9mrEl+Ob+M7PFvWQCQ0zhi30OhCB5KFYwNFL0oUFcZXHcFL0IPgqGLx+Ip4ntzIoVoi
LUZba2kPzfxI3O6yG6PCq0uMCTdt/UeOd2y6R65SId55/ieMb++xmAkeOMH3hVJwmTGnFPOGuc4u
ZZcDbm/8daYTd+SbiNyOI3zA97Y6VSS2m0o7kITyD2h9gnoujE5R3zDdXgmqIyDtUy4wtT0Zogqz
19Lybw8ufU5JJqRY/F7HHFQjdGUosIw4sI1AE2LXYmhhicFk7VNGAUF+GTCsa1AjOUUzM0rYVAJQ
qLPfqQJm5odMOPSXts7mGddVDvSV7W+9UIj/xuSeuuk5qQJ8zRG9QiD9dL/xoAwp5yOVEtXBRkWM
eV1OnK9jmIxeCjDzC6fd2qEE0qBUwGFDHKB/kq7QtJU848FEjyRroLRVpzNew3t68/28OWVo0pOr
KY175MGGXxYivlxVLjHQ4eBqk8dEmwLUy1ZegYNbE/Oyof6WWiop8DOa83kob02U4U3nmO/JYwRr
MbyRJ0aGdKqiANpeEeB2hiU0F/2fpoXoFfDkxEXML1iRwCS3F45HtP7yYhFayeruTJZ07iTrUh2d
at5JLkVKAkET2LXZpDjl1fX5f8qTqjqRXnO0tQnpkEaaTOmizqugZf+zx1knZGwMz4TAnwn8Jt4s
3zIqvrdvemtg731Ptg0TY1jMDVwWMMF9w8UtKxWnjcw+mCHX4v4l865159O6ZlAjRLMz0nKMrViV
KztNaJMuBsg8Y9y+rh5jC2L3fpixTxSycAdeZMyNM3yoov/v43U8JGc04gnmFXz+u7z8QYpKKZWp
PpCVEfYUvC4kPkbkA8qv6a56GVOHbFLQ2upaEg8her7pH3q8awo8tHUb0/KA7oYjmm51iscPiv5Q
yyKb1nFUkyWlDXQu0u2cLWeaQVqWHUO/W78OLXEmeYt+4FfJO77YK8bx+in6JJ78zu1QTknFO+iQ
0QuwQZJzAPkSXPlav+HeAsPVti26NJl1yuXx1uo3r4u0z/mxWq8C8MEx2U9xT3L2d8w2dfzhNBjV
8mExCUpFeWcXPNfOSu6MRiQA6zs/c9t/pXfxyZBRu642a0cLrk5J4TgdvxLQBZgXl82LZWeOYjmr
Fgcd6npZH4P7Lx8vomhWFvYYv47QHjBywuOpvPNZsTEfK9nOcG7AuAfGw93I9KvjcKqnFykhzsLp
qCpvfkESppGDvll21oKFv+Od4IIABzi+QJoBUSgg8jCdLhKoKnd4QL6S/7JtH0DsLsSDLz2DLmQz
RRAfeMg8X7BtYPMzncHQefQGUWnoeRCG3ZqQQQjkH7vJF3nnxJWEXJMvq/dPKJcY4WiHcbzulLUT
iH8QIrgVbaN955VdA4A/YLW5YJI/adQdFfXhGFKLe6pLP4L50rHuGLa2aimusdVVKH5EM9PlRsvE
Nmwh9h6oqHqjeVK0OuImt4xuZzJzKimMi8F79KZTQT01FN/c/c6K1eP6dgj3K0KYWf0KiROtxtpo
C4vidW5uAwXb+zI55bQZBQjMc2gXsbdN8bWoWJYrwNfM8BQ1uGNOFB5ioOMQ//qVwpYu0EjVRtyM
aCjGMo+v0PqU/LZbXoPXOWuAP0SamOosl5IHv5gvDBxDyPaJ1acKCsUNOspYf1IJ/Gla20i3gL9N
y3d22BVhQl/fibXgOWsf4qMSc7M0O8p23LitSRvTCDK+/+4UKvwtUgEq9U7OSXrmJcLd4Lrmzamo
+96q0jj8WVza6pCWZ7KDmPsasZ4mlzj+W67X3/Pd4CHIrjSFS09oLuxUvPgRGdsJwx+k7653kFsK
M4u7iPil1teRZLZoZ7W/kixod9sRiaHx1R0+X0C/0zFICFlGo4zXGNTthHDImDYhOmak7Y8YeNHy
ZOcGx8LmrswwF3Rt0qe9L396n8x+jmFtw2H4SU2jQwev7x4ZVGBQvRtz8DzX+GXfVxLkeHxqGBcN
cHqq/imdxo+/zInzSVwiG89tAfo55THAZuCESkvvBUJwJgs4c3sQ64yzKAgei6FePNxlrFLLKjYW
7YlHcJS5NaXvDUjwTw6qnf0R+oXq7KiXqchuNv4cPa4/Z/Y1DVKYbeqaxX6dUxBnEd54Zkyo0yx2
rEc2BMqKGf/bOJsfA+2kOv6F9eid0bOtP+fRUyMhMFvbsHBS0Bkw9tJF195VGZnqjCzldR3UUviX
gYS3qqaTPHFfdWeGjV8vsiTLMGONL0GvyZE1Hv6QVy9rENmXKcKoMsu4KqaMy6nwNG5sVK1jsa47
NxtiS6RnztK26sxPuP6kU4husx/jJYJXvqq/57lMBnTZ0WmYYYciG1+U30cAXyjxKdICgeSMyAfo
cYo3/SIeOi8MIw9XeEaBI6kFyw8lsgHXWx7pm7HXMmGsZfEu0e88qPmgKyuabNn++yLnLSuu3ZMQ
BDxn4GKfyLyZ/p33ogOD3c4HsYHtZFnSzOrBZtMw9sSBb2AtLdPsHscX3gYsb3KDj9ItLGlo71dq
mctPfqKQU0tGLXir4AIn+v6yrXPLk+nowRHDjmb+aYXNrZrhWxSUo1bxlSer0g07YCk1WhalAvXV
YnALMI8PE99/0bJxe9Vp9g/v4vJXvU4KIZbsRtRHfzfNVEFzxM6owQ+w1BzURlqqo1lN2LSL3oSn
vB119o5+ZjctyOigUpGdyaSOviTJ216UkWzySXuRXBSLbSohW46d9zK+POdFh0b9Z3k7JIO1tjmB
7ApyXPUZPgLG4IPa/C030D75JMey2hXut5MacE54S9ZXehBEc71jNGhzu0l1d0+tVGIfCrP+cYNJ
hJ6PfMb3nuPogPQZCyLpWSTk6jJ0WpOCJsHJg3slSi1F8vNnthg2YxrvTOHTeO7wKSg8xucWNd8R
w49QSg3yqDUz2P774dwmu0uvzz4gBobLSlgtKprzzukioIjj6TAUjDnHguddPb+hiEgmOOx7g3bA
DIOt/LXDyrATuKVaktklnhpctAJ/ceGNyI/FUVlPi0p5giD9kQ6GikXwV3Dep1P9n/GiaVvNvYYT
MmYuVbevwSKXIeZinqDF0lXWWNAg5F3Yjc/OXJWdsEnG8aufuRbKZNaFjEbj2nZ3kTZuEm+BiUnl
qnKNOF+vnNJdG46CgXdtee7HGtWLRM0kRKoEF0bhpweSB9pPsvGQ/ImTPdlTgAfBwJpyDOLTprmH
BfKqDyPcN9mCEUJRR3n0TUpD9lgYviGAdq+zTsxdCLXDL+tg432j0/HkYP8vWIYKE49WeuKLXYQ1
v3yslHCwwFivW3yV1sDqSGZSL0YI7dtOkwlaY7Nuu6vq9kcymXOF2ZyxFaK4e5ZnlpKl4AAhKw3J
+XGqglvpbhOOcv9T/38Hsb4aVH/8KnFZabWLWhgYrF+2LUtnAzbY+o5iqgAOpvLVOGIwyeNyd4NK
fp/3noz4FPTiD9sVleRLuErZSdkVrS/nKvGE0ALHu6XwelAcMntIhH3fpyfnmkzyjJ89rUvRQduR
3L6CRNdgNpm+iLCdrs3uk81ImZSjpDk2RvUR3urqVJVBPfTV8EX2OrfMyGreOJhh6MXcTte1VYxh
HBLb2TZRmtvUxP9UfZD5gdoIJ76OH7Iy7T7xmNQbh/wsIZSxm35l947PKIBJm3uzIuopGMkgPK1h
HxsWm6UQS8CYYo0RtW4eY4rIn5bQBzO5XhDfERO5wUGV3vzWSi6BQou4XvybF/8x7nsFQBU3yn9e
UVx5XOtAnFxQjNZbG2R9m0VQqjCCQ5PIIN0WUl9nQon/YAop0H+t8G820Xnh6umnOhxAc+1XPLGv
eyZTor1lZvK0mxMCjqDPWjskmqh/teAUwga+HayyGuuSkX0ZHNl9X+TvJS6KEaAFO+kF+cFxkblj
EG17ErEgXE/4TisYBYPBiQ7xDVtGTSn8TAmkIokXa5vCRXpZC7xMjUhG94FvmG+mKXJihCzxcr1q
3mQaaMjiMOO0MzQedxtHg/PL2fj6nlscLlbcKcmhJb/2IbjL8NxRlMjJ/13ftmVdNGXKp7ldJ9Fu
HfkByXe6FfZe6s26NDsovyleOLGjdIEAfrhX4OkIW2hL7SMkKqx0aP5W1vsfZtkO9xv04i8Ksokd
buR7DLRyFU5NBPB1+alO/U06N/JqlN60W5dhjMDthpXOHq4xoGgD66wJr9Vy9aBJvrDSoHLQniaK
S+tCr6UWVq1MVeZk9Dao7wi/0bTFRVd3jH7Pnss/70HNJ0r+HWfACbA8hlb0hGJxIC4mD0G3dOz8
0LbLWT6JmqMrvBuGgvFatsxGn989YMrc1yQQaOvDX+XT4HnMi5w8bsuPIcGqAYHgiYJ4zrnYkDOk
JnHkzNY34DV07ahuJYmiRrIze1KylxczMX0EpkktT6mmNdLhiY89w3sqwvjQLdXVXY8libRMLiXH
bKmkMNqC6GEgidyh4FCm58e/RJtEZmgiHXlQd6FOcS5TPWCFGCska3HskdWk5KLivVo+sGoK4fFK
qQbTt/YdhCHVBa69/rOzGlCMseRavOcF/EPj5zI31Y/881MLoeSN55q87W/SsAnMG0vMR9IcFPe9
upPGZlivNxAie02pk7hHOqtThH7Fd5U9od5emF+MHqzfHBtpxbY5/WCrjM9iwViahJgOLXMQB3vJ
Z8CWDFyoMP+VPlowyNtDU8b2tDqO5dXQm73sRa7QPKKPCvK8fTQ7HaeIP4FtQ1ffQJ9xrBLaUnBU
BVG7ud+InVVxkHSBynrnFEbwpibuUpbib1KaMC6sl8FNVw+wTsSigrf+9VWGYqIRyKwN4A/pckLM
DS2j6UpU9ULQb08izGOndNnBb+ySvtddhe4QgCwLmI9sX+NlSzxirllAHKZTEV2iCOD6CEdtqF4B
6rkkX8b8gHr9Hd1moZzgBNJDxY21WdbMUSgckmoahouyMo7LDBaMX/oPpHklVhxqjcax4MwMf8VS
Fuv+4t2+/RC0NdBDi2qm9DsATSvdq/s3370iLLHlvs14C1oWNuV3ykt6DOGIrw7Pg682Xa3mzmEW
lEwVsO94niZvrRcD/BQas4QC4Wm2CoRH1s2kYVMs10rk8Df50naISbmWqLpPy4PUleYXwhXzt7iQ
h5tZQMps/qoVEgrHbDoCbcCvrLBkzRE/eahy/MvGiuodFgq8UrcieeIkFIoOCeHkYjgvhUR3IZVO
N0i/oWJNyQJlpJAtODPIh0SotKN2g+OKA/TsTHKwQQvuJXxzeCK85LVxUt1OR08/i2XoMgjTyBUl
sXa91rtZ2Jko7TE1njdHUKqQZkxZBZ2KjTIE9BSWUjVWw8p7voiZpKeAcTVoPM5WhROnVIfWqTQm
5EghQ7eL5sv6yhJr8FkX5Dbq6XskG/Vjic2rnBInchV/9sMF1XXZw/ZOFhOw1RC6wZCWnrfGc7Nn
OucsuM9qZOzd+utclYDdbDynvD6PNmPTqtrAONi0YJu7XiLVsGB3caW5xO+NlwmTOYJmIL8KArUi
Ye32q9BuzDwJJ1PwWHqZtJmMtNTSJfOtLdPXBo3UruFtTa4YgCC9ucLzx80aAxI9Qi3eVG3CQOZx
bdMplttxKHAXbj0PP3yQMoRJu+quKVDjiAjLeyRLOQbZOZt5bGlsZbVuASM4tKOPPBJKhCS19W1z
9go2JTHssQOjgQiv6f3PNc8jqnJu85HG521TOPC3q7fQofeehVtrxkDl/u12pc5xlT4M6iSn7+Qg
ukfYvCB455kAv4Wc4nmLAzwtBkQf99/TM9S528BUzuOKAYplFTrK7jRiE5h+MC6KrrjfTeVfu61E
m1e93pLjoeHPm6pzTU5v9II83M/Aaa+Y9ifSdrjqKY0pEMH1eVYSM3x8mYxj4XlCZwSWLsGHi87h
xVQ/eP3jJ9gVgC/kXvRw4fXkKAhfKMrAWOS6OUWQ5XG7BQbJY/uA1mjmha2GxCstSgCnQtBsx22o
CGwldTQragP+kHyu60+eu8QJ8EJCPYHoI+IwpfUoWUq8PlpKfqxjHPkLgiQlz7ez7V9PsoHEfswg
2tJy2OsCn9cGp7Hi3YZlCSkLC81sMlfxtttOwf64GmAt/lyzDkft5rM0eBkpxQyFLQaFR628QQn4
MoOTXgNnuChzvVJ356rncg1llzQNKQpYkA7sqA3P9VmDlGFeNz4hXVP77USlnG+e5otjzmEbkM5c
A8lcgiZeZ4TPUbpco9U8UvD4kOZfKxpqM5+Q3CRb+C94k62w7R1cz0XmFyAIKZsSInrGenOaVyNw
q0lz/hH0juMWXIja8DrR/d7925Ud+5OrLJsydHPEVjWGzdwVWIGKP1ndN0VmL8ODK41te21KcuYq
iIzLYFjmD1waGWt7ClTI69Mv1Ar5hwJluTW4lt70pUJ2mpaaMDlQrfriZWsiTNHWaxA0hgjtq0rF
YoYBP6aDQ8zrqRPT+tFTyCJCb/0bPOhBBO03yBVsY4ML662SfS6/A/Lk93ZWfAhO5uJF53m7jc7e
2apBbtjCBkt4Sjh8ZXpwwW3okoqatrGfWc+mXIARSxNI03xuE7skQsWSp4C6yXxYPPBEmzh3iqrv
bCekYlyvqNd90dT+5whOJVy1B/nt+LcKMckGvaX1efYPXdYT2pK4RWT62nT5B+WtEYuNZvb6tJAg
8pLT4FASofd+vNCtKphuNBcy25yJdMjOmw4H07YWEcgVdoIHBYs6h58DyRQUYuNCl3OwTdC6l4ou
G1ylcY7qgk9QdnC6vXbbtY07wAStitNCldz2w0cl5XwcfQKzQ5LPHq3WwxwxjvPRuebGLHfRabzd
eODJ6eAok4anB8Emw0KauxpE8CPp3dbtwhlTGL5bS63w7L16ZRpTdXnGLUATtd5BTVCWx8kxEBg3
43MkFTr9M7Nu2iCp+lN7L1ExDb1az08s+dZrAwpV/VNlimgVpeQ8PLCTJM1audBh6vGlk2yVrRBJ
4Vn6lGGgqnLY9o9ycXRpfklyEk+GR7o5SAnlTLfNJ08rK3k2mFK+DFGJpTw6+AxAQ8/pW0qcZ5bY
F5PCeJgFgrvZxQlM5Jmr//neYyWfkODrIdBMKp5/cldpe0WPehDXPmefHzbPSo9EWvfO5Z1xaEnG
fpSWR6IrRI0zScpnawkMT2Sr2qlfwlSyCDsJiIzL8rXEHpTp/au510z3xefeSULVtedpE4ZZ8FFL
zKjnJGGtHBfa7oHz8rO5Mc0VaXeeApZa5I0xcRoROKNW82WHZjbdNeV6o06Ti0W0UuklQNwgSv44
31JBFzYKUmn/rY4eLcYIO2aSmywxMsB/pYW3ZX44IIbZoPdTCkhhcN0ErlrRkAv5CL98ehwUdxWX
eEab37JOc6YVChDzk27041pmIgjOY59Hhy7Iz3HFn31mvLg/Q4jisOynuAgpUcX/q7qXgsilRryu
0Azp9ac+75tsbFQbCbfV5+FPMD1l5oZUrF/GUWleLfs+mQvbl43pkxZ2lGOcYTsNuga7lur8SSre
J2qCf9IY31ZHbFjcqsX0XGeFq4Brid28Jzfmq3hpDue3PQutF4KoXWnf7E/HkEkNF4PxuOJEf+Kz
IJTNyqU9fBt4DlXOo6Q2Wv8xHVlc2obXPbblX9rO713A0Z+IlxNfL3yRK7W0er5pNeBEgwq0VS7/
rqNlfuKEaTln5WUUMz3JRW9NePHTJBYKaOQoVvYfwvBjFG+i4lUWAsBgPYfe8iWSgP7qT8pYuPBH
KlSXK3sw9e69XIsXsoINPS0515LhY6MqQ6fyhmETE9Ma6AFtcw86cMm4CZU0+yh4ouDhmEr43pvq
aaK4L2Z6G5Peievk5WfaTrcLxq49sBakIcp/3Uey1WnHl+CS98rerknx+EgwrypnhIvPmKBC4lDQ
4Qy9tkUYYxUSU+3Zx5wBmHoGsOwvHiQ6wjW9g4Dy7oe/KcxiHoVPsQYMB1JAwSEDlPFCNWF1LJGe
JWco3ZMypfxmITOqE1ndsYJXKYJn6xmQty5UcENEmeUZW1e1yADPvk2FrGmA1reIdUQGC6wAZluH
7T5ge43jou+XmXyu47i71j0/rQa/O41dGxPlnoOFqgupk1KC/7Vq9BG34+WaIhe5LYsxHUEhnJM7
iwYAAfusPCk6VHhzahxjWwWJlN7QBL4z81isMTMJeNsjepoWOk6bCgnKM2OzWwnzuHrOMm7/Lp0l
IQ7VsX2mqv/3981tEyKn3MKihaUkfX0MrgiHoLr+1tjrw1Plk9+PZuHbVN+7QXGeg51rz28hOmRo
GNciKYu9wQq49t1YuNbdkPI1HTlJG65yM69o2+67F0t5I1UlXj5Of7710p7zwa96LGLkymn63QEj
vOVAUYnuzr4kazvH9Ua/aGxapq5RHNiGrGUHbOZI7Co4HVfAu2PsmGoRKs46qgypMH4ez1h/PX4p
4IkP7//kJkNtBzi5DzP8nTjySZSZ9XyoG017iHndHQibRSWUiaNzi2+oWYT45s5NjFXWmpEPFStH
pHlt6h10PfCI2/s8+8j4L0z5Oa1OP7t2yDlXPnzvmr7ErVuaMAqHo3/ijZeC4LW8J8aGskMUovQE
ugxIQK53WA+Qqu0suauHCBbCYCUUtbzc2UwrB3QVLR6MsDrqJQKR+84p/uMXQ52YvF15+E0RQ/Xg
YEJWRXBmTcQ2Zrx9Cr3go989whtq7VITxF82Yan4I+yoiV4TU/e2gmL97ROSWBDqt2PvgxmNzu2M
54/5dLnSfT1Q9BVq7K9D9N5Y8cmVVFbZv2nWYhh9FfVwluh+dXiOZzLV+TWZbd+3pFQNtUU+5rZf
YLbRPvnoqmRSxYwmAFtLV9ExO6LC4oWUaQW5kzX5+rq2lLRB+cTtG7yMWWk0DsTPZ6WTNZMjkw3F
QmVFi6bEIcaZnz1MdPlxPJZi4rVdrXtGhYJ/FLSfeQDKhW3EeSCkacfynv3iDHZ/PSSMeD7A86mg
ZjfrI+6wTGweZISbL2wzxaRR151kHpxuuLmb9n7xiKEN+IFLKUI9KnmIlAdAmDqk/G7L/XawaDyg
ksk4IORBygT7AdTSFGGXCP5U4sP7HIi+xg7YrXSlhcJ5c8dBtwI7bMP85YECL/VRMOrNK9KJ9gOA
KHLUsHWusq39nE7YgU9GVYnz2jqkB4slh+fAiMus2LJOSXKD5Pu3KAt8KolCGiBfdnnLi9D+lbUz
GxQnC+ghkgPrYPGuhZapBXX2aMJl/UZSVhec4JKotGk1KgfnSdS29r0Brpz2cxcymn8WICIq9rJy
TveMcX6lM7qFBIi7uUZhPqjufZsqs36fDemeHWPRIye2RWFPbuWpHmpbkmWkUI9nBq2omnqvWcSb
bIuilXAR1cTA1ADzJIPaZ16cVZkgK7uYMnzRNX87n31oG6c6uiOUnheVYCAhKItO/c9+99Rez3o0
KKnQ2rtXofwDuUgyYdarse9sqLDnGeJZ1LXeno8Ra7nF9JcJhyJ5cRfjji4nEKc0nbjxoPDjEj1c
/PyOF2nzKPm0G3JuEJTA3KdvKnAP/r96ASbItQ48NtseSdaNMl68jk1rK/jnXQoC+c5DptXOlHH6
1csjDXTY5OJ+i6gS27Z+lJlS7HM1UW21DXaMmrr5AKoFqoljF2lKDlPdIxTF6ABchLIr4K7ZwrTI
1OIP374zvRECPaCLKxGZKlY4KvYZALl8hC/o1Wx8Qu54/elRk9SFv3TJ2poUBIbR4oAhH49NSlRU
/LZsmR0wLFhjm0koPZ5sTHghUdn7zrJmnaqMAk9in5bysMvHHgBQWXP50BmCJeuCvY/cHg/UAL0l
k/YzLS1Alk3sZ+Ya6DYjZDFai6LSZXmq4VWFeC5KUQ2yKmYHo51lNPrFdECJJwnApie66UgcxjWB
1wtEzw+EK4F8cCljVtC8T+Y5LbOVqLUwNEWr5sP9NJRwNjxWim0QN+2Xa4iIJxrIqdQFTGGAzE7R
sNRPIlnkbB8gxh5UFfjQnvwqBSPOYThOpI4hx2yX3NOsjiVA2E9Uyqx+MVhvWmtH7/tcRF79bL68
PfBODmnhSYYxpJZDCrX+Uq1xdlbiCT0aqWAmk+O2o9Rb1K4jMpehvh8zC/+th9Wd61ln3knNrNoW
XfQFHkBL2QKglWl7ljPiujKw9yZNbPQBi5IV5VrmThHhl2E5LYCxr1S7B/uOrft7eoBmlcsgkUx5
DD7PN8RP5eDl26vim6HOmf42ifkjWQ3skdwwgFq8QLiAOQbrK+xEwdb1EqJiKzrzRNvmo4bKlNtO
h3mRqAX1cLsTnJoy2kYqj1pgTT4SRElxLj0//zHefXUBsny3Kd3E9BdJ4K3eO/vWtEX7A4IkRuOO
KXTusl/XWrYdi0mnCXtSCxCYjJuLFcKWLcP3dqB3Er0TMirWX/ajGa73omRh62lh6wr1UKpTjaEF
kmx1LgjKFSIZ5SNr4ACuqX5irkvD9yCV3LBW3drr++aM29lJlFrm85dFp4g8DL+KrIebE2GQmQna
zuS9hYiK3PQv3Vofy7oaSpP5PYQFV5QnnNQ1UPvEMtICbNHWFHoVNnEIxObXSgdc0B7AyqnZvfwu
COzRoP0eoj1Jbq9uvvyDbK21vPnOgUZIdWDngK6BNxZgwRR2iCbpur3wl+97UpQefMF1dcqnMdEG
StFLp+GL5l85nGXNhPE+I6sKuSm4pB1P1cL9KIHm0WtzlVCDqKI+le4pbt/DkYxb+phveSuWwBsY
ecgf62YTTYr75Sb90YnizwvGZi5ho1FKhPAKPs8U/AwFAzv36oTkOnbJ1p2e4GGS2mMODTFY5cbl
jJVMt6TwJBTsrDV4OGOZhJeS0yfzUAhU2EfUkhQztbRKVc4qJKOi6IjzOETeSoNXBkr6mdIx2Ipp
2vwSuuptTK9QQtJhyC1igXXVuVHMgF5NclC6z1pg3uRHoLBhPUC2B1vB0Jc5hVuGFg9w/ZGQhy36
03ykYm7el9S1ru42X3JCZKnKYG/1GopACXNDtYbunupvYfK4hSOe3hkqVNEZarmAhDB7wEfEwq+E
5FHgP/llgHJL0HlaxvlC6+ZVGvMGz3cFua/xud2BB7LwIsxPgCyIjv122D+eKy0My3/cYsryGfIr
LfJ/MXsPHlk8EZmKM0Ao0sOEj9sSZ3jUW2IngH5eZa8Ldun/kIvPAmUNqnbgmEy30jMvhnD2i3xs
cUj1QcD696XT3/XGG+4aoYcqiYv68MTA8xvLTYWIJ11JxUAu2iPInpqNECXJRVDj6h9wJNnNW+z5
K8jOU/ehfFzbV/Pxqtp0OP+kbSmRNaJDGLaj1mEYG0ap2okXr19CDRiVyAq9E1TBY35tJ71I4eQv
YEHS8fSvIN9hCRYmm68YeHDWVbsgocfjVyIJ54DgXh/JL1nF1fbUaEm3q6YS2st2nuJX7LYHXsXB
PVtQuwum38wDBi9m8q8P3wGIS5jtHAnRlVJM0trpGe7HL1Z+RGJWyvk+ylQJ/jUB0c+k6cQKiPDh
F5Wc53v7T3j75KN1cBl7tzvGpZMfFP6M/MCclMHkJVIciix+L0aTQteWmC9gAdWGQlcGFaNLVGU+
caBk/bNWarpZQiwRHpGVUv+wFQcX+CLuY+tYMH6vjNllb2lRTgUp7yMH3grPS8UbZapdKt/l0x3K
dC+vc1Y06FWBBlmrw2dHj3KTQ9jtgNyE1vA74BjSaU6e1ubqdblkCdMHw5qgZ73A02SeZh/D6lNt
Q+qTfrTdtEh0H010zgN4FWvL+eECUPvNvTVHUsyKSNR3V7eNNC1dJs/ALdRDw9a12VkLJMhL5JBk
7aGPrsLBS73h8cP89VZsGhSCJYNW2gmdcSC+90qDYz6fTxs9vDYfTKUYjL2UslHuxb3brwEC0akr
fqQG9EzvD/+CFtQYZV5lMoVMOJtFsl5OINjTdYTtfYcmFzAi8araDSbQ1fWpl1yRn610wAUWE504
0mqYi6+pFRz8wEw+Rk/Qh37YlwjLB2Zq1wbr9maK2VJEqQvOvznjHuj4nwSkXLxywu7BcRlL6lEx
QpLma4pUx4Oqi6dV+EpQ1f8s120Txe+wbiIiu9foH3RktiIpPXwzjtqyI+E8fu1hJfndT4H1GELb
bziXiZG3hcBoBb2MT9kuzIACNppUPjuUwsuvPATgEKB5LPWPHsd6wy96yXRZ013fd9lby2UR7L75
aaYHWRMlLFGqmQClz86t32MFNU2l5NgcjdWz0P0e6eQ7Hv6p4Ce4n+eiFLR9UU4pcfdy2vijaQFF
yJoc9fW9d/O80bYnUCKFIVBkggMk1hjcP2XUbdQQeikAwLicWGACdy97o1aSbFoujEVaqrkTEclG
GFc+nYErs3SfXvOKDo/UQuVoR8lQBG/D/AopenrPcCy1ELBcogG64Wh+LKUMirvRbkJpvRCLF+mK
Q9S8NsKMTe/YNfSPcy9+rmophPbrbHjZOOEadjiG+4Ai3Z8klghwX7P2WxKOjfimc+xuJV50rtUn
hj0BHewNlDjPe9SMk5lLRvuSOBO6AjBY5Tb4okZQ3wdXzTkHSs6ckVV728y1uqRL3Uty+X/w4Bjm
Zmc+cQ6xEufEwPXoTBO+A3PVkwcZmgYZpqdaWiMXWnrROWz8aGhdPMHFlSgeP9HykNYVZfIcIF8e
gyKF4ariYWvMEqKlknKvUvxsmjy23ZzEyBKga8JbfmNh5DZgy4TQX/aTNWV9Ug9YlisDqniv7Zh+
4LnOEB83rFdVUuK7LYLEuKhDyvUO3oqpDsskcrwFW6a7zC0rRAHcKRmQ/fynxRE3fLvdQHkYujj2
E7uhla1/DZCxnW49UzNEsOXe02oXzE9pBxZfc0ZYlk/8gu9wdLEiGCgRxrsi8SsXOCmXeievCTXV
OfZRc44eiKLf8F1ICFx7o7/kHgtdFSUdvUfi2jSuVyVYdydLg5tNSXKQv2BQQr4PJv+46HVVplmc
AW/x4kVCho1hA15mYJ2yr40+niVav1+Sq6lYF0h1SVzqoft6YsqiVpnlK5TXT5YDxIGi5PVljJLS
ruZ6u46y0ogshRxHM+UWgnqv2RMmaX0aPEKSiODufFcC9b9oEpcjshie5vHEi8gwQyN9iyYhb0le
tl6olyyPEnBb/nyPIn7IO1esG8iEQylL4ZErKDv10sdyXGk9EVpH7oBUNjGw9ApCvo1/BK706pC4
OGrH5tMn+0b7BI9wtpKfoJUTUdqF6HVJMqjWxEqKKI3MtSeNtCx01xBvKiLKIsPvJoI9pBrjJacb
ciwWvXmO+S1CrkjOHwDM/R4jtj5qlohi9Up2q0oWjWptj7A7AqK8Ly7jWYZrcrUWryjxNn8IzrQ0
crDJ6cBH9WEka48mKRHOa1MmMvn86jPufxLswDLTLeLCmtDeJZy+W+yOCmzPQ9dHANRE3fQGL3UE
cdrO8QsCoyQO5JZV4FodIPOsNcAC4FL/daCPtOn/8KV7PA5PSjLRdubvEgvrShosSW+CUjf+KYjG
cTT7LLr7tLf2PVVp5Mq5PYk2NxpcRp354EyfZ2qAvPV3QEj5cR8rqhF1G+SfWrgU/ReBxBXQfxNG
J3MeVrjL5t2AK/ttFnsR6i6d9tl8bgPUM4HCxwPa1Q/l+ZdSUPoDtaiXr3VZotFh18ECaHfb129Q
Q65g9T8Hat+tubHJ9YzVTUJTOl1YlAUnzdgtZleyqy7MCZhf+KnoZRpzhxDpfhM7izMcXgbxknmg
xNPXUqAHldS25bbt6X7cuIepxu+LY5uxUwYFsmBV12IzvZoL50WkhNpN/8kZYHt9x4W23BxTIzCM
ZHTI6RAzO3sSFfI7BAgJ6hpTUvVT6k/vjtZweiSehKenc2UwWQ6q6If0AqhszTtEI7C7tPiDFbQK
Jmw2+9D7TWlOhG9uqYY2d7UoeYFNm77dvJsfngE2uWlM8PByP8gjSbuDHNBr0AP1kKgMtUqN3XJ2
IFcZLGAKkH4SbUklIgFFXPoo79xUxRPvGij3HBrU9tweoHKUKI0Cp7cQBLOSxa70sgOM/dkIV80y
Yl5IcblmCkuBaXkqlGPA/rx+CphmBLBf/OAVvNeESa8xza9hhweJvBDiGDg4VjnLAsF22GXNgy3X
2skoFlKipAff6L+vhe1yg7ROqRBxwx0DvqixrGDlv6EaJVXiBy3zT4FnVdwOWT3L1jEpuEqImYd0
EYPv95HGwrzInwQ8EN0vOwrrRlOR/wj8JlN3xjvXqfcriW33U0BCIixv8A9bbCIYUawxa1DBxoyL
SIiMH9+/aVeZkGVQlo5e02S4R+wnSkqSBfYPjfyhz0RwAM/tXw9IScEqtpVh5LqrzNG1M7aUnPTJ
ptlV0CLJ36ARmPK0ENIy8O/6ET2c1CRBc4WyaYdsF40T9lppSa2J7SLqXdFPDL3eQVgEogYx93Ap
EsCc+PYQh8UMXbVb4sVWXyAQ9JULhxKc+IyJiCXRagA5BhMsJv7m731chqyVuP3q9B/IlHyjBtbg
C9SDuZcyZSGkMeZOIAdQ6afqwIh04eHBL2/6fJFHVlh7TPyBmDjydCo6knb6z8hnzxJ4jhsz9VuT
U86RqKcYMqriPF5LXUglNjlN06ZmzHQgIjrXwOuf7d+SNWHcL9Or0CylrHok9ZnVmcnbrj5EX1jc
QDtop6NAWnkR6Sa9/mp6T5N4jliHMUSYrEQFBF399wEqbqxK63PkiJVXjcnptDZQz+nBXWxVGkum
7GplflUDcWkQLfqw+jN1GMt+iZJLzElU3IZ6QPCAO1+wKYiWxrjNSpo6HJnzuoy06XTcQOVZ6fC+
3C6fXXZQH92q2BEXhfNZPxZ4C3rvJIUkx4Cv2w2k+M4AaAvt3T63VRS1VUbuS3Y/DS4TSI8kLtjP
eJNcQH7JF3NsaPsHTA6y49uxdN0tKlORxTUa0aXh23qa19yda7SdJ2jejUgnaUy609E4SRaOo2GO
dS2Gro8uZ9ryhj7ts9CjZhDf1i9P5BWeKlslwaAOCN9uOE8ZVNVSZ++c2g0pLfe1LReA816v2jw9
Hm83UwjZuFv2pbJYNy8c6e1y56ZnXFvJI/pAR5JuhsdCZo7BjyB6ET4jBEO45qqLFF5UByNbPvA8
149e+vkRdKPyFVwKTyOCS/awF1s5VfXE+moKocLKAn2ZFcO1Uohm1raaMZHg+/C+INBejg+206Gd
uKLfTA4bvJBPP+a5qlfNKaKe0q6eXnvKRmjRVK1FbZMcp2xSakB8kr6O72HoJXSTHwlTGkAq5kIT
Yj8jtAFHYDOahnWH+m+ZJ7Vux+jGvMWlwkFvcne2svkp37op+mYx1+mHMwirwQdrPv8UWfxg1HDJ
7PC63KX6dR94JXmV3wOOgbbkZqUnBmYVzm1UFwVX8opTnOXlpM1DswHV85CASUq+VAstR2Eh0Zhw
djIthE6eFMTl2BQU8Cxj2ESq1JRMyzSBcr7N4uDOiANJ65meBxjYeLwBzi4gE7tQPwWer8NvoUAn
vt6bhKTNmaAYnWVY57pN9IBQrYuypMOjeOV+2zi19nvpr6IdTvuPelQhpvu3yPrnogpkVN0EukcP
2kwu9WERMnVVmUwchsn9nUv08ZXveav7LWJ8C4HgRsBNLsNtl0IwSKud8k8jc7iRYzUzYUda0WFS
eXTMV4HW6TNf2HZZ3NXHMdEZrYagz5f3qhtDjSN5syvGTVzfb4YSEqfzGEdpFoeMbk2UvsmXKGWp
0pLhAoYxn/mNnNBl5w3vQ13Q8E+ioJdnmqgy5PkPnbIlg/iVosNPKoUC2CqG7yAChY+QyECzn4ot
L+fcSQEUhBkJIh5It03LsExdzyo3iyS1p28Uf6vwXG9boHbbxAwO8IH8bOlrLoLtPEG0duVmeZUU
6lJb+2NZV2ku7NpB4cYDAstLPy5HAVmNrnRv7C2/MBY9vTM0rqkW1t/numY2v1HYDsdfRVLY5Yjs
Xg1D6cEKRhjAThUNGSYdIvznOPsNwa+Wy4fj4/SIyYFEGS/XLyQUU6PiOurVUocD1eA2PMhudpwv
QcVDpIWKCn+itkYVgdYAPsfiopqXd7UDEEZv2zQzKw7q4eZyHcB3EfQ/oTCn/oHlIdTS+9TgljsS
UcV6qoMsg9+na+hstZO0HAcSWgNZ+DKomhgMs+cvVn5vCeSkvlCuzOhUIvSm3/qME7iWKZauUabU
uOrAEktXUOGyP2S15Z87X2RZUTsD4fhwFwZ5+DO5uXJb2pnDJ1UlbtPsxE/9x4PBP3oywk0JStaB
/QeWz2Vk18gV8f8881kLv7vSrDzq6qBXjPJrIvEt7Mj775zi9lpBCjOpxzl4TpnbZWcLkQGdV0hB
KjkFcfWAlLSUEvmIXOsYl7m2yYR9WsjfiOecrGmiM5MvHsivz6utmrdxHS5yYJ+f6j5+FZIUg+i7
5KoRQTLwQhOwAzMFNon+ELoaLwM6OvCaINh+ACpWOpQavou+Ao1Zp/An5WJP0DqZIRwh9YZbC9Ra
jBVT61hVB5O1Jkf0K+fdIbmZ4ORR9s4oA+DTjW8MkwLaBP5Ufmfg8tztJOabE2mU7AYIEOEuAbfH
PLi58LDrbTm9GFRn1lF15DHJ5CDnYVZ3CAxCA5pJ+7j2QWFlGanoCBJfN1GmIGi4IlzXYu7v3She
vTa4zpgr84/nciyAHVcDqUeEwUBL874uXerI1Td2I8TlSUxmN3J7q62kps/PjmpG/VxDiDzMSGwS
pQeYHUxnLz+Aop9AIf/bwLb68Rrwzk5dDHiZS8Tj8twK4fiy8tLZ3ydKAHedfOfUeIMdVjHA0K5D
Ks7X3mPxVr++7Diu+5RqU9mINSYt9MGsU76snIF0b5HfvQwuEgHdkSsje2isLYx/72fLa22QMu/B
trQT0mie+xwvTlQRN/NeaCK8Fwztj/hpP6I5msM4R+Qz4aCGTegHzkFIycTHZqcFDDrJIR+H2Lie
zOV6uFVCQY9MPqPkeT0kMREMK58+YILKA8MUeW5Kw7lksyV+F4jUaUMD19rIv2n1qdwpP+yzrVsv
1ODfQGQ69L0amq3QPox1dL57GriUNwdBsE3JbRnidRzWkBnWihP0GOA8UBGDtHOJItxniPM2/2n6
/aGUvtk7k+IlBm0bnoldMtqjhl3MB1djA7wh9ZVGiuBVNt8DyGmChaLbgMZcE4eKdGsyZ5hUGehe
ODW8jp817t5NRErEruZund64c1hm9RLV7YqsLSDyUnQHU9IMNnUQ7361Rsf7VobgXeuviLZFEpog
/G7UJnVdV2lwNRFOY9seByTmisNVoz55jgnROFFna8oOEWjNGNxj0eaGLSU3xeT94W7j9/9frXwg
trVYj9qrno5Bvlq/CJnMmbyq7RnYxutm6tL0EvTk42jBQg/HnM8klbg0JY98e7rfkAttrPZkT7rX
e7wLeBWcZRDvSxEvj8cB9FnXdGIfE2hxjGbzmmI2C39BJvzo3GAl1QSV780bImCJSXGoEQ+fSlII
JH4qmdQu4d5nLZpoJHcfv3HOeYtEuCI11AH4tEW1VAdHE6eNMmA38Jjikugg5KpXIGb5a7xQPauY
qYs4R0hZpIbVOCHKfQg3QPmlQfvHV6IVDy/fFar4bk792OveaVtkrPbibWpef8fe+02JkwEGtCmK
Vml10h24PT5rfeGXSWFbZAqicKI06nYKEreb10yuxVj8kGjMB3g/gNRQ14MU5G34VtYrRngtQiLq
I+sA2/+C9AX1TaGxX6XK8jxgqYI50TftKFIIlqZiYV4UnuC+h25zerpeb9YZC23QBcl+vCWKDjS/
VDbn5r1V6mYAvrifZmD7brCh9lPCRrP//3gPDTXXRJj3Y4RZtmG2bV3mDGj+WpsPW8xv1chwgpBF
Ot69+9jk0OKNcNEmKCA6kAFubXFAF8Z0yCkIvk0WsAEV2/g5g2xfWJSA37CW7qVgD0MSfJY+sdnv
Pavq4p4JMiFbt9OXE5qdqKFw/a1mRCgkTq4MvlanNWHGQsaaK0VHbg9zN/MWCUIB+rQqv25pad9H
phXBgAPYdoaX/gMLFHDtNM2tZsNdg5oL+MHcM/7BnxJY4LoTOu7cxcO7pbrnRIpzOJnYijliP7Kt
Q/YKutYClonLfxJzY8QWuRJxNScHQa9B4SpI7hCdscdEXMqJTx+TUp5AC5+mjTmQToHdUBrRH7ap
P5QIu12omOJFm+ySxckq7Q6nVn7TQkADjG2wtU/L6KOSY//o2xC7zM8mUL2IbfnE+Oz/xm7+vZkH
EXdFj16lTjGngHdnqEjBElbdHgRE+vGHYoQz+HplV5J40i/5LLtREUKznvwQHcUOWONnC3VfJTKQ
jara6OaTlKwLmsbjDtuvbFOxOsEAgX7pgf9CbYYPUI0DnIfQiFo/PX2lF0oUehtyppDiaxFpVcny
8zPEOGiG/JLmzcZrQKqFWdbQkEQfKDzzdVBIN6ggDR+XaHaNHUUFtIj53amkqTdcpZ+qjTaMCheR
pcnNYUun7fAHpS4iYOVKQTGcY8RsSfDv54TR3iRh2C8wgzyEdC61Dbd//naQtvdc+a7h9/z4vnXF
oCB4rYmN7sJvwgybx7rX3mhLH7vGesXsvSU2F6EzlbxyFfgPoDlyejBRXKZwWmAvjxzTo0qd4QI5
2nexhWJWrVRqsaAFEY54NFyeMmD9Liaxqsp2dcI+KP+TyEHCkXby1bxjtr4lajAjCuaVhb3qN+jf
4jjzt5NJpAyTuOL7Ajzdw25knvEaUvoslNFohpP29IIgzCBsQEl81lkwnRCZUYb/L6NgZVkSmSVL
YQXlXJYIum/a6FAoZTdXnjQDq1aki5z+jq1U+TkkvCKjYTnIPkVe9s13GmC4CLXbu3u/o4SndTV2
V3VwBzimxOzpPE8dGtHYmqBdAicKxdyZOIo/djbErv6AozfgaVOkp1Qr1ykzclSTlX2MxNRYIVdU
M9tauph1n7XkdvnE4vFNTnRo6rNfLonAr80nYm3+AHi15JmGoedPmOxokvgxJk7ZtDfui3/TRSG4
0G1HV7HBTbdZ+olIf3h2KeEWJ2zvBo6xA31ntwF5dvRk/PzZXHXpkMi8uHVnzv7Jzd7+zMQIHami
w5cVO7aDlo+3OxwK0GBgqGh/4HWuyGxHb8KIvN/DYVaZVbr+RuSj/+DnoTJEzWoFogZU2jwOKz3T
UWFp8ZhdgE844RloxSx14G8mqknuGc64Th3KqwxURY6vMv20lczPqvfhYnLfXktoVzPK4Meh0Oaj
73jLjmVKCpv4dyAPSqjSOxKk4jLVVqXowsk46yo6TiMvXwPmzTmdsl26SMsNIiWk8YOzUVYgNuq8
OxtwLSVfFic6GiCgcPg6caicjoysCDxxGbU4sVO1dU2ef+Rye+cWejo8rDlMGScMTC/nRxADfI/v
9XsJXEyf2fZ0sjpRIR6ntyNgAJY85hYGU31+EmgnnIIQZnIy2NpwHdMooPm0mIrnIea35d4cTSkW
3+odOHMSnFqFm7qou9/P9jAoLKnTI+iPBfICn12khC+CrwdxqMVjvEpKpMeTpMH4EDRobE/Ww5l/
GHHcHVvey/4pZAwxf6AOI5ocjtRgx9lCkIce7AEfGvV+YQZ9HYZFYah50s8XPaSTYYqhzcZRbfec
0FfGgveS+3/tePC83UZdwo7Uekkb5txvhniVvUOia8CTf+4F3Pz0H+HZ6fzifSmQyaZESqWHGI/I
xUnaKB26/KkCldCuZdBV81lWB3xu6F/U2tNuq0+NuzVRFOqnHXwR40ACwKqzMdure9rMtVFTXPPt
5I8VmQEO8AhdU/qK18d9GRs9xa+AIv5medLkCTzphgv5g+/HS5Zl6MxFPPaWnlQJvprkancJk3QZ
jreIx/9PuDTw+/BFbJQEKxR1HgF9g3jZ+3b7yHoMImoVZUo2UbynRuG62EmKzO3ILgIXiUgBAWQG
B0SGSf5Hj6umZ+0Ly4gWVM7lp1iX11M9gxVXk/GVbrZoQDPwGomYAEq/fKxzHHcEQ3L/OSJV5z8C
Wht3ZBN/K7ks4TXRrHEq7AhMiXWir4YMeWy2HAZmRYk9HJUcF0qb5NAXWoppIhu3HIJZPHNB+vbj
+SuIfn8sSSyLlkl75MuNm8pQjaGaedqAt6yHmiV6pQuEBX5qgO2lnDf4GE++VeVHPEJVS5idK3nd
K2wyiQ/VMPNV3yZwlbjX41TjJEINlK1WQzITtTX22+wPM+LWJ2NsBiT987JYbZZQ3+NrawMtCUfh
yu9NU7BEERYcSwGoJVXdydTpLetu8JrKv1jJJK5TLaaRT0kEUx6+epll5xDsXCdJKTLHFnJ848a2
vUT86crWZkOZC1BFlA8FKDllTQr6voIBUfOpB8RSYld6MbtVkYFfHg5bLVtxgJwekT88o9JKjvM7
/I/2m+racX/PPEVQXs06bkQ8F2o2w9SUagwDujtUYdQhsbC1/rfkAX19wMDdeXmIBzw8zrfXdI73
oT88RBtcogw5vpRE4jEA5xNSMIxT7bbCe7V6YzA79jgNd+MOgzcFK+ywNkEDoPZmyZ2lvAx13ck9
OKpMuKZg1ntido+GD/PguahRtXYmbFZ86tlssEG2fP6aR+t3IIXUUvGKEM0YCsq43qXDCNYMmxMK
Efzpizx7k0v8YjGj/oFFSMifX0lFpz2H27c2klaEVl+rDsvA8jHx02yuJL3Q1qg1iR0HwrKbyLxG
OG/NSC0EIPeAqxR69qpaJh+PHItWw90I20W/jg1yvpD4lCFR6wj7RV0AlLH8TPKwtGvLr0ZJiaTr
GladdnPumUcpepJIAqYsSrkck/tp8sNzL2cSEfDWx5QV6zi9Fbpm62VZO1P1BgEOagPUWF+pEtA/
7b2jz3AsydSvKlX8IDWUSBwCXa7wRwvegU0TKcUqX60gJZQoO8V9nhzdmiUHrw8uYVOPKqlWJb/u
bfgj2JonX/cMvw3KDf2sxdyLQ0kbJC91zeGL0LdXmJdpm8Bc9mWaxpiwHNLsxAwSKQIA988L0l8C
Nzrn7yKbLsVKaMlUFGjfRHWsYK3Kkr78Jtk+4Cw1EMx409ifL0PsEmmQ2+GQoFLu/2bPWktTLaRI
tiC80PyMKWN8dNyBZx+56dPdUnFP1ArbSykcjv9F2xyq3O9XAqKwf7ZUetoF4DY2m3kTzu/pSQLd
g4SISd0dFSfwFFBNrgNrqER6dB90y1QKnVKUahsyvOaUi66bCV5kyTevtTY0pVO7Azwl5PMxuv/a
g6f2ouosK8bJfx6EzwXDBpbMlqFtMnvcU+/j6GKs86V6i7MODIC09RCFhrC2V5I0Hjr+fLEWfcJt
pUlQLUhi1kGyvJxatV+fk/jyM518Weoyq1uGObCCLPN5DwOg2iNBW7fVVjD5oXmE8kwVAWGA7iYJ
jLZYZMCCnxpSPuUmyjhd85aBtm7nKeCZLfAMjOe2YIyiV2tABrWVNg0p/dIsb2GLfj53en5P65GR
N4A1r9e22zK4MtErppus0COKGU/3zf76QphOCi1qOm4gLSrAVToklNXpW4J21zVyJ7f4bnT+O6TM
Ipo5+GpGO9bymjvMjofzvSnk4VP6fqo9W6HV0eOrLulDpn27w9hPcaIIH3HuxR4CqbKeqBMpQERV
x9h74q5y3Mn1CHjL0CajG7ahocunpkWS8RiBAmsmWt9DrvAWSRTi0pmLVR1aJlfujrvYspY4m6yE
zm11gho7j9yIhCiLL6bnmKxMFxaQYlTqlSzRiy6BBVlW2qgBWFPJJwr3ArzDa7EqN1iAor+AWo8E
qvHwU5M8QtNe54eepvV74+BNSiDO7wcPGFyuOHrQAI3NsXSiQ1hq7BdGdol1qhVk+JgrUU7VZZWO
b8mDEOHJGAb6vDZ+e6LykNcuXadZsAUebEIS7itma3CIyXxxk+ej0nlK2RT4RjA7lP9tZJMde+GR
1c/tlEX1rDCMGhIo/XWrAAtlSapkkw18gDSgRV4i39tkUt0T2GxSo7q5zyZTR6xfe/PRFtEViYTa
GfGb1K/vc3eug8MlpeoRzK4Dfg1qS83axITwNxU0BOOaCDqc3/sCKvqh40CbM68VLmqG/UIBeCJV
XnMcxRWIOaGdK4o6TsbBmsIiJ98Cj0cUgoxyx5MNcErVuJqEJnHC5nYL8Zr3oBC2q5N6jIbkl5MT
4SG+AC7LkYpbo/Sw4ohFCc7nzVvfCEtdYf9aqUC8IBRVBTdW8BFxbipoxuE02UX73x5XKvudlqiX
99uo88jg50F7JSF1n5VSHizvnNrl/ZooVG3WmZZJF4RCbNvjwEZd9+GQohdSQ81oGIpoi8peIGyC
nwBXvHgZ5lL173eA3xgMjhPEgojcOPbncJ1Pj3LNgUd76wXVAMx1004Ku+jD8sL0sD8Fd4jO+UPo
rlD8XARb2rR7218AFRAUPg73z831SHUmX7eWND3WSMmplwRJzzZWxpFSoKyaPqoNfhUErzKgW8BI
akBk6IRP3YNdbFjnBMKa5sA62Cl1RKAsfIuwea4tnEoaPS1RELwZaZomImSSI6vLw0ColGrVwgBa
foLCOEyubv/wXfC0huO8fStiDMJYriEzhcXeFc264S82VcIIQXra7aYildD6nS8wNNwWDxk8AlQq
83ujcVdUxInK7hOgr2INTJSUkf2DAkx3PuZcqvKFa/v/3i4Aq8LOGey8MniFxQFqYXLTBeglid7Y
FWgMjWuELC+ieB/M+JpC9p71pFmVZm0vUOd1mmyzh3ujhfl9R3s5gnT+zJp17JslxGnTSIRqIjDV
Go/ldKVNiG/R4mO2cU92jN71U63CkPRVKl7YQP277miPtovi62hHkqCIQza3VPDqJoOoX94usp8L
g9KRd7TaDKCfOsmSvTUxuK7nmGyteDo5nj77JBtKdNWlwOk0dAa05KAERyNY9177wqa/lVYZM7Yn
6VrKSG5tUZRoSsEKfOcU4yS4Lb86S4N2wAsB3YZNxhkRnazhB8LOOe/Wl3cnewta6+uyxxNN3jVz
Hr6q5EkQ8htHmSl64g9hY8mlpnVqZ9KK1IDfJ35Mu3wv7x4ywjDuK6DObUItIsY/KzeCZvDgIMkI
CdX8J+hph8qrO2HUj1tN00oWdrK82T68sux6Vxd/2AAzl3pw5+S7ztgBjH+OmezmktDZzBRVrGIQ
KgPAyFk1rLDlqHfKdsi7A69+uV2kgJOYQ3rD5M0YFa139M/9RMzbOQ3TRZsPZOOL73K+bNZQ5DEy
wvdYEBIcrTRmW5hjKXum4TFQA5Y4URZghNROIyqrG3MHgrqBNkATTHQGjYtkb/WWNhLEllwsB1hE
wkdrOntKzRDiKkEQp6siNmg3Tn+09rOpgcIO83GeH1gwpGA4C8DMyCkHb8MYm1otsqt1yYIbYCo6
jpRoa49c8GDkV/EKKWMFiEBOnchd9O8549mXPNcwhPfvVtgl79RRhPyVQ/IQyFeYjSwE+etCP9Z0
PMsaEJ8RwentQNVVX8KmQUAiol9saXEsOHChFgSA3V4oTyihogsmLUCP6H0tgOpwlSZZuo990RES
mmEheS2oryIWjuK6R1Z14zgufIx9tWtbm+Zn4IFhMdtCA/2bvRZG5t8ch3medWbaeIEgF/TCpCUv
ZJGHqasamaZ0vVzbZtPjIMzQNIQxQrv1Ml3nq4ePCYPYqnH5bqa4j//83+g8B3RFN6LqZu5+2+x9
YDtskNtvGlxpdYspxsgqeTRfWSLCsFfYs5FH3AAp9+i9VT+gysPEolyBBZGmurv/NKqEmD9dzhIQ
iRzM+3WlCTGdkf+GO30tUyw78LzKJWC5Ilw1RCTN0EUe8ObG55gGu0xyMbOTaZhFgUVJ1fB0970X
6Qu/4HJCJwvwiyOcX0CJQZ6vVvEA4IqHAW1UP+DXeutyJPm72Ml1cmW27WATkgzdBzoDxsFIGR+J
8SpsGPP26OWI7JNuPLT+PTQQ/AiEi02t07qZ6UW00PGEt9Z2+EAG5VjDkXcOfEjkay+3CVrqyT++
8CpOht2tyeTluS9iAq/ovBttg7STVYADnQ4HqygFvPUC97PstdV+xb0Jrv+11NW3MHkoVV3uW91+
UbeuWvk2rPUFRNQPoUiv2UGyt4L6w/Ju5N7fQYMbM2JlJCPtz/Pn47JM+cbRLosoWCHhLe6JUPx1
cSFzn7HrOVdHFaNyvXKf5jfU6CaPoA8pf/5e4iIEAEo1E8XSic7Ft7jljTV3LEnlXSvDBfGRmzhV
l29svn5443lMvV5mKZUCD8qh+tXVXNua7n4dhWI3Ei5N4pFtMWrm2OLxL0GSXrr2/F5k0wtjvNJU
BINeDj5cPvS+kmBk2vK/rUlWs9rQP5daHMjc8aWcVFilz+BseGXp/A36g8y9CTplwmRDeEZnWqBI
v8bo++MjqAQjlz4tw+MwFX+9COyM7NsiQVcyBEBjp43MRynBq+RrNpQPCRVCP8k+Dx82ox6RxOGI
bDxvivha/OGk7ftlBvzpk+EVrbakCTjD4Kl0z53JWZOpdmCi7NK4tgIEkFeC8dgKVg3sSWq+5/Yi
hi5Tiynz+2aCFX2qbXZz+NUWadcYeEoqlWx/NpLWh7Eu9D51RDqGQyBtbqL90ROylmEC4h2Hzguk
ZwDNfzNq+EXa6bzQ0eHqWQVpmBF4TdsLbzuMgtVYxkmRHTYHlR1ZGQgejA9PD8WC1L84sD2A75S/
Kp1nu6jcNhX5ZODUO9a1iHGImhSJu55X7YmN3SaSlwWC4f/DceEGvHyipJa99p3BHqCwjReJXpGW
gnm/nYXOGfOHwUA8FQYoxzYyUMhygETWgG1ULNrs7qZL4ajOTQthd9bGkD0CrlvAIfD4i2+xR3z0
HiM0hccFsK5q3upIx+3UnlU7dAFQwQ10sIeXkno/8zCaCrfii6Pt59Ehu+NgZHo7959OczqYh0ot
i6qH+uFiayRxOQd5DiKBu0pr1hZ3UyQJuxiiiSChtWkRfUYgEGVQC0gDXhs3w8aRTucGcWNEcXLS
ivk2bqEI6OQT1JHUCdIHqEXYBAnoWPV72BdiEZ6nqqvP5c2oEgzrrT3H+y+TPCkF5CWWQJlVWZrT
msd+3bucV4D6p3GGV2aIBsk3H0j55Sw3D9geQveHi7Ae89ZWUynNFwZNlGq0Om3nWJXptpbZGsyX
sOd51WTDrJ6IKCe1/swjB1ravd6vlrbQ1pX3j0hQsy0kXqvCZzgT2AyoBeqfhZNr4yEm89QLyFEE
hPN0ds7BQDvPGBAxtzwaDRuMnP0UU+i4c/GnmLtyyuawrycyb7eqC8POgF1WYB4KB3yWoXjK5zJ+
w8Yrs/CeBz8sqCFueg1hqjdtbOBNsww8ConAW39DeXdh1Svm4F/Bsh1KCyse3Pl7AdY8dhTuFw5o
ewe6Zk1a9lyTh/zwOw+cr9yBhzIZ9NKqEKN2RXbJGe5jw2CzlgGoLr008pav94Ev169mIEJ2VLCA
NZwAJrVWRNAjZ/SNxMDq9rOapH3iql+Mu/fo9R1z9m4lp0ClHdebvlp+R8lI/Vh0AnP5AHz7ubzw
E+VP6YyT4BWP+8hDezVPd5uWisbYBz4agBApPVQb9t+QyxCD8H2FF8HxxyUUvQFmCI/Xd7sLnyj9
W289Nj8RX3PnLzEi4LyqRWyHPTcd2BNiUobzYn+HQdOBi52SpNxJrvrBwNlzQAjXNS8VBPLO3ma3
J+M/AtnihyoNBEv4cuSFcVw48CtozTIQmQk5oARlM6DZUhfvDaE+cS0IMlQ3hk4jMFR5NeZjSXJ/
cB+ZCNT+BN5sxY/cCTG2CYdliGMITlN1qzXHSQPs5Q5yyD4nNYd2zlIZmAQ31Xnrn7F/pV2oxQhg
ic40+B1T9IbMMCdeyvubWyuVCPykgnFvsOHb//ny3qgU/1fs9L4yRvaRqrgju3t9UdFCNLw2CjHF
g5iVdS7zEeC79auz2NrHd06sJvqCRRgNa/aGf2kUnZDKnvJ+k3fXjQ+OkLAAIMVbC0PqEyiuryOS
nWg+uIpvN2xn/vdGLEu9VvFrnBtGu9nyP3gZ86NOJ/PGKZ4GEJJN52MfbXIEDqGD9LeTGohLRRdq
mZftKTdJFoLM/NTnSBeT3QRpr+oZzfTJ9iUgYQoSOZ7XDc8oOHOf7cPyF5hMiP+mNbXD6vagHY5Z
hKs3WQ5xA/iZNt2TKFqMW17d8I1zOvJng2Kw9IYqkxEybrNhqvbioBdJ+pVeVLgTvf54irTcKHpY
9mfPbFLa9HK1avLcEO19VGSiEN/n4JVDVgyhYZFyijGx/ioXXWjxDieX+ukSwC6n4J31MsD1+b91
irLY9NmWd2Ca42cMp8O7Y0LU0MO62oiltv7aH9h5IXJbCgDFRL/vgHW7OmatEV27degqOG2kR3By
8I6n8BXiFVwVS3eU2TtUyVXV0T9ycVeorJV3Wf0s+p0CcMgH4NoN/f2yDyUnpGEJtJKpf5Q+zjRu
a0kDSne0+BNbnGsLt52A04tlV8rIfnm7Fb47w00vtKWRfRQQMO7APmzQzS7yHiN3JnKiIJ/bDjQH
JsX5mSGAj3XG/tbR8Eplq75tq9iPhmmO5Jn/mmJn2kaTvSIwibT1KngORBo3HkCqz9sVt/30XcUh
dfzrATfS4XrWHFougSjPHM8rpm5yppw+OZNlM2bJZYyQStCSMFx112nBlkdL4Ys8BPeeN7ulM28J
UJiWrtmwkjqQ/sp+Td/HV5kW9mDwkyNkVmi/3t6taIUOLnDGe1tV99uLDvXTF0DofxnBtmdvnkPq
PqfCv/e5W3TU/PF6rnmur5jrcejrU3Af9MCZxddeGJoqRdmh+YLZY5y3h7YBC14R9ErOmkviN/bx
LIrYFinTspYrMAbwJMewR1wG2847C7hFthEQTxXlvZ36YziYIVcVoXfCPJ49t+/yRlVcHjAt/tao
gaAegNSFLo9xD+AyMM2RV4FMJnjY1/znwZ4Q+AZ0g3xr6TV2X24dLCWsj5d8Y4rmxQbGIcNGUDvk
mwNP4Z+EHbJrOxUkoOd64SsLsmOKDTre8MvnURZt++ryLKJ6UtaHVnEXXcS9NgJDtThIe2PMzMVG
z0Ojt/xWipSZPwMsqvs7pVfpVMgUecFOtHcb8ZmCIKoqCpzaQYYAu4Y4i0zR+djiZYRQbgC9/LIM
47zqSDses4FbW3d+3vQP+ZOrcGeG90iA4zeXqCm9r15FdhAQDCcWvQnj3Yy5IY5wBX+2uqUnma7F
3rQTC0Sef51OGEgpyiWNn3Z8WGWpLDvKwPl5kP/R4AN/1/+aG3JEdQ5gGBUs4h0O0DH9z7UIMT3Q
xpkW0fDIJxJQQD7HyrQPUGkl3QkZ7uAmvCTW/2TFWaqiGJgJ4w2zsKCYL2O4T516CzqihRBggnrt
TFn5V5kr9p/oJT/wD0xTeSis3Sj7eDG4sfWXdc4aWvA038vuYhFaImxj1qtpPyn+D8kcoQK3ueJu
Vn7cIDztIBS1V0jNKcG7HDVkMs+2mt9Bd8eohnKNPZS0m7BXS2UlnQV0ctQKPE8OXwl3o/m6dtne
VYjiqU8PEwHWBiuHreJKCYrqBEg0DqALb96LtYJCTmrcRyZ/rLSMD6OBkq7nJz2EmBf4rkZunvtR
ibDNIFFI7m++zhVTjXtihnCa6CXmc7lkjlyagv6Eoy6k8Ohih8LKex/g1ZzjVpzZjWqosXts0Tcc
V27UoUwo6KeqRoWlkRiVqZxS0cdU/rUHntvSXw/o+L+DjloeTQMa/HzOfeZHsHa5VvVVwbm6KF68
Yv1cb3AoI9YGkHtBq+A9shu47d9SfOvomtZXbKW1UQTjc2T5YLAszSQ+CBEDh4niMkpTiBO7JRKf
cBUW1LoQ+gvdam4j775lPS/K5IS71Gf9d0RTBeVwHmz7X1NJXXqcgCP39w5Ad5ZdVCw05GVFT67/
BQ6miLQJKKnHmCbAfEM5LQ2dT8SlxvawiLnX0GcYKBHKjDaLP+8W4Sm1babXwF5ybfSMHmjCaEzk
zbxARaHaXGZlQeYWvu0lrsqvdC0qb7ooLiBShVMO4dsgV7ghLmOH0bu9DnSQ8mKshbNGqLpLdh7+
4KwsCAT01j/He1LJd/UpxRzbse/MBxaMd86oahHfrfgDXz7x3NuUlLNR4jRJVX8sHSCy2UVptaQE
cWPbW+xDn/m1FMfQyU9I5CRRHOklNH0171JG2W0UaYyg3WwDh7uutzulyOMDiJfKq1wR4q2LSjFP
d7IozYFdtMFGaccVt54tyOXq9nveBWrikXYmOHQkyeCbFpr7q/Bnf0ngNWUTL9PcgBOgFOaftBNc
FvmtkBavSFIQ2oyinOhS3nDXT2jNUmEPjPyJSu3bm714Yoe+KEzd8SUNitasFt4KRVcr53so8nIz
yFzGW6CNGra+itQyfFcHokoAwdLpUlf7XmwZGAMq6M39nWRfpOuXWKTUXrlbK7C/8SHYySavIpSM
CoNT8CeYLo2EOvUKd+twL9OkSBZvWVrJ4Xl49FUgLUnnJJV86vim2fFTXphmmbswkCzTFQaF7cUA
ffBuLj9gI7Y8cMfbreo/xX8aZ/iX4JZhdcogvcU0uLdNoe7UCBB9DYv7yaNco57KJ4IK9ff3hSNK
KL4lyOdyguDjDdKOOmVER8QewZ2gssRNY0yDAbgEcz3ej1aQLRIsTElsnMzjpBjqmWJgJVU0vFoi
fqG1CzhjrJvS/aAB33QIecUPoSw4/cDqiHYlVvQcvrnCVY7uDrCcIfnao+KtzH5HjcASz1mvhjgJ
bRN1zsqpmJcbKLgRSCyfVg0OpOrevgjPOes/dg7EW6zVpWPFr25m2qQZ6Dh0wi7rxyXDFv1LQI3o
1y5AkPtIPzRK/lMjOHNicKvtYqOUHjQn0zd6ckvrGIkRNJYz4mrneLMkwhaVtWJi8Cdmm+nWHbx9
MwiN24sshK4UtWk0XtV9Bu5bheLDU8z6GZ2oMVhpTyZhZaHoGhwEgQMk+B7SSFiprrUds8PN1P1F
9/Ku3MwJbuxZXpymYpSFt2987W6/ij0tEMez6b9MzwGRTFWbVATI2SY4PFXmOTzmZ1FwXNTdvQer
Bai/mnerNwJ0lk8mclQI3MB/TSNhAlCqS2zgSXGCbqsd13S/BgvM5twd+lboB25dYvIf3A71IWk4
vmchkK96r1IYRVJGPk38h0cnySV4/IzC+y1Mh5j5fq8AP7LeFr7zy1cWGMyY32j910HQCiH5ML5T
gcLm69vuh2UWGNRucXELuUgFBdqBcvGDnysvQJsyUNMGMDsH5rZOrh1ax3qEHUz6rrtluPeG8oYU
yS7ZM2z5/Gp06QSXCbWKF93Hby7BPlKtcc1KwTDh3mCi8Q8NepLyA8wEuOHiSocMjAOU4u22zfbX
rWPKQuB3MBbKcHeNNiZJWaFHm/m5mHHdnpwFeAG2SwuEK07VIHAAbzpme1B99UnfUWOaXTShpU/M
sbK9VApJSEBbqJmqmgy1ddWaFboCDYDjVU8PHfHzRWWMbQyMu6M7GD9HNy4lAEZcjtYyHSxyOA4Z
dt5rHm8wextjrbDks8U6GDJyOBMhHxF5X/wuGIMDdOcZd0wI38FpKSVMhKxXHvJ4F8MYDPps99XE
FlpXV73WvjIeLJILReI6i2aiCLpcpXUfj4wKB2IN7OkVGtyfM4AlR01nnMuKNUALeGlo2Ethv/rE
VydadlCdktNKsPk/LlfztdeZJQZul5EqR4E4a/izYfyy18FM9xbfKR3KapZs562KGRAvoMHDSj9g
y4uR5z1/mSudZVFVw5jMan1qEW0SBSi0bxkPPek8oix0zGSPctLQCdlwUJDVXVaf6XJ0ZR6FkvWF
++Yx1NTUIbRxVeiw5LQD7zIlArAd+tZXD42arPJ0qADXQ+ZZS03pKPxRAfYsFs4sEFI+TrGrLGww
q3tdxnjCN9wwXMciAbZq3SAPTxaSkjxoKmJaeLIcTgTmmOfgkh5gfLk1MVlH+/6EuDMaICxqbIPj
wk5c15mSVz4BK4WZkPKR7L1nN8Pqfv5mCnB3K4gxpw8ihTtEINj6Z49w6YCfY2/7dpIrTlNpF6Vr
+srxXwnWSg0Seq8bPuml88jcih9AyachxLCb/GiyDwkDT4rNesCnGYGKLeYmPYfeXisyrMzNGCLi
ka4c6W0oSiLlF7pc5NjDzj2m6UACKtek7HUxkPXPxwDE9vPPrUdGceSCVFJjHHfm5K9YGuPgXrIF
Dhg764Im5yjx19Ih2nSO4a1muPY8043jvLQp3Q9aWitIe++HxMp22laADgQQOgvXuxyw4QDmMe2+
IvJgN0RYcAZBuZ1ITh2D2uRuG8jNd1w3XS8krTDMQzBfUgUgPHHZWXZ+mCisK/uDEE9vhMPUe/iP
OWeB8boa9Nk1zfL7eMp+2+SFuQ5+YwimiD9ILBuT6K5A4igSP/QnbwriQQvaPs8TbsvZrqNvtidS
tbkIb6p9vSXN/YsmCyRrPyRrtWmzMKsMlhOGgAvCqdOJ2EjPH3ejVAm/+Nrf0pO7d5J+JUrIxo8L
k/q9+bnNfXPOrSqHWvTYTPgj8Ltach9w9fpfbkvWOx9CTMghoHpym5XhQEzyBNrNFd9WrUG1JDhu
whdJE8hHSFn4ACSIxEd+7BY5eEmd+R3OcXWK6BuWwRJRGkCuIaiFZwauIsadChlUH2vPus/PBKeC
CX3YuIISIyldsXpZgIoYPWhIbZSdAc7KnK5pnOTPRCqDdyAcJFkQm9/QDuHefzkBIdOLM92h71nI
C1atao6d8wSewdbKt/4zdkN0xjjta646RXEPDeIzAmZK8RJadyVKDVXZ3TVYl4cZQq6+g38kzvH3
aj7kxojlNFLj+WhlAVldwxmIwB8IvWqQGfksd/FDrzvLOwO6U29RHP0QnC0kZ2DuwTB/bW03TDVA
ylHOfVeLYrfZ6Cc1+OnHCQtL1+RnmwBHqvWkUyLx0GI5LlvwLnvtgBFIYH67063FBkNzF4yNx76W
BkcKoKY1LTh5S+kAis77ApQ2YcLG41Q1RUbzUobTh5yNhXmDdnMPRW69dDJVHKafCc/cGR7LWUlg
GLa4NF+K0t8CK+Gfo2KBXv2I9bm9S9+Q1vzuSFmyKEPRtYD5BqSkF6QL/OctsAKFKjWTM0yjW/QD
EVBTku0uiyk0MmHVRXliWfWwg2OmONNsxdy+NJ//EQL6JGbiKln9LByVzeuHXChtLRRCOwen3uCM
GCD6vcHGsblVhLjIq/kFEwbGDtB10q/+mNDA4cvO/AtHAb2yiKcEfkcO9zExcCrn33gn9M7TWaqV
M46/xqhYNbRJX1FiRpnqoNxREGNnMbOqOQr7TO3rTfQ9Q65PS6gSpkndZNakpgbHS7cSB5NKm4mj
5kzGnrUIcBDD9unYPOFiyIXyBZ2VzyVrXCl8A9dRo8fmhxddsk9um2HHGwKJPNvgW1dUKcCq1qkx
6LeiQmZY/qxGgkE23HT7D++WpiW6OGpEYvQNPmULXhpDY1KlSvfD3PgKTpVipVAbSmAO8AgWHZc2
D/Wsv3Zi8rZ9M6ltghxGjMJ4jxbSgxixNv0Cgkl8x4A8IGb9HY7YAhg3kV7LOm2N/Lqsxc+x3kVr
DNugo8hF7Wd1rEhhUjKRXIqT9GpgiUy5BRbiYnkU1D6SoqAMwiWc+KuU5/sZG8CXiLwP0o3AzNgW
WPpib5fMkC3A6EEMMF6+/SQpYJSV6ABt72eR1i0/NDKmLkx60S0sj197o3r0Ow1SX+dXSgYa7kV3
UbIBdTdTR10NsbdRgEd5o7qygaDE+m99ZNY0eOo9vFvWTsuvL8H/DU/g7vw/JvEOROZ/jRA2PwiN
vGI7wX2tdJi9PFGC4yCBLgfK7ihOoYWzDXR9dDKslWT5jLi6bkMzVMCjyZPIKWGh47oat3vRRHSD
QlWdvGKMn/E223cy0FHAgHJ2ZpAaLclAE2dTE5kv2JFVQCHE24z9osLT10Md6x0or3bhF451yG7w
URnxbNR8RlddkwniyuxJzHa/VUj2E8nLeIfT0fOXDW5F/iAC7hD4/RZ+lPU2/KU2pZ/kukk2B1ui
F8XA4aMRVnct/kM5K96GWJJ63L5XeUWT3Eq8LaEdZs/lGwWF2q94OWjhTJFaaQCywRiSylY3Jznx
IzCl7ky4/XoPd15tYcFVK4N9NCCJ0+kvhBs1RpUwc0DvCDoxqNpoKDBJXTjasp7jhRnvRMqmB+KV
Sn2ePVRWA8v4Y1ZdLMgAWjNM2SbveHu1HqvaYmq/XL5+8HeyRRcvl+OBKpxf5YNHL5eSJA1V3syj
JNJx3jZGbu/4hgtizGuESj7NGHqtPtkx8l3SqE3biqz6Sb47sPxA3wkhemUjcbLU58jAYyGoQJnJ
ce7EArNyJtCC+PDVx48mriGZ9QhgIRVoqx/uW8D8agi7Qkt1B/jO86EJne7Zde+vOAHM7IkxB7qy
nhiV2gztWNpVZSJKvwtkoXtoG5KdKNnAVCBkvHTvHAbcNFVwakk/6eKNGZxOOdku9q68dBYoI+TY
fA1Rcmh8HXGNON2Y/evC88243E+IDBnskrpe9DSYrO/tN674X90fYjqaa8p2MXHDkXnKrprkmrSj
ipEeXs9Vcu4AikTlT1LFij3ydquJg4RMRGEs12Md4A2f1ubKy07nnCyyrpWHZQFDbzcK5MjXqSFL
ItZW4ecB15+OIr8B2EP6l+e0oq811mjaQjU40E13+RTeDDnkjDE1qMcQ1WbjRhmAYK1DQF/y/3Bz
x/ztoesL5I5nBaD3NBcYvvd4/vduf9SYuwKTLtePCeyq8vjXS/YThzXgoycDa5cc+0yBuuxqRG9C
uuHh7SxE3TQqZXKGOyiPXpTz3CpGebg96GWTU7m1P/X2K2QJ24KNXm48ULFzldSF6nj/qe8NL70K
rrpg1n6BtvN+06M0fV5UZiJkTDI7PBo4IVBnAMP7M1sT5Tor2znBGnyMWNsyuCh3BDuIQ4b8CaF1
D4Wpy8W9nH9LqCpvYiSdpVxWcIEdrwR2yoYFFiDUllMsU8M3yQAJ3SN1HAMmk7ZuVLlrDdOYvKqQ
9VzQYYht0YfOz+/rnEVJILXMn/unuHmU7DzphvFPjWLPx7PpCVvBrk/RwXEz7g9l6uyr5Jv6Dy0x
aaw9R7uxs9tK2q3ZS74dT5w/OC9kQJXbyftR1Gv/Z8bCJvsyIHZM8IzN99by/TTWURWXaW4ILARJ
M1rCECa68dU8LIlZpEfYsAKiwLWh8AQZ9cl1uLgVjdpoAh0bL7pdbtIfHSx4OyNpG4H1+wKAs0kF
IRtIrc7/cVCaY8dp+xTVIZRDiw69paFuj1ItXWEgTeOij9y0vZH4iftsLiHI0OGjEnkDC+tXCvhh
tQGild8Gmh7ePMOgsgI6R+IzMUMoQxhYhqEUiNVpL+uGWiXwpRPFkU5rLSRHyzsNJPemanUzJJXZ
+02cWSGruba67hdk2W4E+h8oaXzevyZfIJma6sB1grcFAzSjN/34Cof5aaGErKu7xda6Ohwur/Q0
8ZoDFASGASn59QtrwBgYCirkQCZIlpxqWVouEtIFHqOlhrdMP0vf7VFm7AZlkFrNN6vRr3gJzZbI
uUEVA1oEiyBcsvflFYmK4e158VRsVuiMbCwxY8c/DSUa/lnl5CvPxKYIBNmTHnr/37W0S0AfUpSQ
TSAIbCZXOREa0znA26JRoUNFsAVz6lDmUO2CDcs6rBZ8gjVpjWEmuy7tm9x5aknJnslV+qdOxYst
3vD1Pcuw7DHvSgyim70gukmvjhkMOwJ9wzEJUGSCndpH/vkzIMTYLja4lejxdcaKs13lpiyOsiEC
hlr07AAB8gq4gHAsDbVrxKzi+5oI2p0QiR664qzT3bM278HVRz6ZLL8jMGAjlPa3Ypbi9y3P0Qt+
CVg/mpJ/dTxHXB4UzxcIA/jEGix4j/DtV4v23EouEPNZ8WwMnzaxWeJNXQkU8/lSN8ein9y2X5RI
LRw59FqrHQ3eNIn+he0hGagEBMYroLdlc86QynJrdGSxiRdVwU6R38BZ09S/l33wktjtpWX+Dk2b
+i+cVAJsUiS8fnSAu89fvMuGkyGCT3RZC4hWueuEwEVI6PmQa91KJVmzKqULHkEy9k51IRqaIUme
vsTkJEZAmzwcGxvsf/K0yjgBrIoC3veZ/mR1YuPQFRpjwyoAcejmqSwL0u2UnAlaYnh+ZNsSz4w2
o34rIkIJCs4vEcHdUVlkITTsqQPqvXHd+GFn1ZCNUoe7AqWMqr5f34RZqknPYSFDgTziQjoEWtz1
ZvUKhaHf81CwMUImwI2F1w1DS2sg/aiTVlZCzwe0r4Bxeg+NVRdGtum1N36Qy0YGTIjT+6gZs+j9
EQQ69Y8ZMy+yamra4iI7uN1RIUk4T0AdnhGAgJJTbQzEfjG3981otlr7Qy0weGKSFwozhrk44ZdP
30p9E9WmyOvqCban4rkVci3gJovdjT7Zur7HJep33rt4pZU6/GKdKP+zVBHXJksndYGBLYBHbbbC
nIsKYwkWG4RP9DO6K8SUzhYhUzogMIifhq565fWge7vdL3N+S/Mhc0VSt/TRwYPyWrwUOCzfTeRK
4LETMjNRomxvFmW9NUULvpjpYUntxkVUBF1ZmPEP2bJ2xRyFBEtOV6Cky36Mg2zaeK+gHQwQhqb5
Ggizf94+jUjY0H/IPfCjpGdOave6oip6YzIRgT4Ycs0sXSFI/gY2cULeP9hzN2wScQkr+1nddzu2
PaDfk8pEqn5Rk9Wtzt5bie9ihQVVJijas5xMa1dUX28l2gYbpyKy3Usr6hLFk44UJZM+dg8RseVK
hsRvY2H38cmfh71VzhxTKkY1zAxwyW+s6attjubK7gJpbvHjvlNtYIiBM4a5u+h7JiLR2y6aW2v+
/e9nm8QMysILWUtms8WweOZ+VQPAUDkUZXG5w6B6yx4qcZb/4NVF9LPfXfpj9xN51H7pAn1Nd9Tf
ehlsLaBkKfNtTeHXqrwhqAme+vpnXLzi+2ZWkmzM6vI6k90G9srFwkfL1SSi6XLbEq3C8Ja0TZLl
3BpO5owLv86u+1j+qOEMnje3ST1fWJSYHBR1Aii+i0ZR9+L8AccHj2DgJoABbym65S5a2oKPwX1R
aJTAeV1UNM+pKWWsEz4TKMPs6taF3nElmaN4tZ/Oh4RqpB+wdthnLgzY3em+eUDwTPTkSXhgIYPd
jYAMadITtOri1eNb9uaUss+Ts/5yzRi3pLQJboi33btFRT6ZpBVXAFEWOx8bPU/1D2qQEwFdcdNI
CcVGXGYLQncnf6iCqST/cVFgSosG0U6Z6rvrEvRmog3GxAIO5tn6UjAHxHFzkwt3iPBV3UZ7KBxR
3E4O7O5LkgVIwuQhqvjKhydYe5fkH5JmBFREmYw8d7LOQLWuF2zfrPoMEFjdOm59XoRESLaaMs9P
11QqHR8eVhSCiu/MuzAECTgdL/+3lFqo0iWzaIqp3Rg9anwMFmKe8+xQeo6kMIMXCHx2F7m08uDR
GcF3dPdgKXpyDw/ThBDmj5wJhhcCFwHRn5m+V88GSe7NbgL3T1sIfEgixU7U+fuRJy9Q34DOzvhz
0OajN5mtZ2odRGKmmkTkvoR13inPUxmi/qonljtTiSa6zKNZW1pQCigoH/iL7Wx6XjMcCtosbDu6
pja84DxlASyazPDbSUxZWvxycIXGDnbK4fZopnb4khHqQHXVvY94xlVIZBegDRfGKDdIUqKu99MZ
19usKeNkJrlMlN62KcFoSUybC/cB5sQXHxuuw8lkXmu0/Cz35NmGqKO3XPHHxOMtKDO7wtc1/6sv
iSbta0yJbLRGHf9IpZE6Ayp0c1KnTre3wSFN08AfTb/zy6QFxMULIQU/5iFQWD+701DRm4JpVoPE
MnKFXtEXsLx48mV/mdCjVxFeh/gMgys8HZh3gnqfYIoqpEsHG4ejbHJo69sVYUHBYo7in/CgG5M/
J2YBgVJEj/0AMR8w0yoYOQkCWlXERAJiIWkIK80y54/wqEG7ypkEaRb4+B2uCqLlImdm2hnQqMuY
tgsoxzuH2lkDFwH4iyj7ntbPyECVljkNmTOBjEsGo0gYmLfBaEF/FDUerw6KEWLstHAdunIetOHE
6GouneSrQRLB2qx177mZ6DPTehaZPzEBvzPv4xS0SGNbeFX5kptp5G0Xh+4YuF2r9knYCNJpfEit
Zwnteyxsklqe+DzihBsSvN0/wb98E0Oc4omsz1pXdpXM3LELelIXSybrCokKeJ6TV/UqKOXYPkoi
Y/te04a6GetjPPAchmI8O6HBPuqKGVOjTj0/JHnIrFPVJBDPISRYq4WdxiRpE+a5PrydnPefVti8
QPdJ8L94RThfuynwYuhVXtYqgJ6Ax4k2BSWZXJvIZFQi6hJjCds9bApPQDBFf+1NKGE3Z9/Qhogy
OV7M99OaXcWpIAKw/AApqwkMXlz4tDsDIBHe8/20FjjALGhv0f60tAI+j0CQhFeMDm48/n8m+hZ9
gBvcBUEgdJC8WqDf258pJxD+8AEFS5MPFAc73FgnocQDCIjyxhx8dFbuBwJyfeTrJKUk9/sbm6mK
Fm6fFHIfAadr4zVuXSKQ2S8uJUnF/2xwQIuUwihbBV2Gsf1E6E5pqrs05wTOvwKHG7sp2ZSrf/Zz
M1HbvSTLcKug8umV9Io2ZYiYqHk1mBcH78klxISdLmZwiEZiG3SVElWAFt0IjUms4s6V8ugfHUvb
gJEXSmRpJgsgbZrtERurnVMusvmCNOfF2HevdnNhLEhQcpK3D04WIgX7pFlad7zdPeQvzKrAK7lY
NkH1yOByEVmu1gH6CEbeQeUMoZUXenwvcWbpQCnjK8cgdtwy0j8PgOWY2DKWWA0M6wNNNkpXw4js
fnem2c8pEGok7wcH7VUC7qy01tTUpiy71NUZwzCOW5k4Zl7mbOnyik01tgxJqcDe1impys7RrgYY
eHWb78SHfcIxUBGdNTXmXJRkx2cC8qmf1PS+kacp0NNkAsZNc70LRzpNaCSrbRjrbeim5lWbBfJC
j8S/unqOoeDpPUmBlwIkVEk8YMTAP6WnzAewL1ee+cpJ27C4fCWgPddU+TOkP4A7tQKJD6EvJNrz
6Czkx79adXxr5QqDDIOUUoypkLOZJZZwySyrpLTPaCj3FFBf/fW0naI96ddvUDTfOBPzVKHcct+v
swR6hPzmVX3eYduYhWG6m4bYh8nvaXc0VghLddYxhhsPTCQCtVBRhcLIwKa3jZm1TD1/XAutZuNg
Z7X4CnEJzIUguUwjsXFQF/Z3geSt5dDJywfWSa8b5sx5M80LkDJapU/d3EVy7iRpoqrruU5akHw1
EQ1wxrcVRCGTnC3jjQ+iEUaNyTU8sG7xdlje5CVsMnTn0WiYoC01OfKTFCu6YZWep2LEM3PNVJDr
9bXx+E4SmOLd9xMZ6H87lFzVAr3YKfj9BopJN+eGvTze0R/r+N4O7KwP8VOxoChWlqAVtHsEKjsJ
Ksj20cDd92D0fBAdwP3eAnYZ4pNOAGXndKMBDjoqq9P5QLTUf0rcsEIlomQnEYGA7fmTiJMg67rW
yYz6vpXYecTu6aHlmQSU3YUiUw+vqzvDfH0jYcWSRizvgxsPQARjz/9twEAiUAM7YV7KSdQGJOZo
7QV1JJYg5m4ZWSu84qA91jVjZy64/5A5i14r8bQ42aA2MVL+L24swLDhICJLjpNWuAPBWxurffhK
BV/t6VSyAlh9g38SP9u8ChlLeHrjJxzRMrdgljjzPpQc7+fBpp1bkkV1mS/9U0aBGD9paIf7R1+r
TQWutkXBewGK0wV1lIXGasHORpQtIMyeHUklFVMtIA6jC0PBRsXYBl1EZx/CHZIMOwrP5M5f06v8
LVEcw8k8Igb08uvVJFZ+M2tJ06tALTP8uH64vPHZW0AtYrn7RtW49HJVsB5y1Qs19HeXFKUBTS24
Ak6ZWOELqXJes0iXl9qIEch+ASUz9WcAp4vmiugA5osM8kdJOHvXLxkFcRSuMvVk9d3QDwD6S+4o
tohoWqLRSsSWWgUkzibC3A/BrFkFN4OpMcqUPZ1Dg3lht2s85nqdfs5lAFNoh5TbOFB35snYluN2
oE6U8jxtrccg/cRnu6izzci0bcnTwaBNzEsuyWgBQtol77o8E2AO8RTroRhzC/IloURQaFMa0e2b
/sSfGWzPqs2RFC9PgXHvSVl38Z3bOIVA/hJr9YAZJVnTSBAATx3Mfv997q2JHTiQNU387iDbVoJP
DN9g9Fr2NLL0VfoG+RWcJEw9uYr0coAO2s+cjNTxFavE3S2uDvs8ExjjiO7ENEqL3HcIoY67xbLE
i4sHo2SuHJ6yQ5BzUmk4rorkN/bz0gxPN5DhMQBky8DWLMFkn/uwF1spE1rLdBiuMJjLAzUCQooz
GV0kkT9fpD6bZriwKIilwt9L0Z0n0J8CRaKaxYa16IhECAEP/55CBL6p1aeZaJeor3465DOdldrf
1RlB4jtIJ7RW8nec/1zAJTk1K2bUsizB+ir/W7ohFCo1oL//yxXO6q1UdknA8AKOs1HlUhYr8oPY
nMftb73ihg7Jj6tANCuVGSil8BoTRSAW24GEDrA/9u4+fymN8q93AkgnBCiOo5qL/PJcM3YO/Dw9
ZQty9MjbwPlNFXQFVzVrkA8ZSwatOo9iqR/4r4pvmzm+oSKoV70xlDI6zCKBSctksVbmxS2w9ny2
d0lXBgSbd/+iLG3a/gfJTQd33gHV0G8Nb2ORVwxm8aKqEvKQAGkGFtgjes+zqqpxWGT2gG5AgnS3
W9CdIFsgH9QxydTHcGSx++LtDN2WeN8fK2WkD5jr/M1tB1k/mUtPgoFh1ZLUrnS/RdYlIYVNkOmI
ESGSMgjjurz4MbShn6yZy4gK2cPFer55gvKHceYIZmoVOWFCEcMA/bQFZprOBN5FM+xUoWOZF6S/
hMWEAETZ14lXiONdztjjCfC2T986lvhb3Pmz+fNcJeJ8DD8Q55C9B8cZN6fGkxR/tr8hjWCceGGe
VCh67RDfmiKQTvvbux5mZBKJpHBEf+ClelhRA6IAqhU6qoLyw4JAfyEFQYZACdWANhugeN4qT0dK
uuMaJ+XsY/kVitRG2dbQ52Xc4/lcW9UEDsMa0cOv0PNgyqYAG0eAa1fQMPb14CSm8SqtjD29yB7X
r+mYe1eWxxACdFmrq/+poS3sWBnbOnGxzxpKJWFppMyr9fSmBd6vt83z209RyeE45Lc9Cr1G9bkR
RW/ZKXetIKDF4r0NJA8+4cupgiRQE9Ng8BLiHUMyZAJHvHQK94wnA+P4lQ2ZqtcyMdGC3BK+FUg5
PQmWUnnF2KuHIsMMzqJdPSF2p0M8/VFQikBHLWgqfap5UoyOQJ5EwUCCamjrwBX4ruvi33iBTTpg
2AoGm2sGcxhWlVvgCZNHek+f7mvJ9muCWOW3Zj5JbkipwDBFOIziGNOkEz9mNvp5vZrev5944nV/
nmDzhvh8jaOiSTDtY13hAfvjjaQqSLu1m/knPK9pr9rZtbQ30AN8JlO+gnARcow9GXbDQEJROGpe
Yu7qA7KfTaX9jxWoartbvrPttabDVnQV09DvDiLbsZBnhn8DMLW8Eu6JIguCP15G/WxtsJlE6lgl
Qz1qXtesI82vkaJHcOIZ00KMgnR8/+SR46oZFgZYAe8F2ladW/s/cXRjfq/kAcILhjWssi7WMXOc
PacZ6T6t2kmC4C/FY8HqPhjyJsqQX05eKANuc4cEp10q8w3UjaHmUZJrBQczWyR8pQ1ME0aOHL5l
Eyte4NZFdw9HAZy71yTg5NsTATtwAlnNn5jZ9na41yzjOSPZ8WJ0LSJet7NoS+EkYNE5Ps6M4yxf
FsgK77NE9Y5Xep15pYqztTSUCY1utlI4bvazNBBruh0qHbCayoCmJRIk7XkjW12mUpopqVtxX/75
tIKKU0PGcKahLzp99+6MXxVh/x6V5ozC8RKfUZZhSk5T5k4soV6i9KAsxsWX+iYREq0qQcRpGsV2
TNTOArEYNGzCfGt2yqKNT74HPWf4zJHbshwxmd5QD0pRGIodK62DSDoglanOPSURIkShtDF9Ush6
iR7ftRcKT/Uylnn4ElZqlI2hZ9a4ZbfTGg0b3nwGj3BVmYb1DKqimQ2o5j+SUHJI9TM/mDgpoIui
WsQtFtGwvQ56boc0MZ72/t3bPUWvVmNNYT+mQHoNoMqNhF7euI0oB3o7v8WIN9KqoEpShdfKsFA9
ZpWTGzci1MaEDtw5eaTtugDuuq1nDAvABhm6vucCyQfaXSmM4PeOdNYsTjGWIpeZwKkxNJdPzcUX
bZvJDXgAOFuNIwFkaeAoVd/WRxiy34kP9ZUShY1Id2sxbGIAlW5X9VjKrywnO2PMnzf7l0/7bXKJ
SO5NYGVr+3zo4txPWEyrZzqvFxQBzFOwTzPfoB/yVgNO6olkbKfPIH2Cxh+k+trv/8ClInqVf6eq
QTo1D6dYDa6dQYexYmjeQKekDgdgkK9PZCQJCYh+yGKC5Y/Gu4MQ3hu5DyqY9+OxxrsrNzlbY37a
J1x56F1HrNffNq1IKAfF9b8v3smyiplIe3d+19B7/SWdCuswv8FiDXlRpLInbVN4qvFOiaKH5blS
jQaNGps8gbsDFnqsH4B7S0LDBOkDuJX1LJG8Zjd5nIrySYiWOhgrPDlvAJX3YzV0eWUDcRy9pnzO
sTEVhSi/OOSpn0Kxnyhmvc+J5aMYxBl2LD6P1P8k3XSWLbmHOyMOHCbFxjMiWILaB8oaC0XpsvSK
YQ3jZBQ3kJ0JlqnDXxU1AW4rkdaJjTDjx3Cuiyn+yHGb3Suj4NzbEPQCagR3MO5lKfxmkI9d8TAp
HgeItLksxyr4psxe8Cc+d/kI3h2/EB5dMUcoW514cT5YgGlagW6mzlNJHuXPvxfz8KS0U4h6/WRg
9wOmHKFYjovbKGlEmgig9a11/Crwdc3Ud/ofq81vb7Ey2J7u7SyTGlPR7aKiX5xWuvBoV8Qu9tOw
8N28g+sxwiCmFiZX0ghF4nGTMpQYzmpUcS+emV44LayQCWM6M3YWfbxz2CytTEtC/WUmzXK60GVI
I+FvZjsfqJHOMNb/YQ7zNf9KFyT1SwGRD9FhFYrxNrqFHqgD9nr6EzDtS6rqf0cVW9SfwYa5JpJS
EdoWluqnyWsGablLDqDgIzyDxcq0XzeKqGdS1mWM+ZGlw8wruQy8spfmJWCcpB7UAEa/yExYHa3r
TP43SaRJWqnzwXUaic3tuqoMG7z/xN9dSwpK3I1cgjsrQWI6xhm9ihX2UZjPkjpPWXZa3g29/d/U
aTXIzMj8yr26oYKmQuah2mb0wGS1XhNkaJSKc2i5I0oSd2Hez7JcuYovhWwjC5eenvbMp0LADgyS
/zpRly0sgo3dNxuorntMstzJVkxtEoSrOPex+g8JCr3uolBxbp8Hm73WUIzWPakvLa2JuHfCP8dK
tbww1kwJ12gDlR6eMsrv8RALv7Q3lfaI5oA/kIC4ELsT/ZJtVblTvzWwBv6iErb1ifyVkL/L+NwV
/40coIsrGwr2pz4ktxLk8hdHFIADTK/yl0/yo7TRVZH+igwIwT/SX/pr2qN6avSA0XOiFMMT8HNn
t1KnTmIG0iHKQQb0mjq7+BbqKb5Kamsm0HZ0LnDL3kl3cbjmqRUBKMLStn0IYrPVVKEsR3V3Hx/z
N+BlN6F09TFQz6K8imQvHpaIAmnKcHF+xpz6dLFzQY9yzrT+R864YJuk+wp2bvgzspDfxRGSg2CA
fwd2175KmGiIZtRzjCVMY77ivjj1/hNuy5rZefqiCrxviu4bs4OSf1tTjuvXxbVzV5VS+gHJEtGH
l5OM1p9FkR41Hf0Njv3hyZAHJyXJN4cAg2Md9LRNhynZ7IxhTQisHLW/tUGX0wNqpq/isC8cgr60
uwOFVW8vtY/HnB59lrWizGTkW0Z66+A4g5T7c/UUktuTCZvMwRFle8EpMJXl+qNGpRhmL9C6MCJ5
qAKXNZmWOdGgMxj6jb0lsK7/IjzdJTaC11LfmmCEhTaVQkZ3Hd08Ksh8WUmY8ctdB/z/khxZilkL
w0/MG0tWO4XB1vJTrW27dCJNyAqsWfJ+iDOOFnSouVFzU13A6mBbK+ZSntE4imUgWUt7VOTmYFGh
HTFKB0SQw/6HDSAbGCnW+BubKfZef+lF0TqSbV9HrgGizJo0zB2+HnTKjH1U+LRjREf55s0LUyg4
7WcBM4kc+rkVyzYCQSh9f7yk9iM45nIPR+kbNo37pLL5KRDHRXklVfsIfiEO4EYQlGHhAbM9qt+D
GSl0HvpOQ1HdQe9XwKc+X0mRyKUrP0sHyb3g+Yt2uLQiIaHB1IGvFf1gYJ+ArL9VALnSuQz2RNN6
YbRfGw+/i3vecNuAl2LxuR6W2vM112KAontp5zye7ptjsXEReZ4d1t4ILVz2e+qaLCD61HDNL7ln
WwBmPI/IHBkmA2Hc8K+SWBRbq2wDhN5al1Su8ns2BcrNfajCtB9UaRZGfSDyaZ3W2pnabaSg74wl
InibKPyetIKadcAk+jPkapt7+c7r+Yak/iu6o082wVzmw5pYh49cgsGyNrPMNFzFtmEF3ZqxZ2eE
lPJAmCuRgQP9qVTUhqBdqW90kjgTL1YmRjJLbCMApJQWTeR8k/WfWplXbS8Vl0cSOecFn6r+R5QZ
BqoaYUJ3NXoaV+hSBZO5LTvaXyFu0/zHStGS1e9BIU9GDVyFplFWFz98Y0YrraO/dt36KTAywgZj
oAxmCHi08Nby8fX4OXyGEn7CDjGgwSmULV/HlbkWo7aGwScCOsqeoH0Qh6C7Hhi1OqZAVQnEWb7x
I4fXhZDDzmN81rCTXY7egCwjnH0/2UGxA1KeccW3wM0AMCmzYxi21iBxG9aQki1vo/4ECntabRJ8
GP5t/oZNG0sZj9SaO1+RtElORJGXE5JS4pLx4+RVUDDnreK+usj0yyV3oKnkINmZarhxNyN8ahg5
VGrF4ulFs5CNT9Mwx4VvLYOnjw+1pvM2iNP9Tgd0jidoUK+CCavxifMPIYE9XPOaOTn0Q+AR+f2e
yAZNCZICWAEUqxZnu9VyTEclOtim8lIjGJcUgxDZqHcO80qTaRNfVtgB3r0XT2PpFj5zmG2bwfKe
s3gksJJkR+EE/PYZZ/NG/WaKnEJpN3W27Cw8mWV5k7G9ltfr6yZoWkd3vyazmfeRQM09b0tp2tEj
oNBR/VoRqpGPJWF38QqlUixaBmcMe7JMqCh45dqVi5cMShch7iQdOlVpixjr3VB8Ki/MvUB6DL79
HWDtykKligBWJy7OsZIZ6UYvyUiHkd18IRVSQ/fPI2XrYKR5m/nuNwD3tLj9Q0ViXOdWtHOWLNHy
7RxQhF8BM8vbNeK2TqgdFX6TycHHdkuVdh7ZQoSNBmFTPidjOaEz0ApsvqA9aR0BJflPqpxvgX/h
fYHTkAhbXNt4tYHURcZDIz/it0q6o0+qvnlDIPN5C0ZRDBbW5k55n1qkQixPPtcuXLE/bI4iYLdE
LJ5rPHpu4Z5nbB5+kvoYIXtvWC0WYUoLa9VgJgZLECzVL/t7kcnIX120+Ur5kzJ0uOAUysAMqoo+
riCadAsVFtvuqa7lgRPaVwZBW4Lr3h0oAPEDay7D6prKNhvwcpMhjLUDpNmfw50zhJMBdsZZKOPd
cnYf/eeXI4x8VJo4n/QCKvh9GmiYuf/iriWOtyRBW6ftdURdV49W43VY0xcIenh8awhMBthMSFcN
J/DmZr4PwAnHlH8NZcmbJI6yIIToKDSZJjtoS4HZXtha37MVdoMRvnfQndzn2DdEAeNJBqZ4YAlY
k3Swl/vJKRCKTszCIrCt+RDdzEA1+PGJ+pnLTXlwyixqKq6caZUlY2O2nozuPDHDgMeOVZZ3K3Os
VU5uc72dXFp48+WBjAy9qWRLVyftb7yqdyu4Rt4Tuto7xDiOvgmJR72jPaQLxjtCVRFNjYAJXALf
6f/recRtagOWly0Tb//jwVlHc75Ccb4So6n6VIiOXi9e1uNfQb5F9kbKqwJh+FWqr6oGQwqOvZbu
npHmaxEX9JyFabG8i8uNtWToh2ESypOoBrpYAGE8lAxxHvkn76a0Iwkf2HqDsnaxQeYM1OKZA8GP
AX1QxiFwz49fKTsZP5DO9BmTyna8EUJadax7x/1kNyWGL3Su7UltFNc1fp9zLbNs3z85CAb2oxkS
Fvwwh6T0KyhA1T6uN9SeGxJU5QXWCiTSk/LqIZEVN752/b/o5hcG+xfa0XiJEYJjOH8D8mpyi+EV
mta3j6pXA0soRNY5JVszYK4ZyTYJ4g4gZ2+hTZKnvUTG2sRaGcGxzoa470y0Hi3ub1zaRfB4lCdS
YElaz5SRTFIvzQKgX5UAFm/cUaP8ohTaRvtW8F3N9fmUl9tSZpycYzHSbJJEHq3WKJuOAdvTBRgL
fhPYmWDAphNPBhAN0IwQ4A2SX+FAzzRe/pzslBRwPYM2XznVGm5ClFBwd1wDUuwVDbsLGPnuluMJ
ibvOfporOcAZPHvUnfSKEmt8U0VFAMM2KwOaE3nx0uikhUCVfM0ooNNglYQofzDaICsX+Dbcu2zi
Y85WK+s4CZ/kujJFySHPqpwLKpbfNTPETomaE5bcrXE5lz8Iy6lMJGo0WN+tar/gIdd5+gxAkBTX
YumDs0cPQChBNs+GkC3AeRQXvUA7ADRSrp5yXYMvImAJ6JiAvhAi2EhNXiziPdp/h44CleHikZIq
S+l9GemU3bCOGqJ8/Qhu5H6NSpQn9S6g1EFPZt5/dtIECrz2JlLaeaBYwETIk4Fde4BLMeMdSmwl
/YHNUUuTaOszTXzKqkxJn/sIh5yENklYXJQylGvd+Cw2ykcnpmh0rFtic44HY5r6FyWFPUL782Mm
/bEVCS0y+849K2ws3GHLoUcsjy/Igh1+J0wziTGsutghdeXL4eo9zZ69ljiEOkC6HSH4rTe+pmSg
ABSj+1RgTYBYZKaaCd/12dLV8hp3kbN9STlnUJdZX0PjY3PBibwhBQj6HkJswsO1nz+yhnHnGH/f
NI7JROXFqaIlOeaRiCaXDUem8lny+2GJNiBpLLQaPRDql2cT5uiYs0PVgpl9T0K0ZySJamqoH8Cl
l93DxMdexA9Y06n5LbvmLfxdPaCQQqezQ9ckBwPynBY8J7voOEF3rMoE5rk/oSMl3dzF+vFP7Olp
KcLABJaV2UupdcyFeEWdL87UvZLZJ6qxSB/OTDwmPgFzowEXeCGGhpOot3IIDW8uNwb3nYXIElWm
dNoNdgdaVI3IdDEv+ahK7eZ6O2/6P2eFwm+ldPE+CUWpm9uiBjN/6rLckOngrTD+DhNkFX8Syjxx
QRNsvAlfxvdUr/pwcbVixN2pp2T481s8cPS3Tur+sUa8IzbycBcyF6QCx7XzMH+zXPZQJP61WIrP
sOC7FppdmaNjLc2nZaRxJMRKk4M3Crr34T2/c9yuLH21ObmF5XIduKdlnTl2UoB586QGBzQop6em
z+oobdLUwbPQoxLnLSWs9o3o6cb4PlQ/AAtJpg9PE3/MX81WTiUDoqd3vwvkWjpprHyIkZb9y48k
48NpjDzHvLvK1n8CgNDPSDe/qHHM0W0CD+cVR6kT5aG8mGTEnWPhIO22sizbMveMBzFvSxtyiSG/
56fDc3LjCpd/gz6WN4Wj3i/4iRxsSiDLIF6UyOPSj+66c3fyqJY6xGuZ/Y1JLnpVpe3BxB0Pf+wD
1St5ImoDP/U1yIDjw8sIMTRVnTdl369DDu558B9BLAlZYiubjqChxuiLXYEkbMA5Tzy0/3Os3DZw
gEWp7JDpvuIuJrEfELYeJvC31c/USFWdRyKd49eJ4MqmmvHNUEE1enG6tiOw7DBxH6Z7OBF1do96
++/TtyuFFfkDtV23aV6oQOaCcXINQfl5w3C2VgAIlCY54OizqmSoAZdaX+TZHHYXRurkEn2Lal81
5NrrQ14JRvDAtcaFZJjiwP4GOlgmM/6dRrf/EgBN603BPOvN/JcbenXIiWlnM++1egjuOENphdA0
83st4DpA+PlmCTS5MohJ+EungEcpWNgW4qs5b8nSPyzY77ekNKBToQ61mqxbXeBeIi5X14MoJbxR
AlrMez++zPfQCJ19bSBeXhdik4Fv5XrtUqiLrzILnbC+fRmUcysxl5jcqmfjcTFQ/1M1o4V1iOaq
2gbsQ1Z42ZO8WXNTfE2BNnmaLtHzjYiF72iu9QXl31rCb6Z/0ttIj1oEHPZ28qNaPNigBOoRwCLq
OMunwBaJvrVEBl6n4311HLixCrWuFrY7nBUXuO+E02FYYpfzB3x1frX80MHtT8tf9Ax3YOdFNTn3
MGRdKfaSB1kPFK/4PeFAx7onWxd/IOmJ2z7ijcKJbk1resAwWnGzDJMBfq3S4hVQHUDT6RQRRJ1F
o8V9bEhu2YyJNIrLTrS2CFtax2HHEWEHim4esFxRG+PTHPY4Wc86XGaX3qtPeFfjSauNpGdVIwiI
ejClJYyIMZ6/few2atZKcyTs2CI1Lp4jTHv64jjH2guH6JouzvMilNIzg8Z3ecH4M9xRVbL90khQ
Wb53bQr1+aKXM6pvam/Iq/D4kXTm/lklHDvpIPTqMtY8FOssMZtrnfD8e1yw7AS2NE4jq7heJlpL
MvCYITSS2MIpp3086yA/Vudfylni9Qa5CiVqcuMMLYQcC7Qlz7tV0izyQABoUEdRFWKJGT21zrhr
CBJaJgiPRabwfPW9z7mOMl1KBo80tJ+yz2zElymZeiJCvQOwjhsG6mmV4YRD0ynb0EETVNkYoDnf
/VOF0E+dxxl+T2udoYWDBdUqhQybEJzVHT9VkY01QCCBWADrbYuHDs6C3tMVSQSd/RpSAapzeGeJ
1l89tA4SXZuKxYSN1T7Fasy7pVZqXY2g3lA4N2Eosc1Der0ntEkjXcbhbE4QBozwj8wP4fWkqun1
0MH2aOYoXO+4ARM4QbzopXCTEuybfvE9/bELcDLfBGcbA5Fy4CaCghEgvyYM/SJatgr4f91TzyYM
xriUTmyt4kvhQwRTJLPdpsiByefQxhJX9OQZS3ZfbZtEfqbC9JZkbRoFFTJROAk7HSkJ+LI/ZesY
rKAB4Y8ktkdp/mKC9A/R4cxe6kGQWmCoq1NEWvQoF3ytBxqgqzIA6D3LD3AdeTLrKAMowN+tD9mh
8KoGHmf74Jr8MXHujdMZXov73nx8scx0aIo1pEY3N4MX8ZyLnuMkh67Ec7g4LPrPKWHJcs3F9iZr
07Xv0Nng8pNEgAZusZEkXvLfWL3JkCkWweBPnUzTTNTSOni8DiJ1PRbOgn5YSDSJfhaBjeJMwnq7
12O2wuhHIURQ/gVBsgJ7idx4LtKfSTbZE+2MqXyMYgwPNIaLKmv/wGRf0BlV0GYPLwbJ0UFslObi
LfG+8Fryg25MPwTv9sY80lW4Hq3c7g7HVi4Jh1lLQ7Zg82Lf3wZ8ff33tkBy0J+P6vGtl2MUqiLL
2fy0fxs730zOn1DmKzZKQkoV8XTysF3ZkjqNtbTKiYg9kyUK9COyoFJn+D4BQt1OKJVT8wtO8v2s
GIlp917nLn6xdnX3V9s8qgrYqpsuxbh+30ZFpTQO3NLBPe+FDM3zrH1onhOVGoBlFMMbfrlD2mmB
iKfNM8u0N5e3cvASEQcjPljWVexV2fnDWEenf5M+IlaeaLbyvq3Du9txNh2sCJIhW3g4ppqmRLTK
4Zd2muhGHTl8NVmbddOrFroBuIu3Ad/clUoLeibQyP655nBo9H6q9UFr9fyKqy4BQFf0/tMOGpB+
EncgScanvJok6M15VInzaIbeGYZPZIU4q7o5BHQbrDOY8ypMQFf3kOU41pGJoUBOJ/IR99Y6wuW2
un7eBRw0S63dXpvxrN9IdTl029P5WcZRWgWXbj6eJgbJYyCVMGPcIpnwqalIZO5OiNf0GPAeM035
4dkivaI5D1ECbTKaDwguH5Vf/BL9qSk1WpzQgjBbxG7vHYiZMZaU3HxPxb/NAAeRX1s+xHHMR0I8
BZI497JsqU0l2XS88gmu7s7GVb4Dq/F+F4ALnF481Zdkk7017uL6cvfu/Yo2B2GW+iz94PsWgMX+
nsHHvJgXun+gRBSt4e5etXCDOGeVYGDnGybTBWnx9Xtt++023dC3MHUC0vXfwLIkkg2CdLmJcmhX
ec3n95LvDf20V44WMmjhRk2pPKYvXR6bX6wTBHWmhF9UeuWkKfrnAb+Zj0CTXzNSTAfEbzZCrOyY
KQckgLXDWmpmf0ZUjUh3prQQbXK1luCEKJJeXU49JhYj8tgrhOvUm6KXYkwF7vO4phYo2zjzu+O8
UR9dR3r6DBCe+C6HRgaBaewn5Cq26cf5uudfa0NvbSxm6USNVewPGr8SLduT24bHGOkmuyKGibX7
Yyr+DxKK0GoR6QKSlL1D3RdqqtTFn5lAykyrPdWMzD3FL6eGX3AIw0DOSigqXBX5gi0+0AjvaHd2
DeR5iBcKlzymm9Y8Uo4fwH3ImauKPwxMpER29j9IZVQ2hUDXxLuABMe0+h5jDOMCrejFlxW/i7qB
v7DD6/YBDvvr48DIyCom18r+NBTWG25IqeuOXVNS+j+3lUtoGfueX2clrVxkdJqRoT3vrzKtwePe
XA3e0kh9lY/ryj/9HZUbNv5Q0rY1vAnuxlkSsy5+ePsYyZPbvg6vMd4VE5lJ1wXcuibGpAy3VId9
NSEog7SxhKRYyN9F+7gZM6G7DVqL5/BznbS+B/s3EFLBE0X8xkklktIZ5Z8Je44JSIvrjfMoY9KK
czVodmynqKZpKN++V8HmTHEFZyZj+qlnYU1DY9FAgl/TOklWlAs91GSmkIRfyVrnTSDP8Vo/D8hA
io7Nx3pnz1GHVyf7dGavZpz169vpXYfoFq42JJR3rAXdMAg+SkM39ingxTn233rZofvepiGkPL+y
o5ITO8qDk0Br2Oj+mpCk5NM88FpaJ/IVrNODtJ65qU6xKHQvtkGBCXmX2JXBeudL3j5CAsx+Ybfj
Z6FVjRAiaYT4G+CpFU8RobFFwH7EfuI5TAuXKm4d39BPuL/6FBRcaM92YK4Hz7/FYMxhsoRCel59
6isjU7RytmJ4i+wk+C0fYZcVLGo+D+nC9mPByajgxt66PURhYExD74uABHsF8YOnoOy35Spp6trz
vu+ugyXHd+trFksgOAuyJ3QbpQ0dCbPG+iGD05BfZR4eu4JwYNoKpab2X5tg38202TEP9of7QnYr
lRz7Qske4Z6lAweApQEgjq0pN8uuPL390CeZ2gjhap6ZiTZ/YgyvnYUEPYJ6AkckZr3xn5t7/52p
RgvYvGITvGhO4h5gadqVUeTR3C5uFAkKPX2KSo3sibwy2euL4X+M+HDyZ1OW769GdNBZch1TJzf4
xwvG1/KX2EoOYQZi3exxAmaJKs43AGUV+Y83qIkte36tuBbcNvudQcobXUbGCe4aYK/wSl7L7nUE
GG803JCtljGUo0UcfiQkiffR0iYCbOvCQC5fiJFfPc+2Qq5CgOACVeKdqcF50JyIufrhqS/DAiDr
At3t4cN+3eLGg13LJM7Mc8R0e/IJFTQ0FfQwm6Z25eY+9OvvvMRuQ6cbN+zqAuL0GuZde30pN9gs
Lkgcn+PbANxfuSqRbJjtAtZ5Vf6obRoCQdsdE9XdYfXmDG3LKomAuf4zvEPAs2rVOE0+pYXZD4mr
nhXKko8mSWIeD/1oz015nToXn8fzfB/SrjHtmSnEMLUvyjDrJDEFssRtocHuH0lzebcIDBjpkovb
ZLpidf7XaPbuBj8MpxYES7cokvjlvJPeeP+djtYp8/TsIguMgSd20f/sE3Iz6Cnrjkf5jBwCQanm
RCCAR0TJ6ALqq+3uocQwzfdvDua8uienOMOtcfOMm/S5njnvyHvrKBW60eztQ0ixh73k3LEwKWiz
bfh6DDAkrhNDkDzK0tCbYy/XLtxGOnKMOxLBV8+ErAcBuS4GiF5+4dD5wcy3ubatz7Ym0ODzQezv
tnEUTsAnV120LKYynSOCTSGYHB9d0pMPm3PV+cBos+98c8t0rXwQTUATK0FJiIAwcx8uFYuQann/
UZSu0l3xluy4AHe94LImLLUH4EkXnSA/74eugIVIYmSnedQzimDCIHEh9g2QOKKWWVI4F2BgNpUF
QwAT6/cl1EcS6bCdMC0uvUDEo9luQUqNYWmE2jHTapvAxsmU3gkacGVA+6FBRIgifvBXAa94PKs4
4LnMdNVVPuVmkxL81QGSLyHOnn8BDIiNxWKU2sw3nR+jnR5psBXXkh77dWbtMw2cfbI3Rdwbn8Ia
tKCly3uY+T5tBRUiF6rmNkMU2s5phHOzF/End1BxFFTwWsQOfLf70mRPQI07DPDs5oDZmMKVReyW
aBq9ZCvKkEoxF4Kj6od8rAvzKBRpLyG3NETXOvmGPmibzK4/dEZ/rXi72ddw44/b6+XN5NWTvkqr
Wk11aFk3t1RB3LchU2FUvGqIZTLJM3PyXxtSkzcHEz2jbAXWl0raBkos6OcHakPJStANXfYm4Hxn
e7ykpmxMqpqhA6BRT0UyPveKJg22a46y5IRAUV56S1BmkYEfIx2i6P/aLeff9gczRkP7nlJXdgcL
E8XzKKM+GZYSIIEwyy8IPoGvBnqVvyfOjhbp34MSCc3/f81cVyAkKn2GZO8t25Ci1kLXg/LrClsY
ciL5rBMFzc68O+t7sD0W3WZmoKVtDN1Kpd+WLlXXXejblOZA3tw1WNWv4Sgjs5pfKy/zDdzFwu0Q
jw/gJK/UMaoiE8hy4wNUrVxqUoaF/61KJngb0a3thrPWUr/Iap61TIZzgozeiq6gGUAF9epSV7wX
py0lrPHHYSPXqySHBOeGbQFe6owUko1NHkrVsLBnQXp3PbZdzJ57ZdQqfgOmzg7OpbzW953OdrKZ
qAc6Q3xbgmaETXCthTJsG6510FPc4fuguQOH3Iuuij9iIRQgoTh1UxJLtuHtUtHO3bOMPvvCZgm2
pLt0fMXVfzi2JQwf5gGboy5KZIm/YVAZryKzDzgsjl8ag2ARX5XmUIQ+jIJTMDkAKD32ViKVbzde
W/x/+kWiWuvJAug8JOVMTQu0BYmNCsi/thluaf80qRn/UQ1ArFBhwSuc+vOVUQVK0ozXbL7NJTVa
ifuC6XdrQ49JR016uLR0TmfPq+9xNiZEaq/jSYC2pjKVraG0bO/7Ins4OHA11gQVTkF8co9+YEGp
0yAFAiPbopjnfyhwmyFzFRoDmaAkaOgomPkvSXv3kHgrVngMFa4tRZmgxvdWgwIsHo0dQvRARgD9
1JQ/uJiXvluu/vsygKy9PFCi2+gcWiRiCUWTdWyJ/3TtBmi90mwSDWagofTFjUaIGfPATC+Cgdq3
jXxgquqdwYf/KP6rpRfLm/RRpD0RZc+PLfUB+Mry2a0k0EgMVZqWzIQot5XtGkQv5HNrl58oPiV8
7k2t2i2RYzCWcp1IjP5ZE4piVEuVH3czBSE01h18SIqXB9MO9B49RaYSbnedCYenXP0JQQFwD9Nc
gTx+H3/O8qrhVdlXXufOzgNjDP/JT9sZyeaNE7yFq8Af9GTHWds9SE4BMGzqMIVCfvwywOwrthN3
7+KxfmFCaqTg6IDxoeT99ERHLPtE6a6bFF10AfUhsSiIRGSNInNxjvmPawux7jVkMDuDb11jXueF
brHkjrOfqQuyizgLcsxiD4fU5uaP/M0nkvSv892/SonzTuaCfF6YRdn9I1r+ahvj+vH0sPxB3VDy
3mX3K72LW128pn8nZubw1cEMxA6tklTNKfFz2uraA525ZYdBstjPN0H0YAfLyx67/cEtHg1c3GmW
W9ZriKKRNKPxCfmPkrbJQqlnjwN7gIKsr2QJWfqZE6A4a/zvfvcrbezQBuI9zCUie77A6qupTSxo
eBueLFkcRBgjslPlHLXAFfRmnyvBKxFYU5Vxj4nFROYQvb2WQFMIFbVCBrDw528ZvinJTFi7OlO6
RIvrEwnbzSvrFzMVC2WDK4V/szmQFCbGoVNxoviq2/d6SH7LhC0O5MTlyAuy3TuvEdBk3AUhhh6F
KJWzBcRXDK4gxJWQN+NA9LgXp0tIDoXOnbnIL7WfFC6Hl1L12deNu49i/R2qauDd0hIh5nEM1xKJ
3FnubRCc0XrLdnjeh+Fw1JaKTGlB4njd5DmvcX32chTD6XZhIxC0/6WqXFtFNQOJn9kOfIha30Ow
04EaN9dEEE2yPhGmR39E/nsnsPjLYQpHWnlKhUo+WARRvsLk3T6L1VjxI1q5J/WVY1gBqc9aIz28
tuKqNVbRwzkY6pOlTdcjj1P04V5GQTAppJNVJVfCThMledpd6dNpit/AZnIWh543ZH9qPAALNcfZ
kDmb6vA26ubqFRkcGihO7HHMxxUPd3YSHY7jiTHotC8PeonxCDBI60zglxTOsu572DtjYlVhLILT
U+nNv1d1a1ib4xg1UFhioFOWOtnm+TYj6F9LEv7YqjNYXsVAiFXIitXH30OZSF31Td4pcE2a7+Rc
yPnTIspIWqfiPDOUfJIDkX3R5SckriELGz0P+HzMZvHqEjo0DjgFJs1XryBwgCAhgArFceghbRZf
yQvoAU7/RmgfWiHzyQEbAsctU3JxNndqumXL7wmqPQ8hkZa2v4JeKgMrsZ4sm2gATqAzI1MqBpre
cmBdc6ad3ibcaTMEMuGF5QkLJ7FGnh7bSDhPqbjUCYTyxkmyi8bNEmYiwo6iG/VW+9s2QbEwBhJy
fNkKKjBcjyAZp7TVYRnmaHcmNlvGhs74MWuhRiiWYb1d6w9q+m8yFisVXwRUsu9w8bwuiHHSHtw6
SDXqngw7yT9JWUw6u2pGN7TAqZNbFN098VDuPeaEnFKcm5UAREoJjd9hch5ChP0W9onlOmRna4iy
IZbLCQSZ0NyPoqHIwcCA5Bvkg+wUKwBNYqnNxQD7qm9Y+fUIdaurXRjxW6HYWDNon6u80iXx5mN2
E+wxtwhjLcTxNYs7YiCNEa+XxujMyYu/U1hNE4oRHR7pzJOMyU7wNCZraZsfPArOob7SZAWwUdzQ
u+cHpAudXPqFGkfnjFGar4z2arTnzrvWhdw29CehrqD2H6+oe6rluhy/jFuMYcm9hxIiezvc5EN8
vuSSUGeXzbd/0GwiNvARKIJQIPvTLDDypdfbKIElQKXuSrA9aerl5MqZmXRrooHke3d6Rp30b9RM
KmxN5kGhd3xUsqvEEHlH7grXmddOz8SInUF8d53AjO5fiWKBcojNdtoK7ZMAj8x7s2lkIc8GM78H
0Nko1FJenbZdzIfIOf1LiiDTFE+pGYr+HUCh/D0gIypU2lhQP1HrhbmVVIBI9OW1TBCjzahwC1UU
zv6PMOMaMdfc8WSJBlW2mZepNn00m2tK1knV/DJ6kDdshmqQTzDHk8k+ml9en+EcHNawBOkHNmIh
jwHQ1Y99a4p3gsGjNJUM7ybo6eBpAVTEcQp4OCqiKQgGKXGf6gXmTscPaQ/APecVPQZwvzp+F7v5
edyg77SBk/BpTMBD7tS41t9sYAgI0XUDnxScZWfHgLLrB8oyMLKxG864ro957AYz2Rv6zec60xGQ
PPPmkYaw/76bq7YwTiWs7I5coiEheB0f1sz5QjGuu6iND+bMlKUAlLM5YQYsBq/BnuOqKHbavMIX
G/gw4fKjPOui3GgyosS3KH6KwrG2GrIi8i/xCAkRy+MKvEcnHItOvZHS1LCJ966qw+8MAb92VXHX
jYykzbxkJqOLI3kFzYbyin25kOiqh4eMxtN6pmnwVOh0evOvEDYM7PVPLZC6gFviHahYBIPF2XBC
CIloY/v7980VzhefvDpvfSgjBWGbh8AB1xRv/XqabECAmkJ5967p40yd0eXRTfOYkNiUOYLC429h
uY2vz4M42oO2gs89D2YcsnAtUtcs6y3aEkehdhd658/gVpJX+ipDhkzLLshOTlzHsXhAOHQRSTmg
mh9AIan81dgzooIeZvAN4Up23zd7kKaeQ48MGiGXWOjXunf5pv6rkuYrdTlt6Ar5fR5fnZcZGPao
7jji81y5mEAejHOCxHifb7T80fJjNKEqIRki99FSsQbYfyouVw++lO4FIoDNeMq3jk2I8djVHr2I
6UCMVRoo+8Vj75z1wEE1OYPod8eIBIAP9izxkcZJrFZ9AaGDyK8JqCK0ytLjU0NR/9AAyyR6rCwh
+5ADHrsyKesd8+l4OHsw1rjm4EQKtg7bIzBspgxQQxZhMKSVzatxUI+R8f6x1wprgdm9951UrGeA
+YR4V03FnoHQ2aFK30wpEYVZDpy2GD8A9MGKyZsfnBF6pTgr6lONeKK6Q3RgBQQ5YIl462SDBR7u
EP4i3X7PdzCrzx3Qj7nNYcn5nlsqG4S5/Vf55A20Vd81CcsOgyVNlgHaX8pIewNGEan0jVTZUQxN
zKWrMs9rSjxopjZ7s9/Xb+1VJYS90P/0lz3zYualdnhgi/dnJX5nyOKHWvc/YAm9KquQzh7DniWU
2ldfAw2KjZpiT1VPqnw1ze5BkxnPC7UyYV1Ts2gixkBNCthXemtcSjycI3ZQRbhtaS0KWFD0iO++
1IwfLHZgBqGRl7KPvbHQr0qN81ZuN47EmgTMONykETfM5LAvhXp0tYavKygCu2zj0yqR4jTmKRxt
IZg1XjhHNZKbDXXn0YMXD94x/YjN460KXqFV2cEs9m8B80HgMDC/FSNMyDTZMCyhwLgxuAFILI5b
UoBvsu3Iw/es0TE03pyHoshpAFBvbPfvqswM/aKI5QBS7bwp2SaDR7PKPwl0jgd89m9aO7VKud3y
xqj8MTodR8lIKPt6QAM69H7rIYtn3PJVzoUoYODz3fmzDgZsMUv2ynpSHTqSSJX3rO6c2AxBDswe
hKv8btK6cUQOYm9EqW5Qc2aIfIV9TtvsofHOP7O922i1jsNC5C7H+iHFr0QfEIfVTIJugB0l9xyb
hcgP9FgrdCjeXFCdvidazEni0H3Z5PcI1eWGogQ7BXq4sfGgRIm4o5VuAZZ+Q7RQ76tamD0k1QKk
QMSZF2TO8najqDYqAfxj1KCS9PhVSISx+5/G5pPNsmJVTVXJAmAfhIgS2Gtwz1I6+fvBS4dg5Ui7
upq9kTA/w5k11IYpjoQfmejXdBRpFj9+TIxZ3wX4InIgAV7UZhsbTc2Uqk9LxmTK2h0ik5wjOfu+
qQwmMW0VfbuMoTq94BCeBg29rx9oVSb+JHZLZmpSb3tRH3s4MW6KdQfVDy3NLiWISjvILHUDbb2C
dRoELFtnMFGxq/GVYgs0H4LKj/vxUBL/md5H89IqGMtXVmmyCkAbTmGKF9ZDJ4HsMOfTuwmj8EJr
E9p+feCVeq6vLhmWt+F05IX8zOlogC52/GZfdpWDSJgKE3wyH8lKbu2Ou9SxQ01+Yy2Wr36FHCvn
S7G+CG3wBW3yTQ1Ho8q/ZcDC9BIOt84cP7a6hnDc3OpE7eLPD++Y1P6nQM5eU3ifT4wQmWY+3cj9
x/LrKCH1TbuuNY2ujxQE2xB78Rz2q801h9GH1o7qITe6VJz//6bjXL7uILqk/1QHXJ8oSOjxkH5i
RPmHr7IouOuzMpuBxztFWfBngqSKodzWdaI6KE/pwL9KfBnUKtAc7G6EH9qJOri67Qn2E2Nci+Sa
v4YHlS1bSX1/NpgPTZ7rOaKNEbAzTqQ0dR2Y2S9d/RnqTM8lZ3vq7nhm1qdalia+X92m6h9TewVw
Cdy7lMLZpKJ6SubBXXvzvIyNTsyrQKb+MjC8VFVjZEOMLGCrwUSIJhjVApoEsfVTIH+NMV/WN/71
qqULTSLnt5J0Oos7y8bqT9QEN2PE3aJPK+EAgh1Ol3uthJnEwNDRHH9JLww/yJinC5LUkoE4mTEM
1yP8kaNvhivOjXJ7c6aKFu9Z8fsaV4rhsJSyZoRUGD4RuZAtR41MPU1YBVnuOnpVgk1SOQQ540nR
EXMv1nq1Yqwo0MDYbMp+1+m7uDYr4zeIl5E30R7NU/cSUV2dRDTSZ5uyb/expKL1sA6bthdJbDwP
5zlM1O4khcvr6/pKt99Di0DFWaAys78qOOfJ8urD95tLo/kEqZC5Q+cLDcwerEjWTFi3I9lc4TuL
fQ40z+ITRPkCFtv0pa/jAL7bmxidiwNZQW50zdm2xt3vbm6IuwuulmSZdmB+mz4QLOWA5x7Awe4x
PKf8SDEAadODo3mdyIfVYJHS4dH4sd+8g7zZgcCd4KeGAiQQDSdtSPFm9WL0cqIZIMJ4U6/Do4vA
RknzTWTkwVvlMZxCr6gxNf6MvVlbuOD3IQUn7w876c3t47on26FPfOJDPL/QRsWQeNxYwvloGso8
MBx3dmxIY5NFKp5h/8niQea1dIbzFRwfy8ghjskk9qGmkW9/UFKrXjkz8a4+s84ccODfUf5FeitK
CjaOdldSq1YVftoQoWzXNgXR1waP1I5j7W4FA6Bt9FsZtZZsByP5UlrJcDpkovmi426dmrfSjnA4
j7K9Uf9aZJs4ppvWiVGYiKGT+2ysX0StnDJC/kvIo320noLPq9AQVphCVesAEXN6DJYdV8oxQDxZ
9M0hcZzwkq02n+I5WtLekGfsFwKKYvq7Rdd0mQaTNWk6jTFUMr3d80wPMcfcZk2ypnv7sdPliKKt
BtvMwxgw5ZnHSoxIP4q75MZdxgiKR846NglQDcrJ+3KX0ZXYcgIs7ywQNHcTChE3R5OMjHK153/l
Wr4cur0vqVIxGFTFz5OkjSaNKoM2O3VhGMPCZoVZQvQb6+A/RAy948NZ4dRVrbB5q47xCAgfwG41
676Beg5kfAIVkQMvuzLCRr+c/J2CQaeZX1VjOjIiTUYtGNxqr2F87XlKDhFdfQzVwXggy77lrnqv
6k3qXRBOzW8sltBiw2UMeQaNJ5ok4zkRWPqHFZF6X3fefSAgKSLi2HrjoIHDoCUko5NTrVoOEvqc
IWViDrT3oyUAHsS9R0z2N4wuT9LureWOilUwhJzvaKIE+U3q12V1MurUuHnDrvblCAWwDZqjlxUx
OMIcBXoH1v0UFx+8uqSb0WyG37vPIetzdQddp9kZfl0sEgO1NZAgkeGW2t/MXe/awxb2fuhUR1Jm
Bjt23kpY48qpehsS/EQTAeAeqN0ADTHIRTeIbrpubqyAyZxFwCcxj1DO1m6F2v+FV1eqKO3jJc99
qKsOqYPmb9VfGKno80TOWrX6QfIneV1xfV6DwsWS7wy/nJU8PrUtpeKdaf86W8LhNDtLyVk39fp0
VN6131vC3PYn1OSMk8NoTlnhfGVYWRH/rvU1lYL/WIlOOPxATXx29SBixpX1aMT90wcjCCg1pmze
8jvbCsMe5Y54QJhXL669p3AOAUyO6iK1xvxOj+gMbG0Xj9ii0I/6zterNmDgML+cj89/iaVZ1ump
EDUyrt1qE/ufvEIHco4G8L47aYd2okK7hS/HFtRO+uqqodDfbq5uFkHC9Zdc0/+6uLuD1Eu37/UP
gyEoaNjZQgVA5KHOjsssSw97TTR9C2uwqsLKqULqQUFy7HbJCZ78SmdCcfJJrtRXpa591aB9M1/C
y18Ji+uWNvn92rrkdmJy1yFCMZNui3sjaM8o+a/XLDILT7MZsnYFRByZSiMIbMoyPEXmB5FFw+BW
4jmFT3V8UKga8Gja2pHGruAEerrH2bvZ3GgGjI1GUoyyggzsUpv9tusKmduhlUEbKfor4Tz1ZPKD
/vOXUFZTMVk2vJDsKHYEmjyxEDNQLP1GuYLNeqOST5ipx0URqZHZC6Y+TDQOtjlGkxoLqkYZRuBV
Y/0aOk2IOCwSlvpN4Iw0xbfNT843zBh2fOhnpBeXR4/M2q+mE/nsinFFIPDpCSAQdQ5V65olS5ls
ALVuHtvOMEf57/6AVcMZsxwACprgkILNiLGx3sN32CyxZR5xeKW/bBCFiox6GNYTsItnEpF7BrLr
kD575lqnebr60j66iDY3QqGT0dlkPPfrk+uSOngCVLQdBsSkecAuIIa6FhDLHHUG+XewdQ4IYYCv
4Bm2QVUyd1k5UvNygyeW0xORdfxHemM+YRZfIlIRRnnMNtBzQym/mKe2PiTS2pfvs4QjZiY9ouyU
N073Gr8oW/H1pbTnnfllyHklN0YHqLj3CiJvEQyK/n+366V9LXzAa7Nb2d54uanOLEiTJTB969a+
iRVl6y4pC8sxrcJjtlJ3BgCDgPHvBaDq4K9vyjqHjrPYx9tz077T+E5zmR7sxRXXE71Fb7vmxrKA
QIkqnhBZpBQPKKq16Ey7MUWuBkCYe+/X+v8KqTKVavjfkz0E2K4XdOEWEiFV5nQugHQTNyWBbp9J
oE8MOBqKoUShOiNHGdiUmDHCKI9svBnzPU49wS3GEsqTdww0JaIv2yhc2dr4U+V+cUNQSWeVZ/IM
zv2nUdg7mFYTWzpLt1xEtOHPuYh8MLtLYwNC8yjp+Oj8NmMxjcDg9EUiripERKUxW05IS/ROf/RB
mwliPkzkPbJHd17R8bNWvOmeAQthtv+WWiLuQ8kG8V+tXhZWyAjBbrSNW6Bokbfk++1wujNtOIcD
L052+f3mY4po37/07pGWY6oBw4kWqwYU2zZVw4Vk/2fl5IOzbtN8E1+iSSb1YnWswFMmC+5ZlSe3
h3rY5SvW74BwR2BghFTVLUl20nl4LvZu1pEBkq39awmPqb8DLRN/HHTKpJCQI932sFuEGRmGzXQ2
dYOkF5uLeO7FCDMkh55Tw6khYCWLPzeJSgVocEza8bEbYqb7CxbJA4aI/Yd7CfBCZGZrEWfc/WRr
cqAihWC1FrGMfsHrB2XwwaKeAPdiDLhiDBqCigq0XOP0d9f+59atUCL/A07hmXCVXVAVUFSfWYx7
dvcUVmZRhqj/YsQFTSPCjiwV9IvukIDbIsNuBsCR+vXyeejgqBLG3T1z3/VpAxGfP7jbM651NjFd
pfax4VfGqkborWlbUrTbAizG4+vdH9cQgtT42sQOgbvQtZGDZsnq5RL59dXp1Rj/0UbHAwSefq/v
3XC7pr1mtgvrCIvcCv/d3zo3EGvg9o5VQGCx1apibKzwHGqkQxBYik1a1OA8FlfMAix2+pseNxfz
uky2ikSEpXbBL5rsU8xjkPw2KBi5Xu0aPU2TL+sjQeQpvVr7fCUUkjhMbV1L+TUCvL0fKXQ2mWL5
7JCAV67kt1kULGxbveOgr8T0OGZNiusGp94dRoiZNjLEGdZAPSTf9WMtlKHCDTApLlGF0c2ChnFp
hG/RO/3sDZJsT9qFFdJPvNPVDj19xkK830VDbqfLW7Elnm+pvKar5h/HamatsDet9GfIEtOVEppb
PfaOJk+UJSFA2cYNcHlD3zHJM+WeyNSKW6gtzjqydIxQu9yGALpgfFbr4FYzUPCNUZqnan+Z04Rd
snZgjl8kXNOfMbsrRpru08gFhveh81LUDYDDll8KwNHV2ueae2+KbvaAmFBWG7VbOX0GL83L8ypx
APb4XlzI484MF9+KZIzIEP2qtu1/nsMTIQrD8P3vz66TNoL5I3bEYlfC7Qw9q57ivJuVp0Hyd+tx
pEqG6VVnOhNdM75bqnp3TldKF4C318wLzRqNpFCheaDx52aZYFT/Vo03rRqzxE0YYsW3J/uTKKtB
zkstiS4r2OEeUCVwMPWBH798EAPVsQXwvPQ9RLHjy2diDXOyCqe0pbIobyj9E3i1TEkPMu6Pps8c
gDLjU5PjPHDnpO5fmt3PSBBvWM4DVhpCBCZamJynabVfZoe0Hcuf15Y2peZ3gDxBDCvPkxDJ/Dcq
L/osaiBzzU/Ytlbxrrz54sJd3/43xl7A1OhqYtsil5NiMsHRkNDEZs0B884C0iUUfxRJaPe4e+17
Wq6oqCS8NBNefTl6UZ+jt8LhsJj4R0u/UuPKp8U1EC7QUa4ohbYamwWPzSmUZ3iSphte1hjafJGL
ElWanL69qitnrzgASvsFtjMqaxFkRU6PttTGt43bBKqKHkiY0esil15vl5t0TSzh84UkfpSU2IQk
wYaiLPxJ0Pk9+Tq/jMEPZ9WygglwAoFNOMVCzrh15tYbsUlysdZ+Ewn4VgEp+OP8iReHps3/hOSo
e4NmOntaVon5GNfs94TsuLfbWpna5RizTT4pVvdtl1FN2CgV+PRWfUSfUNvhdx7G5J7+GArIObfz
C97YdY8K9NRBDzpMWIdQVNsOx9oB5kPl01ZsfQeFv2H70vixC+9kTLid60AmtSA4mDxQSwZY2keF
Fos3fjILMMg686veQ8mbgvCs8bbIlYip+34eNEJMX5jeWJk8ZAvynCyXSm6u5SMH+ibDmGJQAuM2
pkcbcRMcqqfzGtr2v0ziRXY6CHzAz1l4Kpy3XmELDoIxQCym/JMA0cCk6YWYcS6PdjdZP8EBu5SF
fQqpKVQtqAlDfv+kakPHoS+gWOHAXlYkzBGdaQI+gjPF5O/2zdPs/mr36HKWsxCkzWWVwPED2Hsb
ozQvBlvpZLeXWG0ybTfWO268QMjvh9g/+mdUQE6o7WBwgpqSJn/+DjRf3ogkPVy6BowrO9rWd2pl
JGQG16GDlU3u8QkXPgUXoQtw9Upsdeqr1rfyKod6UuShao3fId23+1IK/iSPQXvNiktaXO7oeYaA
Ixd8IypCuJUVte3Zu8KN3sKf8P8OdL4cqImsVlfHCrxNOtdmviqVp5mNmm/QhIIir0mxe3RW3xbg
rNwB7RH7iun93pMEJEXgo1u803IdmAPqTC/e/MV7YIfbxzfgN3g0o0MMNzJ2cEz3QrK5ZeJgVtVq
tX/clBL3YwnUrRnQcwCZAz19ZVC5tpfz9A1o6cKa2ZL1G7ZWqFwADY87v0rcD264aRBVxfVu3sTK
PAYAsrqnbxGwDpGiq+9IQynXjqpsPg8bQ94gsgmE91ksPVPL61ysQDUeJGIwxMdsjAG/5ow4AGO9
19Jv58fI2NBb+/3YlbKscsCZRn4aAbYZsDJS6/kMsQH2nu6nHEzHUHanAy57m5kGlBKQ+rAZtm8d
7tJSuRzBgHOSW9zZWGbXWNBg/jnVH90zjGB3Qk/ZuM+BnQWz0EWSS2wbv7Q5BzOJEdbOPigHSoby
aOdwItFtOo2aiqXKQ7c4T9cFSWXAshPr5uewKLRwc+4ySBCRYBnyWgdFKVMj1oqPXlJ2aYkS8U/m
x0Y0+ifv/MfdSvuYD30qUa3G+BJIqnYclKUtcLnlQTQsFJrd9q1rdqA8YgJBceav2o93Uupf7i1J
xpzfXHa3Np4EcSeYjH9pKbUTfxa0ot8UbElf4lsGB3B1co8+ci+rQ2S8S/N92oI6ZHvW87qTfXQE
Nr0GvmRgqjFSx3kRDVjP53wBrx/s1kqAS1cVCWIPQ+nxPDeySCiWccKxMbZeWBVOvfaZkO6s1c51
83ZwxrWKtrLOPPaTtY65KlmYBbqhDqP1HitKHi1r+d4EXZpqwXW5tIOFHFN7ZN/9NILxCE8OWzUG
uV6PqQ62jiLtwpadhWg3LleNlJXUKNpwYEToVVzTt9rNcknQQYBW/Z/zZ6z82Ae8n0cvnEsMaIJK
1YbF0rmU/k8T7iCKchGL8/+nLICP3/CXPHUP1NobeTRNLPN08DljrIuqE9v7Nd0wPiqbe18bYn5F
FwfiHet1lLl1CiOs12XW5AY5qby4QlSfFhlti/8n9KH+aGAh2BfDNt120Kjhx5DgAvaibFUzmgPZ
2HILrBfOTMFOkMvzEIiL9D2+eVCu/Gsa8V5rOcCA6ZOEeQMsFo2aEelTrqwTivAS9P5eXS+Qp7JI
8ygd/6gOapo4kwEwVugR9Z/CoNeOf/GRkI7FHy3rcgqkSO5nYs2V91zdkaJWVASHiGtISarfbLpc
kJ0uh8svhZ9mfqZ5JzhW7wDxJoHIvbK5OfBgwsq6AIBX8dwjPVLww+9pyTwt8vZNjQqL6moSM+xK
5zO2ukitUA/YH7TbDSTcVuTv+c+D6/F/gJOuhT0OWK//FihCADPFlexH9aEwG7Xkc5BVpGHDPseA
pgK5JdAXYALF7RSjt1kj0p0oVxtEuEEi2H5Pwc1Qai2rGQuuU6PIqN2UpcMT6mmdZY70lRLElUKd
wAb04BVv4+ppuj7ExM0CKtCZUdet8ZiVnEVKHrfWr6PkG/I7ErgbxPNhL7sulaj9CA2WYygRIer+
1w9bAQsAHp9gd+XkmNfnhoRvcA8OX78ozZKpyh9rInctty87DP9YGSqzlGoOpQh/qat7TnWejg7e
6QzF1pbn35RrbwrEHPY0bywRYboz0rUEe2Zy7gNhky/4Met4NGU7+zvYc1WioEfomO+ScnsqzDi6
yGv2AigoEf74qOdhJDkK6O1xvUInffIe1UKN+ZQkTDH3Yc5i7P30i7UN9sKcPOUyLC05oV7sORDJ
iur4jfPweIK/QzyjSokxdiHfJb4iBkx7yOyWMOQOn11QB14bAFSKnvAk/lLPIvbu6Fv5ISlt9OGV
cgx9Qs0tTg49q3KwbHCEZ1ZC9Sy1uNZknoVymREBt9YrkGc9+td3XeNLCdoxrAPTU6Lu1xfnbvAq
b0TRcNsYYDvT09MpIV5BnPM2lxNbGQWv+u/HteQy4IUL3XrTQyRk7m0cltGdhQnsfriLWYKlm9S9
r8zsobmEBJhC9ax2GFfh6qm2O2NupheBWFsGWnEQyP4BYCbAtiNuCm+PW1dDlmqHcR6T8wt4Esur
NhYDsrYiEBoi9NxLb7enWYQYNhyELoKCOT6tylTkN2RYoLN6gPhDFkRpMzeySO+rWjqjm6QztStf
B//vxQF45LxQ699w2qvA+a202eBGgT0bG12SLqn17JCTXASjJdNwnU2MzYWoqRrz7fuL3GMEya3J
T6Enb6jf9NFjUg137CzEjBieFP3gLXFHLi7xyOayhyJDqUbxn0Ln8yzfxNFXdYbash/GEkvesbne
WJZ5SkNKdGroLmm7ZvyYZrZaCVz9lNtfWnQjyg1KBYzQ3OMYvFHnJG6WZMbWgKQm7K1v/gzHvw3O
2I7L7MZN5Y7Z+kp91/gCmL1dzAFYH6DvTFF2MKATYzjRjf0Og7O8oRDChDUZo7Z50Fz9V7C52rcr
5hPK+PehuM/tOZ9fN/h8F9Ns9+VEXMt5PJZzvFu21os8o4BDzqla28mm3So4sKgit78s4/36YKBh
bCT8OANXbj9mUZRVwAQoDwboVJ7XNsuOuJkliZq30Yy2KuEVk6cdsjqJNL1iOfd5Lq+Iawq+Tyin
naTu02dq1JgKYcp+zpbgbbEz62DkhFaDFLMpr3hFv99/NdK+5cgHNRonhvUrAz3iYwVt97OM7lmb
QImwpQuaePsSCiS5fRivjcBmJuUZGNyp38Y3+27+6rsLMs54xOYSgNlK6QyRQH6sQi9a+yPELKQv
mo6XqnKdYfgAJQA8BGrvfFOVysNfXb12hTIYJV06Joe/tQcO7XYBn236AhGdxrzxl3FaH/IHh1JD
LDSNV/sAyuUI7PhTegXRi/6X7plbWhCsvTitHOEpje5fMBlK2imTDlKGCC8JA53X5911v3acnvKR
epR6QPsAhY9XDM/pA5FXc3ZfQDVaDBk9g+1ikxgVbjhMkqBp9G6qPhqOd1wqek/3JnCLhpFPO9mf
D9y7+BnkQDYHcwAz9zE4wceX58XBV82PQJoH0s0n+gmLJdL0T/XJNx5y/QEXR6ocRnQNzxMN6JEe
nKxKhiagxEXcmzaoeNJkFxUNHA6BDF7JJ2Z1THioUR/Y5BZfnqBJG2Ibge74Hqf6Jy0Tn31HoJWT
4NKOdtmbkBFO1r3muCxSYRVqRMQAwW9qunpNEWE4YwCFQlCMovHpSl+M52HRsA5zXP1ZVqKEF1QJ
1Sk0BTQXNVE+TavQmE6IG6IjTaldoYJzXmDM1z5CpT5lja5ByWzrSp0ewkGBMNLnQY9cLds1m/as
FyM8lgfhagdof+Zlk2l4qhgL6qfFcbKivtdmOJnshWf3qvQHu0Y2VyhFRGinpk62Cdf32STPFkIl
r9aRHSkfhRtiQ313VBq6idxPaDQ/FSQsWk4R8CMgl0IyhlCKDl8SWernYbnBrlp12+lhscidIDua
50/AkibK3TyMr3WUQBG93ElaP9pjIf2JdnzzWYXWmh8L2J5djpfrOyP4/W/bHYpkW3CrFD+1DMLj
qMegf+VbtfWxiO2fmXTW5XIVmj63qDOIYZVN6gMpem2OJwrv67URqAcVVzzpvhyFW44P4X74YQa+
dAUFqsELW6eKnn446EpNRJGIjrPcrdEPdw89LjhM7XrDu8ufUBiD1EKJ4rwpuJ2wAgdfqujBPSZd
eqLwYnirHiEZHkNN9sRzrutluKFYxZO1plAQO2z9G5jPthcrSTru/YY7fGO27AMG+/p1or889etL
bbMCt/jrRuqw1/w8o9ng6NWmPGZk0FNf65+s7fLqfK1/EWxrb93pAyQu7ltkG36/39oZuxZtcpTv
cioIEiw2Y0oCzH8BkYFRP9wPIygXjxdgQNF6yXJWfNGarJ6DjHdYFEq09o/Y/oSClGuFyMFxeNtD
M9B1a8X+gW2QfzRB1XCZjPvYw4TpaA/ifRBDzJJt2Gdj+EbiFoHtzqEbsXM5Ii0j4Pt9ex52MbR7
09p5Sl0bHzvyPHjk1lCDuPg+06RDa43Kte23XiIuaV4cDpIiValA1cwFjgkJWo4i5vWgeIEIBgDm
80OaxbJvekRGB0MLNikzNo1W04kQELf6kR+8l7Ffjp6fwzGDHaLMqBbUPw/6qHcgL0/4pR2uCaN/
GAELAYFKkJrcR8T9AOilTdClhb+n950Sn/6EOzZmLyBY4fx9aQQ5ePizLpyVb9Aomf04+M8ZRy8u
wbMmHPpQs3UW0j81JR21jL2gQILcG+yxc+d7W/T+PPgbZGGsRZhQdAwNPluxiBLCoZwWpeY8X46G
XiR+ZEY+VU9Pdxx4sRPt6G8sLGyEv2ZqNi5KE8K96t4lRiP9hUp4bnTNVBP6UxnZF5ldkulc8oGG
2k/0mFwrASU5rgwV3YIOUVca4KgEEv1Wb6oh5niUUoLfDXJSiqCp1tcZoaqkXmFzwpgxgA0I/7lW
0x0xg9cylUoHRK4Hnhf65eevaA6LFtRAG9Q5VfINBox+YnUhsGj78+A6Fj6N8K7sk3eFircZNCKJ
OEYyQ3ctrLmLMQA4Mze3kwoh3A1Ca20vH7DCicpX5xR1DSyMpue6H7oRpjLfJEzzwPYC52dj23Td
hoXHpQ0jo9wSW+xA10uedDbFAg1Iry1sfYM88QzxShp7KP51ANYGatGniH4zuR1po9tPzXq4jmMQ
NsnFX9ZqoYz0r/u4HuakSV17uHj/RRbcmnWoVZWZQDYsEk2b41cdENiqaJvkbkizRgAihqGBl28l
lizFnZYJ/5rCEXi/tu89hnLmi/cpQc0nP4xZvCwsavLDyN/J13x0SFOyBzr1zsB9De3qolkp4hgq
xHaWijsgl0gF6HYNb0wrI/BC62sQ52JN5M6HWxbuOoE4i1ua24k0kOJrd2pMLDwVO5ynKmMfiQBm
nvQC1YQSrmg3G186Sa6GrYudjJv0DelJAQy7ZGYuOsXT8o59n6T0L8bekToTxD8cnq149FAzx4oF
K6v3zH4me1D99af4rqKCgdSiKvYm0Ivcc9s57dJ9KGyyxiLebiSoaxwG6Tq6o/f40GfzQ93uXjyB
6yuXaZPoZYWRel5eng6YpUp9MLOny+rIqbmlstf3BhjEagvBhszaMlRp2ZojPsQSYil5tWPZZ6r8
E4AuSndSafKgL089ZSXdQa0UoYnu8P7cVFkxygngZ1pZ1ZpjAhwolecPAyHwcCbKgZRMXdF+NtkY
yc5sf6/g/86D1oj89yYMzhAvwp7j9Q/hzTRCJwkkd09dD75KlXG0D0UGKCY6Kc73C0yGWQPovbCs
gQCur0UygRSPelF6lBucY61Wk9uAN+k25A+rgiyCA/159R1krt14Y+D4rU9UOo4IgkWheCWBYfvA
Fj03ZUTSMSM+USkRz+KyLVCY2Wvb5hvRYyFgVYmlV/Jojhk/3uRkai6mRUN54OybSAwBnZrcfvXV
rkhqHBCDds+lZbr7sQ1D523JPaxdzWMbmhD4nT7/on8Io9n0TcITfP3hqve/B6ipzU73ZwAdPy4f
nnP6nBUDMoWdppbB3NvoiEdJOMcDEEHTXUpsjvoc1S91HVuY3jJzG3SuSFKvsqWnlmySkZhJYwhw
FU7kQQFJo7yPwl0IpeorsO6RKhRVfRPsHei9CuLZ4mYKegQGcEDZuy0pGGvUZmdGcwwPTW7zNOY6
kpaRUQeT5oVAyHT+eL2Uk/qJneDyiiR50mdW3v/SyY/4dg6+in9LdfCJpLbmEq+4/gp3NCH38QCG
k1fg33LMuG71YzCwgMsFYHNSMXwsF2MuX/9e0njEp4pqGRxiaQYkbj7MaL1Wkj9Sc0JE/u+fa1/3
hpWcURh7KCXMMcQE/2S5aW+yg+5KBmu9/RgmmBj4jcry1m7tVyXH2rm6bXACtnVzTy22JIk9kI/Q
d6edrhBhtBcLllul+MVWONyyfBM+dbfi+xISl5rRY3zLQLVMfFIK/+pmnTboF7d+mT4NCx86dPIF
rMLMwQMRywIuxjWEYw0d3UzQ9NH+260hV9GzM0fgy7u+pDldyI4atUSEhWnrbArsTRfGM3jasK5b
NZs9fyjdjtYI63hXNCB8qql1w41BBFfpoKAZe6qLClO8Ax4hFaeVVtZrp34TZpL85sQzkaiybyf8
wBE/hXqqf8Af3PoTAXlsQLoLl5laSHNxtf+WFusVG7yd7PYtoQlhDFbNWA6oQwznmEBFkPcrY/+2
CxL6L6SM9ILsMfN+gGY3BnYaK+2VQRAz4rMWe9/SJmbpLT2sVrtmZhabdwhotWVw12rAb5M+LPUW
z2AFuzHFEdb7NHVP2NjsfXEActTSuM3p6/Wk7mSFLScNfVz1Ijwg2Y4ivdMXjYHFzOoCdScXMfR2
UfQyGssC8vkv83wd7yWbbMzojuiawR5M0vf1Dq4h1YMhnJXTo+f7+P45z2Oe71EiJdNvXOArrK4S
RDFh9caX5ZdiymzdYM+S02P21131onwvWwN8ZFltOaOwZCtURqvwSniD0KoFVf2QQxlcHutbjCRs
vnTzdTUIIW38LsNOUxZSBfoCXMLLDJuUF4j69c9ozLct6/HJ71chktraqq816wCaJ9z+ltFMHa9w
MqRnw/MaUlA6MkA+TIk+vk9nRLRxpLW8/ow6oUSSRqVVJ3O2cdImfEkksFBdRVok8or6RoGKAa/8
jKnPCGC/xsT9TOqHLnSH01kaO90S63Yp+dffd40deXN5QIeuTrozIgRh+BOdEhvLMY6ARvhLLKV9
FjS2M/9TW1+F6Npdd/nzL2Pq8HIP1+e8BjW6dOU9/v+RSvi0DMt64gJZk+krFQlKV/JEZ0c02+aq
PlVUUI2FxdBxsY3yykqgv9iysyafp1Zzb4/u0Wj3NUP5ra4zHXGDC+jnWsgi8UqpY/B6SOGqVHGB
CZn7W+ecdMEt9nEZSX01ejoOZZYJ17CMd3hOA24eeaz1RMC5XXmqQTlA1k7YJkTQP3+zNIcWejRm
vR7s5zCfJm4pzlQSggg0Fmgskj7hJORwrFFG6xpWvJAqEEYpOw0yI6aWP8OQXfjX5SZtJPigcwkF
XqilispsZgIxO2OPYHzHGboQzfhXodm2CWEexLO9J91sq2ldDqO89xU62OwWe1z8ovtOblfdUBit
SSMaLQZaX6OY/wDCVLv7Tvwlc950iVTdWpm/oNxjrqDg+ztW/F5xdQqBLNt5RTH2Vyn6megLJIEJ
DH2GEfozq6iTjCOaXQw1bcBhg/B3LCipZdOmmy8tpJwxde2sqyTOTeNyfN2z0RWE38KoTTNPSoJe
BvFFSEZ5WzgLoEQQ38xuss0je5F5DLlQbWiedzJgYB1giOIrVyjxJ9j0rO7wtzmFNVU1Wxe0Xxhe
0Wkdlk0hlQyPqsVG1+nJooQhj+xqG7gGdQaA6oKA0GhA29JoQUbXTZUdi4UsQi9unVWIt9qZBiXc
CC95tNhyevr44QucbdxkB2Y5IgiEtZeNxcza/AcAP81PQDprMrL67BIZEDDKcMyzJ1/S4+Jg2A75
Th52MID4VO/lM/CRPooBkbe6fqwojPkIiV+n1t1VMrm9s6kt+BhdWuSmIQH7/g5jOojKred55TYz
Zcl6RZ/SNBooTehshPswwP8geW/FTQhiX0838irQQ7LSd8css7lcraCPsj99eG9OyLcS1nZpa4og
BtDhqv0gwwHmYVE4Rd34hNlaa0oy2Eu/qvdvt2qFSk2PyFjxCPVVMlRqfCBvUuusar7syXg/RZHI
eX27+OAYOw92IJpNiEef7OIbemF3pAgdCuErSYUmXFCBfpqjEpSY7taHKFGYVuej5RASUz3PcrFL
YoshA7IxmkT9EnYVo44Rq8wkmAcLYmiyucjd8sTszobaBu6eE4j+k/6qEN6K/fP5xBU+5t5NC8Zb
h1P23HgXBsUR4lt/CPIqS6Pj52JwfWxoDYH1bNYZkCNbozaWQv3LBDSptDck2eEzKsXPgV8sGp37
oQvsl5UePVYlCBEPG7zRa+xUKTcL10glr2oADmLgq9YvQPfHN3/NTpdKjqu+3hLKTzTtfN5uTofx
wFejdOMNkYE7Z2P5MJs33rH2D48eczeHtPk4LE9Ay/jEOyM4cw75mAxyZJxJr3pFAzPPxavhguOx
71DP8+fQ/2MEV0AlKrzKYod+/o6KYr/qebfI1yRmdTLvb0koc+lPTwAOcQgnL4kNTc8n3Eejciij
y2hTJXqq2USEGRd95lmC5lYWYC0M5sY6TdJdvMpXrEs34J8Rr8XE9WQdCCzhK1MJxBAkMqQEUQTN
1/DQIWt/RlNsS3zXep0LQt+AgIs95LEZpymuxjm+DRt6QYefq8p5QzR/fiklhVT7alylyOum1eQ2
fNDh8FJRi723DYMipHk1zFgE0oZgxRMDAiftERXDCvdPTZG4qk6Y03349btd4+LlDQdESjnqbh2z
D1mfCkv6mJ0pQ0jL9VdU5DPlnBPH3BRtByks/mGR/qehoy2nXsGx1j09fSIG8KZ3QLe/hUKwp4aM
f9w9ewMr4yHiDjd0lpE26VlD/GjkqFN5gmapQhcdL+EWxdrneVwTpFwIi1A0kNX0DL9B/JXuxaPY
HUX7Z7l+qUQUv6fxhWaMv8Hrr9J1jPZObXLu2J8AsWmf85Gxfd8YL/AAP+2YFHoimP5/zTbdWEyf
PxbQU215znTNwSJi2olRtC/eowTWeVtH2AxEmFd0E5Vama52ONZRBeehWa61SaaCOopUGox7YRH8
D5gqQQ8i/+rLZfdw80/hKVJkr5stuLmTWadjSrPaMBsIZNLTMbGUKbznh4zVywQ/tn1wpAukylfh
H7OYcwHHVpbB+cFc2Ajyo5p9TdkKt1REN810o6dnTkBAR2qEghZbrfhMDz9UlGUd8Qu6F8q4h/Ht
2qiW9P4iM34jhz/LmgL3I+/YoxgzHJC+Uv3HUq1PkSlDLWdXswNB/10ovq8trnLtuwgp421R9E27
EsgeBrarm6KxO+4r+8MitjiFWGC6KM08vsvCdxFJXwLtw4meR/oUTRU2HTLmyWAGweffWWI2lwP3
N4NTjwAdpSZTCSmY9khaWODso1XtN0ixRHKMNS6gG9BD4bs811k4RPGC8IeY+YxeTpPVUZS84Jta
4zQD/CvWvT1ODf13gOJEY4rh7o/L+6H0UGE5uHnp1pZyuIZAd9Q7CWxtaYLZRvXfNWwcisK93MfD
jbBdIUWR2C9w0dLgCBGYOQoPO5ZOMJgcK0cvO4rM+FEvLt8R7r+BC62ySrAPHArg0GnhA4W3OL+p
67xmJQw9P2mFZrP8PWLyZ2J6dvk5igvZJ51lzBqHZLCBcR5BIy9Gr1whUHBZ1N8MlKnyg0Oi5xP1
tz4l3IeUo/Li7EJ+WOUI1xmj2ZxHMsB/cFO5EbRo9DgyQh8G1tjELFSR4toMo8WNXE4zlnrh29hw
hY4Vr9NvZs2DYr31KhSM8GXgs1nbnGM659CsNXjknBkGkvLo6EuXrJmtijh6qO8C6o8w+L0V0ehU
dVqDv5CMfBtTWAxqciGID6hD1aJ1qFGl/SLH8bHkWVsHM8W8qYQIZv4PgK7hGlsnO/PewskcmzS2
z29QFlJYyYwT1UN3a+27ZOxqpRe/UrE+WhdKhjjvSswxc9NEl2VGktSH5o9DFZykd6rrR6HRExX+
szVABtIrsipFjIRySZVhtoP5i1EEC1U5gH5tFwMZegrO8vxVyMtTF/fVNGiSGp4HiKXgrKKmLCF4
PjrdxPN4IjV1HLEgG4+DWzFWbLYZXUoDlTRr8plpF5HuSNuGDdVC3Dzj0ppTiw9aTvuhU+G7X+//
5NwVX3ayIcLShbobpSCQ7omlTsmKilU2gDKuJRC4XzrdSfD8f4fLEhS2IU3i6xKd52LylhLvG6Wa
e35a1feWmMM3VdutWUcgx06Zf5WMF5sqcF8xZ/UgWzWX69vwM3U8mZX4rcKNdb/HEVLfrQVshcIU
JGriyP1D2jerWEWhctuYmklCbrFaPqv0biNZnmaXj5C/TZE0M/VB9jISopXLI1BTHlSBEgGP0H8x
e49fhZbxLSNNBLnoXsgqOPjVLrpgUmPfFOt7P2Qx7cClMNWZKe4DKr/+fDccX82thgEPaAr6fVJQ
XbyCpcbcV7oNLTkSdxVIubcYXAQNWBDQm/LrlRl4ISwVJt2e+hZQcc8PESACsA0ymU25ep0uhG++
0Y09POxxG4J9m1fIv1NdixaJk7Rg12TNZeISb0gC1KSOLGb+V7iZ8+UoqnZz8gtHC0/KU6awzT5w
bkPniix/Xe8YF5nKpT/0sL6rNAZJuR83qvfUIG4qfSI7tEWgKJY8X6U3Bo0KChCVPrIJC2FCJGQR
/eLYuAYOx4JmReCgSTWzvSn6exd0xvYCNLV34FXrx6Ja4pTwz+45/itgt04LgfHcSY3NJj00IlzZ
VjRkJVfwlsJw2wW6HZC1p4zo9NitkCWaGWylrJ80q1ZoQUx8xptmqFIFEA3g5FiyrSwhsk81sQ0R
Sirwcx+4zwJqPoWGYhSY4BVTVo5L+NHUCNS1ndSnZLoQaem1iEsmIU2m8J/+31o/xSnNV4VyWrR9
vi5egM/E8TKciKXJsCS/Dp0/Oz8K671gjnK5yUH719pKSWavZzob2ikOXwk0kT+DnWxodNu9KRSV
YBBM49pMf9w6LBn340ZGwF5GZ9ItTo4LNlKIdu2Melk4phQe3Lgcy6WLgF5e8YqIj4e+BMSKnpF3
AIGieuBLhvSgJnH1ag7CDwXfafQd0Tgbrhyfzan4XsBxw+lE5/HkSzuzkLSODyp0m2iiyfKTDHN4
rI7lQpoSly9iKgL2VNM5Y7uWCO5G/uWvxHPdfjuOmzlwveN/n1rnh4LJOJxbLHlhLmzohTTI60yO
KRMbbJbPmkgmRErczNgPrnMzLzpiEaW7yrp5ASBuNgoxKwbwzEKrWvtGC5k7RwYJmIhMFhZ10IPn
iumAPGKPJCnlDDNGdeEskk20sP9lLlodEOUdzBhhdFhhloLBXMd54wavLCTZQ8b/que8RRBnTsqi
F7nkVHRipXJ/uIgvlLouRhJOd7vTuIFhShIO+r5EFy5z8/S3PLuZau+MyCESWerY7RcR2vYwwUch
aaYBSbLW0jfItNZZx8syVhPfX6uNzdGONwVChb2kCYtn/DvCdltyQiNBlRCe0460x3ofBtDphM4+
VoqYcmPQTLLK6c6JpRUxmHd9tWCC1g+r3oiJdCEE8njyzL++vLNx1M7Ba+TgMMmZ96K6nv+trhiS
hhz7v3hzGpEr3xe7WZnzyFhvKZebEdkQUM1JI2mgWnbdlwhTZ2rVlshDR4fkfS8M5kviWhn+qEhC
uCbTYFvFjde7Zy0y/eGMvqYuS8hJg0jnv4WSJJv00V2AkItJvkcfM6OCTilN/qsa0F8AZyUJ7/f3
pIW5t90nT3VFUGdzX1KxnWvwbggMqTxqoBaSGO2JJNtdl1SMk1+exTDXmrz4TcI3eJP2DynA1wpb
8S2R3sO3Z3WUqRbK3GMl1TsK5979oOwaeFNaoUjm0ePN+gacXYtBuyLEz5FcNVwUlfMzfEw8gzhp
0H728Hr3HZvu3xz8ClGzCQc3aLHYFM7t4SMRqCXhiT74ZXsCdFhNar+ctkXC8P30tOQUSj2V8/WC
KYbFkHN4IjKWieyIWYPf+gRo1zZMP86WgYAw0KjUs12Vha7IC0uj8qLbvsUhx1QZ3TDWbXIBKuEz
ZLH7W+C8OQe/GMCCyMXgeoHo7rZP+dXqPAAOnTK+H4vm7KiDyrEpArxdBoYodulh3kS1G+e6mPP1
lK4Cy+wTVuE77J/eXiTA7oIdVQK8DUn9ijwr6cFSvwrmizzZ612cISe3WmIkKux7aYFbMaSmVzwk
+t3iwWCCoPo0uxkAAyHt8lKIwUMdITR8VzqZJ5ZO5ZIs3dst9Emqa0ocIuTUUdhf31ZbD2EwrJdB
FqaQw/T5p7nFgc+H8wtauI3oqVkx1Siz3SZI1MpvuUC+xR9zjNncLRtBqiWrf0NbSNR+uqMfnIDa
gW32IkJHz4U2UIkM8uGHP1ARlgEuSJ1BPXWdIOQOjRw3P9vb9NZsZcqeyIjYloHRmjtfaylvAhoP
B1CyFCwhZUAGfbzK0COkjixxiqQki8a1PBaNqQOzmvATtn/eztXcjfQhTf0/fP2sXmY42a+4ic+s
4zeG5RNxHocRsc9XR80lgv7rqUdhmNEQSsHVhSCiuoWX7qpnnWO9eGFXtbLPsU9IwLslG/Lla9vq
c7CJ9+JCEmOf2uVddQbrelen46uyPXGnUf4ADIdaiBU/by8drzw07YLSzCQxbwidqh+QXkPFmhDl
LxBKbK56XH/I+c8icX33XRhLWoACGKLeCOpE42HSPtmZiXdDx6aST+n+Zu4GMnORJmwtkZnqDieQ
Z7oPXxxN8F+KmurjpSbN/K5MYFu8pQF8UgSkkrhnGz1vxPB8MlkC59a9aRAOAtvSJumQdVFyBYk/
JH9agk6dG6RxCOByYc59yy/PJXSyksr9VJqaF1jB2wEt0FATNU2KuN3rqtWoqidDHdrj1BQiK5xG
dIjPrwiEeI940PIk1uqh659vYwmoVQ+4txNEISmS+c0YexZVvxfFj5CyFiiaxS1QkFYV4ubS4p2H
I/zVatO0i542B4zfPLEyu32S7MxGyPlwb74iMWlFUFQ8vqvtgxhCeBkrikspTOpjPDgmKok0k4di
mcrg2R+b9UNhX9KtHN5IdvAaVqg6FbNeZyDRzyqAJ5/h23pjG7EM28AWbg3Emox9OcttMKy0iY3j
6Gjw153dMiqsCD5vZ6InSbv7dz3CPUZbr6WPrebHshzESJnFrSjm6ng9QZ/TgT1MR9HrS01Z8pOn
0bTt9ikxOUVX9HUbZuIzWYIWoblCFYsC0dUeaqIeipWI86LWzva6oiZDLEQiGhFUHBle3YECRNyy
4u23yW3HsDWZjcvliWdDF2VQh41CPTtkmBXQQaTf9kZ6ohH7hCY7iOTlB0cccVD4GRld/3T5zfqf
ug4jq69YWFnDR4LeJzDZZXyzzB0urT45aTbC0sYRN38mByFpIeXE3KSlfHSZXvUzWyTGAV6dNE0U
3FjZCpS9fkLsbhnwnzKsQC2oblesfU7qkLDkAMS8Ra3LFh0YaFgAFnwTFcSicNkMH72ihUfdQdzs
GMKxxnbOKeJGf7Q4ErM3pmfnmpo1YFFfuoAncUL+ujb7EhOzYtZcpTzbun2hpqIdVM5J06bXq+2i
o25YQxtD9Us+c89AuAYSK1OColmZyVOP1/CH2UykXUGwgkOXZ1sFGhHvoi0Z6q5//mSi4YqzYOez
Ahv7mLw7E4RyXGLTkATTeKLowdgJMcPSOxq86itaIb8aqLyG7F3WiBr8ul2q+qtugpg88GXnckbT
bgsGDA7Ozh9Ipku1CRfWH/vKDT7DiyKnCT3cYK+c9wP+ciJkFZtnRp1gf1xH49zn5K8rh8itjeyV
QYr4lT3azlvnK6aWnQXB3VqMdar6Vh+G9Dg1p+gdZ9Iw6vzItWxyETS3saN7GuoH/mzVQ63ru0oo
wOZrEF3OvHExfA87m/5WkahSKwX55Msdnd6BmuPX2Pw+rCKpg50LwFijmgfKk5jnHxoP6tpWyRp5
E5zbeiibpZS3KgLBfanN794t5ovR0UqMyYGNSGK8DJxHeBGybkQFyi0wV4FzeR51C5/e1Un+Uioz
7Zi0ZOvhh6qQI69Zaxr1gNmwaPEUpO9X47O8AppPzWDMJgD8KT+7J7DpztukZBhQNx8EUGJIDnsY
dp53HgV117uaIT6f0DNYiu5DFoCs1vPlw3gWUKvVuj8I+uAhkHuvrClhCyRYCH4l5AbyLGXb8vzJ
xaYe3zDL8Hhoh6vQL5G7zsY6JQU/od8WfwFmrS9I9eGS6mo8LClGY87RsbN/weK0chp+7JsEuWSM
dev4wGJ3Fel8OlEEmbCvc7DNPvC4W9+IcqzGu9SI2h9m5Rheg4yL5AjmbHKTFIr8rdQOdeXH68nx
KdjB5qysDb6xRBO+yC1rxrk6Hml+Cd7uwTbC60X+52Y6mtHy7NSIvGC7rZmXtvXEiWQcl3iY+vv5
vZZr/dcyoQRPT0nkstwSuFiX+yGIqTbEGYpt31AbuZw/WZ3iCaw9bwhu17lTHGoOq8xeQ76tXEGJ
uCeRH3IU2QCtM8FIJS6lKustAdRcNf1YRgfavWhynwe+dzh21iseXvuJW6coyTV3/uzs1kzIKwSq
f8T8vzeONglnAPwnCenlhaPh2B+PgXWiUXPV1PfQW/fDkhirCBxj3wS0hpmbrgh40B8DP8KHWjL7
jh+DgoxsneHKMVVS9tbhxdCIGfH4uxj47sY44vin1DzhIxpzQ+povtYZUU4yY1AB1u4EAHZYrqdE
IMd/Mx5iV82VrctNcAsvjttbSg1e+2ad+or1WnljOAz4nZl/CfrOQxEtqoABXAWT+KyuoqjPkToc
JPrnpN/A7uSOjAvAbZiPGKucE0C9+7gNRv7nK/fEgpN+tICHI94sNP3/4wcsYDfenDmjNUPHPXU4
3m6CSzH3MecWyDokWwDQAEae4+bKnpkkTQTa0wWqDwCI99Ak76Heim7BdHLI6Nk6+S+Hwr6rHpYp
CXcqiZWAmiwWR0GQnP1LCEiiJGdLfqNi3lGTQN2I1dHvcAtCTip+PQsS9a4Bv9xAGhvh5lsfqRxW
JOmDUebg+TQL2YoDxqxeVFegbZL/G1RCNKU1FYdEhrNs+aW8/ilfvcLy0B8kjy1tCfjfAfXnkNeF
KUfBGobKA922TRlvwwu5sep3wP3YH5WaMv4Ur1725empYnx2ukgFsC1azsbdvcDcFiDpmCrQyHFP
0vS+GyIeT1PNNMKRdpQ0+Hlzo36QVFFcAJHBbWnl2VkkcoxdRBKe7Tsm+li4xBGr5hDpIMcuwr9a
N9Zg6Fw70acU8Ph/NJJYRix5nJPvlcJX5ucbK/xU740oXYufyn2aclGafMljwYhjhKkPm48qMwmb
wZAkDJDX5YENUN2RHNPzxD8hZQO19ezFQxT+jMm8FMFsZwuYLV+o54FcsllKEMdUT6eLm8UYtc2r
dImJzP3dpT2E1na53RHymu+96mBOtPAqb5wfwiaATSYV3GPLpwa+e46/a3UBsY+qCj9jthWZHN1f
dpqXy7a+29DLPvmEKUsd2COC9PWIBnPr8E8/HXuCteRvhLZ2vPcOhE3P8p7CE0y97cQOYvyJ0n7I
3PxjCr7emPz8cPPQvqNqzMssJbFvOr+docBgvnzYBjR1THzMwT51RPWXYfuYGeslxB3cSzWMW8Eh
91R2mKUBX9VrpYa7gicGMRetXwgWtWNkjbAZ/XsJhuoUZwJgr4PhUJpfI+as0bRs11GkwNtQl4yy
QUGPNlcE1u/Z4d5WihuOoKLCKp0ZzYgCtc81twFBsYn1XwydFTDkM03oLlh6Va6l1cZV0SGOOwvU
iq1lCoE3nqL9VHNO0r3c3QqZrcaFoy7Iaqux/OaFJsDlH8XtNtmvDVAqDZ7eo3p1QZwGx4UHFVyY
EuRu0IiXoMfBUr2hsPacgWFC2XPlF8oFf7CD5v8ZTRWtRrJdWrsSBeKf4G4Coj80y++JyMHypSSk
v1cnimpsq3T9zXDOb/kGJjwwsI3UaJLkD95ZXcg9IUoXYxhWxj8ugO+8EV01Y9XTS+sCC2JQbNJH
/8fjWDHdipXVRe7LJ1C1T2A3jqZhix/xg2BS6e+qw2Uqo+Zs/kkkdUY+xpx/OMUw76EiJeELZXvT
1OXUlZK38+6bZlCKvnyw3ArIKyNPKABeLmJWB/3Y2CkIZMXZ2fOQg0w+FL/J6B6MbeyefSy3NXPr
WHR4FSStO7Tya1ciTJ2HbQsJklTIqILLeEa+zFseRlCr0obBua4Wh09mGFTPOOUsx1CsNtU3wgun
cRmoiNZrbkD5swY44QpNpgEguXnY2UEKg3zRoNk5m1oboWBfIXePhzAZPAh6Gr0Xd7tvrgYVMN2r
qbqNQWEqlpX8oz/rZaqT1nu5zjGFubDi/Yqd1qT7MwoBGk14B8xTJ+ZYf3lZoq6w2JAnrD8M+sB5
dBdxBwqbsLpvV8rLARIOMBRiX5/sXLAR4VjbIfzaSI39wzNsse3ywye4RmHprei4c4zUOp0J/FDT
ymTweAo+6Jf68Zn4QHP0oPD6XFgIWqddrouFVyMxwmqAzV45FMlvr0u0b2LOw1eAUNd3WUB8Ns0K
JHqZRO9qd59Z+u5UBUrkB3rQV/vxcfH8IEm88nHq00f6J7+5ahGV/LJsRfRTRmVmoScejDccWnxp
GKtgDYMSCad9+CeHDJt92iwSr33NIM4dIE4tTdAStRKIGpN/Wjtl4gntTEMBNkFXGARForuTd2Ss
sG39RmPra+BlwrGC8tuv689ctdEQ6cLDYj7azVodEbrT2aAOzHF7HB8GUnHe8txqaoywvVUJJRj4
E/RNKSG0I4BONla9hBksf9V/pl1Pld1eMMNiL5lt2ouywm4reN8tiYNTc2EeSgiL+mv+bDxAwYbG
e9dO7H3JlkdjlPBbizOsPK60Sn5JCVjZCwWWSRFhlF6r/Gl6ua2UVQkC09o0KNV7gHaIYzCrM8YM
3DUADgwnpJa5+kaCmmsf6m4p9mzx0BlJQZZtVxlDPFj5tiLTUB1tgEN5710oSrq1fv1jjmRAas+F
nborp8VXTHWBKHc1bmzBkguv1Ads7macPr/YCo0AORBD/SgXcEzVBsTVfGIgbOEfo2i31N3L2YO1
ORXV8aXFXRV/5x9qv754QX5Dx8BoAmjaKY+xd9i9mSIi8OUMY8lQwVrPUjA40u/nLQH4HeFBltxu
xfhdvOYCwx4ll6G6WVUhepwJNtDbecvaGfqC2wRfWzNBirlqIAWTW2p1cNbwOpwXZIIud5zWK8Aa
klCGTf2xS3T6HSfACI6s4AwVmAJibOM5xnB90rEKxkSiFDLLT2umw5CgPny7hvIfTOqxPBT9jg6n
W313hbn+azYtyxOgHtpYHQvxXuax59T1AQZbNQ9aOwABfplu0klB+0BA1lXnmGVRE9XRo2oGH0Hm
dUQSf0nAE2Lu6N0PI3HXblNZqdrrphzWLNCFGh6sL7AB7B0GPAvHoyH2eK1IaZfkesiOUfvKcXY7
n89XXLek+DIwpX/o4gPuv+XIGUzQIf1nUQBNB7Nm1HxxEV9lEIfJB8EImO6xiPYIMFcvkR7LFEvs
UWnYf9ArcrHYakRH6IY/nZU4dh5lGYL0t5/hmjZZqEG2Z7Bo0RgSYU5XUQmj1TOyXDK0z/oxk0j+
QF1na0hJ0EhbvPZJty4F8PmyY/6cTCtbrjBxggS03RtpE5wHcHnyGSe0hqjLDhoak7ImTE+YVHRn
Y407zkQf8IwVuF+Armh7iSA4poBwVg6iJbaihg6IHaMEWfrcwmSCIGkAk49Lfw9auFgTMpbI/juQ
ZvO0kOUL7C08ydbWtVWjgSqShJpAcV7ALLoF81rqILnAJgWwQhG4kz+/a10EMQrtvAOLvsH/i1o9
eaDVGorRYXPjyHnsOXrcf0R875pWBpLKV14EIN5jEoQpuLBD5eM05+QCGzgAQBgsOirJruXL72dz
ioEFuYemlDZtsUIPRzVojLPioUuOeXfqPJpRoE+QGVZkPGa5GKQPy8BMYJJfLkb5sPePZiyWBT0M
q9wMxdkhdY3A7mnsfZRFwsAyOLexk1TMJcUPILDXBeE3F76xrHnbSMs43EYVjVP0vEO24QUCVwBj
bVmPX7X/wq0kfna/vGmGUFT2vzYAxJrVcZzzbyFc3H90rQHaGpRnnR5UmuV3eOsH/bTZ6NhgeWpG
AW5EGeCZj9B+BPagKXGyUpNss9Vy/4zZygePCQJIX0WcWAhVUavrJVumJXj8TGhlUIlgrIZC4+EU
vF6xwT9tTEbwR8A4avJS+BkIcabjnySBUxcol2skeR6AzEWA1lek7jloIOtP7FHHFKrfb1Da85Mq
Ckp2TzclkbZCTYb4suvJGUadr1I+kY2iXC5d682cTk57APPzBak0ihUBdDMi1Q8FCczu1hYipVzf
WmBs4zvi2oPEgalTFOkPTtcNpO/fJZ5RI1jTpdmR67Z9N7IfrQgU8E6UPLl8J4Z1AZoxELqDLu7w
g4RBxGaq3Z7e70BvpzYV8Y7Gyt1vzCUbVMQPlLk3fdQtjpK8pEAYRUZm4trwim033oa2v00rbd6N
O3TDFGJ1cB3vR8fP2ooyIhqyqPsr1SDB8s/05A/4b+aceR6x7Wz9MLqElJowzgp7lsd7AUjCknkO
seZ3gv8PFbBwlZJwVtg+bFxAYWuQeWxLLpT0df/deE2iGjrxnRlarpFT+3T3Bc8BHlA0rBhu/jeY
3VyrLPOWDsJZCX9o8QyK+w8m8aQTZE/hnZn4u9unoCt5GezOIIUWTkg1UVJIgBqjoh8RJgutWDI9
nWsRzpn/CSiefSVLQwpdtYvwUkd6kOtd7CraRlfv9k+JJ/bvQJxWopsxIxMAWRHUsoFsfGUqs/Xs
pAKJnyjSiIudPJUyTHqdM+ytCExbIISr5UljOSMOS1xKUQUAuGf8N7pmflzBRy/xBqAh4IuTIXgy
CHCh+4u+8mtIPQqpxZclQyWaYBGH5HKcvXm+7cRzhHHQDceIaOnmx2Zp3Q2k7qRdXkk39nY5+37v
eN94Cd4pgAN4jEAUApy2GGQakdW+I4gB/XGnQOAySgoE4ovzmhQ7G1otFT37U1xik+uCjwRUT5ex
v221TTht1p8u5BV+s3KK+HOJaPwkGYMAr0CE+2faMp8qurb8bTBBrNDuGYI/drAL20eJks4wLTLu
wqUIrnZWDSHhdWyqDuxTC4R2iIyeXRFDDtcrRvSebRvgH1B1MT3XrkhslEZm7yaQ/9hEieso/Ibr
M+CxoBhUn5m9xmJ7k9UMxNrUzSeS5pOlq6rYHEc/1J3Wb9cm59ZSkjbrms072JRIKMg5Un5WYTVO
MV2uHMYY/aXPg35vBBTOXL6eA7EN1T1Q1UiIFJiVnw3KjSYJuOMpmcNMMA5nMwAPSOhijOPpuZTP
8ZUhNFtf9tmEka5vFQOpDXDDAbNj82w2OSHz5N6kDW/9dR8VN4L6Az6Z/Vx5ENC+HUe3yayNt9nh
5c7Ml9VcvpBsISaur1kglDTBuI259JkUktWwr3ydIw+42a0pFiXzLV9JizE9Us8EfR4zqSaiMWEd
FkYOIa1ZM/8yvy1enTxRkzODke3dNsGOguOHeEoSmh4YyrMKJE2AHmCQ7nZSBuHcUDzMDmAvh2tJ
3dKAUv8rqtGs2wRS4GNzHjdKz16fw249rXoBvhTj3y/5DVowqjdAUnTWWb7B6Gxitbtpid2DS563
vH3VKwF/+ehzL2Ioz8MPUeW/sIXcGbLf6A5jpeFgwvBCofVvc2iXb5A6eEXX34NF626qXw+3rhOP
tLqrtZCZH1mnMMS96pASkN3nma9rIfjdVPwjAKGBAJK4rYi9xK5GJSxbAAyYN2JzsZ18wjPF26rL
8Gd8vgRySDkvvKhWvz9hti4qecpI/Det/DbqDrZ+nS4bBCc6xfPKUOp+7kwnst82nGKY9/1Hscmn
VcPOOWBvqLKjFtnm6OlqmFwDjTMqo/8i/NdGh4muBkJJ6GmBocFQnq1Yg7n1Kl5FF+el/dPlrc9r
4wVVE/nfOyxCaueETf+EzUCHQYeGOOGvTpbfK9Yk3HKDjXrlDKNdKcBlF49bEvqhDjlkSygT3tXL
gh8AIZ7lXeJE2qlbuPjXIRixLiSlsvX1BHqivAsuBV6gPrWKWqXNvf9YJvixRRNz9aB4IfNjCCSs
1q2q5r6+yiOqo1TGAQHyMcKkp4Q82JEuZFb/EjH+qJFfoPfnVgzPJcfszSIXufQHC+G5Zl+dAeeq
rjxKaDl0w6my5bmulJJ1lhFtKzrHnzl3tqRiB6CfdyQtZ7LAKnFGBiywbMLbIL5Dgsd0KvjjH5S3
Br/+8kEEv2hmtzQ/mIoIr2jb5AGZYXyO7z9sfjtSwrBPWelD52Z/jf7ApMYarz92hdQZVZLyovKQ
JlZPE8Z3DifIBblrN6YQ+QjJmuK0o9HfZECX4cQS2MfB+TDIIMNybMHZ8iZWtUPRSPeOmv/TmUdI
W44NN+r3aQjPLQzJL4OSvjqri6pBkzY24WyVVCpT+M54qeZJDGHtUCROsBvfFrNfgaZpcfd5qI+6
kXqh+3lUp6qgFC32Ny+zgV+lkMSdEotnEkDRGcTClTu0MXmH10PXgrBGzxJnIGJrwdAWwqtmqllv
Jm+nE2aaNSVuoebPClQgRXbhOYwytBZkszTqOt4C8c/GwgRCJ+Tlp3UwHmWM12NyFWX/ORn8Q4RE
BDxFiLafxgNiVMWG6WB9PYozURUnyRmqR5y+5GjfRgLDctjKdQaeNYizPPmzXb2S1E52MhHLk8kj
tqjixFi3S9eLKEuPEm9qUYRux1ZDjW9GuIqJE8nvliLe3QnA2aWnttXCnuLTSrDpp22ypeNGN7m8
/zVtidC2FO4QfgWKQfpx/tLes29qSZwjc3GOXC9rAId1wqMQ1B0P32wwExWupRHu+zOxXKSaXELe
7uTzIN3zf02O1PgxXvePgLY2T2t4i4fjeCWFbCW54QrfBNNjiELVvD9eEP10KSw1BUsuwWZD8u+Z
8TQ7eF8U9KJzsZTneBvXi+3tko91ErPAgEOqjWTT/xnD1KkZR4DTMaufNUMoIaTeFedlb+FAaMiM
1ZMx+epMx2TZV34qqtxWIZnujRZm2h2n2nPqkeSFb6gk3tuFzI2k7k5BbCnoeZiYFdbN/grd366E
PLto2cgfKYN8Qz9/eB1xukVjiKDvVCcTzXnAV3obFCZ70/GmmKCTXdafcQyE/MLWIz+zh7DgIFHB
fMqJArOywuHJqWDGsJUwxTqRedoQcmOYnU5eP3g+TeWYTYgMGHFU1dHPJoHFlbinxouhUkJsDbCk
wFinJbAkZnWSTECEGOZh3nDH2xfMlQjJ8DXvJO/3FP4qSU1aMxsa82djYIy5n9H7hZKq+yEPrOeJ
rOazIpoBEFiyl2okkRzqfpRA+2p48/UFG0wVc1amoSAkDVVUEkxXU7SJHGjq5xLQ4PjriD9LIuwQ
ddfXAQ9paZLuxm6d41dFutFa01tMrRPObcs2ZZF/Tgfz7m8obE372j0YiTKlrdtvzIgCjgywpPWQ
gXQmbUI4Xtu3pWMkA/RXPTlSPhhFBJgxLTQ7ybXG99w30PCdnw/ekYZ6wwSMrE7yx5vwK3enKSJL
hqyKIAeqO5hsgS94k7yrL0cN3l4qvUnk05u6hYTeh3w0nbabu+Id4oYR72/R05+Qh2FjXB7SA6+T
pWLNmhh18Q/iCNb5XPS6gx5SuafRf7GRbq+C7xi3WQKNl7crITp+MGgsRjAKaqkJpTtjkxP9hb0i
FE5EF1CIUT53M9UWJW5s1zgrOhE1eBrnpjyJMnTSC9tVjzrmYX+y1K98O9S+ZTzjl8Ze9YP3hNJ6
lbAlqdG2CnW5WKHAM/tFP0NmEBxf9PEFPqswEoheZL1B0Feno+vZv+g5qRBLSzlrkLRyxhgbZQyT
PN4e1sYPWYl+nSPDwM/ksELWQd6a7Zqs+jQCohZzRM1GD6VjY6HhIh2xHlqgjNQ2NsqvKIBZsikx
DayZK9vQ6RGIsWgjwmViRsx52PfxCs1DDNmmFpgvxg7Q0HKCIAQmqNDQ1dxA968v1AI1viFsQs0Q
KK7K8YdnzQ8nId7Rpx0WEZifzvRRY3AlmgWrhsNmYDmN0KQt4ffJTQtxarNCf6AxgkRFpDa2BS26
b4krKzONEias4N5Gao7pFCG6bhoC6O0LJzKlSJUonAvkaNj3YJtbzT0C7TPDNFFc0wz4nvynUQqS
1x1gnrG9AOIzAFM4MMMDo7tSi+PXc+74OVxCfdwDSEHosXSbK3r3Py3FlxaRUfGsd91fmx3VEE8A
u6npD91xh60LTaya6c2PFKK73RMj0S4GUJXp3fQZsYbRTh4FFywni/r5nFZO7m2iY7k2as+/vYkP
3Bivinbg9xkalHxL/tDMWkIVkFHToR/+aTx1DmLjGGJNgIu4UIeF32T9aYATl5EwYIDzVUL+CRZd
If3zeixhuePSVpZVh/uorYDIgqnbA0+RgO09xP6beYjeeBcMfsf1aEPdXYO/zCZqMBM7pvw4kREP
ZYd2kdDpOVyC1seiurSHsVvVqMnxZnOWf3Kr8UH2TGDnrclnajDdvaE8tWDSehzwkPLiarfZFX6l
H+EhcA2b6vqMhl/7i9dVHrAyJtHZmj8lxpqmDdc4oazR2Xi/4P0InshxnEATjq9UcnKkV3nNuRuz
454fXuns7vOnCcYPf90tK42ZGQ5Wc62Vb1S7e1EV7RH+gS0T+wB0TPimhII0NDn4OwRmXAfiNXIw
mwo2ivMu/Y74HNaK5uZGm0SxR1VaxWh1UIufy4Znk4cpy0BiduVLxu5MFL4n9oSfHuVBQJj0bCJC
SsfKmRk7TJdDsy5yxPiQw3Fi4Ng2NYoqxDg+yNatvAnh30P9Lu1egUHjOKqpvXfpxyESAqqdo3AH
w29d15bToZ3eH1WNNSQN6/QUv6HecKJ815qQvFq4qjBPJiijhQHE6vMGQF2b3XiB5Ec4nivBYDDc
sPl7TqxILfrH9yZEOi/vvXSPTGpqSPmz4JbuBWuugwPSuSr8aU6ySbF2Y0qErF99D035FriS8mQs
zVGTP+U8Dh7cuyRHxPq61w7ifPrb1V2+vR/voxpAZZ2hZtMfzMcQYUVlV0zTIRML6wGVW/d6R3Ky
wXDMv1NLotMzzhCZhf12rq+7hSs7ryIbhrh0H1LPAa4woBsUWWpWInA5usq81P7RIuk6JqPDB6Ym
xBba9bM7X7wdiJ4oEs3whGAfq+khKapqnX9wkKQJgRlcH+kdfbBAZ+8WpNASdUCNeoqcsTnFd2RC
7+uyek7DK0+fBKttfc/IweyUsjHFd7JMiGMIisxpf1qB5Sid+hXjAFx6O/+d8wXHkoRddnqxTJvj
SKRY8YpiEyfntalwmsiVM4zFVcrNN22IjyrvlbU4HJZ7ozkwRdPCqeJRLTdOaBf5zTznuKCamsow
z+jpaSmbGTpWmhDczDahwD4yRNTO+urDoVhfhTC+6UGm6YGmLgo6hwBzMcr6hD8VKW/6SzqXOpcm
u1PQpg+4rP4kHIp080fubDrvuGiN14EiA4zjkx85t2q52ZUo5usQzARbdcW8/FVQFwb3YVw68BEz
hJ0SrANm4mq1KwkZTvS4iGKAvON/Hx/riXLHjJgipjFouqP3TR6k1/OSFjQz1X6CK2KqR69U9QGD
5gyv4SjiRRMdiESlKbujNH074GoZPiHR208n5n2XLWRGubZgKFyviVd3OON3ipBlTUORoWCSExNl
zhGdOsuLZPWBVZF1yYrYLHRG/qC1PUX2kZ93x9pqSjgrO1URMbjxTkx8kTdwRtzG3OD8D/zeqsOO
2wI4TYTlFl8HtyYNS24eGDIYrHWxD84CtNaRHK8GGGSjNDdXEIPl/MvA605j8ITI7kIQPwOGy3QY
YA0Xa9rQINn/3JY+2DivI75ciTrFghs5XGeSRuSaqbL7cEw2D8NY2WPKvMROdlhuTRDw1xzW2iHX
4EaFfgDDjJctpXeRNhI1t6S/WnxXosu326w36fPFALWHkrWCO4Nj/Nq8DQ5B2G8/LOniwFud/2AS
8UvxqnIpAOZuA3iUJZaGlSYF7TksMD/1SEvG0/YexEYMA0O69dUb5uTrq7Y3cMNgAjEP61UUf703
FUr1GHOLB1SV6ayFoPznh7dD4TnEZkoMhnwq+n6dkpsbLDqM36I3EdCTFzvSKB+K98NB2u+0FK0g
pP3nHPhqfnksfFsxKHLJglPhziMVRxE/DDMKxE9Fgoqu2/w6QHSXcXplDWKCN/R7RfZmmW4wSeOX
3hKKCUJ7rRlLTAVYPMKIiDxKBJ3oRj+FesTZDuCvE1fmdRWq2AXiw3HmiAvvo/RFNI9eTFVvAXYZ
f0DujRsaZqSaesXWBmGxj0GstuOQZ/U59e8jtayk+/DWe+ncNAhKNf1HGqug5jXEeEA8D7UnkAWN
Y0tReRYNsT779w65KWp/4XR2WstIP/up8THc3hzgmlKXaJeV/e+qhQ4+9KbRzblL7nwE+Mga54Td
PzDtNud7etspZ0c1H7eHl1778U7hW7ZYRyVco65Nqpe1yDc6uXsMb2Vuvhp0bczAUpsJWrswbV96
dJleWFCkqP37BmPouaFlHu/nBC53z1Ip679c0uIu6Y6n8gXAbsFbcYMdczcwmLgTxc8HAqYYcvyB
ja82NWT3bNMBFyXTDyiesrHgfMy8QUu03NC3FafqO8JgQ+2ys80GLXDlDyah539/KxtyYw+5CFsd
G6nCNZ/blMWiGM9eV/UzJvtWYyKCWeBDhsamDnIzfhrJ9hTMvE2cG+NpN/nyVy9bfwPXfEA+Z02z
IfTsRxHh87clUzt79Wa74OB+RiX8obt/ermR7ITtWFhd8RSeGq6a5dir1HVrpnQk2wzURh61CUqw
pDDtnUEXrUlVUTcarRNtrIysGDwU5f4aHfNPSZZtV+yxCWYK/3LCtOhlafcxC7je80x6iLfVqagv
BmTzRFzFoYpJ6Y4pwWTUXzTJHVFhVksRXujwg9lW/3HKOA4Ho9g1Ke+2QhD0zf2LMwJftEw0iYof
LorbSP0g/8bLgUsRbrA20ynXcu1XY7ZpGCErR2CVU/vbXgt9i8m/85aKg00tIvVR4vjEj4qGKk2R
SEOd4f6rHV0oSLr5WPaV03MMzQMuwMpLC0LqbEDLf8d/drKSNgd8Cm5PnKwTMw33/VCrUorgXIPI
iKY48iDGnN66jbG5QV4GcedpMxGEgxMV5vSMUG8EEXq+0dRwddSxNXxaOAnZlcrV8KIiYAMdh+qZ
+vklc3fQPckyfbrRGOIW4FZpqAx6l1dLqGiuQiwAAGDwNIB8NDt7GfVEf111PRAvfldK/lYb3aIC
F232XI0tVDWPpbKZJiGt8T4FSlvem25C5+NJUgvKAchYUV6NOol5Y8DiOnaZxJgtRc9WnW38Z5rO
zU0KDusvip1g3lcdXxlpkhVFM+6/AVDg8WzjyhsYmXfNhFW/X4Ggq5oQ1QCOuExfHixsBAcjAhmZ
QS6ieY7hXWb7NXF3yWt5kf2rnCwWHjFtXv6XD5I1yfex+3YZMZuSrqeLS9HxlQLq0JaObFDXgliG
2FQ9DvkvoBZrBdQLoXmSUzB4BACiRJJjCQnDwfK09K0mIukdC5R1A6o101CsuuBV3/d7isZtSuYB
O8XOf98uRQJFfWwSB1wn0NigmQVOSfJd+L9y/iEkPC0l8YEvs79b7QpcguVr0WeS7O1LoEzLeHpr
oRapeuh/SXlVu/hcKBtyuJnmR03PhBBAy7z5/26+0yGdXdgvbP82/QwjkH+JVHdlHIouGAc1b+fx
PSVOSEW3vKLJNOqu6n0ATz4YgWe/KdVq4cjrSlmbtAXIS0qubNO6j1eGHA4cnvDVFFMqvEF9vLEs
QX/ls7O6C23ZKzWiAMeERDYBYgPn7GgqMK+nUfX5vr2h9vT40gRyBzvI57sWfMILBU0HnzQ+Uk5H
e5Co06qK6FGkeFDE28e2iGFtKH33zxyjERL2W//bOu+i0hpx6/Y0m8skABW+bBpzO73CAUjNPBmg
d7zX0Pjl+pxk8EUyfr/yPxPRKJGNFrtBJi05tsdFFjBYMBH0tJtzZD3N378e/x9OhdghVqx0YQKH
5KZnMlgQUoQTRfCCDcBAnb6uskN7caCAmFLExlf6jDeN077EvMJgyRsT9rhdogfcVhBG027hSvqp
+vxW/f2heUcBPAu0lg71tCXNo6N+S5DHssPtDdtaXHKt/UPEe6EvYGKMXnFNJXHmfvwF4lSF+Ox7
otZrlPNuLPy6j0HWhe3pEbk+vthI8Tho0phqnb40PD21+H+7xSnCHRLiDFuNBPVy8iokr6U5ms7P
F1kx0mzXdmq2vDbMpnqTN5rLrIWl5vkD38q/1eoeumsKcyyyQOe5oycPODZhQWlg02pxOAnJAvUi
LWzZh72GcrJyMIg4PwuG3HTq4lbeEBaQdw8+RlXK0lXPnTLWBKf1Cdhi45yG89A+Ul1BEov49AfP
4y3VQBoug9IN2vQ1PLwy8EZAwIRydH+lxkcYsCxFqzHfwFVinGHSDj9uOJjIhcdT2o9e6gOn88h5
NIksTEKMT0UUNmAs4HRsZHOxB0JuyK6k6aXm+fUEjjY8q+9P3JKAyjIher+Gf7YbvufwC8Z2AYMn
13E7i81YzXTwMMylhlJ/egk/0/wUE5hCNyYZtIRNt/jXoBe/NTUNV+50rRvG3x2tzXianEYySnpb
ovAe5A/nzxeyk83O3XULMyxWyVIPmP4GxkEUY8z9NHM5GccQLh36XvmaWy0FgHG4dD2ln7lGXfvU
pqXJhdW4fQrdPuSIRI5fU4J7wece6Hn35CWzfQlF+hf5XWXjLkY6eD9DqtKPWH0j7OPR2CbbCaYk
oX3aafLsWOPRTvdYaODwvElsNW2bH8LAF8hn1aZ9fV+ifec10I91yZHq2+99opD1kw96cswG0GyM
xERuup8L122F0mVUWSWJEJ0zHJyTUHtZ2dg56qpOTfB2zIiLDwR47uk1HZfvdy2MNznZD+4tjAc0
L9Yc4yyzDCoUgS6l3e9WYZVgoUPAIMEM5MMQAaQb7yl5grz3AOrY1Hl2n/PbLE/eJG5ph9AJPjrH
enm0qyCzWFu1bbDhn8WEew0/TI7kJZZoiPTizKqRxkKKiIa+uBqQ8k5gU703FyVBpNO6hnaSeowh
ExwOxycew+3zoTLRPRFtG3Yzza3zDKBVQsJAXwWr766Ygu4dnSUyy4aiSyVD6PdBD1Yn8svTHzKf
qw7sCU2/bUrLtDGPohXGCDhAV9tvPR0d2YiwKJaEj7Oxh9PqnudUJb6A/Eg8wD9TX7MktwO4izBD
8vCCkhsopdjhqfohRnGkcLjL59OxJ+Dvqxpigt5z5yQ3cThNkCqEgPhO0d5TGYlvVNz2IEMAcJgG
u4us4kwUbTUiQWyXAZWHYmrWFwAQVymhPYpIZ8mxFLFqMYe2qfoOFsoNx43sUIQ8j47+YPvbckcu
QbeXBXPr8MPwX/RuUSFCcqahh/3zz3uINGc3a2AA2e9OzZemdRdIDfDtCdio+F75fdlchTzmCmqe
eeWoXPKICW9eGjgbGmvJeVot49l6oXVEhIFbYpbxk+Ci73yJrGd29v6mHC7ftKf2X3Wo8q/IrCnD
fNHqmu5CNm/qHsVKnptsLshdsQLfFUd0osefNRyxhItjFvfkWuDgB8FxDH1iH0R+ccHZLgjdooL5
vuNVahLUr3TV/4IrKT+F/VDC8Ygj4R7Tdma36LXcklO56zYvvdvz4GUJTtADDOLqZtFFzmOADLPU
bdQv+9CCHZgeGxCYiZHM3JYxa3rs+pr35SWjahqHx0ky0G96V50cYGgxdoJqUMeovr9IbTX4R+bv
6K3K+jzZxKwG/j06ZKxPiWTXMii1UGOIg8tRqOeZlSn51W83KMw69oIJ+VfVLZaBOyz570dJ4dzx
TugQgaiWWcT0+dpBNUpEjDuuRpREg9YYmt3ifBcDEJeUPZkFFnZt0SqgZ9Z5ugdJ3Fre79xjdmFx
6C5hFMMpvMT3JVPDCGjMFI/K+NetvekIEe01n2iIzeCA8fzH6AEf6pGP3lrAp4nmcTnKRhgagi7/
QGnkU9dQfXbN80gvhInxVyO0FyHDvKtOBbBM5bHbUZKJS435N/RlNa4W+SbrwgbZ5t5/ingMZzYY
4j9hfMm1fG6mRj6c9hMbdYdj+dN1EMSjK/ZE7pHT/2fs3ikJcCMyfaPVkgwaRSSRkJFOX3EaWEWz
nAevJd8MHEuBT2vbY5+404yKpmbvslmCGsdU/+LhCfTSOTh5zrIuIoYuEJnucx9O7xYYJ9I3Jraa
jHKJk76p3Mv/fCDmR1F8osVyxy/NejruYt7hxMSEA6IWeW62/RW7pWb17KVyDbD5qFstSFCeY7wM
2OSwURW2OOMaCt/QOXzvLy+XXv+xHbdzkJTe4GsVQhULPhlLMucRxG5jBdbcOTn+2pdVjeAJF/rj
ZuEnsFzu8aWpQ4G9MTgQpBmne2XXVSpvGwfsaJjkOlV+i34sOGmqPrJGxlA9jtc+ewxNJiEXjjMT
vlkcXeUvrtGARORnIBkorWBslZe+ohec7mFmOCrwM3WzQk8kZ+LUnVvFZK8qBiqMD9zuJnKfyf3V
9vUtTA4gMiBFbKm6zxWoVILd+ZZF3chJvIC1N8PWJ0cDaVkk8SEQYj2lyzgpk1d9Bke9VZia8lsS
5meo5To8rOIOnqG1ZXT0RNykHqNh091/HBxIbCmh12ikqjYbBB8jtFKeUKed+2IEVdcgNJinGLtE
jQHPaYRHqkOEeUwyoTPi6EURF5PenzTF9qohjkzQoCUGE5pEPiU5/Ge0N9AeFtgupPHMr+v18w3J
Wpb9qWtE/W41azETzZqjM9F36SocJ13P6B+mHpB6VNzDWWeGqnMT9tDjZcrigaxFKA991oPa4xDP
XqzTYDVmm4cL7DB+3Y69LWOE4+8+YOC4GuCVPe2V4GiBT8+N9a7c+n2OM5UAfyKw1hNNWCitDSOK
Bs+MdveI2VvWN8rIkaAmQ/p0ODBWB6olQqvmREu0RWxwVmOzhgPIMQC6eBWZ4EjhQJh7k3zH7u1s
w3t4y/WKDnxUFzaPJbAu+IoOz1Xnpv1oFMan4OKjHVloUbrFI+Sif1DqwB+yQPSBweksr5lBToYR
JoVO/aHnjClZWDazQrmFYWHpxrBb8+2jou/rzX37xJJQCnnIEFjVFX0eAlF9mqeHSpjL5qUt78fZ
cgfdH5udZJHPsNAdx0Tkvk7TKz0TryjSqOPWo0MToYg9dcg4nJvpZCoGL3P4Ub2HsVX+bTH6lj0T
j9db7dOF3MOe9ANzDffp3frFC3K6MaCEB75XwrsgBXy0Hg8KaltxbXdce9kBIZDRKqh/fd9oRozh
kOVSypjhZHNLXDtpAmJL9CSI9xcvF1fNAgAV3upZXs+mQjVNDbWhuyNa4DSy+m2Q7KsIlWoSyn5i
CISJmslknwcj3WtzekfR+ahzwyduX2z3vRvZ8q/URZHwMlRZFXML+9MLa2j6m6oM1BxfIEqy6K9d
DmUEhYCqaA5iWLpvOfVtK0LhLp/cc70E1+up+tKz/SOTXx/8xMYXiWOrIRYs9fCuB6QHrU6K7XfS
RmOb03g+r8irXIoZps1rmH/ShzTK2c3Yxc91tp3ANojwm+8HgGY/8uuz0gtS+KwzyaB7z3ouS3nl
FJo86JC9mX2+NV6MW+CtNFWYc9F5qSrDq5fYJta2kYSA7A9O5xZVfbD1kBzGGeRu9Y2pzxTtPua+
e/gqRg4Z+FKbXAfn4HEiJvcf2rkrMsjkMAoDK5ecObhNpnpeAaav/8cEzCI+fH+n2ZiKqpaNS7a3
yaUf89uhszNpZfVlNPCFJAYaWdmPg6xn8KMqEX+q30zOfal8rYrFOQojZcxqg6RXm0Ljd9oA2Rjg
S+CgvWtpdcmJXDbcSjQg2ivWXGdUk2fx3KfrgJqYHwzIUlLRlYgq89wykjEtOX6tKw/9o4ZnW8+W
5Yon9GZel7F5K3MkffM0SUn2Z+yvrjM2xRVXgDQ/sf00K7an253bLJsIzHev5sOKMHJWNZC4ZiKZ
BrbMmdf5egTfIVP14QwxHRH2IHOSMolmliI3WeQq+ZYIpc6xwTg3ANuJLsb0sIXRtLMYpSkgVeiO
/yoRWYWxzwlNOm0N0wMH5piz5v3DHxPmZaH5ZVYIU04DjbG9USYP83QO9K26rK1YfmbMP7uv4bE1
fR8NvWyqWc3TN04PWxneOvaZARxl5N6wFcEkWD54WhUYNQQWZstux5Mn0xs6xe8illUx/XTlunDd
BT1eGlvVxOmCcouy+qNVyPeEaUZpH0hUSUNTM7R7TXJanNRFl7e44kjJ75KwmGLXuUjqFp3CLLp0
ZW5z7CDkL2NaOODSqGDvXThe0pmziD9bbDN6g140bX/FwPNsnQtPBn0tNBxsNmmS72z0eb5O9IrJ
9eAW+f6oRkQaSyqb7X0GuQ4NC5vHwX0S1F+g3Wjuil5rEoRX1OXIvOJdIlgx8GpFbl1TOET2t9+e
O6Pam2YdUHhfDWbpyz5cCyvlMIWG7f3BQJmZtBv9oAo5e57X78Yud45ApEMcA3m1/La6sey904d3
7pYhqqN+Yd5MfPQRwGrx197epX+fwgcm4qs2PzlHHNgJyDMMal0x+HCQh9/uEjepI5reh5InNSIH
9Lmgj42uxpWJULiDfkf9CAqRe7imaFZ0hprpH1ak/tANVFUAQWdtT1XQqeQDf1VGBRO00AeLRkvG
OVzcQO6VAUM6MsWtwqd7hw/6oR8tqFNsnRLIGXn7lrl6AGrg0aTd5ImF1VnFe+Y+nH5pZ+vNuJ8C
BFY0bdb4btI18Euu1R9Zpw1egTl5ICntnu8swVBD1PxPdBFxIoO8LnJt5M2IOwEiiUKWGpBYwFK4
nPMCsuU+ufbj5rk91A3Ddpa0ZUmU1cWlPX9j9xYyHMaqchakjnugCH1awS+H+n76nOKNKoPqPLY1
AmAxYNN1mNrQvW03NxnNOOEKJAB9DAwInB4pKWXanla51w0zQGxD6vudHNgZYmByXSY7o7WW6icy
2EbH1CKUJkNNEwp148BpqvGVBH2sc3peX0XsIaMiQ6m6BVy3p7qxd8B+Nwwy6vND6sfAKC0cP4sf
XIEk+0dbQ19oy5wZRk1ezthaKj+ooTkdefPL36xuuT7eHj7fqYtDHDJt5dEgk2xZjO42/IZ7Cxb+
/qONrad7A5oTXJTG1IUjZBernuUBwwFPdxu9X3WtQ7lI9k1i2Xruj+ShFKygeJ7Xa59Vn8pHJODA
eKJ6hvbSbi/s3aX3m47M9m0EOlIq0VF5XwPKgzfgfs1LIzzM+W3X5K5othFU6Ihy4xmDr/3kr59M
4z17GvkC94Nm+QhiP2RsXsD0rURlFE5WDXf9DiJib2myOV1al5iEk+q4ZUcFhYLaw9aFu2PPU/eR
wHUUBhuSE7jQlFlnQPOWrZRLoiPIrm3XlfL7iuj0ibXt12cn8D85vyqG54aE/FQv9cvcm93ZUMCr
xHd2fSNnO/IuYoluCKEG29M77mDsMZcUkdBhU67kjJgpceCq02JDfGBGdeyRxDJ61iFSY256kvql
pHPMwuQN2QDwijDpz8MeB+3oifuGR1XTlzaPTS4XcOSt52IWUs5ip4vGfiTtJIiGyqjrH+D+A2bV
rnLAMDpiq0/2RjrNRePcYHQwHMNfneEqull4xFnbnXxpTMBToELgnTWrYzU0HPmyOWYhLVhez1F+
0v8QCsgjhEUyksWXqyHQlRF/1Zukuy9pAHPCkICFZ0B1RTCvdCDjYUgpAXvjoHzin6rnrbVpnQRy
hUKzi1BZFzU9o6CEK561JaSr4keaQ8joJJ7Z4lz5G92CeM+oGJrONky+gz5LnrC0+J68yf6x/bmi
fAgQEnXSScu8xvpVI7y3WsaYOFvCk++YwgsRGXejpXRbdDGL3ORFFWFycQXfo3FCDyAXjuPepDA6
rTLhRiBCN9zVtd4W/uy8xlgISB+06gCZOpCJr2XPrA3zenQQLz2idUlxi24Zqe27YqPnEAMma3Wd
Icz/LXhFQ1mXPZ7/RxJaNC32kNk7k9hRM/ZnrMKC5g0zqyhull+kpA0Nl+O64iubcHudB/cQALe4
3Pj4vfgQkrbkTJr8LU/1uNxkpFHaJdUp+rVswY5/aKluC3EySmaXYCqEpNRTYjDBq9fbnUt683xm
WY8ZbmpGNcf85h1TfG54leHKHYJ8LeldLaCPCWIF6jQLfsOBwkoWBQvjq1IMra8th68YD1kfzDH/
FCYfiw854tNwKmDbjv7Xh37ao+PAILiSTCiACHYiGabQwyEK2DWIXi9tyxgv9BxcOPGb4f0NE3mZ
LcoSpiC0IgnJoVKrbQuhpd5gNI0Rf/uWq9bFw2f/Kbb5ct/6lhATHtaa2SRNySBqM7TlzFGI1gfV
iUwhBKDvrze6SwQaE3Th3NKDhNz8WObmtcpZOllKxQ0chgAMw/c6ASHYshQkksGS1wgw65LnA0SU
4yT8W4rFVrRq5ilbSRh+YSylmkIHdNy8vq1VN9z2yrFvZTQgXrPzaiSWPXTeskVSVUpXYnkKkC9q
KBclgoRnk+FShKQQSMOm5/oNlvpWB8k+utLnGKjDMDNjJu3sq5zQPQ3YqTFTSfXzkEfRTIXyBa9X
y3ZLDIsJZjd0/Xxcx+rRUCY1YJ2+Bany7GcvYpHCftJG9Xe6qyGrcdfD7yNjK8UrshtX0FXWs5pD
jRzU/J98XOmtwV3bq9AAdYdTNnH/XbQ2NcqW3kpm0y6ifwO8kKOQIAo69dJw7G3WWppFjCn7bLLO
j5g/mCopD2nenGq/MS+VjkgxX/hP/Okl8vDcCmJwdxv/z+1h640pKP06pscaRlDL8tUvGB1FlxaO
+OBIbyylB5rXo5/U+q4GIbWb18KWB+jAUw2Da8YGzBADu+mdyYEEsxclA6uqPnTb98beAZy/pHxD
QZOaRwQNLXBW2wrDv5k6LCz5m0CN4mo+LbxONgQdd2RKdu9ZhyD50eTDjJYgbfP91+si3Q2rXnJM
MykLpWcQbsfrsAKoWpVirfd6mNC9MavyJsogwLVN0+ZKfwISIhaZldmvNc2o8Jv+GQVsMEL5SQcs
Ep9A0NbI5jLUK+FuUVfpx79dad/bCd0NurDJ0I+RAsLPDhqS82o9Vlg7oAB99yjnrUCBlRajN202
/bhirugUbuPFyL/mZkI0HNeZvv7xB4GGHMTk4LYoyC+uKAvTQz4m2bMiLrFqPMfrm8/XQmkmWr0d
CU5nTRrrvVaQUfyHEQm5C08jVgitZxddxq8hxq2PRQlbEjx+moV0/aPJ1a2TkMgapiT90Vw2Ygcz
WdlXJksKKsd1eXMA6dllIqLo6EadqgDaTQvl3RJOH/1RTApKd7JVIg4zKIpESTuYSVAbNTsN8MwZ
rJ85hkBowlaMLkboayD4jOKetPIt64XDdcwyFNkpeSZZ6SY8ESxZxpaq1tnsOF+yb87S4n1WNO8D
vAaaOpoNe7foPtKs511BfK03SmEU/LU089267c6y95NXJB7C71CJhg+EOqNznVF3nuMBy3+Xnta/
6EBwbKECgaNninclXHbxKpXqecZRxv9owvTkMIMuDfLmhOXoxWchKE5Qow1zhNsgWoWXXIffHteR
kQ34JT1RkGTE8MkmAVtlFu3I/juwNIrxsjb25Zikkse9VW0UCvLb3ajIiG1uTQ4RLA0hgIbewXU+
tNR+Tw7QPmvjoLgsIO7ChM7U5dCbrX47oL3NJJiA+FUWnsYblmWDZB0+7+GR5tRKj8eUL9C1ZgYj
zH4yNC9crTpMfWaE09Ny4gx1vsCJYdsQv4l1ro4eGF+FGdrxxHNMzd9no7Rhj4rDQMkQ1yLeE46Q
5RH9OwmaYO59IjPKx2ZD5tGsTFodKBAZaFE1unec9VV9GdBJpJ0omkV2tju1BYP4cZ4fxjz0JzZM
Rt6Kp7Wa91lkeKT5VrGP00Tp6p9sjFOMAtCY8oF7bmIGQYlf+Yu1BqLJUiQNRhYyPKR6MjcLh49l
J/RS426fDaqbdtrU0K7dUjCjlOUXc9EobOjehwxDad2YtXfNP+TThPOka2l/2LCs15GW4eqmaIqs
F+/8W9K3dA1F3zE3JCOlowRyxFXj68ejZ5djACXuVcOj+eWDaX0u4LuTV+ce4ueSuq9QoHbACOaA
fJGYthe2l4wVE/tfHzNyi03EwwuMolFnlvWeaJP2FLolHu9roXOzTsKIUWCM2+rt9UpuLMqsYuRg
Vk0oKSIZLFrI2gdwYz/Ds6cHjX0x9Ru0bYva6y3P4jF4ldoqzwmWlZ22rA2xe5e+uGQ6V1LMZthf
/Nq51lTFF28gHyyBUfUvlgnRdZMbuHRzjbTH+WqisSHZU72ELjaebbzNQnxGhRvYxx/X6CTZFYLL
ajq4X74o385RLP5b0PhiskZhKa5BHLNDfKdRniQ1/kzYfctd8AnYAnZfsxdQMu4zrDqMCPu7htFv
YXn+1qXjieqGj3wjATROF+UKhlJuLrX0JTwruoNXjmMXH2Mkth0kDzjMvwGqEsamo8UX3c1sAQK1
wZ3thLnYWAhLUELRtDYvy8Zdvu8Mnzq9TEydppjOOSSdo+mm7yZhdM2LmchlKjQLY064MyEI6i/I
sATLSPEDpS2/xIg6Fd/64ZEgn1gcER1TR98DxogA6NGEEXIz/pnnfc1dY4rmmK0Nr6jwCxXJ1+Ob
aKgKR3pNBT2vVmn9px+T+wnfoZTdHeMJipu7KPeejTLI+tNp3NQihIDWZl+DJzlYOBLXBeebfsBR
ThEiw/CfTWOtr7y+30uXnKjkmiWv9OVKTJHO5I+FvoF7jK0JZlI1+47VnY3+V7PlxiTepTve141n
H37FT3HRuxZ5OwXWusxiV7Ti6OzZrFsoqT8BkXwhMTqeLPLob0J9E73XKheufzbp3Z6FEYcgKe2W
P4D+B5ml5/6u4ywRihP+hLFVWsWUw0MJLdF5co8pDXJLEkTwWgjZGw2/iIDp6kQSf5Igr5ZSBvV1
5tqdxH13OSVhZ0wPQvVsDNbt2IRm+mXafq4SNd2M0MwpMwwwZq4xgrrslrsFE8PhbFUXHoGUbbYf
c8H552X0UAVK9e75CAkC4YatyXyhszu22gsawXe+BEDRQJyUHoFL7TxGk2Yu6HctoM6WmBLCC67w
3z6TzgNVDsR1gkiMJ4bJY4tRkjr1/Lwb7iAEJ+0e3Z2jGqW5ldo3H7aC7lz5HIGXRoliD25JJE0H
OJiWJ47kZYKr21GUdkBwFSzZSGrx4xal/DMayOmzbX92KaJPWhEaRCXsGZ9/Njd5ZOY379idIT91
L/gkVlaWTG6HizpCDG97FKRNql7yFk3e/P28sC1Djskn0Ket2Xi1Pgy+TowlRVzDYkYivCxLOJVp
Oius20k7vTWR1F63/JCGNx+Kym/gHpbYCRhsLkM05yi62xX+VOsT1cIyOiT43goz69kSDUFQcKfp
e/ePbEPwprssqtE2ld89ea6NxVzY1JLlGlpnxDVMm3LSR1d7ZtLzKoIA6v8y7eXt/A35TK/HC6iA
ydPK1o54EogeWqvDwu7it5cfTL1P70Y/GeC3L5s4wCzd9TL534n+ORYhHbxDKfdcPI4WrkpbYFux
yc/UujfQVJdrH1s+VLhbb89FbCMupdAm2RPPT1jR5/zUqOqnOSTaWAIkrjYyw8fVUHI9MNyAJlNd
Lt48i0pXx4gDVbqg7Rn7bJ3IP/6cO0IE+ct+xDeFZNCOAzFFHLegOWgZ1ToLD+aEzE82T4qcWiih
knvg3rBJiqGNNxSNPn4ZFiOeivtPwpkTXRUmnI0ZBwWx7NCueSPhpfXx9ZJJ8JabOnY6+sklQ8JD
VauKta0KiD/1+mdPdmEoDPaN6UGMlw1gHWRvitmgLlBMRS0VAdzZBk2ZvMYDfaaGyzu/vaAInLlq
xWoh5rRcajXLaYYTTmynswxngjNu7YnoeXm2mgjp4lNpA6qoGmqaN7zxxqgsd6wE8KUFaEVmd/do
LNwNMS2gXgocmyyLuCQ/2CiskyNzTCJE2S36T7oZj0koR+mzFdb5EQJzcqu6FoyFGHu1/qiMcxdc
YJNRON1C53fyVSiY4P1715fXYuhJ7OszgBnlFAAo+qAxBEwTP3KB5qqjPsodzp6ueFqj0Lz8Dwqf
+bnv9TxuC8sNXd0RnkLiokT6yUnOCbRz4mp1qDRDpC8gxa5rD1cVPVAxizE5q1cchoBV/g/5oGQG
nCnImja76m2gfD/8SN9qBzMhAIx3fIKeWajn/f35G1qANWnsX1LFs29wbGxiFyaCjrwCvVY3E38n
sz4IgaJi29UUy1tRVUZLcknsU7mAIYgdgFFoomWZYvF2LB9JOGu/7PDa92pyL6vvknvU8pZKgkU/
QWfrOdy6lJP1gZUootwMaYna1LD6vhBpzeEChr/O9pND76GHvPEyBBbMSD0iUKPq1P8He7lUugPD
Qf9hHPQ7l3LeMvmM+lji0dR7IqJKT5NSnDGA6bR++gs2h8tvubGYTNCQxJ+YkhGWFiiXyaARw09X
OB9LScWrMYBlLbgD0L8XhwCUuDa0khfgWd1UT0QZq5Oh0fFhC9t162fvTlKAwdT7mw748hwbzIao
AiIWqSD7cdHvUgn3FXr20+GyNYRHS/LCOb1Nf8oyJhI2xY8yOFKotIroIcAmrYQ2NR9ziLvwXndd
c2/zYVZ+O9dg3wEMDlcVvDgz3Xf1lVpYgsq2ZamsO+lcGHjU9GDwMImb8vRfaD7yUDWDx91ydKR8
0BuqfQiVvx8Weq5WNAxrxqzSv3VeKa0LV1mh7R/RMpzqE5V0+zAjURwIbU2Czq+VoK7H0P94fYhD
+ufMJ02HaHXPTdUf3hO2V6rmqnE79+9kxMwwWh1OqjP8/sFfIoabdAgO3EFMYBvvskfrRsuPOtrW
fPyHkqskxi3+jn8fVS/zpkXtiHS7QFmrdhpa6TBIRP0eu7dvct/BYbu5UeFqcwydKyWTjDljaBz9
MykcxRJkEXmg/B3lxFXO8dL9N1dnf7dJaBsRodbjK7rDJPGrq9FaaD7mtns8KGosh/hzjYNBBKGZ
m+Pd2PAju6ObOGobLfdXeqotsVu60iYLNuwYiYjXct1TRLbkCY0pTrUf3DXo59migqDMcAWrubbk
0BNWdt7E0yftM/Ys65z9T6reaJKwM7CJw6wSMV3hCY2hXe9it5siE0+4vqWG+/ajfznw4oQknUqn
lZBvG0Sgfeb5WpJOUsv020MQQr4lDJITm+SJNaozGeVaXA/3aL38mR3MTDlWKkXggSZobw3W2vFg
akM5vFpGXkzIpW8doLbp7qtbM86ovbIKlqfDlGIkk3EXpj121nBj0kYA2n61LpYioo7cBlkq22eD
zjkvpub9xIeAUsGyyLjFwSe1D1kq46sreSLK73PyPFNLZd6hACB5KHCe/3rT6orTwMa7rT+8sTmL
GzS8dGPMfKuLiwhEL7ngcSkJ3Bo7aRzgZYY5Yun+VRhO0gWumsia/tcV5LNSTOEFDTz+AsXwfyiZ
3Dx17ISTI83Sf4NukoN+vL4EseVsqj8nhFSLYcWgD6lXFGWEzJdbEypu/K/Taw9ObroZ9pZh/LwP
YZ6B9l/bjsSZiRQhkKulZZnO138dlE5g8cyXhSpVjEybKLLxqvMmAPHg66IE0XzOr+JstN8SDNog
fSdVOR2zk1DPa5+3jeW/BM7huHn8XbTp5Qr3uWSx195K4GT5sswlIxzdp+dtZ5zGRkurCtO8HIk9
LHqMF2gJc3cKX2xxRN4ujgAHVHVtSzpkv0lKfN3wmO2Dx0O2y1dP7v+pZuOcdzy8y4R0bNfvx3FC
LCpSkRgkMOSMjbe3MNdqRRYMPhCUaQkeTF13d2gB+ALP6hGltGBdU/5TGU0HIRNmF4/CE2mBfjyT
nsPY3o1oMKuqG9aUfDXnVY6Vu0vRLMRfk0xIMIW6PtEktiJ5YH/vCqD83T0q+ouy7WiDaytnExao
LJqdGv952IDtsdewrRKWh803j9aE6rMnjfVT3gR925L1wOnUDhENKvKHrnoSNuL3v2YzQF7C4jH8
5kh7BVTTlrhnLt5/hhvPu1oBEOLQtmFw0spr3YN3Vs1rAeOiSZKioA1Mcuerk9N+o/2TP3TxATMU
x9WOidxni2RcM9V4oR7Gb+tS5juLstbIbTKxOjC8mhQRaEODh7wEi3g7dbzrDqDLeLlJlZI/v7cq
3oyTZ4ichT9i8rSNeSsjgV4Nfix5zc7ZhhBMlzhNUaWzflxCeb/74dgyzNL8OXo8LcC5oj5Upu3W
2O1ZEA2c1id+qPxlny7srFB7LT1dR6LGjUZthCc9fMWhyeC8XIZUr/M+fe8FIkOHYdf/VzWiYEFF
dogLooj9Z6DKRf1R2ivqxuJgasE+7Kcy/E+7zKv1UGMN8YterAZPYsoCdzUYnLfqdBSu97yfExu4
z/bFRZsSzMdAxfdBLx63sk/fmk2dubPhudsytvq+iGxGnosHwbBCIHSYZEDEf2ZlTDiQb7igZdOL
hDju5nhRHhb9ia+oQCqgvGY2mN9S9e+szaWBrY/dWcOzm5Eneljh58mlHNG63w2PREnQFi0TYJsA
5+6g5URHkiMD3dNqTchwUdPq1Qr8/ejF82V03vgBgzoNaR+UiasTR1TpiISmfTcWpuX4pMBZJ22/
ziHL2PjoZuAbRw/WH3bGW4Kp9XoGyvtDRqAzRsDi3yIDq+jj5i4MZkVoPJlH5Mb2LaztI90fqLgM
MnX3BuJk1vWMTePYy5B6bnLe2qWAzzRwPXG197Zfc4yd1M5mdK3Z8sFJ7KJ9GZwODZfsHk5fygvI
TYuxRtCuG0/AtgBT82A20gc3O4cDiiFqaHhkLCoP3bxtu49O13XjCT2xYRDGN+kVdyjDS5mDDpUR
npSwoE/BnHTPzjSZQcszJRcIwrTA9EjZP30RXxf9t4x4ZKgC70KBtiPiMXzbkTt3bXNASgCGuZpF
NU8JjT6lpPmMiVYAdKk2EdoTxoigSSt/QH4NekDhVy/HAhCpcgyodTQ/kob6pe0covnVYwmEh9W/
oFr9/zVJEe3HRqbk8JWpRzxAdiwh925i4O5V+L86jTQcHNUSy8g1i4kIXtMYEwc9kefNTzYsZdsH
4F+Myf742+KZLnlI1NArpfro8+7ipnSS96V2M1TRMlGSjyB5ajkNNPe9Rdoyl+5lHRfo02//sa7z
FTH/7gLPjfiZIjZfmRPKfXzioXaocClKciwRmDxdxNqDZ2O6QOYfPfW3quqRPK7h0+f+GY763MUk
e2kD/Y0VvFQKleKMIzGZbgjMT2A7WOZ2Sm3ILSSQFtDTIhM4737tCB47cBZiEvIcb2YJ2pcFoIOY
7RBi2Twm+hUGPoRDYNLdjA2TiIlfAD6LliNeAr39lovZFdA2V8xSIRg+hIftLPrhA3jz3v0LK0oA
nGN8fPHnU0S5db5Ycpxt0EovJMq33+hcPJ/T3vi+eEejC5box32WQxxabZ3GeaqzxEs4ucIKuMy5
vTmytdcz8ES6wubAnCakH0dGkMhPw9ZFZB3IKX2C1BkdDH1dS1AQrNlCZl1vUlZmOvb9mIvuyEz7
ItGcgp79uT53zSO0dAcZj4rNROdJ1P9zID9pawqSl5DvP4Wcvp+uQ27/sPcIZb5iOOatT08LiUd9
WvKz3YG7B7YT57TqrstMwR2Q/662Up80BZtcVAhkgnOna7Vki/tROvUSYfffQ5cyAqRo/0UtvCx4
EnJXIH6xY38te4PvI73mMwmGhnGJyYrrdID8dGRkjJf+4a0zExnfomOA9cZJc1xOYUHaeva8/52l
D0O+sC3vHGWpMJOD6466XWDVlw8cc44ppyvZv5YDY155RWzhi9A19C7Q7VQAkhKQr9nAobO9+cQ5
UGiLlJnjqhMplyGTFPpZ5wwgPcYojy90rZJ/r/bYEzt3k0KC99MBo/xJX4Q8YicbfpyhvWt3WF+s
PTcJktkKQrFPs/SDHPi2wlybt+A/nIzQCbW7EjIBHm1eQSgtl2FkacKgw65EdsqEQ4bLKIgRMMhM
lMJZNIUvFlhnFRj3/o5D16K7mauC4WcOb6+lFbZHhIWU4esDav90OS7i/a6mOJGO/d9r7y0IWHPo
wm4ZUIG/jGUt78rPPsR5YyArm5iIKsAJYdL7FD7uVe+4Drw3UbpjpJ75haXBkVP5ldKHZbsfIoFy
PqKuUU26FbtwPDBeVw9fT1xznqNxjyUP9x2exWhrOj+RvCvHGQDqgsP4IF4ztyrC8QGLt3TequZR
x5j6TgTJmMmk0DYU6NdWnd4Hm1i+OGQ/AYc+51IX5EYkJKBUovEPRn8xq1V8rD7D5OOHERKZ6V5a
SjhU2Ni+y/l8/QIM7zYfRS5+lqmWPnI7IV15PtoJYPP+rsIKx+9JPHaS592A9w03muHasS0iluVw
nDRBDb3v03+mRT3rtLeyEP88uSg2Q1+oWL3ZSvbvjkD7C2crJ8LVq/Px0eAtBRHucPaV/+W870dK
903uFzthVJa+60yGQ5oQ99wrs96qvoQGobsEzi35XO3z1jgj/6WN+TTKEkpkOP5FhjD5bnNR+Lvd
1DBQH9+N/5TRqLDaIlk9NSpMD9xTp6Pcjq6VREJwTXPyBhtqCdneU9n1AENjU2U2Wo4d9N/2L99u
4pE2ZZVORgRUykrGlLc8WhXAgY6G1NUyc1Dp5fPW02JcK53XfY4oadVsErEpzbQbCxyj8bJE4r+L
BFNbpwBKy+lGIOuXOM4g98kCJvmTAUjTdKWxNjWw9R5pSde2NiVDGh7iUhKb2iFpDdgwc+7Wt+5m
pGikXMY5T3W22Tv7zvAWQYc/vbKWIWbbZXr5UY7uFHMHRy30EHMvtyxqoW94ICPzT53koF0TWPX6
HKv73bi7X+tUCtRktyLjK3Gij/CS6BRJGxyksTwlJwar/oPJxi5kBTwoGxEIR27GcFMbdAwCQNb6
OILR4KfhaX3QUEoFRrL+fwcATmSr4/PPMtrD4Rbt9uS8ZQ2EZFuG+0rcX6K7H1sMHKhXZV0Tz+BC
FDSzCkPg07gENB417XDJ+fBoQGLOkwe/ftPGAMr7Hodul0+d/G4QmrMB5q+owrsw0c9Wi/fFUVbf
FRnxb6RaxL+BrY2dDmgm2bGQgs0tQp24siHLREwDupP4h2WxPIhqWIfs3oQZW6m02PwybR6OenfK
jb1ad7lvn4ePKNUizD6GkfBQ3MUZolKg/US2qQctCMOlXMe6H/hzKDkdBOZYg1PeryiWYgJxGHdX
OO+UVvNlfPPI62QV7OnMxmEnRP4sMecQUZv9hwzzbWDuMaNiG9M6iWYUdnX3yxcfRAS8aVm6OhCK
7ToHCj4Uq2347d9VqYR7W04FDe3PiQa3dN3MhX6JQ2KV2pioyITH9aUKeWLUmH9d44NiVJzpJVof
sWaqP1hPppHkvWl0OaWfBxR2+gW05MfD4ow1xU1QP8DLsLaRO5K8lSeLzkSYdz5Jp4I7sWH3HtHb
Hm2c9ujhn5GYgYo1UcJD1Rwl3KXbKAiY+Wd14gOuevPLKxz11HgJnv3imECqI1IOJXEp3VUKnMP6
85yZrwAJ4k7thqQriHMgGen5kgfM4j8hRCPAjyBw+XY2dbI4qs2HZQ20rE6eEdcbJKH4m9P2hwVo
zoyZNc4H9P9wkLROe+vse5oLivAuPqGyIGX6yaj/r58zyAXiBHf1lG645TvOvGEdxZnbCAyVletn
50m2miNFEZeXEx67Faa7/0ji+37YMEW1PK6M61H7YZAFzwUylFHqcG1fGL8+mupayX+VMWN6YMIw
8Kyg8h2vuWojHFgPTJwtSYQrWo7A7yIl3yxf0gis3IsZWBlYpOcSccY/ngIuSyZ/U3pkNwIEEaT8
z0My4NiwMWx+EMCUh7ZICL2P1bU2hdQJdxIQIQpPf1szS7Q/6GwTtjGsAAa6ahMrHU848zr3O/IL
lfUzQV5xAZiEdwSDhFsCDLI53CcnKLeqG5mGNcFz/iFC7mH2nOnHKm/s3XfKKjN4jpAvcWBzefFv
yUOEAuSiWtXq7vWwbf1iFBJE1evl7aYsMRsoc0CSfjbtD8hJoiNQshvDQzbEsusT/AMRjkoSmsJI
5TAqAypNel9DKwWQGmjbEHCRFzhUhi6DXvqfn6FXHx53EXceFGGWDQyfdgid7s0E46mcaPmcWRgW
vQq4bh/atfgCBm2hHjCvMMoihBnkCzX+D4dHwLfSPVEAbPxdtlgVkIDPKOLPGLGDv2NBpw+9fMpW
NFy2x3ZBT0Y6n2mj8m3XUOxsxEB0jZMhsKctz/Ajgjxshe5G/WLDEM7Rv7lzWLjzd1WYTWknf2CP
Smwqfc5e7wWwnxCwLfr3sEpQuk7DwsYubFlp+27zrWj0lgx2u0huH0jdU5vev5QlQKg2gAbyp1QF
alIndI4dfWOaIv+ZFM38U3y4CxMLqCL8tE+CjIIwSmsFpOMhd5rBaU6LoLYqVhv9nkTS87fCgmPz
yAR0X8N1b6yemMwLfBhVt+LzINc2Lwlbc52vaKBAqP4i9NkZREkSUEWZK2BN1CGaVWktdZCbPltF
xGoFJ7zEH/thAaCJVDL+1A2QYHHx//PFvkH2L4GlHNwncb8e/Wb3TPdKu+n9nUgXGjJLECdL7oiv
lGh25D2INj2PnD1yHzG0x2vuEwpvfLVEeQBKwAwFapkt4mavHVm9FSZBVdbkD0ncMm8dByQgCFSf
Gius8qBFYRIJvhPzEbu/V5FYfZhnvJaAwFKYcttiGiXEeGh6pBxBomyF481e7NfW4Fton/Q1o6gt
YhnLm068TcO7LsAgw6vsN1a2UIpqfD1T6CDppto1OxOIaNvnPGChPJkLKwYI1uKHgFd/c4fdrxt/
3dzMog37ZTxIYiRtnuVROh1Pp1xN3pRospyo9hhvTvmDNIHkDGANjkjzd5ZZib30to1FdSIoprXN
4gipmAuFq1CK77XhVGRMDRfq1AERD+9Lfbb9rP7OM9JhmPOiVkbVibbjWGDMHsBZjd2bIJqGfdDr
ADOT2uDPf344lqFjSWG9Dp7qydFUBxEDY9JrkbBHEsNlhufp88ohwvNmSfD4VxYFTUakwa9S5M7t
32qgaq+EUTeftVS2g8VEXiNUZg9FKO5tNs3MJQPHaUIqcTThRTG1mXph02U1c/PuEhyIlX6vXFAt
otPeeKtlt/9buglIM2GYvfPW+R67ioTXmiHsxixwLzcIAPGiuy1HYZlxXsT2TXqkzKUbsCuplvOf
8JvIsFvEjxtdYrdiOsaofAft2Ol/u03NIPrmxYOID5YAzKzbncq4zvG6oYQzd16jP1zb+SXDqnia
5BrsvdGSEhrwcuG6G3OZncsTmz+tnFVb3MKG218USAOsUG5yaQIw+v22C1bP+0KnKw1uq3jFyu9g
4OoUb0JmSHUVj9Mc4D048TZoMNp/YZ/L0jF6tAZYJ/jGCDsaH58my8aZYL6SKHfcoX6hAy1btzkr
5VWkLN4zx5FqdSMxAxHNVZ3ExXV9aAE4+pHk1SOTylnxpPw1poKzw5/SxNVsuWcLBqbuZNQAXmXs
vMCf+NKzD2igjOr+u0KGUeLcFw2wWcO7LdULFz9eXdIxl4iE5tJ7lKjJ7stQStv4Ds/sN2Nrkgo8
aR7A7UuYcCLtbBMCAKHZKikKgO64jRcWuQTjmwxrndbm+AW+aKp1W8VN5x79d8k+daY6Vf7C/q3j
PB2liDGVZQhj6osn+mmNi7PocsBe3v/a4JF/bMsR9YG36PSQhYIIv9jq1hMrK3QQ3bRBtiwSQKRl
Lw5brlH4mDBBF/QhJhh5shl/n4NM1Y+ZftFgdK6R4pQHO2tKtADusmXQ6rhmV8BNeOwwr56us9QI
KjZ34u6PzUCV/78TK5fsWAbgTx7H8Astc1RiQJGnICV4OysOtparD84AvVupZjW8eJP5k4AAmSnb
GyKrY8XamfsY1SEvb0fiJLVs9t6bB4BSJHtASRRkVG0BC5kyZsxAjxhNpGhNKQgxvhFOsylE+nnL
NiDjDKHNhu/G73mdtSBw2wByKMmefVZmVWNraxW3t0DnijIC+9KX4gyjqq42bXIJRwPadGZICfNA
FNoib9eA/7AP0GbS1b5D0erh+lFWN4TrN01uV8lSwG+tbBmEj/V2u/KQTbVp20C+xEq/D1aOAvne
hD5PHqdg7pqgPlVI+R6wfAHk1Jl19yFHH9tSkwcUEKTRCxUaDZjLWDM61fLHwRhIvu4SvFR78qEa
pXBchuhwNyKc5f2J2ZCTu7FRtFK6nxepEPrADvqUNyRPpzQGANeM8FGUg8XTQyzeULpb/qotZZ4J
CbvVrELC7dHvoja+WQ6sXp9ovVSBqnlGhV9ZOGGA992KZB5mLCl7iKmliZe6tWtvqVw6YsixJPKt
dlz1vORF6TgDxDacBiwpFJxG+SJ7c0ki/iEjuFYcuJROZPhu+4w+LoU7jnkwn0pygKzpUUXzCBWf
du0j2fAqFDYrl9jLTzbMfV97+Ye+ZVmRvDnKWebidTRW7aeOeEjQcavb/C0FT2JNIHBjERAAWG3r
gwsHdf4MqEnU2PmxPSfjL163X75yEbc87uDYaH5yNz7+fJOdXRDD33pggDjCoX1rWBZgyschWZ3r
EhheXXZeg1lSFXJMsOE+58T7qLnrCgPyYryHx/3bR1fl4SGnVyryhzBL2+FTSDyWwtJDin6tx5QX
scwoOkDJkE2LDo8+Lk01XzDf2kkC9S2A6tqRsucYfF+jlXxfVXs7PUgxAqMVrK3qOLehhJmoF3bg
mN3TMvKggO5HYUtICJz4zk1I0LC100rYqojVmRd0Y5OEo2CK2OFdJHCdo9v5ug2+ttk7ighg9fv9
Upu3egniRDtLSw7W9L1o1mX5XjotDzBVjID+aAwQdJuzukpL66KAy4jVk/tVyrPugVNt8hyCjOFB
RwoKTKNAhzs84kCl5UOciWZhNXKALpA/Yt0O8kVBAxPQmBJApYWaPiXWV4UOjX2MJG+JNJkSE0CS
JMZQtTwwZaFDkJcX5wN+fv9BhCfZL+f3Whd2clhLdyimbukKm0vM0nxDtDNSw43AZ3XNyoDDUFqC
Ax2piT67Y85l1pFRnc7rRHbkp9ND+OM26Z9Ez9CTg3bX+rz68unAljws1cwyosH1q7o0bv2255Cm
N338ctDTuzhYUZdANs6LEi0b/lIWN9uJh1CrK59PTwrFsY6eND0/jYT3nNYJ3HWf61nuY44IG8zK
kJliPq41dP3Rp+/Y0hVHzqnV2XHwMXh5Y41UXLSjlbpCVTsmVmZ1Qewh5xp91e1x0RJ37NVgnhwA
nzAAMz7BEt1hpQOrwX/eVxdrOKUfvGjoTdISQWJGmeiP87BhXH2teEum74PEXrO+h/QWg4qTmHvY
WjIpKPVma5qLWf0xSdZFLKXttNCp4WOBKJK0ZT41WxooaOyOclwil0wlLpys8syZp9ERsgTTHJwZ
IkNmTktC2FlpluAzwB5UiyQoFzKf4O8OJDOYHYZgzegXtoSPGDIxQsYep1RH3rmHNgdYsK60mS7n
oqwakoiS+iotamuZ9m+LhP1xfnZ/ZyxX65Ouk1IPziQssQX+sdOAZC5zG9rp9ZqI384uM0QEFdL3
4pxI3dS5pac4r0QHWEVBC2dBsMKXq3vrTQ3G2wZjlKAqcIP0eI1CLRucJOZ9HOP1llteF+LWxso1
77KS/b2Mvj2K7kLBcX9XDq1Zt9FmAonbywtv2BNmZfVZdcn08MR5/+LrvJS/vyRc5q5ODSkmX/z1
KUpR8okxD0sLQXNcgECyphRujjcPBZB3347KPnfYgTj8O54Zg9va0t8QM5IL3sRXzMIyTC8h50iu
fx6qcm6T1vY7Heb6P3Pdd/rHC981LrYENGFLmYp/FJIB+xkYClMUHIDv02eRcHX2dLnOsg+nJ8WW
One7XIUWK1tmA1cDbrPghHpVa4U5Idk4b+jG2CUtxB6hlaLF04q0FXV7M48Ay+D4nfKe/fL8nrTq
+H07v/3RyHhppAneii59nKzfcQ2cb/IzOja3/XFYWaKnvH3mr7oWgBWgxsslR3Z2qU8A01xvSOCa
Lz5V4H2eyJu+jfRAIq98773xy8q0+p3piqSh6cnsn9ichn+cPHT/nlOQEtODrRfCQIdtRaQi2IfZ
pyMbnZznNWnYm8CCqZo4a5SyHYJqt7WqXSQaE0HGjG0GjznM8MfbQSaz4rFACQajI6OkRZkJ2FYu
prTB5OUiBfAG62ZrYeHB+rlW6x1t2v0VaO1pPUSUvXhW/II87mJwUkQlAIfRukIBDsdet9S1VM/I
9y4+rY7mlqC+1g5Nnp6hhOapYtPJia3UrFIGC4JLMkjVtwx/Uq1CJEiJ8cwNUBRnjsqm+yPug1JS
nkmmirYMqwT0DEIELil+NWiH3XdqZjm3PkgK0S+os7nag5zVBZZIvswRAkmXcu4N/PwTp1LlwOTU
YnQ+Lg7gpOb0Z20fz4wq+OMvey/ZnX9se53Jy0TOaFkn3qpJwthR2BO4BXSjyJk/VKu+AqaX96iU
Fl+u5wlheDEqfS08oDflA37lR+gLxAaFeh1U2wK7QHyCMYUiyO6wWkmmIfXQLPSDewmZYUdwsb/W
0dgWKTPJmFLoqWFhPTLd//1JpFGkI8IqSFy23xeri/UkZ3QVGquyzKINKjyKyPBzV/5ktaEB3LRP
p6h5qzJPJrLPLUpJqK4FvybcmC4hhlgo2y7VFEGtDg459qipCOBFjpfJYIAUMvak4/QgluXegyjY
9Inv87S/07TQPYRRcR+mhmru7+IfXMQCxKwRy6ilDDq6bBZcDYa5tRx+9Xl29tH53tgPju71uGgP
Dg63zk/mPhsRGIVcSGJ/ZL8+H7RMphTCXI5l0oPxhVeXGD2YamClh8dZBc+fnc13JYOwNHSVbeKV
6xhqAxn95w8uZBRQbc87FYgI9Av2HxhFz9Be5lPiuMhcI25IWkTrTjwTP2Zey2gHLezhTyon7d7D
dUOMTp+qIJp6FoaHF1TIwkVO0lwfXT9rh9i0VVojVhdftL1uGaZWpKuoYhdyCr4wYv3pvusq7toK
FxTf7N0tEi1JrlITDkPsjZVU8FBeZpekn2/+2H3QyRMXo5CNLQe9t6knvwh065o9bjVvvqOuyGug
1bevhheTBKJ9j94cyneLmuZYpWLo/r357rr4LO41c/lqv3jqaydLhUmKL/5AjWlOh/ln7uQkuBuV
AgCbV0WzZNNeVkiZPYOw0CIEc3O/dARdW1qmQqnW0y0nctwog/xg/+m8WgsXdxziISsfgqgRauYB
+CH4e80okgTzZF+9gtH3RjY/2omJEpt5BGtxoHtmxsO9WYBgRye+tiHFxwATVBVqlrHfaW0aoVJM
m0g9rCnqY+FoUt/d1sFkyaiN3va+1B8KpAeAaX7UpHZJ/Y/bIg5cxHMfgrz3tmvfanRZhKGlFZB1
oByd2bUXjsMrxSvF+m8Znali0DYapWMNXWBCRkge79seuGtmtrWsdRachS/PevlVSt2Pyjc8r/j8
J1BKbdYJX975PSBCWOWQ9eJc6FdJgkbq69Mu+rTz0Q38OKY2ZP/E/Bat7iB44ryTOXiXxS37/t8x
dObs6wPkykHST20+faO/7+Gkqopqwx5/pPnqP8zOpMy/nZevRRnHPk8u2LdG+F+6B7FalA/Rawy+
nWVFlDVM5Z60WtLDIgXc04I9YZWKN4T4C//PHgX/XM2kyTzOsgaTpmNVIYABUDDJbeUcXO+gDpx8
NCw6OUY6ESkHEEC+H9G6HIOtdNal0p2UcAL1/JZgjtCBIL+00zrSFTvs+gH+jJyfr3rMPBU2TeNW
si1CNZZbf9V8MfATlzJ5RVsC+HgC+Wg6KI8drIBWhxBiWPkd8gXKuLVzhOhpR1cwyqDJbtgYw1bE
B0tZmcMdsZdPlfbSXFYcvCW1RGGCJTv6cgY7im0BcZEPYhvxKe4YzfiYZLpfuBPMNm9VrRvqN+u4
Wc23n9vKiAf/SQAZKm1n8KBI0nY3XujbKDcnQRE+qKlb2RF1oy2sQr1cThU9QoEWFoTmyycg2W62
PhIxWlRR1GaiQ0VU8in9PlGPGNBfIwn75IYLXZitW2ylh9EdLI9ZVGW0q91cey1eY4Fn73TQJKZb
dELQ0CYqcsYO4F954yLPIVwxdqk9lRPzI4qsyP3qwLITT76pv78AT9U0YA4bao3mJXqo3Rm5atv4
6IPseAoDq5ayY6S/WH5VTLUCXyIlGTuYCdzhtnEkIhMmo52oWNYev4I+rBwOJX3JPtkQCUyRUutP
ooDHrjKaRxWo8WbtJ+mrB0iojBQJnZk4llEQgxeJ/Xmin36+mwjXFKkJelH0Dul/SpRAzpWBium0
tgY7rjKETwn6Y+v8EPSdhHvNf6U68hJ3zNKYqlqMEAvbey1FM3n/1F9oMyhZGWB7Rkc7QPhf7rVx
VUWuQS0yyWBnoiXbyFcIOpGjnLW4L2SLFBhPidWGmcncCiafrt+KNp1pHBi/K0YlFt5+fOW6uDhD
RpZutqFIFLwP7FZt3mLEfLE3ANhk6sJkUINheRpuAJ7prniDQZS8m+F8zjog8ht/p1o6BmdKLkFx
VVCp5M1rgD99oeGd+sr6qAoNBUpxXArEDFf9kA9bnP6Zl59a7J+2gKXXIyQrx074Mk9msW0Wf4Rc
0hkO9GqzQ1SxA0F8+e0H+VH2Bq4w3o2J0jd17H3/0jxp7OUWdCG6nXRc1+5xh+zeAAwi+nnzUrI7
EXGomQgicLds3X8IMG6pfLv8BwdLT1aMFmyDwObHfKHN1fPR7H0yNOl5dCF8wzNIMb5xRlM0uJ43
OMDrAHCdkrkppEPoyPb1Y89zWxrLsXK0pFOC2CrMfTjCnRRlMhZ/PuwxJF5hhWOq3hZaFHpSJN17
pFCqwXwLvsFoCV4WJZ3zeeXUl2+XlLXVPLX5vk9JsY/iyKqaUQio+wb1eUAdGGcD18NhR+Y3Z6U/
lwk/iSasxwsnbccgubCMhxBZ0uN3+Rlkr957dFN22SNPsqHlYgOe8QS4ihMihS0IySIv7kNYHgrw
ZXSsKlfC+YNSpk1E8FjIkhb75nyZEb8Xllm2Tc73+B0vieqrEzdM16LwMRDsIj40UUHDgqZI31zD
KiIx3fNB8gKDz/8q3r7DOwSOqukRTZb9rev/qu0IqLUGULMCBOuCMS6QER5vQ4SWU1iSh/6hukdI
6VpyVO77RcdD/14Mzury/dJbNZx1cL0e7zhSsn6ZvixXs+7e+skTtnzsPr3ImP7D2fbz+CdG70yA
D+PeGMoamUm2+RkR/6Sx/ftmHTF33a5Z0tPyWZg4H2yoFu0ySSCbKpAKI/Vm2gzLEMSyJNb4FPu9
ZUB0TKPNv0sVDac8INzUf0SoMrRTfWG3fZzMrndxYE01x9EYm9pHv7nw21KBAeH+4eajSOqIf7k8
tU24ktpvQYoOPfh9Vouq1P5wg/HNMSmNzTUaI1BDO8A/4iGhMzmZ4iGP6vByAAwJFdS0ipC/v2ZX
Cmqx7IV39wbgz9NFA0b8ewYru6C4siJ/x7xg7a0G77ZF5ovF+YAWPAj3E/T4c4ZSrV/SvsGZjn/P
874AYBT3yGonF/ytedVkaCuk5plDGM5FzSv0rD16l+8gkeI0UwugFYQk2K7wxCZr7BlgBQrf8uxI
leiTfBiKLbQv8ApUdlZ6gXob6utf+FGhrN70qkQVATg7FzkBSnRUu3+iahBhztcbql8S9vyRCfff
56ADjCay3xxPWMDyy3GIv5icYPcnXSZjmXdwd3A0WhErDEUPhYPJzxm3fmg1J9IKRjJvGRPVsrNI
eTYpKJzZ5UDW/+DuSC/6Q+KGoeksVXVoJvkUlA+rq2Wch+sIL9GQeJ3/7BS6b/UsrVTQJ3yUv63U
aYwMKFG76qGBDDZaB484wQBGRIChG/NyvcXMsUFnxr4yi3vqq1e6N+PYp9+6zX6v1n48BSi73wYX
7vPWlmpMjp//Z46ujW1JKdBx5h8SLs2XqDG/MS/UolUEbkpHgjVHqDzYJdVOBFQZ3Y68jYxeB16z
HdvD+kc3VH6ajCrxh3E2HdSp/QTmMlNqFstNyPh2NbkhztODDgDI7n5EVaOTB8sp0PXFkTd2ykJf
hrwky1n7MbSUkO//0AZG4HFIS48gqR7WTGdsfSfO9X/9NWnd4f1wECHXzSMEJrC+58MjCt2J/Y64
VzWN3gIcG4Sa/KrzMtRnNwIUOBWiTKorRA5hpBENS/I0PEAamhKmE4FRDcPBDlFU0owoR0hhVVzP
MfxJLBnQ254ybCr7kuQm4Q3PwDWsgSV5vz+IB5WfzujtfOBKcm2yAo93LeCdWxGfrQ+gWuxgBJ9m
lcusL8GG30FD4fvSGgF4783psPrqFghfgq9yLsV/I1HQlKQQLiiSAX+FoGxOSfJ3RJsYSSQOTK97
nHx2hwDQQr+Ntt1rqAbBDqZxn35blEpqrC40nNKrLaTd8b6t7lKHuFBGm/HTpvhH4qeHv64aaTZ2
F2fjQ/+fZWD9XRQmaBmu6KmsS7GpahjHt5FeQZIXiAjYZ8hhPaDJQli11GjCVVMBWouonFbNsdnj
BlmojZWKfsShSColWuc4Mm59J7MvyaoQXtxl+XEWIDmS++mp9EASTZ6KHMPDTMFpQ/l/kMlTNuwC
NwwMiHrVq0PR1VDm2FNAETCvhdEAcF5N1KRrYAG+l1koh5LIHUDv500ap7B3ePSo3eHFqJiezpxe
CUsCVf6Nevuf0eBGI3yVEKsz1l+BA+Rp/1GsUtj6sC/U4Qi1czknHwqFLMUVtKKmZyLvYO4dZ2bx
2B7KvI6lk+8QLPsnFxiZolYTNWiVSAqlIgsrsH3avihG9rI3mmNZkXq75M+f0vxHJwOlETlMj3GJ
KaJnMqMgZ1nLDpKNuKYf5tHFCI8Xr2xo4e8W5IcOQm8CQEKrsK7IwOFwJk+0I/tnbpCIRiqgAfI2
OnDPivGdVLBz2NMip8K7jneHIzxaeNql0xVYPUNlnO5Bkl80bLAs/SNhXmkQ9Oxza0n2zvTvyGYr
WJOCKYDqFYKIe03a+3JLvKXzGfqAvIg3onXd6KNw9gjRRFYYED6cGsyc9zv7/8+whGrRORuZzTl3
5LqWE/kqviLjDP4UDitSaP51o97LZyDOtLPgT2XGOWUSwCaBGUuyuNiOUsNTBTGjmyGt5MO6g+ee
9i1H7Ad/0MD9/aYP/Kwn+mei+rmn19c78f/q0Qq0W4/w/33ruXJdPZHWj7qwYeZwabQS8xk6fQkz
LVmcVX5VLOullQmnhPZd1JeKVZ1ay3LA/B1cKaGKt/6Psz2Ulhf3KYnzOhohkleRcTekyj7gD3LY
LkZYTPOsAYUMA4uT/ZFYnsyyz5d/m7n/6Ifty/ylam3+1Jf8lyNeT8eBUGWWHMRGaYL7JFloeovR
mbjRq9X5WIu/lKUBE+OiiCwKxCEfvrnSS38NqR/Jhwd8W9Xj91sNSysYa6ejal+x8WrXVy5K+RdX
gaw4YmQTIl4+e9k1kxLLNLkVtVWtzNv6avpfThCOkY97eabycGqcrAN3oTCnlyV121XINNk5kROS
+RVMhYgi9XHgzuuIV44A3cISnzqhcjVx1NVHvAbYe9F42Rcmv28wRpddGpqx2Wq1P8AHtf/L0Csv
nqpvGYEWWhMykT1najBjOEiECg+y+6VEQ0DwibN88T1lYcvAt6PVm6PfU1nfTfVmnGko/1L0+8dG
ijB6Ekt6/oPAfLj/YgRic2qHqCJAdJ5V4kLGwXjiKkalZ9szrD7NLVgN7WYf07+fkXpH+z0B1VVM
PwXGTJKUPeIf4f6YrLi8nwrC66iY+Vk7aw9uwnbswVD+8hZSIFq36QKKnTHS2svuz9DyiN1wyM36
CA2+JhFg7F0NeMUcxUyHb6FIETh/AltYSM18KJ7V6Uc3yY/5yKoxec2YqLb3x9LNLpUJnSY7Ar0S
7PT91JIA5IUSdB/93JxKu6pn2IQbD8gy/2snErNbMokfq7NCHYBS0V/nwxKw4+izA6XnV2xUcQRQ
aEJO77F7haGy2cyJmRhc1/+Ye4sRqF5dSbnDMryu+BViaOhpt4/XKoGEsPHt3V0gWqVZiG4peFZ0
cLTHsoHTVYX42MrU8xlZOtW4iWmXUxkYPp9iXh77Hekz7TNGcRnplE+L/qeQQKCN50VUS6nqGnk0
V8xCblFvzwXiLO62wIXXA/myO4ugSBvINZdtqEK+phhuZC9DXfmgfbXbs8ZUtCvYl47AwCXHyrK5
kmwxAnnAbzFraTiRtucO3/Xosl3yui7GtL7H+RO5pCJPHQqwtWvN+x0hQF1Of17WpsA8h+zOV82A
5rOcR2i5Ao/gGSX+Jj2vOVqDj09PsJNvhoAmqT+G8P4uXD9VeRbiKBwEelYZJOumtOi1v865mjTv
n2eiX22fAK6OCxAX/ei5YMqlbFIMNATsY3ZzpQtsJkVoFRNW5auehyytKORggebuQ/b2GLycoa0a
zLuGe/+SVi/gf4jhEIw5KtUgK89PTQ+wJ5PSEEToaSRC45WoK2+s5Z9svr/Js6NDHLnEBshEE66V
av+BRhbtCwQabMc7v0PwA9VwII6KGlNJ7Js9B9P1hNlSQuhKn8SgHjSAOpeIWxmU5TW9QpV3//FU
rqMEnhiDChj302jTJyBfk/GRiMVYturWLLc9sdux3ds67hywGTovsKjDW//wxecJviFs0C9KtAdy
GF2WlHZHxHdFwIQHUNg+sXd5HzxQcuJX/6UPPC00lAXCAQMrb+UL5XZhWrwvxVwPnALQItQBoO3w
IegX72T26TTyBJMzeEwIZ1Yn/QY+72XTBKRY+cTBcOvdO6unBbUWemwPBzad5NLGBngkKQcZS5xX
f+JPn3vxV4PDkc1lRG1kqdxrKevOyrGx1iAHHtwGrxKlKcGzj36bF329U1ZL/vGbJoda1lPlCpY4
1KTJ5h7lWulQRENg+oNaLa/8cfltMUoN2QmL9nAXKA4c9mNUgAfNex5RGqPqsdFJqyaR2bYY7nOD
Cs1Rg/ai0VTnVHrCFhbloguI1UkBaxiQSHcgNvsWs/6W2WCtmUfDjmQC6vr4Fu00KIG8CyXHDD4E
2HqdEpeAcJyO/Up30ldqcKI8876zKah8QuDqg9H6zXXIw5FIwVzSC1xvZnpdW1Z4BByNruVR+fAX
YoI/geWMQrQMAAfDN79WPxi9w6j8p/Qpedpq2Kj6jKslBGXjYE4OQzUWXozF2BTHwZavFQYeQh/2
anHYgjkvKnFS0/IqR4Jf9H9GpZkdcAOwczuB1m70PZvUkbZiv3AN4iAtGB5uSU/RPPU4jIlbVKuh
YAZXVKOSiAm+wW3nr8z9+g+EfvLHXH9MhsUQTqMFR5YiOUfphkzfTWW8gD3YCz6BRd/EEbyeX2Yd
71uPpQlbgT6a4avx1T+lM8ObTqPvzGoXiIuwsd5DJY4fabd2wMeiL2teN58HkvHjfdXRyscaqcmd
xVwnA31okW13AJ6u3+iRrdz4KpvKrTRS2nHUNGjZktF1vqIWlQdyloC+G1wRjYJMdb1HQzAPe4Wd
C+5fXXKYPeJTHl4RtfcLWe74l9crn/qjxzE0TbjFdScHVDaZSqqZYod4hoU2OXHmEXwN7y52VnX0
Etrd66AkhhY7Drnhtxd4rAsHl7KnbbZruUFRuQhoVoPdBnM+n2Ba/NiL4WmbS1jgfCb/tEd5lZS2
jlW095Orl3/hHeYv+x4Bxiy6yO/f4UmWGs7hQD7siyAIs2N9yl+PohGCesnHkrZZ7BaCcG1oI3r8
6AG4SNAolgA1m/XLmuaIRiWbcR/b7jz+NyOy/UMBRpOst9axJUfXxBs60+MXyNGZ4x/DqvPJSxw7
/cX9eBV1ngZfU9PmWycD0P8SIhdVnEJhfdOV1iO1DVkDrqHIg05zO+rwszuQCxYzPJz5NfSj3Edv
aIroEd5dXbKg96mbkcr/+Y2tzh86OwLONeXN2YEluTnJoeg79sfVGhir4dYq4L2WX8oj08msbUmE
xSjOzhjOk2VuPBlW+4zJe9YiqFCKvW1b9MJHrrE8n3ixW1RP1prs1qS0lpRZzZZdTppbmmeEwdBS
6oTBC6/W4csLBpo60ACjxbtDDAkSCOXmzPOqX3LreTAphjqL6N11UbWUmBPmsBAZ/uYjvkrfhQEu
dovyLx1VuVPwM4SuoptAfdFH7yFAeuk6OjVQ5263frXpmD6PCv7PVOHreTbq8rffx5IjsxIhDqRj
PSWFI8z1mTyFCLDneZulo5M0pcFqLe2ogwNSi38pQx2urX7C3JGFGdAAGPAz3aVLtWJM6ONPqq9+
UcimgXlGNAVuB/R7hKcSmQDr7rusaHzK7d4xfyg/tqJCAoRXnpOjO/ATMVW/H7YqKpsC5h5oEyto
In0r6Ufdq3Ue8LwjVTL2WpjWf90fSE0s/WflcvYPhYJnZauan+uahVCvtkAnRMgrWnzz7nPoOVIZ
Dn7LlKilnXquSWtwNxzNtHak0hivygDjAK4zyokAEqQdNHBNz9KBhQJX3znE270VZyDuEhf/wl36
VMlS0iZDtvA6w6u8DraJ5GXNQicN/xHxP/SZ6kfk7VF5vWM88sEH8HJBnEMaF0HIDN5egD12l98y
Ry+V8HFe/+wBwvih1BQhTy1eKcEV+2RwQuUserotd0PVynsKj3RUGAMo7zOQfLb0LvKvvbj+ohiu
nsmpuIN97IkCEDkMNGJj+Nzw2/XVF8h6bzktbaCLHm4SSXHJt/7PwkY4ZAN7q4hLv3VE46twAnZL
YUxpvCpFPYNcWRiWLAfyVHVKqZHxLSlksLj3KgfSulNGmrp/IXk3pYAke/KV+d3MiHxtHqibstle
w7fLg4ZeGxtrrX09+KAcGyjjgGLhd6blhQYDUQRy9LEGKL2eiJyg+dQvjwbjWdHPr/TXvu4oGwTb
gma+0rTPTzdR/J+xJlofTLswrGMEEnawrnaY5SMq4YvS4np38uAztEOl6VZyL11zizSK3YtluzmW
hXmeKqWQjqkysVxPMovROPVjkCzK1Fmwn6tBz7rmMw36Lgn+ApSAf6ttP60J5U6wFEoQ/QXGhDbq
L4Pve83kOcirkWd/ZvvF+y8TJkZgn7O81BVL1xJwW/TwebJH54GTUri40tBl64fQjfKnX37Rvsd5
6RqZjFm0RT2OiWTttUtxVqcedALPKohE+aHNN8tsh8im9GGAw9wpCHB1BjYqSecvTRls1fP/7xly
Fky6VbYU28/cDA49YgJ6NG39hwFmI71gURXdCyQIRBZ6oIEwAjxVFIguOYiCNMBEMgZckKNVsDDc
+6rFxUrRUsVF81DMo0sx2NpGk0z5P9e502altD2rhkOB/6XycrnDn3IxB7rwGSQ6V9bHK2oVKv/5
HVQUE2O6Z7UrJU00RMEk5Ya/4xdedKypUCvMEVq1o+ahkwXLKcOuTqJtln5hKKXp16yWZ6jar6/k
T/aLBIdxzAsQKr6zA+GooFXeAHTLf4RrxDdI47QEiur38UUpCJyZfelOcSJeBFgY403Gl8IRpu76
flpsEn91/uefN/QQ5DoXMwAUxIP6xSK9r8+vosNPJ60q13Ckauk2iyk6jjnUftju6KLqKEwaHUTH
gH9z/+Yie2lACYESYHmN2DK3fg2PWzVvBXYrd2t5q7VRPA1ycYMp1pJPfwUmXzZdETBe845rhkWW
wLTJK+RLrc7jPZAhEANxChYAAoW/95B2Y0vrajob8Ddk+Y0L4wX7qkcfKWQUZu3gR0x1BxROWUlB
Fa4AKLzutAU/c3dm5MZWM7nt5hbIXrEMxRQb7gGAixJtvpI2WYSo3Yn18rKAUwhVBV2D5heft66H
3znJANbZEwhhTPOoZ6eP9Xe7XeO3yvvgBnTAmIrDXSRSX1pxIkIMcXBilPC2epxKt2udkyxUxo4q
uKmmgJ7t80PIZ4xXgA4kY7/h4IpPJMf+Ld5+n6KFUKMwl/UhYLswVBkAL1kYjKZ0QdErc/n09DHo
p9mUJCDjr2mkPS1mMJ+HagM2XEh8X13Kohol5AgBMGpAjP/axFryCONTOek+ZQk4LhQYsGjmXGfl
roEnEeEHw8uoqif9xGQ34J+ZmNqyUp7NUsua5SS+18oP65kINi22ydzdbS86Jq4wl/7HkbuM4gWm
HCw4SzagA9X1KXsnLWL3myKqJvqmX15UEkZSjyf+sjWeR8O6gjbWfVUnmc7aByp/Q5+O89n/+wSk
trEDnpOdg8rb87ncUSFUAQuzfNHa78MlfeWHODkx7j+sDSRCRbR+x4tSHil5CvIgCPJ5aR61EpcJ
tcdD7MuSxrQCRelQm/TW91EJmij/K3tv7kHvrb0OtRVQ4OxduknSd5R/tZfjOyU/WmOvoUQE+XD4
LPK6mPWM3F+uI0bKu9aV0E0ILlJQz1E07SFKuLqQkD2t1XuAuRkNEoCE0jCKkvcrU6uk4Luba3mm
ojB4x2nbFKIt43cYAd6xNx6MwdLOGD7ATyJDtNFizit0O2+FL+cwPgElWYh9xDaSyV7nIQl85nex
aGRWnIy+Da4H6b6/CqbnpVMDvGwp9emmt5B4VdoWyJAnwG/PfdfYde3R/xkF09vg4qpewsrVXiO9
wwMZgwxEHcQcT3Yej+8C3H1AH/bJMY5j0aUkb1MUzxyST5TlBoXxf5Ynr2C/jSTKlJ7CX7keajps
Xq1Q2jmwWkZJXXje1l/ho0gTM/ZFa+iSI/g6FAT/pzQnrXODD9N5YRTGCnigYANEWXXvQKZ1mOXB
Y2hoVU+HhA1zaayYc0WYB48bf9GlwkNWJ+D5i+7o9UZgsizVQnh3KRS9N0qKKTr7YOD8T6SkA3qT
FLvzi6YjqWGtWLUbi5ka6mjXrc4isbycYIwKUB4k6Byy50g0Xlru4TATXZ3devVECM/d6BZfIwNN
Hy/J+auioMwVezCkfi8t/XZSCv29i1nqor4LLTU+llpYrRKjSsUglP3OSQPDihOYnskOBrrpOva3
8QFgA06DCCiUrkaPWJhO4uoRW6h/S78SOxslexd+6sgKgs+WMaWjQZtIlg+ZLTOFdWwGp+gKEMvs
LsdclcSoO4hIrtgs5OQKKscnzZ4tsNcznOGzOYs3mBUSpobtMUEXwLw7vgmjQEX0opzEy5OvKL45
ZVJ9VPv4vTmBXNtPDVSzQOhrCgpBRgmfOxBNXRNPFm/9JkTeizCW14WzFxI+5lhvJ2z9AkSSnMVP
KWkZ3N5QcGnrLopxr+A7iJVqqXl3py2hf8Lvugy0Ba7s5KQAVl4+dFb7iGN1a390pTdfo+5+cEr8
Bt1w6XuijhYOa25LjbPrJ50Z1hUflD78jMYxuTlhPbiXooy1lE6w2N8V+V4BxdVPVsCrBuyKkmrF
cHElpSA+ohgxSvTFiOo7oBjfqm5Gu1zU2dfkaitiMeJ31jryO5Rz2oFWQvCwdqFd2LKH3zcdDy9E
JIBqWvMzH724z+GVQxP15E/hGNudK0HD0GUK/lRT+b4ClhIyOoaptc5rb+uv3ff6OdVp58jpIagw
8W2ON09OBHnujxfycYjE5RKgZl77JSgbQMx+bii5/k1Qxdb8EzaOR5biewzlTwUlf255LEDfqLaR
I+lurU27UOihHzxSjYys+se6qocd2MWv/lBh2WR3TtpcEtvnYJzu0pG9UcofKv6w7mIFmpLb3UfT
+fwNhfuBq+kjrWNKacl6b6/MVRiiLnvh1vJuoVfqJsEE0LSRWt1OnZZSH6oX0dmX3St86upgwWtP
ZioQMElgfrjep+bdFY+nX378yOOk9npGYtP6a0Wi5/sqjWNDdauCFt9EEbmYQgwnsHY1uaR+jz4d
92QWtKfjuP4XCa1G4C8O8BVnpUKcPCGMMZ9pCsMI+eu331O5G2Lem90rMZuuNn/VsYzMBSTYSMPQ
KvpRi3HlCI24Pz6MacW+pPHWNZh+z6xAcE5w4VY0qnrPo2mCW5ruwL0M8vi3oQ50CjA3nbSV9GTi
mlPj1D/Kcf7vd3rNz5vvIyT2rzFqKXyHE5HJ0ZN1RxuxwAt5x256Bw8rnveHw80I8mhhG6tJkv90
SmmZKDE9KGmfKMMM5rKgOFgvmCBObpzP6zenFqqPi5ga1FN+D/I3HVruP0cB+wBgJhZD1B9lbHx+
vPbyAhxmxLAYBUWtqWwIXMxY5lJhLP7oFBeTEb4ixgy2qgefJDBTlZo5m/N4L6yuPoXUSIN7YE0X
w4ZdUr27MhTZkjYop2WpI978w7nuMOLVbO8YPP5iCzujTPHABbI/IAwpJv2i2wEqZJow12H5GGxQ
tDyAHG5yOto6D7uixc8q8ZsL8QDd+qYtO+/CNxMN6CkZmaQRb4FY6aj++MTCIrALkruwWZm1NRqC
Z2oYDqsmBpHegfytYNpOAnzGt8JoqNJ8MLDJUKAlAj9+yr75nfiVk2m9KoQWYr9AqbJxK4Mpiw1j
Z36q6dMOjigb0VR2CiSq3DL1BnU9XufUujNFzmI4m1wH9t+tUiu9a/gsgyv7qrllr3lLFHFl/dIN
9fKGwsIEEJuZ+Xoy5HcEVihvEUAs9x5S+525VW+NZU0p8D7WM494kVvxgdggfC7Bzb+UIwL3ax9C
VmO6BmzD+tKV1taasLGVtP7eqtRzkBDspeNHpt0zHF8wJvY+y6p5Ojwm5leUp0kEIfypEreAGeUx
m5TduJN9OAPXv/WntdexizifWDcfs8xUlllTAMOyTA4pkoIIgt3P2cX+9Y4oNL3EZATyPXeqBhiE
cYMFS/nVZekRDPktu7Okdp5uZNrzdPnhemxSMZY2Y6G4P3iNSbZxicFu3EYtxqPJb2U2xlzBpJ4H
8IAvizfW1wdjnnmsl0+vmO0s2+cnuHqe9K1JsS+1Np/C/3VRJzUGDfkeZde3fevhwHOnMYm1QPlZ
M9iGingsmsjLsLDO6SH65prvLQ5TCaP1zu5eru1fzfsV2zY6Dv5vZmQhDuWs41+vDPsMV3Bvmnpe
z71ujshYhclMBG0jsWM4AdlhQsCf4hbQz0AzpBhl1DU9Y8kJAvJ+UxnO2Is4Bv7ThKK/B235QuWW
Sh8cgmPmbwADsBqBn+kVWzT0zlUttIsA0cmhcb69MCBQvio2akV9IioO3wN8E4+LquGz91ts0+tl
7M7Hl+6uYjNkGxEOqkECeXemZ5uRJY1t8P38oN2kSJEVD6F6awdEpOZkNGqUHjk/XhnyaBMn9GCW
Bfr19unQWvJi7RJmM4pfYBplT94iTbE1ZCOQQ3cR+zgu1lpMnGAYkLp3rbJRQ6rZB6ysZjoO7cxI
Q2q9Uzw68P0LXhfZBpwi6oz+VqM1Gm2933czuxe0u5feNR93KNEiQdX2O6fbSXzFbzGJsenvQL42
lPLxKBR+IsRuksW8TPXp+qUpcWO7aGKRWSMexvB4Z97OIyZf1hrzrfvGSze2wKUiM3dz0WtU1uDW
JH3NLZrHcrD/l7sCyFLXbAgOVbRJiuA7rnZThDdTY58nOKqoG7kr+meE6psm2oT/r4p/nVvV4ybX
T52C+I+VtThcjq4CsMP7Bl12qFKwa5JlQlJB2BEisogy8MH3I4vh07AfKzjxFwdgGdya3XlAgd7X
GLG49wgMsgojf4sClkGiXojqBbllRrlCe1S3PGH65AHkh31NVXt8tTcuodJDSLAFRv7w1BV6CbH0
zlFpTzrGADABx+Ot4gO3ypdxAcyRyACoYE0PmFF118fqmpaEYx104Zte+EctVcS0AygpozqUXpXq
3zQMi01CA7zo5b3GO/xjbHt7iwTnwn1tApXjyyUYrLPxyfPk6jdHvSXzCopHIJ0El0GIqvl+vnrT
Ns+fijI2mNfnTxpGTRD816gQqh1hpxbTtCQDtnzIvDnNV37v41ofTbSft3zPHlnE1kDQWELpDP6G
XDi1LrPRt7rn+eboF4Fdh85sRVjGBEJSXtzi66F6UNvgrwxMZEu38W8iWzyj9AsJjSQupxCqpTb6
tuXVRaBCODKqRK5ZFRknZcvEHQTICMT/xQ3VE2ROnRKs6xdfPBfsERV2KfujvcqJ9ciM7FMvMx0E
W8nXIiU/i16XYwQXgxQTnMXM90qGwew9UZ8hNVYbni532RMCKIrzYp9acxuMgrXnP+9yCO5iSG+2
+l/A60zZ+6Y6BCz8gnezWst5FCn9Sa7V5KfCuk2vhNmmN0BPHfUVBVwrAeHQ134wvoB0hrGJZmsN
NZIq3fH2CpA4V5gLkB90yrgUVRXln9AH8+JVcVAZP3CVV51RDyRnSwmhdZR/fOZNUSc+E+fpc+6d
yfggu+CBAyWtDnMA/lI+gitd30WAfSN7aUf5tt7YnVFlYO+z2zzptF5KEbSUDmVXiby/MIGce1vc
L2DNCjeorDyizmrbGY+kHQGkLyaJam6WKS1KOruqUSS3sS6cMQKJCndvAk7C05mb7GUVgv5dmheD
AX1Lv7q6D60JEbJwiSlx8K7jyy3VlMAeMshfvhsTRBpIyIlbXj3cZwBYYuVqmzmvFDcyviuQRxZv
0rXTGEO47zPovb0glLVR0b3Jhf6h3s9S5g/0Umg1SZCN6eM8pV7Ey6TmIG8MfYr+ZsVZaIxvCrmX
Z0Q/BrCU1Cw7WTZ8i7lUkaowYF4RhqyDYTqwTMcn45Mh1avSwuSK6NEtSzWjclgTAtV1+yxmONu9
lV9jkZYh7/e6uqjHMTkH+EvXcMs1IucevnLl5SFC/qvnS1Er6yYQs1tquJ3mpSgkHo+7IH2A3nbo
O2ANsXmI56/JoDZ3+hgITsoDQ7RwxGKbs5iu4Fbix9QwmjoeHc8uMGKjpQCbkRzUuaS49D+724yx
HZMYlB9ZKxG05zIJBYlvkgSkpp/8yovoV9hmIDNCaCnhYjh3YCGvVql9djaKcMIXF7nQc/i4SK26
df4QZgETl08e1xtitMPE/W4Dv3TMPCgshFIQ4WXAZWrRdqnhevG/AFL4TupHYp2O+aw7sAkbqmaC
o/Yh2HpC0zDMQNs8g/jdo3M45RNR1RMuddYgdMRjrFSb9HBShUa63koo+m+ErmTYBbgd6bVnXBDp
+HkYANP6VcNcD2WGAqKAtlICALy6xsJauoyAFB9Jj8dAtm9Mc5P43fiwhWexpyustkd8Lmce86Fv
+8YG/RoyBEsaOHzh5fQIjjnzzByomKA6U9yMAju62Y+yDT+B/FL6B88kRbwEsbzf3TSS/1VNjnL/
wGrRTgG8MGhRBfZPYngApMj3Vq/NkfE9ZfKTLwAWXgacbevgvcpaDHMlm/VlpwITk/Y0xYvT4avP
sXEg4o4v/hZMjmb4hzw/qbtxTGAWakPM3gF9KNXbrZLPWo595cnyf/gtOyxlyXlSadaKkFaC6sFi
Gb0qcF1w21l77QKNu94RliCkIQvi0yB3gE30oAnp3LupoNs5vj1sLXRA/s71rEQckFWu5a4fmEDF
p1eTyS6MQEsta/tPiiO0oqMCW5FQGjtqs9loAzHInIxcObqFwZlvaFanTnq/2v3cMm1h0yGRfq9y
Hd2DsjAxT2yOHIcfCsHOayqZ85os6oDQOQpvob59wKpLjovxiR9vr13dOIDcGK1lGNkOAXEAt+BC
OpF5QmE6QtZULnJokkOvahmUGKYt8so91yOCjoyawvFbJd00MTh4cgAuXbn9771+pEYeXVKx5oG4
7y5pxm6VA4gjDJL8ZQ6tCTa4V5fds/uSlrZkDEnW5QMIxcS7npSg06DQurQu0J2nBMpwbugIfNIX
8zbA9TFEBd87gsxZJsZ6/YkIiwqzOtvT2CP7kwdTaJ92mBxkNSYw9/9RhxkXrlTco6hc9rBA2iH5
FhB51kkfhqkB6oNqS0i2ZR09Jp7c3p2RAW6btpjLIKisAzEVnQZOi71+Q5pYvVFtvWLMZwHHIKhH
Gpq6g3r95yym+1ftM8LRPtBB0TzQJMlnXmMq97Ab4PoMzN1wNMJ7vfDqW3U3xtLA1/n49LfbYO1i
u7XMB+/f5uBCS+n9JhKdE1nr1fknXTY7gSdnZ7YcT1q6UQx1l6xmy+frOJGE01KV6TEjPZBHvIKK
rPaBiafZIFpUkLs55Jjx8qejAo70oqwvLdBJlDlUJXIlMXu/xa6TTWrJrYKbctBQ7+hzX178FG0A
HwWgAPJVyQQK9k29Kd5gy6aNSlKQqWxF9whaY72UHNHF2zjZnV+Mkws+OBH7qRZaHuCPRddpJd1t
U7fpUfKuPAWh4V8lEkN5sPytMz9V1vf4glbiUn+4UK8qlE6yVULbOLAd9qy2Uu/q8eff2boIp84G
BHcMfH0dSDzUJUV1cSn1haJOvjbOyBy9DpS+i6ToLp6KUMDvMo5E5yQ9Qsx6vOtVP36pNuuzr3KD
TEfjVr98mDhAch5cDfE5fovWTZ2VUCz0KhQE8G9Lg1l5CpfAb/11xam9Ny5rWk20/rSVFTuJ+ATf
7ZJi16UjWTaXyHY5yA/vwKM+Vjc0SeQWoQljqz/fyOq9vfm4TP7E8o+ItzOtVtTmIUkhOhZxonmY
g1pE4/0QjF6YuNjjnuNGT1GrE00fgmdLRNdmWZxMbTIxdgJAbNY/d84jfQx0D0ASLc2BwbAG3C/a
TsFcC6Ah+bkeHB9e6V96xLTvJNu30VlQoB2R57nd26FVdcZXxFk7FNq72HHgZpzgdtjT7t4jMBod
hP3xRdI+oOO4gXAf7U8bJ0hDeflJgCIAIlMjfbaBquTDo1j0ElkWtbhHJlwJ5gZRMNVxCSIB669m
wwIV97WZCo0Wb8KRCNchZtA8yz5mjq94sh942YxFrR1sK4sU7WzUas/3tlTnjPTdNuHWo4gG5vi0
Dy6WGmYkflpSdMyfnWbH8l8QqFoWmJYpbcibCrT4QA5Ap9Veqm9gxsJ6plJVGQNKNdwTQWNP0P9Q
+rkiFXwp2+2S2ulsQNDpiVClhZcM9NyFKHRRRd8wr4AqkLiJBsxjRtsByU8ByzUFbCkNqTWsswPq
LN7DOzVZuCtkYyqMPDRzFesfy3ZnZYCl2T9xuEaBZxH3h0XqBbykWm9yZY9z1BK2RtohziuiD8ht
r/dEwAPWTuCxCxQbU2WTtAG+B3NSYslqs+SGN7s3CMT5lBSyKUun/y4kvSi3f0zh8G93obYjyRcu
Q9elw51kbt0jCxQmLTyYnoQLW4wacC8EFSSPpiSG44lQWP7FdjnbrFlqCZ2YUsn10cjxBABUJbnj
70bCBKEQ8klQOyEZ+OwUefrnGjQFTmYdcRbrP1zlGNQULXi+l33V1pHQyKSHbfUO1UM/27Uq28+O
th5bF9be3mwZV+z3/HKVvNMwGUFgPlcTi7QOWLHQKs562PneY4fLVK/+lAHGJIHbtBe4yuYG/2GD
m0nGm88BYvae27W+yDUjTWKC01u0j044QH0ZfFyjA425qHOPoS5tWruB5pSOZTGKRvEWvATIRtVC
yEf3EHFinrqNh11LuA8WjbZxoEQTQmEQ7PYn8AjJmfOimxGazO0Q1jimBEAT/OxtsmJKBt6pbHIU
yVyL1Fvik9uwBQa5jAd7xtx/h4R92XPk5Y6KKdjgI9CoxEkEvthGz8nbYjNpr4ihH0Seln6TBxWO
IXiK4wa4cF+1W6o8q5QE8eUzgPlkpAtQf4TUHJdQdMs0CxW2JTNVZAd+1bCePYv+eX4rKEfKuI1C
Rbf2o2ZXKlIzU6aMW62XqI1dGUK0sLFQoOv/MU9m7QsEU7phc5m0WfFf+SOTTyVi7kpW/Z0iS7r1
ZdCZMND2GrywwmAyH5vZiThl71HhM2h7OjQ94wSJ9tlhKyntFMG0uUtbXpxaOul05dvs+NF1JHEl
GsvQdJmFQUjaMwkH+kbQXg/pvB+C5EUkCaNz8uw+xqjG+8seX2LlMFwRiTETBXRHXt6Kqml5qEVR
yPA+B1LIL0iF4pBJPcH7YhyIiySQXMfabVUdtG7kyefa8nKBUFfa1t6AIg1rgQp/FFFlYTkEJLPB
a2pQamMXRl5TphmbonIpwb3oszUZP3E5EmY78zfoP8HuO3pzOSTsdFlW4RXWXHB3LzFPWYCys0Af
CYmz/gaBUjX77J4dd9CLREfcmA5SEdD8dJrc9LOBbrN4jcLlHslPP3aSvnjsI7nninQXC21d4YYw
Meb0KLcckYu9RxHF+3rYzut00aCw6uxeH3xYXn8L0z4c779TpwXnnSKgEvHQqN7pmZxowaWcWd9M
B3KvahCsFbA9rBzIILXrMcMAHX+QwD0sca/6TRrzdtgNR1IQkBCCXmu9OFxOgciI4yTZ7osUVirJ
gLz6yGFGHz0v5lMr3T5s6ve0uCEn9fRz87MfqC8MEPy/awfMcxQuOC/wpTHG1uQXDqlnZQwwTc2/
4ICbFkH0+Wz2QKZraOkBMgfs7v8oh1BWRw2oEIXGlHOejekIShmv93oWXH6vBsTBnOXUtH1EG6Sd
9xUY/9XvE7jlL+tySwlFbHcJQdtx6HQV9xE+UvpP+lxd2BSdhnq6wyodUYvROivSx5hzXZIPjSqk
J6mrdefgZ1P7a6INHoq/V5XcxPSEi8v1DaQjtuqJvJaoX45sZroOTcNLBjanGNE3dMpy+Jbuk+/n
X1qSC4jQiUCuJYs/GneTjKNGnuk7F5Lo6UoQRPYxPUbxkgeHGq0HbvHyIQUQo/BkjSuuQym9dYGj
YwkWoFNTosvZ3BNHk0Bwfcd4K0OZIubtiMMlKCUIZKl77skObbV0E7R8jSgS751g6fP5PgPrDIuo
hL40PPmgCoN/unZaGlxxc/0tsTtDOJOMiSgxw3aarLSbNFIMnDpluqCrPLHgVmL5FW2KURUbErvS
5KYMsAE32WyZUrtQfH125pvvGoziBc2GYifcJnWgNsPNCnnlqWlS56kPqgTxJGsTBj4F6ysU2HcK
ghCIkfYI4l3T44cnm6pg1iiPK3nJqMohj3MyCr/xfQRBnMhwuH57NC27MmS5+19/h06gpxUdeXLx
ePYW6W9EOwvT0gSkksuFSJ1PtgNIepHwDky8qfUovNbHGKkdm2vQ0TRwG1tvnhQwWW9GIAqX2Eg2
xBxbwte93aXFzQ1ZbUzhe0c9L5JPSlCqSj33yUHFiD/u4wNui9YCqGpUP2MO39iZu78Uhy8rP9Xe
5LbcHuch9KUYCpFSWF1ErcfCCEwDUYYjTH0qJ1cc5gpnNwgVsaxfD1kpAqYEiRccxlLq5qdwoHf7
n/xNUREOKJN+UiQeIaBRxMx6H8m/phi/rhIr6E1HgQpFC9zbhkYtfvclw7XpsSXRHvKtpW1wEKJN
xbgMIASgR+aoR/HWLgtVkxKXcbgre3QoLPuDRsCc00UPfVfMFuVmWFLllLSLg5sTsb02YSR9Z/la
dzBxD2W4EssrUTY2ZPAorlmFZ0uFL4xpi8bQEOVdBIUVKITP5zqSd2nLZGdzUotRRHFTyUalPM48
CFbZAg9ow4tVy6JmLG1Kp7yspJUKaHhXLap1JgXEZq0JPEfIQhsIBJR7yVBde3JtRW001Ag2WxqB
mu3J3xt8OQC/gGnM1VgQQmHAN7lW0uOnVa5gb00R7fO9OqwGWWbsLnupeLgxkbUVhJVEoiy6jWoj
JhLcr59gGMsG6Rg9oBcAv0i/yHzkW/Xaq8Ol429jk8Wj9qBBi4CDbBfTCkzws2aExAv4cI6cWo+W
l/3RsqtoP9L0vEi7mD+C8eHrJSzA1iP4llTMds39DEbc4DISNOZrmnA2OvqV+9JbGfL6yYyQGEqD
WjFdP+N1jIWHL4cFB0ul4s/3UFnlThhOiK0ZC1PIj9s56CVVGh2bi5iWBFRvSmgSVoRdHTYWYv2e
ddwM7uwyUi+vFi2/0W/q7OB1cNikj5T7ZCRjD8bwfOolobDxPefF1hS4qQEziyhXaxc/tYLsEiNh
uvPfPG5AMgAukKN5dVveOHjxFUMiGPvtBRpvvUpjBtFu+B1ZENFz0RiDzY+wjcNi4+Kg8bwmrcBp
B+20POHyBwlVVhn0pdFKXWubxRmNVz2BDSRA4pGei5yGq/IAN8uzslc3tl+PprtxxD0/k0cYh99s
xU+fpA6yPdwpX0RrAMVlCig4tb3BldmslBGfu68AfGJv3Wv99/40G4K7BEFALgzfHlGVCD/f/ttD
CFEZf5YKlM+9/wIIIRVz9i8yuKogfD0B4WdSbsmyBWCtS12K60PQga037H7gEVirA6iBfoXuCrHC
mlc0jSwiFNU57WV69Q4vnvtjBn9RlvWR0QW+CZHdHg1oAlFfc/H6wbIkyewxpOjW64dK0XMY3vv5
YDbE2V7u+g7jgZBv0vOcSlHTRqj8JPf/kXavwt5pmTD6ljPvtKDeW2gJbRqzGvCVuRUUFTChzTcd
sGWciMztyhYJE9+MpQ8QdrVa6H/umQWy7w0UAtyOmVlUl775dfQP7naeVC6SGdDyqYkqKZq7DDp7
exzId9Qw/HQB4f7NwudgWaUEWEhx7k83t1j3t8ubxo4hbNapMHaz+n9vRSXeXi9T8FaxrEb7ZTa+
llNOYnGAPHPjAEVjy4jNg5gZ7mZk7/iAa9mL2gpYOZlTPLXU0B/8+c/Uiw5Qw271GEjg/5nGs52j
klT6/On+Xm7bRJPKGfMOr/HL1r7YcvqwWWYCSHm0Pv4b2855pwwSJUEoM9SUmlH7M5CLt6dwhTgh
SK4RdGzpWVHZmZpfH8wDC9de69WIia8Nsdp5yZc3P01ZNdizvXnO2oqLFR7nY2sKDZCF4Nr3B37m
JHq6FYhWqHQ0gYFdcQsnIZItvGUlRec+sgb28XwZMN8zgIGK+PE5zHzMkN64QaegTByNcUoHVBI1
S17f6YpnbFx/EV5g/XbEmIzxT4HSBEN60b5iRJVM7m7k37sEJnnMFB01hc+4xGFjo+h6t2Eg8z3q
AGdgbelonZGOrd/eSg3KCev39bNGyviQOhOYAQHpWfcJqloYdOUu0Up/HicRv9o9c+ng80uX69xE
yQVF9ITr90aZu3RBbwhlcwH9Kv9PDfHNlElViuPBrqchDpVa0jyjNPO37IOYTmE/8+a/+drR0+qw
GbigkXvqC+pxnOyulUVxdwJWikjVBMMV77WLz1rh6LS5MIe2FGvvvR2/572Zp2tJppG0xJAXDov9
wbsWPOQG0HY8MrtPiHueUAQ8npJ3gOi6aLxvwaPRli7blCiB7ZaH9YNDDBrd4GqEUDdwVlSfrSp4
nueiqO1AeqMefYeKFQlbfTS8SJxophvPljhNPwaLKjh/y95jji6lKDy5HJBjbWrHOJDaQ4WUT2kn
zv8VX8TEVFDTkU+jjY0v5KnEqkIQtbO7fofeKWs5dacvuyLzDvWMTp7q9aEC1k1mcRmF8vKX8yim
woOH0azg5J3zU0uKmZdAHXDd478n+/PVwJmKQtA+StmMfmWtsxL4ZDV7etXtjrUST1NVPPQ1Liwb
AEs0sH13CdjyLh77OZnBvi0UQMkUxUaNmFNho0X62Ags98lJjCT1OEKllhtuGwhGltWz5/thjpZZ
oUi4V9ZsyI4hLmxoBSGtOIvtYrtzwT8oenuQkQjFWdC6iR06vooYG0FCG1yTr9RLMhk2MKRJWIUW
pvjATO3bZavj/gFDWIZjyPPviD57WeAL8TEelANPmYmhAESxvNci4CxIgKNuvnwBvgMmK/eGMErD
m1xSQjJ5JfL14gt1HdO06zHy0tdDEdZai8q6iEs+LKbW1hfMtipr3z0EdZrFDxRh1ZW1oLytlrbQ
z79JNXg0buwyesDEyz6sY5x36iWud0ZPtl+f0GnNazER3dWiVSkqhrf9n5v1Pc/dGy3cZpwbougg
HgvpiPugQoTOjv0vxrLsaW/eAJbkwoTmOT/IM5M6mlCY440I7YzPfSNb+dS9uT8g+rI+nMytVftL
Eo9b71WbzzxzukwYKX+B6UeCAHAcHza7nL4Uy9Mwu5NhD3A56K/1RYHKrA6ye6oDH6SaNJiP9Q/t
dWWcMdqaqhTAIHeJ9dPYT1g4qmBcgnE3u9REBVtYrq9Yozwxd2h35EPfEAH7/cxF6BDQE2nMMH0W
UPLVBKkF74DN4l2a4YJCkYMxo2zruJMvfz08niyJETIXlOpUR5nMEsBXh0Q8qu0IsOvI+p1faoeV
TpIJpG8UaIqq+0p4JJIsIIsfnOBTyDuUkMvZR6zZSOqraJcPqPmWv78USIm7Ue1MP9So1U1gbN59
ZDAcnD++2zbffT+v1HL8k24rd2Fy05t4zhy/PsX98PnItfFKbGIJHuAr7q5ePl1d8Tfe0eIiptOc
deCctY/bA4ieQ4Xxj9CUxHKI7YyX4W7b880IdWLVlCyY38IBbT6qXiEPdHziW4VJ84Ypw5RU5Hce
1jVR+leLGe/vTlCKjszF7cgAhZ3ws7Oml5GnVVNWtW/h8lp8yyYhKvzRvWwLlNuBEnbTS1SvlOC4
e1t8uFPurDJWklLQSCAGJW59qxksl2JyC501Wa0PPp7AgfnIMXnTBHBVWcBPjmEHqvBGXJPXdcI3
lFhmMDvQhkADRIp2yWrFUYsYImBwYWcPyDBK9obSGKDxEluvDi5+bkHgu7xxODj1VE9+Tq7s2aXS
Lz7wlJ7hGsuAYKcY5X8nHxggYHG3IlM6h8aSypkwJZ4IDW5nwea+Y1WKJy3wmTGONGw842BUGraz
OwIxwTcxRDENSsSI92f3OyCkaHr6OSFZmRwv1/TQr9YRtyzb5rGu2JJatwLnI4JWPo5zFla/IEE5
QGuwrGHD8AgYCVoAaXdyFA7sN417cbBmRBOjfPgo8IJhpxpwG0AaVpYkhiDEIPlMEXPH0Ry2+NfB
qQhXCVOsto1oovZcgMR53pARDE4CgU4bqo9W8oPEpNRUV4hRbNQwa7zXhfGdUHxiwNR0vICCZzqC
wN5HngpBpbyCWtGTGUHBdaBVEjhs9tOM4H2zRJKYzpl+9yNWTxPvM21cFpkCJWol0F3jvv9dN/nb
uyS4BcpPWMV/7/t72jty8OcVum5LtrKAGtFfKrciSfTwJ/l9q7yiIzr+fAHiqbMRHiDcGQDHT0aY
EefuCf9eQru8souOVXeHEabOOn0A8etuxDwPnVKRtiXOL+b9tMKbWApHmjd0n70kMxJyvjwqixh+
28stFBS9snvN239hNfyrRJOyBkVPcF1OctxRe82XgJNyN+7b/VwCzAzHEN6gGBQXiaq2RZGASuDk
7Jn2jtE0HlRUIyVaRFXgo+lTIvNjH5hgIq0ZBXdr3kFm+FY9CsPo1VjbRZC42GHfPStv71b9C3H8
Zoic4ytI2JqPd6t5WlCJZc48G1k0zh7VBsgjYxTvocCilndAfmXf9zKog/jtz2N8PDmNRDF2bcCG
zXvGBphNv0CdE4/goidl/H0hViFfuhL8WrMzX9vuutBWu4BLn3aBYP4dhKAYGywNLAusW472tAwt
j1mpYIf977mU0UkEj0MMhed6xTUgY3Bwt0Seggsj6wRWCm2cSGP9k0i3VjWocTQdeOey1CHx9qRu
t7saHY6yJUQaaCTLryFVmoEihzJzwHixz2QaBt4p6YLSVzJxM82XEVO0BY/WGZJz6y0nA6NMwdkh
D8/r2bFGbMutj24Him3FRH/UePCHHZxGOHfcjUZqqQfGPCuXBHxv6tpKWzz7Oya+0P8EbQmHH+56
+UAILLAq9uZuxG1p4mKMN4dvltJOjEnE/GLfZVdScTKDQhmGtfCaITOn0Wc/7f5yIKzwVVO/f0qP
64Fpjx8BaDWqktEdeVEVt/T60HM08qb6fUg1dZnKLTcg2iYmB5QD+IWp6eKFjaVwzgGwhWkoVfpl
q0TbbayL+97ZRksHB+q6faolyhr/7aUTvSMDHcj9nikOmsnAiE7Z1R1ojcO4WxmUR/LJshFLr3d0
hL8e5b0C+HcRYg3nahZR46uhedmQDtf8f7XGUiEVuvTEXqjdTj+4N6jNiLEP3jAWI2TqzlMSQMWI
odRG6oyeTgRXU3eba3pYsymcPMuElw8CXtlZSfEYH+CQ8tMVaSHOZn6MuQlNgZxM9i/TuLRVuQSj
gXouJBdr9weBu9lKlg9nR9oS80bt+aOmRxvrlGj0o++0CguQj2ZQacfFrb/3ZfZvoJnbFiMnNCV4
uaVKyQQQe3SDHX1gCzqhT53hiYBXQymPRLcjZYFRwGhwHlkfoaO1IoSYXTXIzjUvO2vNw2Qqn3tX
HQoL6ECyjMKPZfJHdGHwn6Z0WmGKpPYzIntADry+J/RLyNtkKN44IOZLMePKkDXuI6SPkVpKH4li
b7xFPG0KoWNmFwukDAOGCra/HqEac+7P2DLlZFoQMcpGnqq4EDaeHOTTa+dqPHyOYRuwVFrldWDw
uSn94B0z2Hr6YTiKUOOYG37DlSb63T0sz5baJX72/F0QikBGhzcJFRanRQYsGBoi2bf+mVfAzPqc
fSBO7n5XufHSMhAmMOSB7hoTkDjSPB47Kf8lLhTOk/+WvzD7nzt9zeNh4m0w8xqTTkvWSdebSDQw
o+bZa4No447EBe/JVjNdA3SuMmVYl7gmvA51pOzF79wC4ak59De6RTZ0KmpPxhE0yB2ToLJ3riVt
IXYstnaukz/FMfBcbnF6ey+bNZu8dkvbdyh8TLjw9xD7OgJdt4+yNdZuYdchuQtO3PpDGtMVnJos
CGtWOZn0+i74R/0hE1YknoYk726GV5BaOcdBzUDT1p7w3jfGwEkC7J5wfwhehdUcf5KxX9ujW98W
uuMRrd6zbyGaYwoN35OZJMOdKSjgzCC5un6AmbBWXlRX5bwlOqeQYZ4Fo2D5xpIGmOaK6unN7gVt
Xdz+mtKdOj/GPdTsxaa/NhSnAvY8x63ek8rvRgtA9ypB6Ovq41HnJjbO38UZLwjThaLPXbCw0Nme
RikJZFpDz5evcOLVGpStXVshs4ZavhWI3gX0bdNVJhiHSJ/0eetVSBhhTw7+rbNVd2AeHFlFTLxF
ihSW8IbM9Nq2WJZB78oLr/8XUTfH6oFMiSGmNhPsj3G3lL5GH6a3Hyw2zZ8Gc6Budds/c8W0Y+Vz
rnWhgzNiU75KddZTU/HPsTEQbyQXu202CLe+dh7lK5IMLKEo1OLHAdQuAKsW8OHejZEQD0ZIahcL
YXuovVoMtmsePr0u2NZKj1GAetsGMzTSMJh3mlzivP8q+tNiEiolwsK60+aRe8/OUp9RGjPB9kn5
p0NkQu7JStc43RnEYN+7+ftcX1LubZwUh3WG1Rre62poEp8s0IXL0TDnvqWAtefj7RsiIC3uxjvl
jcJHURj9bWY63804Ev+wMyUykkQFH8jeTRNflPM3ssG3Ag1OHjC4Zz6sMqdtELVDMv6PhdHkAUvY
vQXrXWeHxbOg0JeCfmaXmV/JbLsylGDBG0YUsQ0tBFcrpqBRtfA5i/LEIW6BaQLHevh2Qq0xp4b4
yeS1Y2ZpjDBt0M7UZs88VLWOBF3k3wiUAVCcDem/RJ93iov2uStA0ZD7lCKn0ws9N2rScHCnEyZp
8NbAuPK4lSurz+CIeRdUXKZX4fKKExcHrJFhdybDaBpKeLvE9xTnTbYeht8HX8FF66IajVGmeG08
L7FLk+pmt0b6rztD+GRnVdnAIj7XLKztGs/6+Ye5UR6xRvGt6ODQBbhPpthx/8o3aXw85fhW773y
0P0Qa/rL1fO4iCxOZg8memg98S6Wq4KGpMEqHYQQ9eAcr9rLuDYXEs87SQl9efw7yYjrTiW6vy6c
DOA+ybKNnBZ0M9O6ppibEGVIs+lOrmKTvFfE8W/5hc227sEvAvbqjTZ6Bw6sY8bmX7wQNvC5FFFe
qfGnK7aibFnA95AC69DXz8UvNJnZzP4m/FMV+FV4UVF9qHV/gSreFTdzmdaBisqAmJFPRQSS6vx5
2gJxRxIzb6AjzhoxsLBTy4/tNXi4bUAroqCR92tfxm23eB/npGhIeezXFP7WnXDpNQXivJvOdD4K
2oP2xD6qmHTsw9S2agWglB1ygCG+UShK2UA/ALqE5kl1F813WEPXi9F5PJUqRA4e5jl+hNbGWo09
KDi6EKYKv8g7Zw8GhiDSehlL39692Qej1lAZPGJXzNIWiX+IRYrAwpl7Z9mJ1XDhzZMX8tIT3Hdo
5rC5+3wGmrB/KuYdJlBBFQQtfNEFiIEaYX8B66FBL9ahrd8nt0efkk22Ov29a9mQvMfHhMFfS0x6
0zq8f8A7zqO4L2lBcsuatwFcCtUJ8FzIINuqga2lQr0mq/A0Urb7jCwru6TZFmPPPnYlPLiXYy3Z
CH57NIPhnts3IYi8nTDnQUBdNRiHyd0Hh4tXUq1fVuemSMGKnvZfmI40+1n2eJ3LjKhbTjqnvp1N
VkwBDk30JqWwPU1PKDwrD1VqV6FfAEMqSR5iE9Q8n82SYX34u7QVrTs3Wc6xJz5Lo11OKJl9ewHy
ts56Ev9Ok9mif1QmBj3SNKGvXRJT+RzFRveoLUgJAuOskWWgY2bF0ZEUbUc5NvsgZC6PEJdu02Rd
1/Ab/sfz1JFTYeg4u6rbr1E9YGjpX1cfkUBqxRT2oQvPfUmkzSjQhnRGoYuGhFJPS44vRczbUa2Z
ajCCuswBIUAglpB9ThTc5JYgAFCOZTCraeQewIVe4/val7iPbpL17Iw/FF2/wumntO25L26OuSgC
5oxJOaq5on4laYticVOK/mEjF6YFeM4TK+XonaGNPq/RNqc6nwXr16gAMxt9rTTlpMEgrNCEf/eI
xx1PM/I09BxeK1cwVNjWnXYc6dfUISiv0TWy+cZUg0SLbrMJ998MLoqF0OsBrbv34ycroRbD0BZ2
6OwgsxgFRTUAsvrhmZlyUV0cUcF+22KhdyyLiY+dT+u1tPVPERxZz8eAEhcPy3d5ASDbFC4Bj8pb
Cb9M0+tIKPrFwDDZ8k6H6urvEcf2aMLpTYO5Wu66Zr4hTNVhaOaTFIIJq8QQVPqFrNWCtI0osglL
LaVHxJjdXbWRdgd0lOkR1Yoc2TtRyLk7ZuPskkzmuhTRbFEz1aDEEwbuGb+DHEDmklKX6ooiHlvR
P6kCj6aCDnnFvtipbIH6WxNOP/77i4vhfY6guhwvGumNG8zAN0Al/wSsaWWHpBdCjoQ3C/V6Z9kd
HAmSo0eCrCPUUDRAt5w4FBzs5/uxytMRRceWJkFZIZUoS2H2QeKEa0g23Fs7GGbzjolx+65Q+ozd
RAsjcvNLvjb0Z/2lA0ioS44gGm1GyUVjWDbOJUM5JrvFwd38T82CLYlQyxSp1j+gPT/lb+3bVYOM
OJLjHBO6VmBUe/dLAZdXwfQhoLAcTrcBObMuB5Jz9S5d5hMThWAK8UarCWtUh3/TIUPzFevWzi0d
8RmdvdXPnTi0WSpguejXLCeGyFUrfGQnr5p8d5K2IPmERyaw9IDmTdtheZEPcrPXUYGbFfPva1UM
xTV2HfBudRO0iJJPZsb92FI95yKhBVcb7cBl65BkCyeuBFFf+AXRg50M+JdJn1Dg6LueMLAysTgy
L0NJCWPoj3/s/tPfnZhpk57Jy3zi8S1R3IDlqQYGVDC+I2nIuKZOa5dI9z4JcUB+v2Nb6ItXQtht
Kn4/VWA1X0Vlc2B+4cKbnq3bdENCjzIZpUNuE3u6+Iw86peTREGf4cTBLxzj/twu9k4N09pwvEAh
rorHpzvaNutro8zTG9Rds6qgD96AK2OHpUJWGVfn0+vAGDcvZBVbXp83923y6P5OZLE7Z3qm/jJM
9rk97pod2rfYBpoqMo+zAcqGwya/myETjuZaHzyOEhUFquHoI0CrUEp79mkTbvvWzk4AP+pw+2yl
FkgBr7NYvpl17imOYZuRpryS7dSwZsb6kwhbsvt7eDk8rzjyH5ktXxFDtBb2Iq7XSg0XMOrNQVPq
6UChEbo6af1pWiOxxvrwYUxRAxFoZsY4FzYb+be/RBz7PpoyakTSsuuDoN2GRcGCpg1eAeBv/eGb
SyA8JMq6HTZyhYAD0aC1XSVdvqBqdxvAluuUKHSGwAQ4jQ+HT8LVP5n0XLBP1PY0hZPQBY1Q2g9o
yK53ROpZeQImRztWz52OFbd6y/YwQz61wcy8rarW4BbyylCBiVQQaDwwxi766sbIuG62N573TV5M
bDAnt+HlxnG90lwIN28o14VeeKj8JCp4RwHWyo/ppmPipmiPDcvI+twsUrx2AQWBlwp3sw+TJpcV
8Pa62icquiP325wGqkOGnxUzgNNt9fNyxpoQouAa5Z0j3acfI9iabdT9lxKpbCTXxdT3J6pd1l9O
6GJFm0H6MSWW1oefhN3SCS93OAvk2JnVtR4euPf8+jdreSNMpsZbq/JqEDJJWhcOxHcK5XsSm03W
8gpjibWyNCt4zxepze0HaDmV+VN5+SSfvSUl1HszRCpaNykP1BUyRjqaeVZ4ohhxuuGslRtnBa0B
c6QNMrQbeySSJuQ+SGtnL0ov82LwW90meCLzeqJ6Tqw7Ee6Atqs4kuzWphrK5LtsmgsqT0FNW3i9
dclQGUG3RJ7IZDCi3qV0Ro8IRHtrGxX+q3+gPz18arTpyDZ3mS/gh0ixAccXihkY2EUpVbguZobS
OldD+uuv0eDTRHAktO+J2zsJ/rn0Dt5SXBIy/bRMu9F1re9MvP+GSDQnA0WagCW44jERLRCwZIlI
U9d82Jzs6MSmPX45qvQGYBqbuXxPr9nqEriY+UhbWm/7gZoPnWURHoImpuvLHS+ZW9zwhTKpAA0O
cBjJ1t6Ag5/wOWTEwLfJ931nSRQr8ommT4nszW9u+rckxEvFT3Izs/FXZfAoO011H4GUEF5EMq2C
vfgGWIu2sKMdLBbeKbJ5FIGYozTeycn4zhQy/YJ3IvOHyiyM2z8kMbTMAqnEuq+ppj8AT+NbqDD3
JTiZ5+QQ53D54ElTAvOL0vkt0swhGOkzA6ht8WpFEw3s2NoxvPntZ2BgflPycvg0LbVEkzJOGpWI
ZvtoQWhlooO+7v2IQfm1pA0RaY27wGGFhSpc0tq79/OpJ44rdX4yBECSPHRlxNWLeSInaIhFdKHe
tFAWO0jYh/A6ufTJJ4RATtBvaaNoEZDdsYomMTLBgfZVVhs/GidejauSvvlfgW2jsFbBLA081D22
xkrem6oVKV7cm6vkRPUZopqkyR52vlYsbVFFMTbOvDbTY+ytbEJfeIynE3265FTKcAyJhL3k7REJ
TPRQYyrdASVqn9rNE0oFzFFg6gLkwLHCvv5VIoQ9unBfq1e2caOh19mvdKXXGAtiG+dJdC9BINxb
SLPa5LUMzS5V83UeqXNhKY+3NZDAsZB7J7wm1PTK5fiaqAUFNm/cafrikLyOAt9u6zCUioViu9N5
qZM+bZJawuJWFOLrESh/r9cnNhu6U18dlHlxci0XzepsLbfRHXDmA4DMbz1P7MZvkw4ekraTV4Z/
/lJHenXG/KumvlHy18Lef2EzfZ0R4vf3hkh0ynBqJ/KT9ifDXKDAAkZoJwkkx/yBNaLQh4oevWq7
BRa9fLXSzjTwYDoncSt1iw2eZVLfn3iRvmIQ03ca2D5wd9z/bVMGFkbSdSZRwuMlzAR7gnalM5m6
quJi69QmqWJ70w/tavKXqDGBwIPJC5eP29cKBMe8dR6aOpOp5tP8aCXlORuw1e+bgD3nZ/3jWvqP
4HlUcU4xhaoLLebtuav4pDqmzh793MqPSuCwle4w3liUKYO6VEnrvugM/fCWFSH6Bob55f1ej1U9
rTENhO9QnwFRJ+qSt//SoKIIGIocbyGyFqmmZV+Rjp3LG/+drcM+Rea4XFLL0+gWabJ8f1X3wcAr
Cx3JBWPrUNG8sWvZo1vvGg8vM1cy0dwyEMyJbN0rMPcf4TWqMXjcwRgCd52zjlke0wEPanVRVxhe
81a/VoGDdriJtIaUFz2JXYNubRozuQA/EcBThmBG2PZrxjcyf3XW1cbR5Oo+ggyUVbNMZ1PYusUX
cLnRoUPZQ4Wrk2HazmR7D+PxA7sGeU2Brf4R30IGgLWvrIJtJRvQTwXhwGxVoTkWh+cSWHv/nSCc
BS+LoclZ/ZhZLKXb61qOVCcMGzst/9WPnUYTPubb0uBaEJMshelYrNNC4hUQulYRcynwuTb2yrTh
eR1E9z25RSD9CYCfDCgTfZqrqkF7T7ARKVEhglpbGt8+ILhj3e6FOWRbyRTsx2olbubbsUX5Ww1Y
9dDx66q0guXoWkUmILsjcgGNQZx0+6dvohNI0buekMgqsNAgWFg1SI4lpgsNZviX77pxBOQZspGp
Kk+EZqz0Ct6iyB0PTaYdUGclPDoReLKwtjUs3/v4VaAk96+ssLmPLUBho5AnqABbAE0JWoBbnNbV
Ug9Vj0eKwEeIBDCDByjUFxcT40zeOJ42nf37Aqj48Ct33arRNcAi8fxKCSwJuW3D1JRW4aVF1A+z
OZ6IE9kyxWinO7aeT/Bhfb5faacRBroDM1sKfijjSAtqqoHsqTLV8J67Zkk3lSgpcLFNEVdf9e4q
tbzQm16opc7/gcUbmrj+gqdtrl4DRhpgb9OEk+Yl2c7phDVcJMX2qviphYxTymmwSpM7wXpv35BN
BnFDgmLFYf+leUk1gQCqS5ypGQhYEqunJxQttJr4QdAHO9oTMuTzd42eeJ5HXk8c+CGeS4r9HC9B
tTGePl3U99S2cb54VUwwdmRA+xPYbIU1vtli/bMCDS7Yy7iIb6hltMsqMevsiZsJPrKY9AUaV/3J
Y7ISHRYPHpEiMz0/xwmlj7+XI5KLTDUQskSVgqBjLzBFxkVWWpNmEIRFMJzFdQTxvX5lAKyp/QCt
nykEAIRUAjhtWOUbL0AKckkpu/L2HIcIX0+BrIVc8bb4A8XtuP8lTDgcNfVFlRa2dwx5o+N/l4hX
+e1VceQqBc31kmi3q8BuFW1AME+2sb6dcp+R9iOfpFYxz1lV2hbRI+jXTDx1ca+we4q0p9l4vxNa
j54aBJgIUBzOsygqdX7cQ/Fa9WCn+0vqjQ48s431ghEjzPna44uwSiHoMCkMrp7Mc8b+0QNXqkfn
JtSb0Qkt+m0HWp4ckNkxhWxIjFXs6IKfqIksA49Ty6ktZclrytG1QZzXIzftreSqj5m2Ge2KPZGT
7ZNcOMwYBslrev5HoD02Mh0nSGAJpQWABZ0aJ13O1lQwnEg8ZctW8Au2IZR8jwz7j/fl6TqWiQHp
WUnWtswdXIBQW9MHp6O4owvNjTlDFvGgtUEEAiptfdf7bDGewYKrOyWEKD0z+WG0hu1s6YPi6Q8V
JsGH+cNAlh90tw65eC6nFJPglpArsQVYCph3HN2NVKoEopXWTvLOzANshR8NJ5dPKH8Dt+8llJQ1
zOuHpMAYfkqqF2Qafz26WKPNQlX1rmByAgOP3m1N9UQ7oEa/BjwWUvLUj2lX6KVpPFkbzXMaIUgA
4uVqoG2eTfZvQB9lNRupHzUxgPq6joLvW+IktSHcNHfH5nkc3D8m3OhuIUpq3PhFSwg/HfN/lmXH
EiYa74Ua2yZAbuKS62tOYXm9kuTmbEQbwg4cZ0EAD/ATTRQ9Qf25jlb9RsjR1qNEjk+Rw2kag8W9
Bo3h/kM0kVFmmlufCZv0LyIkJ0HUUvFIpLotGOM5i2Mc2OV0FKWvEh6V0kz5AAjjkryWIdQDy+bv
t6xntYTCn4305hRrFqAKNbOEzJY4Hq4ssUpm7BNeicESzh03xv3+OsrQspv3UEqz8tQ7E3qGDkT0
GWBReqOerEopB9j3tidHrp3kX2NljiOlpuhhve73ZYtyILxMpDHGs/u3hXiy0raYQoZTN8FnT25a
pYXofUskGL16Mlp7DpajPWHAM+VCzJKWo2GMxGYDU14VFaTZxqCDaWOfMaFgU8bAsgDGpV63oNTZ
JudVI88pYzLubUEkZN5PbqebeDyzL9sM9OaHtPTg/7qWE6IFKGtcCVBxNMO9WabxlfXClfdVJ3fD
qmbMDJ0Zq+MCddLy1ylv4cFwwvYEeK8Qp2CO/9heBVs8p3M5Gsh2GQzrZ39UnB6cAU3yNvUXwDLY
8XcgWhaQD9DhTdTCM+6TEEUVtxUGElnPNyx+swSQnFem9dbCobfq2HOW4JZ0knHFoB7MWcVW7D4c
+Ny+/i/oqpeaCAGXvrMP/9qKpJzNuPaY2B2RGqMxR3742Y43Fcq5VmP6XLJhN0Ah8l8Tk0qun50x
HJKAi692WA2U7qQXVmhLkcO9X2d/rg8h0qoQcGyMGUjkx0M7gvrMwpH4iSm9uc9F125S8kkBvPjz
sU9Lhqx4RXgOn9FqKE8tZAzNMdbrDKBn5wDgYCwREzVb3DAprFIl3liM7m8a74z43QId0DRYxw6m
N2fvn2AyHVp/k+RkkrVJCw2MWAlr0nUUb0Iyd4buX6MeDVdx/Pe5hKDRSFjHQW+dIdqaHHFrOL/u
7CqXk52Ka56rlm5fa9dOTpjP5Wqi6qGxJdu+NO7gvuopRdvnc/qU02ZmDH6a39C1+IDIQ9PjkA+q
H2Tj+sPKplNowzYLGzAvmQjKuNPNRhuaCbHbBBFt1GIQGhSv23K0ZQEvLrTyNsHB5CAGU2Cvd0HN
qHQM7HowH5jT9pP+p3z+xDhcEhoDuhKnItPuTRJ3Bv5huJgVRzovrBaCRU5lF7NvgFxplPnv3EOK
WOQUabWW0bL21ekEC927I8WyPBa+XL/y9oX8D4ftNzVEq4bquOjRuCjztppKlEg2uyW6n5sPCpQG
bL17rgzBR31D/qtc1DZqLiXMbUv+J7w+MIqXjlZAwGZcEosUsWghJift38B9gXYelSE5PRUhDNur
SXaesigKNxxa9SE9lUmw/ltqJB8WsKABQrah37NUz4+rsXZXZUNd0xideIED6mhruqttLdIIAeUp
G98E5pXKsprxAu98pre9srcLo08zTHcp+5vC0/dPBeptgIhZBK4D02vfJpAkfhn2Qsn3rYKZB7uX
j71tQHLI0LKjC8b4s8TvTZJo3AyevK7uSD+SEM8WV2Tk8r/fpcDxJPi/XFseiGO04mb9FTSIVgoD
HUoc07BUz9YeZsqs/iVO2aD+FI7imVV05hhldodkP/44b5fdeKVA94IrfqtBWWq/CU3DEOarE6mZ
5c0B8ya7EEy4tHs32ImWzkBV34VifG7QtTR8qCLIwJ8vXvdjhgCMk4zxgH2q6HtetqrJeFL1Raxi
HLSAF6bh7kqPbV4tnNQ77PWeM5p5bwrJ5DPkj+3fwOhCZD8BQRuiWRANYzsopxkpbNAWq5tscduT
9H75TCcnVFj/1uZ6UoHXH73gy5lRyp0a3WLapmAvD2/AC5zo7/chpPHRLVP3cuWoXyPlHxEEpUmf
FzbYLRpGb1hdp8tL+iRhhTHsug30juK4i++vKnnlSHIfTZGnygJrmalK6+Pub9jzDxTGeI56ejXF
3rVz3Mzm5KEKE+mcaBTJgta8AVeCzTkOfNFUeijIRbqPwR5ljcqmd4DzuT8YcC31oSUjVGSSl6iR
1Lrse7iwU/G9xlQJl+YDH/rePUK3pFacy/fQRE9Qqzp60BXdGYOLfdGGAdUFYkVRtduYUlRNkiC7
bxdqei8FaUZ7VVVVAALWVbtoE0JKe1blrZIyDo2CUvUeMj1e+K8vXO4sS1qehT9gKITbpubKjgmn
XP0AbUcKchEKYY8+CsqvK/44oC5tvuOa26ILVM/V64KyRUdojnLza7fZCSgpmijenzuzmO0ck3Ch
5QZBPPFGZaPrA6mhFMqkv0JyvMbkEHz6fXARrWJ2UdM1nC1GPMnzDL8w4U7UD8lPiuOKBWiq32+k
Rb9HrzT3bsq5WLYLHE1O/fCTMBjVhXNL6u4+KYvmWSybkNvb70OXvxZBWwlmCAxyr6DfdhTUqr/K
42sjZrF1vvokCgMx2vlnnfvqqetF3vcpHTLDuYG7RtydfeUuQMjj11suz4EEDXhELOLsR5ScDa/z
8/Hn9szQzx6I9YIrtW/M3T/dx5xmepXOPa2g1mBcFg8Z7k4Q6TV+JGQKkR8/hTZV1BdmFxz9CB2m
cATJ3uWgQZ10HYf4YHSrpPGKixVGPK/JfZzftzpo4IdLCuFAKeOK1DwKFKG4eYPwUSeFJbgAQTNI
stcMlOSiaCskGv+sEekqJDcJwyvoUZtg42Hs3xQa7/+yStrEXhO2M47eVmcQA6CytQlncjxkr9nb
XfuGPea+EG2FzJmb4zmMZ8Z4yVidYMwuShHVEbPICVbSmQJUniBGlHDPWJaN9p43qUUVb8U2ZkTS
6kNfnpQnZDQ2LJOi8fnJjVi3ZYW7ldT58YYhjGpx452s4v6o447IRLTxD9Ng9kQv8x43m1mMAxHl
cLgB0Osion5qhyQkb5Jyr5xCzP3dMDJbjojvx0AuqwGubvZ+Y8pbS5csD3LG4jSrDSsoP/O5hqI1
+KrTEYWdqsWNd47BUOj42nJYZRS0aLlq2RkKeYxmWZhAl0M+OVcBZJFVGM8qO7edvyGx84jrm4od
HsnCm6SQcN8LvshUXgDnhC8uDmrCvl9DfZCyDeUEHLXxAMcdH1gmLvlc9sFMr9Qv3LlM6iSOGdYp
8SUmqUEy1rtrRZoPoZTbd3iuf8cyFqWXQJiKhpC8ZsTYh4DQ5KITLGulGDVr18nwnhQlwT4kWEgh
6nOG2U7vIIP6qWTWo5fNYwpBcGs9YmPUzwYr4BXvYkvIvF0sICvZ26YWb4kRo4Ye+dKRt4Xi/VAu
XMuVZDOsLcy6pd/vJzr0yUlxUgvIc0bOakx417iZ31akUleTxnOppfMmC0OIlCAhybP8St27W2xF
QDr4XC/7MoSQImpdHKjBO1/Jwh59W/NwziOm07ro5qtIMJ/J9+eNWZT3LBkj6Okge6AArxB+OsBY
2DwbqTtCeacoA+3ad+sCb3Dcf7/ksVbkiocvsGbGkf+s3Z2ezZIRfNRqEnUS2Q7pUNda+Q4wxJTE
tKvxMpfeNjSFS5AuydOFRoKegjZ63Shyc8J8QpgSRh0xc+wbq7l6u63RZLKFaq4joT2h8qDC8IVh
54kTyNsAxSh4T3cx5ug0jd7pQE3v5cxGKKy3c2BmNBh4TitlSVtvswsrmR012N3v3Jvc3iHKjV3x
1vKVzYjfGoYauyrI7+uCMYQ16uLdmaa7pCwJ45dm/sDJPWRwSPNnsK7Aarw+nS2mg/WPch6mW0UH
X+4Y26CxNDQmOTRvCgw6xpAX3s5QS4BEs0mdu9pXC/vlX2xZZXSLyN2+ZoTxX0aBY82Sn7f2hBd2
koSaKcVmp2aMYCzRk8obqYFMj0FSh3je5gBf0kXuxWumcerw7ebNI2yodgqSbR5gQQPXw7si7BqG
gtgQM1HCPt2AdcM0GyKH3yC7C5InwPYiGEgpc/7h/wStF0I3h9cDI4ujxoszjX/kjHgmbBckLfXa
pw35OnRpyTsfZYXktVcUHF24QKTgLLNvYNAu5J8Oi5kRTOP46nlVKBf0ZRcMido9MBMnud6crSx2
9pKaKy7hP0HDPGKfMrzIO2t3SciJidC2zZwHDhUle4hw6pM4hM+jHPzQK3zKP1+vFCSPiao+DCDc
BjjhfIjdbYdrSLJSNrj1X11SA04UUPkj+qhQRj/zkb/sjrFXll+dCCUzyU8XjMZ+/60sb6WTlrCs
Pe6mAC3I505VaoFFMDpD7bH/rvnHuFZM2pEzna3oHVPnJUG29WOYRUNoqI0Ye/E26eFozT1Eea8R
4w1EU6/lljLEo57jVdG7mjithu99OoRV5Ew6HNVSsWBGQznJ9xQmAE6Td438Ib7zcGrzTovVEZ+v
hXMcM5Zx1PUuCyJfkuFkiqjN0BPNR4loOGHc9Zixyj7TM8SA6ZfRpOj2KUJ3Da//lm5V7vxy5lZY
r2yAcYmTlZHX6bvzVWFOHGzl6Q2LSduRPoFmZyc1ePKWDxe3vNm7oop0Xth2Xmn+w+xmtV8zEGVN
NgoxBlTIAj1FaVqUPDl6C01RJIBWRLigjp0mIATqTW9eF+o9hnhdnwWmhmFrAOAD0WH9QoLED+Cx
m76c6WiPtsZ4zTc+rALcYJVIsMf9A24UFVhpsOJ1JDOfwwl90LCTBWtFAwhZd9sCbQF6j8QY1rlr
bMZdHl5aqIXOMuSB9jyj/Wz35JxesCIAotEJGpta6jEqBYZ6EBwwpkulugg+3Bd1HF4CI/03EzCL
m4URqLaeksaB2AQo5cdqLRkWNeLlOLMD0zlRUFMJd6n5C+Qrz3KAH5fqm679XzBjlYRATbeWTGo5
eHuTcJ/o6By7tdGnlpIi/fCoQSa/lAx+SX/Js2T1naVkV1pPT1PqKunXQbt2dcWWeohK8YdTLSaS
suxYv3b0qw3BxH6kc0QTqwvg4IMuMy5Uv+RFvo2fbwgFcRKF2yxVhCP7jxSmF595/1IeqsPaPUUE
v15TXyGVFjRJa92aMUA2XkG4tBuDzY5FU+9wt5bHkqZFa1gkdv8l9cmau3QNkJ3kkiGLmYOdo5me
3HuRQF9GQ3/5vYdrW9oBfkjAdA1Zl+crPSjQWttpvqKNsmQX9A/cccqkUdhlTOB3F/ITBxM57Dxt
i1O9cN+9HgqDz+XzW+hCr30WlOnHwIo3hP9myfBmRm5e1EoYRVc/oxvBu9GW1mB7g3wj2KONWF4U
EGzPmaUEmuX5iAmnRpSkrHmgTn2jh4I+rzVnuu0LiC3/p8OTzMyrTeGcbAHh32XFhEd7XsjZfN2H
PhyRUOnLvuk3zs/yaYeXsu+Mf9scLJ0gZLqKRT2lV6HeGxihgA0CXx2ZPhYkZN7LUKAlPe4RgzWr
O4d1lS+Sb99UNsF1LhGKtGrqaLu8lPAvvNEP9KMMQhmjel/rPNsZXp0vtLtgyWcH8i4iH5MPqcqq
X41sDx1eYXzzkuMkJt3CQjnLP/XTKi9Lyqj4VIbFqBew0PWtXIFJnAOxsvbszLwfGbVSFVIVqwx/
fkpgzT6Zn/1ynaQFM8QUNmOS2dTo+Iu90YPxLhnhu7hmEnvjHcmxbvwA2BTMi6i0CYbBB+hRba4T
3hittldXoSSu1yRynM/iy+VvNbA6i7By6lS4F5t226pcIBVYL0oMllCTuhauq3RT6UmZsDeBQWEV
VTCP3xNvL8g/ngudZ6V0jGjzYr22x/ktLgLFq3bTJRcYjLsrpcHR6zcRW7UxbJlq7NNSjLZ4q5lx
xQegAzzvOqx2K6imIkuS1anSz2lxTX5ITmyvPWUTMp/rVT40xA5LNB44MKV+K9u9voR0j+sASPss
pbcOwsxO88/yOhAbW1SAZruwfASNqgCyR2whBvOZYU2UIUyBrP5xRASvq1nhGpSQrOTKHEOso13R
sF5HVCoV1pre0FhMG6NVmJzp4Dyv+fsjyvziNbJTPESQEmBYHQ8z5d+RG6G5MNjCzI6nLWEVvcTA
wIogl7XV3qoH6hLkZarrtNZMjFyM7CypkrnHmSy/B1SMtOPtoyFfe8tTpDPMMUQeJzNB8SLVSmXn
ZE1DAPau9EbR5pdwcnkcZASLw/88xuksHNkLs4CR+Jl5ghQo8tjsESpUCr4j/h8NO7cTq7GhVCkZ
lreDhORw/hm6AGv8x1PRctEgMbr2ByT+pU1cZVGXHyOg8RXhA11GGANJbQSyqs3+IaLAbUdQxc1r
U6K8irfmqq69pBxFxpO6T2uoxZjkE3aldP6J92zJpVKhAClbgd8D76XcysaGoU8Avibha08wFnUZ
nznNJhoBl0zLyXlKHI2gSTgsc+IjVFpXmUpISiHUyO+OXmNdcRdd6/hK9kFCwaga8oDG2OvSKoIE
nLs25cMDSusj0g/76bntZHr4yeQcyr62BpBK9zonMWIALJR+f3QqaKljOUNBm0/upSzWj2ZnQTb/
O6UrdY5NTtx5zl4MzFqIDYP1vXvyBfWRqO9lcH6fOhJXn3Xb6oUFDAp+qkmXNYUZTVVPqLUVFcpn
JtNGdb4yqeOhIY8kqBNSkTZi5xr9ryPPMlt8H3vpXwfAvu56SFAJWfAqsdqvoh9xCsv1rRroP65x
I2KTyYWwOiZwrXdIvjqjMq9Na2gGz6ST0S4XhgLfvT3sEfmAzdpJcCYVd/fYQBpxE9RHB7fZ2eob
OTnrePrlFRPOWXxTnD9dEjz55brKUh1+F12rVsy1tjHl7MpXT889VIqoMVLlXkUtWCGKvOBRNREl
TEpZ/sdhsF/hsqb72vJqTYKMBCTdDfk4gxASOv6yTNUJRcz6xwvJUJpfkWa0uGqBj90EBPGA4vfi
VVAVpbJd800bCfW7BugymZbzRlJdnWg3ts+LuNhHBqFJZn6sp0V76lTjhsJcD6uhtXvdnv9cRfbJ
x+ReFLdTniACXo9BisQocjj+E/xQECSd/2EMoQh6q99n0TVR1cBChixUeNnI8mSEgvPFi5elLveF
UcTAAB5BTGqJI0G94+/cO9QQ2Nx9tlFrDadpillcRXDg3+tTj4YJp86x93xAd03CF9g0dLAKItgs
/R06x5YE5aTjHthjRtFB9VueNdamNmCCd50isevSt+V/TW6IKqY+eqlBTDOh8/4HK8EDX5iAmHnE
i0Wb9nNzHtgAFcDXAptGQ4TapcrMQS1oRc3qR8fHi4bYqnDSsjB9ZGBIPe16ewrglwXopX72tjUQ
h0SFxKcXnzYQLNYAaMAhVqVBOOK3XTE60K1eufHbQSdEl3GW/You0Pved3j91jn9ZhFgxWKeWGLV
3Ob+SmEP8izpky8Bn9smQ+cxOx5Vf+t4ss8iJy3aD1HzV/o3AviHqdoq0mOT4OGDaE176t93SXrX
+GVxpwC62oufeQrE7yMqcV4kXPvy7U17Ax4P8I3mZXy/xOK4PRu9vONxjlh00fCkp+2zqVOki9aI
zR/tAsQHkEmihzkQbpyVIeBHEw/FnUEBjmUULw1tBjhQluT3j8uYCDzpXRJLN55qZjNXDdAJiv+X
VroIU7HW+URbVE/0qHucPrgPqWDPChWkwz7j23K4wHD7wLBW1YruDgUjDh7mCWz5w+8otaYMtzZk
7inu1gvLx9yb3+MysxVS9eoXracfZ5tmwsxSxmRB4WxIWjCuMg2ZMRRWnSmk4+fhWbaE4U85GdLt
BhAauu3+2K06j5zG+lE8ZbY2nGKvVADUYTe2mivLDTkRNoibOcEPbx0W2y1tzzDap4xIk6F9BtfH
+/oD1WaSnPgrspSiq9OoL0DbrzmtjwiHrBi3MMU18UoiENVc7VM8ExFT2g/lKa09B5ACbvsniO+7
bW6JXmFKP6v3tYUw6h1vRMDwUxta4/MVnYDb1d5E9A2fO47XnXcz4nBJ1fMavfPmiZYtHkn5KfKe
El20cv6x1Qi2UOfyMjCzX0djm0V85vNwJ6bCd1VL6FstVmCw611Maq+G1rYbO58xKj+mRsIoImip
9veyhIhBlc00ZIRPBvHCiI02tYiXq+DhgseUUFKPxiGCkuHQyVAnFUI5gYp4a9mJvBoMQmfxuK0N
wGwzH04FBBRJWGJT6ZPgK+ADwW1h36+K/I3j4w2KWeohPAzHI0kwa65CYHiWdg2IxH0eMvRMJuop
Wvlq3tvZADy4K3qMvdh49gy47TIoUsh+OmnI+LHq6ks7CkYA6l7FkHVvVmzfksltL8mSeg/OaY2R
DE1zsHm/NbM1I5pRVUZ0ZSV5q/nrnk/wObsrRyPVtml22rS6D+1uekJ6rsv/csZG/u/i+h/hpviV
ewJPWQVnGrBF0BWNAFbrRqPXijGfytIftlWWwfV3F+m889la4ExB4MBts7rDYmQzZUdo0vcqgQ6i
08XeY45D4uQHOs7PLrvKeyLXMBBzuUY1/y714PKpCoipdSyoG/QMt/Mqka8lXNk38x5n3FzM5+T4
Q+itSFRq7YXx0IeNm8S7plZ6+TjsOAUHjv2/odGmZJJvL7NxpJNk781HDeJ1R2ErHfXzTVAYzN1d
iiGgSZMmkrUcKjZvC0hT0D/Lgk5YJivIwM8+nh+jbB2k2wu08R8pGP2m7I9kpcB9AlG5GnmFqHS7
wtfDAIzxLvFIY5gbP2JclDN2rQ8/zaCK6h6VWOlTqEnKk77ceu9/LEwW8JweELXBV3ja+q45aq+8
0H9kPmWSngHeTakRQ09/Y9PFFfd/bXyVDtwViQbg67NzipNrDvQklJEih/CkiwtCngy4B/jtNCZ/
40UCSLsVCMMVFxhkZrAOqgVYaW7m+TIKfyUl0n8mHV4I59Pu0MHKNCDmZZxTYLSzDuWU3PbyH8uU
P77FvUNXRU+4H52urXV5erIq9LrMYpEzh7ySdhSkGC6+nUKxi2pwQYYgeQzkAATy8k7G+8roW/Nn
hgxD9HEc4GTPliSYt030/bH9jo96HrUwJ8BByaZbGTnMN3BEPzHKrGLIJ8SmlfHjhe4jvUlQ3J4H
60koQUK2zMuC5O2DBWYUDTkLbOaNI3ZsCypAv6oKc9KfoCbADZhxauRYD9ImXabc7xeD7r8doagL
LNZR0Etwp/rcllRs7phmEkSdt8saQJd/XbJm5wpFDbJiu1o85TXV7bZKYuGjOjSBvZNTLVtFXdDj
XfO3ql/nCW7g50NrJ1HCzWb+2NLDVVzfjqICpPaVPL7uqs3ijrUFQLXbm/4G28WuXKwIguYhZohC
7WTHYPfH8ADlBIaa4QYVlSO+BBWc0+PUGcx6FbCwdyXfbbFUDxEyYDhsaHxo7WFhi/8FDTLtpBvo
GKHzFKbWo9IscoAIhjJUORm4gieqr2Coh8ICbpiy83mXgKMVUCN4BhGkR1RQdGMTtSHh1/oArSnc
n5KR81J+MGq83XibA2yuUyl9+l7i8op2IPqkidP6F4AkTvpFpemju7kqY3dm1Od9ROR+RzCCTWoq
kPeBpLATmgNUJMDVH8AEtqBTQtfcRpgrjSQNKEkvb30XxW7LfQ54yq8+7MHrrbS7ZkPyjsj9K9Np
oZqTXhl1g2lKRvzwCtTGWjjyPTIasIWK70tZc8T85ZiKt3WSyXK8WmLSxdy0Q69AzDJIzUhrclaw
lVinkR2BFFs2bOg0aGCwaZ6cYpzGGvwb9Wnxf8iEoaJTeyAZB/vnGpdw6/UewEWQJTLv6heDkA46
wGkKShMuNINKB9PMHWhmwPGZyBfZDWAhegom+Phncufa3xqJniq/LrJhjpatlw1eRoG01+l16YRq
R+qtE9NKZYQQO5lca+/kXYaqN4dES/jr7hm6SzcWNw52T+lbVcNqf1DiTxjiYhZC4cSAUMFcpAXV
ejPthRz2vqOwH8520M6aa+oAjYWr+lLulj6r0LG+QTvIRh9/XzbRXbV9mt4l+cVp4wKn8JAlV0jR
KQoAYWTiopNieb32tiWVMst6+3SUPAaMcfKgcukb2WPb/9xSXVN7a9BNxu6xksYK/ou/lZvFCqKw
BGfOoev28WipkFhVke5B9MYZnKQ9tCMq8UK0ulVS+PNOQ3yqdoTSSCJryJqUILLoBcYn0ypiHt79
RkqtCK/rhkSfHhQ57gdYCYzcB+kXDviWq4yLm5nwKOkTiU/6eSuwnfpZURRtjttvFBHM0IBhbnAX
vxq7RmPvHhQWP0ZgFYgxrJzrPDJU7cUG5m+NA/6SSbcRfeb5We9+b5gPeh7ntZ/SJ3VRt5aV8rbE
2MtLdFNpT90jIKtUCjZ92LYzIwBMr8tga0iuxrVVH8r+7xITxhduZUL5BMWXLitZ+3sy09knXEfE
NFKnuJulyX7bLG9u4y93aaBL272QeJGHs1XDrErxY/0YFOC9CSsEdHpTumTNKansVLSIAIK7OmH1
GCXSoReNyfNnzZ9cUCy/7gASoK8EL2qHJFFJROHU9UIlHB+QGsSiNykR2zil7r/pJZj63YoUcK45
H9W4i12BylBgYAmklwo5TCLQup3nMyyFC3K69LVfgLtE7PX3Rhbgl92RVTZFuKTbfI3q68aoJ98s
AsReJDYm0UxpneJubE0TXSzaHTcQaXTI/4dCPA38uoR3ErXpM8bmewJl55Cc3Z4LzHk/ZMaak0oA
f2U3RmEAXtlU1dxF4GxYB+YNSOsGcWBPuPr+4iXIY3yV4Uv2Ian48jpKcHJaFZFDH3ynyWQJuBag
LsGryp3imSU6Ipn6QD3i5FZKPeCVS9veoznLogrKmj82q2BntCjBoe8OpdKItl9d8BUtEKTC+ZAk
r3FCE4eLcQOS2ryL00FqinYuoZmkX2iIyPxhKDp0AviHZlpq5jbwcFOdojCR0/mRC5/Nv7C9cWEj
76+8o0EBJ63m1gJrVQt3dYV+t2mFExjwYemA8pDMk4PLQE0RCzzO0MUr2k3hJTIkMy8d1svGXJWZ
X90CbeKvoEewkPitb/UxA5FiRcoUW0ZvUjw64mYlzF2aeXfr+jKVqLkr124lhGvRMdCrOmMcQsq6
FRVWaJAm7Aq+KkP6GZaUum5e6FuAmB6/v/cCLN+tN2KB67c6XSfarhlIsSQyLP1WaThN7W5h8QNi
vfdPPiNi/ZykbKZs4ts7nSIh+ksy3hlurpoUwxw+OsCpGZF0YpnHQllXlAczrR4GvibMGL22g3e/
qrjqD5NCtIpd5JhuPye/4vAi2Qj9qvmv4KHUeRWSDAvLqrM0VQcsXaYJ7fWGaH8hpA2yifCPlQ49
gk2OuptZpZM3cS8A4i0M4acJu3vQKTkMsyT95zwaylyY46YMgorhGrNapXHhaWxdFZK5+UX9JG4n
NGb5nBLpKelj2c9aC1tKvQiA7Uu48ZFN4eFzyxz75KxHoSiRUeKEhH6bt22HJ8DMAMK/ngF/4tY7
m6qUempmbcnXmPQGn7cd/Q+DrTfMl7ZBkwc3ZjfVg/YuD6LqFttm9JZAWq/3H74XJatC4duWAc7+
6hgr2ASEPyQ3lFss1xoa3brOWjypR3GGsrCND3YOm89xczpI0L+5orI7lrk992V6LLyPZTdEwMH8
pcgWyDFLpRKDHmoDJrPgKgY/Jpgj+Pc1CV5kGpLx7wfv9FEj1eMm9TLuWMRJEHAlg0BcIF3SoBCn
Z/wHRecmlnLpSs9Jk3Z9RhZnlEBVBHCo7/2+3F/FcDRrOXY7dMmfF4ehUCYSRJ07LSrYXHwjccGD
V859EtnyPlE0m0/Vi6L6KpnXwnlsP+VRbLp5vtowbmfV6L5NgWxexmvpzlBDBob9ZdkaY0CHpQBt
X++zxKB/Jv0Y2QqauKXPuYdJRCOkVsDU7mjuYJZjQH+Ck2SXYwHQYu8zThLbekfoLNF3MrqZB62C
+iYfkDAExBCScu2dNwz8iMfHPhCLmsJuruG8lH7QjT+TXRGgx+UDnvVpvLw3BFO5OlkxLdWuLdyw
9bbidy4pcr+L2QPJLhrBzBwXv+ksQzB+zz72LkAx8JfKJLNwFCuFw6beV2+De1DkkOpI1TIhol6y
8UlUQJvFpqZr0Gei6utR8K327SeO/H2AJ8qsSvIo8QRUYw1514WYU/sPqDahQqV6NLizzY1FLo5V
pNM9fN1Bcpy/wEnLYJ5nx/StnKettT2rjgwQBTC5HvVkHHILLPNDyLP1PfYE+UaLgMA81n1i1Jd+
4id09NU47kWNYq1CKAUVb/4qeuUHznTi9v7uKP+WlUQXImczLnAz7ByXHn1emHsFAAARASAQItK2
nO2t+UroyxTyMtRojiIhMxLDTrmpMtAEMzj8zQSan716Jf+rgFco7EmSE0TpsjXGxQw8uBwWoYhm
oPamXlQMNTeL+efZis6C9rxReqOFjrkMHZxvLqh8zwBWiM2jnJSByxMe8T14+YLKc7UQRZZ6YZhS
NjhMiQ3oAW6UZ8yepaJ9nP1+GcDNBmC2ehKDDwr2ogAhQfgIwqa4biR+TvUYiwSN/M7YGeusmi5s
zjbLxZ8xeITjdgHpZNCqCcPG0TtTivhYpppHba6n7DRbAX58Y0g9Yls3lpERJAQkKWSW6+Au35sc
1u1Up6aU3DJghEeDF3VoSMrytJHOOiiRAvTla3SYs1pVhOUxeUf+UObVCBsaTs+IaC6pThZDbqnY
1j89Jc9lHlxLwgUiuvdacvoXdcmvv4thX5YAPtHdu9gtBqhHshMEGqMbhxxlkDBsGy22KZEffeQi
4N2vHa/Ni3083M8vAtNibY6qXkjLXJ0+FcQyo8oX+MzGD3L0kAoGmJfuNJUlz/z+Lm7z60Ha2fg2
CcaEKyeIJOmbtRqZu7ahTSNt1bUKwSAFclmnNPlpGPI6de3kMMMjOdaw8E7mKSPf+//L1Vrt6QTV
xSwgvJr5Rk18JaQ1VBDep7ErcwrmlLgxXHv+t5mOw9fY56obqyMEVYjY3U80JhXouFVPZMePRIQt
nlQnUFSwxR5mJ4Xi+/Gm3xk6zhOsWnA5ik6sHsvEla+KsbStzDaeczjn+6u8Ep1OiJgCbjivkVcN
mfsoNBM8HD8iprXu/DcaMJb++LIkvFXMEZShjM6EzSXp5jxxAhkmm+dz9duhy4pqsOiMegCjU0X3
gvQjW2/f4raF1vcEMmPK21OEIol4UvOqzzh4QP0AoEXTTCshTM5PBWEXrOxX3WJSm5MH5MrZtupS
gGhtE8LfzMtwPZQQhBWgDPiqICqguwTaaXJKKCiKyjUuJJAkRkBjn0Grv18SNpouHM4tB8S+ZFWN
ua5a+pH7wDKaIlLVKo85phffZmW6BSDO7ZLjVfSj3u8buk7qMU+EhId+Q6FxEMCnPHfMvxP06yOB
y+Y51JPPO8KmjktEGH7O6A7EFDLz6t/mquI33YIV0hBx3/eUDn5tIQZdw0aqmrVF7Qtw23AC5l+c
jugkXO2wjP8mkTIeIzDVAB++dfzBiC89qDd1Ti8EiAroDgKXqa+PG9nwDpXSxog5BRrny30GvY3G
JnOjM6aZ+Tg4qKcGikIobbdG3TnWOSvRSdp/2u4Jbe2Jmn8NkJJb33Fg8tZI8PVtfnqqr7qEWnBO
akb/pdbVFxasvNxpsk3WbJnWC4G+VTY78p58aep2jKUEN0iJiQWFn9287BTyc8/7vmcozRc5e6Ha
Q9fJlra1pO9+NLtI4GHEcK7vdR8II++MjFp+VJaeJW2h6mjhb60I4YtuKwz0GJtJfBZooCfwD2SP
UndlQ4uhjRKudb+gEqMaW3s8IccCluJYf2FEhzJSkcVnNXLMCCF4rULPCQ936W71AF9Gb6wNY4Pi
asiN7VQOgCpESNIu3S6QY29pBCWf4Me0ehkKOchYi2Y4dVCpUP1FBGVhCF3w4tbFo5YWBd1RYoXu
EbyApZypmgYhawrVpmlw0sFlraQUSf4ktfn+j3Z2QIr8d0g7AkDnd7HBt2HrVGTmN8aqjz5RI25E
vFrRf/HSbvp+dWOPPLyBp4ZoG0IxJq+lHhne40Tresq6Q/eQVMMb6YcjKVN9G8jXpwrLnvDlH2Bm
xVG4aox4nQY6ge90iKHNkEvCyDLD18YcIqdPUGYwzWmXPX+mXI/W4C/EklFvaOsNsnXyPWFox+cS
03LANKmCv2BwxQftZVDst07XgIi1cHuX+DAn80f6S0k0OG7Q/dysIrvnKm5AOYJ8ezFagmXpkEIT
nDvV6NJSg+usDcoN60Q7tkRc+u+7T8olO65gV+PCprQsZHSbp5Pv826DqOyyLOIb128mbAyFCNKH
3dAfIG6DGUI5bCMfN7DRGJeIcdZJwm4WPoRVTXBS++lDih6pBoVCnGjSx40/TXbfxYN6pMKPbw/Y
uTZFwKJCAdj+qQM2QrAKbssdKvNRma0a5rgqM1h8umakmXfiMEGkwP0jqY5owyDNmr0RbD7HSNga
kNPFjl/rWlGyVAKT3rsZ1MENb0RnRDMoaca2IykYQZfVdztxd8z1dXZW/QUFOXgpZgUrqbT7J73H
txRyiGr73aPmTh7sk5Lds4kROqoET/FuM5+UooIsrptfGYeixT5nnD/tUMdBar/bLwJPA8Vfhidt
LfWZf3V4MOwrHHf3HU26pOMAEDZjYwW0Yx0rHlbDoJGiOdBP3+QeY9qLFo5O7BbRMGbtcELF8M8h
bLi50zCnaDpFPnaT9Sqb6mFBLvOQD3UMUtvZk1h2RJZppogESi0EDmJ3EJlGeD0QUZVMCKS7OB1A
tFcT53tn32+zLJ6BwkzqrVtjTL/m2mibX4Vh6l289uecRY/f3PioISnXi6OF5N6l48buPPIiKLr1
syPDlSeYYweP4NWC2T/BnuUhnoefz6ILLatW5hSr77zY+E5UiUDbCDayNDf68M7OXTjCcjCpVqn+
CcCNibJJvflITV+wng4RsUZ3Bna+YPUnoU6+mgk7qA7m8mN0CbkfghYxT1wm47YjyXA6pI0IdlnT
NHjit9W0W3BsVJWR+huWudU6xq+dfP9y4UHw+Yl4axfC6oj58KNlBIm/Uz7bxTACKs7wfO09uwZ1
tyHH5tDiMGZ42p+VAWbRj1dbvhePnyN+bTX1FzA6o7C7nSdzKGh1gpRdZyFbOzRdwRJKVzZRVa9p
mPrTzX+RbIEBUOhl37bHw0asOiA7ShQcIJkswq/w4doMt11/BcsqYxaqkCDi0CqRTszbij4UJw1g
K7KrhCGXP2L6rIFoVW5mGGQ/2F5jH3mvtFZ64gE3YPNpEn3FNbQ3Vnyvtw69EJlBex9vrV5ivxeF
AVZ+qA5xofmTOpKt7RROAUuZfu8zuotkd5e7TuQirbF4XKggszg8+4hhn0rfWnNtSWvipKxIikqP
qTTqMoOD+mqK5tOiDvhHlECLSZ/QxYcFB1af3IgbE98WMmQgmKKB2ZEZ2ah/DXQ5XayomRl2Q5Zw
LiWTvJUvoxTJ0pYkFdK48h5ObnMnEo4aym9sqDQwKmEIY+2rpAlAgJMnzEIEjlXapXh5ZBZCcxqV
i6A8aSKHvLE686ki7e/tClKK1nNT3b6igU2Owh9KCiIPQ/1djpDl8+GUFf3QK8MWbEkY1eAadPeK
iDFO+Na2Vezey74ewepsg74/pN/VMxIjvSkbxkE5x2nwyDIrOQEECC/IfaAxhFO9zpKisrukjis8
8ftX2S5HluPKftUA/uj831uKbt9nHBIzvUmUGafes7974mP316ZsxcRsxtF++La+vG1/x5dvfd4W
uSne+7gpQaFU36REuk17rvKuyEeHuIBOoChZjolmsGZXp9vuYD4pzvPpxlN4oIusGjgxt3ushUic
ZgF7lyMGK5x/lLBBqrSv67OronhZbnSrQVkrbgwH7bJYt/heSJsoQNztXpbLSK/t4zGlvxBXNJBV
ZWDmbnHF71gZT0ya7i8IurqG4Q8tRuo0R1h/2gtK7JOb6vRSBeRE8y+v/dkrx1Dehn1/CCXtySbX
dcT2MgYfe9DyfcALmu/3UmlRxlijWMIpXZEdwQxwtYZE/nz4FDDt3n4OEau4rgOOcea6oDpKjEuE
8ocKHx8HAioHSXZRumjkpgQARpqgqfi+EcDAtEfhc1g6lKPy6HR5jPWXUOCgXcLFQQiqZ8o3PWth
s7MdVxEp2WFffItcbOVKK37TD2vOX0GE8b2evLdOLXV9+mhWT00OAc0W/48cu504ft4cvwDkhgnf
KAvNPzhnvhwRUXq7ahjosV/S6MjR3KMXKWMONwgXr2tfRtOtKSojHcgV8GlToie5LqOSOjSN69is
AmAsTpSAsHPHFL7q/4ovE3F47utEUOXzjoo1Id/cshHZQl7YkctIAueKGTAWnXPHOc1650AfKxb+
KN0NUn1w8OfG4KVwxh5DNYgPikoX1WO44GiMl8hQLT1owL4DsF2EGX9/elXq5d7Fj7KyWuaq1jfz
k1rDLe4/zHJh28KR+qtlzzHTTIPyAJTymuLo94rOq18iYLnLzjyCskFc9QQbqypo7i0kPC9HHcHt
3SiyeV2VEaAuJddya7N2jQepsWJAiw2FsBcfewTP31v5ivqpMs8xan08EUSjdHn/Kf0meDROltCi
ScafjWF3+24k9kdb9yALOOA56RlYHWpQLkSvDU+WsHnZUc2SYWRSgFJS+1zbG17j2jglW8HUb8LA
s8XubySIXXIhunyGA8bDJGBICfgqF/PsC8y7Fmhc1uSltGZMdNDRSTRwP96NSrbYJ8I0A23xQda3
7/ivTx94MuEOhW95cv6tGGdZ7iazDjX2NM9IljXhJKnzs6TYEuucq+MrZJ+iZhej2gyDAwg08cQV
jxVZEAVI9in9RxP4zQlcYXSYZj66wVsZypuz46Cmv5T39swlGPh8cQeA5Lg7zBuF1Sk1rcAd8g6W
O85AwQMSiEGL/x8L6SZsdm2SQo7Hz+57Kqc5af34TKN9WSggmchwmXsJEwMmNYv3O2kqrWaxZWbH
7lDAV/9B1xk3/ZVHA7gk4j2IspHtjcls2VzzP3uSZ+gYMAQjflesFmhCJ0GkO7KpnVkRDAkWfDfS
2Koi5f+JajVyiGy+Km1Zj6UuEUKdNVnRg1WVS7/P0swp8m4OT9xf1fKPBGgnUI6pP8tn/1d19vaF
tzrz9d3qktRxRDr7N5rsM5A5wWzfp6gaHIGGMkACwes+T0pJxVnXNzqxXK8ztuH8gb8hwSYKZbD7
4jV809BVf7qKaD5ljjkJlAa2M75aIoLWvudx29S8IDSQX1BPncQva7bkNjm14i/3yDX6kZutmBU1
912bdyFyKThKhe/UNkcW9MtggXHjo0UipTElfj2k+2wRrZYrJ91yiYE8uJuO+uDj9hL6oQWf/Zx/
9/0wBRfW1TdIyt6y6+sRUJdPArPT7j1eD+wM1NRIdJlwlIWaiSA8QhpkXxaqLnXbYBcw4+TGsn2x
C+MVx68f42mksxtuehSsWLoFjeTYeu2aiBohGMvBPfcLMosSx+t4UCcEl15RyS5jIAJ0ALqD8DCG
HVyX28LRy6kH8YtDDrFJEMi7eIqJLt5SOUhY5GAV7xzkMQNMpp0B0jUKTHga8c7v2eE/EJJZFsCt
z91gomgHZBJW8CFmNIO1DVa+WB64hUsHP6SrwiUYO3f7jXb0ccfd+s5ifZmdVqMvulhUPQz1Xa0W
dd1lo5VL2ImRQb0gsONvasJV9xt5TkiOKoUKRKGwJKcQ2ZWq+cnBlpUg1f6loTy9JISlOswYjvZf
pUae5N91z93JpVySX+Jhhfo+SOUDkgBkDIR6f5cMLjuAmnWUwoWdTMhGMkfNHr28xBCMuk9VgeAg
GCM/VuiRIz08VYXcI+GJ1A8wGUKUVK3S6TcPz9TyjJYRqCsPzAuIPhCzBuTPyLLQ116sK0w3g6fP
w0+gNMg0xEq5zZ2QCsFrQzyasqiYK0m4wLTnzElaH+OOY6LM171rSnv/d7oOAJNQP2oIeMMzG4BO
IM5QSsKE6HcRtiTAz8Lz4GwsGstu04PaRLq7bjN/Tosa9Ewd5UlFxa0mePU69cNGeWWk0RClxXqJ
Jpxi2hnU1pcfiYy4ClA+dwd8Rx1qNChU0FaBgPxUGr7Vq1P7M1RwVy7yczVSnH+/2a3EmCp9+FjS
m3ls+JEISi5Et41XV5lM/Jykj7r5AARpWWqjlI7t9BCPL4lidxEbl127+8ojVnAE8/pG8Zv15OrX
StLnqBwK/vXQjlRNQ6QA1qoX1yvaXP3ikQ6VRfSxveQiRGluejGRcAmRrK7zEDXgY4w0CRhgSZE/
JHl2AizftafEXgRNjkdhiEUHIMlIK5Blpjf2DmxUoPSg+EWJPUCt63U4G0KQ2zySYu2V+1362/yS
7QSDZmDUepLCvDoIFeL+D8T00ZMmHAo8HBUf+sXrKN4e6Go6cUMq/cWEhYA1jyAybxsso1iri84W
oJOaVGi7/ElmbRs7Zo23Xfiw8O9p6fHsMWgEJMW0c3m20qus2Y6i9m6DILc6waNwal7HXmyXa/ZP
fjF6f525J6a0zbqKarrVW2jaCjtUAaG5CevFAVbaDdzyrR7Zhdmlm6dQTJshMYr/Qibgykmv8DPG
AB3FMn0VvPOqbKZ2P6g0ysFQXUzy3KOsfevQHs8IVIGENC1/PewbcqtnYerxUoX8QHU5oPe1WzMO
ZffF0alzGnLhtDz6Y9uoUzzsJBhtzaY21A5Gz5Dr2rrLvaSrHmRLD4qKzyfseyn5+DR4mjlc5QvM
c4GQd36lwo/RoXwPe4lWZQzRIdVhqh22Jbcs+Yx4Xw/cDRQjugvbgiSkWe8y6PJ2DT47446sZ6o4
8q2fLyC6pq3MM1vDy3eACKp96FJmpVd0RVCElgOgWQ19s/hxrfsmGrjMGtlfv6JbkAL5BZCXMNgH
C3GYCJXVQdQjepIsdZcKr9irymNa6ROyH74u0CJYFxH7kykRzeHyL13ilirnLR5uo/jZ4RNeMKGz
SEaNpy3Tu0ys535zbTp6tfgBTnq23Egw42CeL/NBMGNPurn15gWERT2apw9KkCuVX64fbegjL0hy
Bf4h7SP4aZeVB5D8vS2uxpBFVNyIccxz27hreDrQv2WRBy9bgFeaMNc4bQuGi+3/8wPTPKeDfnrm
nsENasDvbkMUSjHrMV6PGbZQZe0oYqbLMRkNbDjKNITxYxrQ9swnD243qt9R8BGgKeNs8wS3aKyc
lPoOG+pKlIJZDYaFvSqqpErfEO8SIfmo9DwZ6KjMG3E8dxF56cqqM1B/bsaQ2HXGGJVgIBH1pmWj
6U2ZBDPyM79SRjDObSoxm9RhZ66rVbXPY15cBcerPUIf5OzCvXNZoAWkhca9M+JPOCrwoR+Il0DN
bsYAbYs+KHw0vRcl1lM8nmjX1qytpb4/iWzbEyiRmeFsf2gFm6H8pnw/RPCYOD4xac/kVrFmJvSj
ldOHVKxxRg26tWd+QJOcPcG523W14BeL0MJUUrOnytvr6NVOxv4PYZvqi6JWVTy0GOEGCZQGWwKe
6kwWxg4ulUw0Xqu/n1G3MZ+7DNG9LQvxSxWYeOaHuiK9DXPqk4fY92zOcc23LCRxkCDq6bLYJ32M
OUWy+cn9e8SN7rajuAEzPOQrRBlToe0gXEmIkD9FsC44ZmlwhJfYLHRCJ8iyzctIlwjoUFlAC1ml
7VML6sxDe6Wn8p0IH1UZJ41ZjFtr35xYDH6FmLJcXz7c/D5BJVyc9HAGQzJJuinO+vuTq8ka9vO8
I07h1sdz9YHNkhSOF9WKvX9lyvP2PG6cfnbzJw0Q2ZnVms5LV8YpcQDnSvFxL+BAqSdFvjufzuPn
fZlZuU7pr1tQ1c4EMRE83LHPGpu7pHV3M/UAutExMIhhHrd1Z55RTSm/IzPIMQC/m2Sp0Uf+AP5b
nZIqgGRSQuDvmQSkcNMsRSJXumoknqZOELny0IhTKAmQHA4WkyvB6jfF4xXl/AzyeCaDs1RP62D9
GK/sYZ27fJOdapRfqXnOeAkUSaJMuH96plQFZbGAK9lUgzrdIEpW3FmhZN4lkzKtK7BG94r3aOZG
yz3Z/jpz4xKibDSYcGpIBK091odaPfDGplVu3WZC0EB0VNVSzIj2kVM4VbIte+41LC56FqLkjDx2
37a8P4egXP7dpFNuPz65PAIpkeB9BfEEgvZ2ZIUIWTVQr3M3geCm7saIKFLXwJgHacmFzrfq/OZb
YCn/zHCDnqy0GafAmDM+tJAS+ZxmwjImkom00k08VuooNc0Tuiu9LrRFxA3yRUO3ZhVKk5QZhhGQ
sJq+fGINyHG12lnE4Kq1wjU8F6ucOMuWLu11SMX+zebBQ1Agl72F+8Xi5cRrrKKTGDn97/tLY5Ih
pvIWNJlBwLRyI80opQCWaLo4NNl0vmyEDRRC0PoeJxoqh8HzUa3lkwkrgE1oEsUKzqad9Z1b7f5p
D6qwbfBPI7eEjuS7LnIOFAWHKmLnmPbufwXW/NWqB/VPt+MjITMHNKMY5JXhHrrF8ENUB8p0XhBm
U40QNw5g52/uMxK7nrEx3SqKMCX/N7lrGH1slYpcHgoNsJWWVJcOmVKhzCphNJlP9itujmwxkPuU
is/zJ8K7rYSwBZ3v9gSJESkA78kht5O5rr3Rp91/oEyUZM4ckLGxF6bUYPWtgukW4cXhfno6Aqxe
0XGZHIKqEsJXN8jxzs0Y+aG2cYSD2lvXIqyLwKxY76ZApOUht6f36uC2PBxQ42cIsXfLChjqX16N
QgJFdCreKv2Wr5MYyDh50HuTRgj7rqJHolmWzgnnsKcYY9fRwLUC9rOfQsP1sAj9SHHFJiJprgl9
q964jXcQezNFDl8klXkUfI8svjVfCDCRMlj5BRmqAAeP1VFf4OgOPsWWcqwEfRBh3YISqIyvnxGD
3naZAl5N+uTGD9xLtzAnqTstdvKPkX1gNWn+1TfVkywuRYTICAISHs1iNLMs6P2C7KvpZm8jHxzi
tytl0sc14ccobGZ3rUBmxi1o/MVJ5EL8CIqsRoaQI8E7x08Bf2RFI9aFbgf0eLTR6vHHDE7X0IoD
QiqiPHVN8Ps/JKYZymf0MoLIkk7SeEPJBaUE5dG/kFk3mbFml5fjs7m0fRs6bCTdCzffXR3tJ7Qu
gWiPicqVHcOsS949ll1OFEyDeJjYY7JiKz6nQY1+luWbJH8mHPBVAafn1r69MET0lpKHFu5g1CQM
hMProzcJVJFLbtU1anZFO4+uRlyOiCZlNPTpuvWn/vzJDYhUyZoGgc+lLXSXkoQd57k/ufiqt8Sa
U9tXZukmrZIi5SB/NeWF7qA9DI1ImY7Rv1jgMVnRkSBtZvXUCjI9yI7ONg780AmeqHogJF8pwYKs
2Gf+F3sqeqmMX68Fx9aC3vlxEfBkd8fXXsW15DDk1Z04TE2xgaWTa7upSG2FRT+rubHon+A3SXJZ
Rcu2l+J8tGYiJsaVEoy2qL6Ohm2WhWqlN+y9uyxElDedHhq2Jso1CoNr6cnEPkN1RizKff1LSMls
IxeVYsSI7rO2ElSFidWNbQAnm2HQX/XIVpMLVqVFnDUCO6mLOlG7fXevPr53+8LOPJpnR//3/ibN
WeE0IRuJh7XPuvSQii50F1/0CIU32PcdrEPn72GUxcB23KXqZifq+QCJrWH1J+eDc3m/d1NzmMwS
DeTvDVMWGgWbNvEscrO7vL8v8mQD7e96jvy+XwGgNNk20DnCHbZB5w3or8y++4WE98KhzRi3+dkZ
74mHrHngzxbVfdx2mrhJjdErvGOVCL8JxphFHw9zealUzxoLw0pw3SvuugX1F4jgXkjwkl/c3TzU
O1j0c6UngrdkwXe6mDUh00fyU8gw7aSHGP+tR/6yNoHhTtf9a1o8ThpPwr6BJLAgvVtNL09exrYj
eebKIy5xBADMXq2Q3Qcz+0ftmHnhOV163/DwLpxJFUW3qbwHe40uHJG7qs6U+DVDsjq2grDnUmuy
HS3fB3y33MzC/xjCT1ApFQX/XN3HlZk991N90lT4mCe2Tf3L8rpku0XDprDTazo1CTS0rC0Cw9/b
dNPxIzqqBTl0f+fj6ONTO63nyw5nT6fuk326ZviIE/MFU/BLWXeOmcosntRvfUGlIAnP/c1XawxW
Obgm3lpeOgSjfjp/F8KZl5S3UPX9sFtzV3QRDGojwHwc5opQ2AsKmiPTl7qrjunDWPzpbJzJ4Mo2
PLZyLdQm2fq63/MZGjfhnK6DOvAcz/XktzcoeGE6GyIe4shgIo2jY/LVsu8NvFWsDIejEKncK5IF
uu3jMZW0TlgevHRIOfs6Q1LZwZogHxuXGuE/mG+gZtFNFypDiIYJzkMCGi1YvgA9ThXvVZ6SL0/Z
jhKc/0U09xkYCovLHVlPJsMvnaHKv/vVVDz/cAZgc4uJ1WHvLNlHncJpZ58o1tGPxg7QmhtoX8RY
mbvzvFX6KkIrmR9UJT/D69LDuCnPpd1Inu2zJ8labeh2LQmyTW1pYTHPe7VCb9xsBIeoY+uI0AG5
X+QAoE0cs6CXq/WqeGWQdA4Jaf9LuLfgwPW3RL6slgU20Lc2Wq5ML9U8NaKAETww76VyhsDePGqc
CnDbchLpICxZq533VlQWX2/aJlPtBPbPpx+47D/CCR73UJCR3iNGR/UU9f0pfIGdrJ8bBQG28PWW
F9JlkMEi5nXBZn3MlkRV7l5QUMnJmueN/AV5GC/2AMTeAAgSOO3eEIV5rFnMlsLTVSNXq0r9bN8v
lvd50NSdN/o8y9jXg0KodiH115vTvlgPGPqD7hdXAlc5sW9E74tc7XEbUbxUBLGl2+E1ENOuuG7f
wycSbx0O2A83aatNO4OcTpqLftKV4oqwUwF1VpN2oB5ICs3Nn6hZDncPq5X46/mkL65teDiNyo78
xxurk6sj4/O3NHEqtSmJ0vOnamSmI9/lXWJ2x1qCWUxsbxn9Ko87Wlj4G8mQ6mjHL8QDOdSSDLfE
Wpp8DLFEEk3bGw9twDhgio3fyo3BjYThu1A606/0pt2pOx00W0DZhJUisYYG9CVtwP6gJ3/p+iNp
pIF/y2hkn4Br50RDgBdFgZxWW8eyMTbjR2wR7urQdFwtU0zdRONs59v/unEflVgCQ7lUwywTBrLm
EjYinEQZlQG6agRmrB7ttJtNgNGvyOvN9AOvKDpTSmXGtH8kK4bpsQK+s7rToqLwGFIJ+gichiEm
1hIb7+yDObehRn/MLJmp/9DC8tGOwL2ZgJ4snvR0xKBY9/kEMfd3qHstVjDioblz3ei16b9NARNq
1iXSIl7/N66qd1Jax9hOswV7Fdm5yu/vIDi3+1QkD49Z0dB36emluHDxzrZBnAKehaGKK7XEwTvL
0YJ3/XVnZVWz6mEMcN3x532IJSMrKyvvEKr/hXEN0Lu+GZLAoE62kEVBiZRfZkZcKRIpbLo8YzHD
xHv7NZ4c+UTH9rDjH5tSzZtoar5PbDf11gxzGy0IrkLIdxAy1a32g7rbZM1fBs3F5naFXEfADAwJ
GyiQTU5MjHIGKHYuYl87zry+q+B8jSp6jHTecATsFPvH5zJBkrdvqdPu+3a9EQRc+xDHuzx+jyXl
FgDIYPmRXljLH+jYVal9mNjI/gPTp9tvBKAei1hnaYtSsZCLrrr/l1WU5LEuHL2dAyT8VeOHi/58
rq3aSr4UXA9CmJ1+tEjMQW5JbMCsJDmesMrVo9fqXbvV3INWnmPKc2J0vOxHlX7cSaGLzFmwJMK8
99p9FnC2sTSCuoMSC94IGfhp4NJCOc8VWMVXUfvZq9mBZ1pge5OmNSco6dlAaWBJe+fD7xJf571p
ymXMSGkcT+0MXUvQUdQLzAf05/CisXnZg0Cd3hrU6fODK8zx/6GMnjfF+LNHpgrH03ZoFQ8iuyd/
8VfBRKFuJ6MIcpLESzSuf1x/JdH43MjL7B1C4jmjnvDmvsrZVXA1kBq2D8LU5NBLm79xp81UGxgY
W/1/kwcsp8ZGjjbBtahkX7hiMO9BNoEM0gRQXhrvgsIzYpVrg0KYw4XlNpzaEbZA0nmFgDAHc/9y
7njrPhgIsWjcXbJB1URu5W5b2pLoS7+iIP3mZ7dQq6x1nibyjXkwbLeYskE9oT/eamyiRtTc/I0t
bGU3PRIwS0gPmLBTeZlmFAFIdH4ytbsihiEA1BBY15iMnKswy9ZsYuK/flYx5xjKPaSlHmtXFGHU
COx8CULHiv+LjCH1bjEGZCpVZg5Y0Ie5Rm0jRGWhBnFwShAU+JP4qTBxus0s0JtUWhEttlZEitld
vYg9inEnXZ9i1M+BcwE/m8H5dCBDHWo0FJR3VIL672Pq1doMpoYALrneWpWP2HFrN1wZRS9eD4wa
9oiQ5cjxjWWXgtQSKr2UYvOAhISL5iMCRxPDrB6CsFypToTR0dgx0Yz2+y1P37flb9lwWHNCh6Dp
SILlgFEgdMtyxyH3Wf7QjGiVT399Mx1Kht9dc4/5UViVBOqcBihsxEumFDNGMLctcBj8qE6PM2px
obPwy2vbbTTKs+6ApAxmVhIEEt8r7xG74bEsjmP0/2V32sbY4GdhnxDuea6xFWjwToh28N0VgUa2
aU5SLtdF/5rlkTdlYoox5gM8ARPPf8mDbs8QLPG+9c37EkZgLeXRo6HjD4D4ImHHQHTH798osY7x
byvc84UKyzCllQYQOVZKZ2A2IVecX+NhUQBVn6u3oD3kajSRHzp+hqagRolZYOhWCcc6a63JdWvB
mjEYANiyerUxajtA9jyHvL32dLpDy9UxFKKxyuzKR3raKWV5KHeXTFA+tblPuJppsMR4btBVgR+F
K0JMz5yEuHu5MHyYBYFcsGDVZRhUTiPqtSPFovrczrwsYwXGcIQmbsX4EKwtnY+gbOpTfVUMi1P6
DOKB3PjZFNA+TJiwc/+dwDYJfL5JRJeFJUL75e27TLViaBd7E9z6pMmPq5NJSH/COjOJ6quzWxmv
lIcRIFa5pRNAP6vjPOrPk0jAgIq8x0Jy44/GhlP83SJ6NiM/DVzIjqIaChs3ELKaCSRN5tqVjPaB
OS8O5aRKVhuPAGb0L/NvvDHKKWu2q+g9RfeZJxw5OBXSMwc0SwTPuJcctnTPht5ddNlr8mK42fXc
HmeDDelpsj2Rcb5bu8mvKxMdLq5UEg+z6fP07Wb4ywIU4Z8vU40d1WmWHUDRoid9W1Ydtt/sIi8r
6gnNL+c9qJ5EslTt9E0NlB/X26Dj04l74avpXG3StK+n6N/ARCowfY4muREn3CgeE/ado57x08PR
usy66ibL7yeM2atNAVBeYuFUBY0qejWjT3C/n2nXNoUyR2vhQ5sAy7XaxITb3FdkYbPJan/rJt8y
ZA9ora9iA2+uEAvBJeK6/uDcw3/CeZqbU+N8JobppDBjPWvsHy5Jd/50BPwFFXyxygCQAv9E4dRn
Iv+kJzDUFVWdQdzMSx6HW6PRcbpN4OaRZoKoGYMlE8ANV1inFZ4xFOFkrUFSAP+ot8LawhRLw7YY
m2DZldcTEgyY1AKCND6FDoPrIAjNnnmEPcA2lm8+WKW/6nejtLw9bktkY0QsQZa5Nomc0jXchsCu
xZnVznRzUZjAPvjHnWkWbBNvSqICZfAHWVvY6fKAEvnt4pEqeniGrWgntmQ0OLbZoTgpz0fGGYkW
7QKgyH17O4BKnd5ppZzLTH72Zu2OXrHKGDLj/9FuYOAieoRDltlzn6PBj/n+QQqCXLv8BFaLzmE7
/8J8CIDo2WxTwwBM4eyoSbnOaJD6IvZEfDuNPdWZMqy24LqbkuYgrkzmwKTSOU2C8wEX3+sLgsrv
0E/7mxTrUvBjn//dytmr2cMQTj4UJi5Lg1lwGcR/lWuhomweuGeIajOg404mDBwgc+2zB7EuKZcG
B9B0pGq8wCKMrGZPWi3c1RiOt4KyeQ2bb6q62an6+fn9NAflOAkUGKBYPiL6ZJqrqpeZE2jYhYJ3
mzz4TxMDjNHVDgfbwsADGRavcIoThOjX0ey/Rc1ABW2o2M236LiuqPKx2Dj96woIwFRNCbzxVoJ8
LZnSP56jQ05VloXX4i32xwa7l1RCNMRIfFr7nl5Zl8+XtJfVBY+cNznAgyqbn96SgD0SY+YKSWM9
9h9yA59i0IMXGwDM0NjomOEV8EPw31RiSRweE/EmHzcx5BErT+u11CctDdj5H7uaqOZeiRVwF90W
Z3QdOug9ogpArHLC1CHius//EcjLM5wC0Q2A4AnhiESLXlsTCgV5EQrnQvtTw4JL1SJIIxDEbumZ
JB1w1o4YifIS9NwukHT/u91H2B1PgKAgI43LxMSgzfQmGtcGFNTLyhLaCWORty2jKDwRcra0FNS6
sxD/ksV/dyX0KvmlCafEz3R6qxEh1Gl12alv9T2riVvoVdHs+JeKHAw0tZxoV5xBxtiN8sR+RWSs
a3Irmn+GeEGmJvl/uuHypbCh5plVn+OThFstDbt9I53mGtCJ121CLRlZt7NtZaXq5TAyu5YIfNM/
cuXPXoxrM0Z8TbJH5BJSsdODrcBuvu8a70hKtcj6TIrE6MvSyM36EPxsvJiTqltYgrSEPlbqVF2O
+ux7hlKFRQpCLmoEFH4ufyhI7U1uRm5kRnmQ0TczvhHBhyb+CdHcOOIEEOb1WkyzcAKQZNTqkMd6
COZ4ikqZMGMUdQvOGp6yg5QTTRYG9x24bQ1W9UE1nTSCWkxt5tayi5WLj6OoiV5HwN8qlAnTImud
gE7C1gsE6nXbLZp2o6SlUHGxwCSG3rsz5fKMwhUiyaCojQz4LgMNpkU9Ig0uFgZijMsWAHN4/T9A
GDiiqgJCibGoawm2Ked8YMRDl0ZJcRBEyMSXrrrPF6NZ9o+dNhwrkzrUpzVEYfcZmVbUGj9K3QVV
oAFYd9oFOkElSLPtiFgl9edj4kKuHojOYynA+cctRJAiwRKySYVZAYbyR2qeSZVItWjeveIjZgWJ
RiClVP23klZNMUGLNKCz8+ZBu7vzePIdHjHsvl8Cs3JbR2xBADeOlOQO+D5uBe1IoX9lrtFlD6q/
2vndMYRueGftZjsbhVPJM5mzEUg3Vag83oguNab1c93OVbFkD/eMiWh1vmxcSdK1sfMc7kkQ+8Dd
uHFsHDslyHcZkLqTVbycOjneLOO/XfWiea/GYjmjuJX6DKDEmYBVbUZS13z7iPJNV5mJXWlRb8Xt
LVWdSa7zxZWQCtdeok1x456mLo6+jAXjPKWceJbKjcMtiAO4n8gUN3Ef1JaoesViISVY24NqDec0
01zVjSX5EK6DIKuApP5+EW2f3qOVYVFNQkRCJcyTOchtl7g0msJKaOKIi8X/cOnXjRB6KbAhAAlh
UMWIPyDX/+lJANBoXwBhxsanKRDqkNtLG7lywuSWCgq+N/Rzum0l078tioBM9oGg4/9x9PAmk3iX
m2uvrGiVikDSrPpu3XGORRZS7MzsyQVg7zN5/NYl0nZpA4Uik+3lIKt+B5J5Cr0Lr0TE/zI0c0Xd
n8tdbj7E6eEOu781+Aau8uoRIq4pEc9hj2wKD5o7xTySgnY3YGsaY0CQoK9rU4SFAoZygSTFYGrQ
nSXZwmIFbEzICHPj4+3w23Ef3oRVKDul+4AVsROpOye4E0WoZ23kFAENCdhNceWxmbXBQtgY2dXr
7IrfrXlMOvR1PoTBGIb0VGGw/cknkElp2xgTidp8cDD/312a0mLp4g8+QGYhtLZVWlmglntIuRjm
DK4NKIkVjmksori3ymcjvvgM5Zc+ps/e5pTsS08ib19kh/rqnKG6tUBPcKg9R3tRyUTW5lOmPY2w
d5Sn2X2udW5kkh7Spt+7P7lAP/yCoU5gCV4XSejnOZJGvEomnD8KF4iDiGEbpJLe8BaqIZP2gvUL
gOpe+vQp8O7CVkUuBADeo7I9xzIgPfwkk6+Z5V8mcJOlfMvihqyHFJwof9PsrkMUAVK+pU8nPHcy
PUnnrUwgqCAVB84ZUy/sIubZvqTN6neMbI4l+6KSvhsGPBqn7STUOLnMRdEwJMQLsL+HTYqVVsL5
HWhqGJfCx+B+rLy9nTd+RcqgvHu7Ac5OKQBjmp2qdVGJZ+jScaH7Qu65Cvc0sMrhJ7HIBVzzUn4f
3lugS2SUiUxrCWjyqcVcvyUYveU9k9W9XL9QveqfDzTEPvsq1OwEXzD9bPUodrBvmOCnz0OX9Kup
pbmP31n7WR9YyNPy5LxHT9UrdJHda8v0JJf0wp7h27OPPPMsujNZMd7DRL+6Ha9QG5KLHy3IzAxY
k6RWlXHUDtb+uIV3YhE+kmWKbVwsb32S+pBFBusZ0pYESoEnWOjTV8duW9sNFeKmR9xP8u2XUxev
yLQdmPhe0msgllA7PStg6iKHzShqUT8qKp46pqD9k2qkI1FEmzo/OEdQacKB/V/DnIZcwk4EPEOo
K70zM7Z+SX7t38sr8PFTCLkJIFTCGzAyMmHCw9xEqqH0r4bAVGIV6MtOdhaSfxE7S04YBqnFEc74
qKB0EbOwyKapqsvy13LPJwooPbQH3iOxVyvTRnj5K3IgXlQht7QJs4ViOVvubLwzuZc3lzzC/OP5
4gD2UM2nA931HMfrt3FR/1+3Ifu6iB0Ld01xiimy+a3eEJFeQv8eeMyAE70EI2t/SJcyAojuP9nS
Zyh6QcKRxY5+ts2BYiRplnSFHSX2u0igSocWlzib5xVgCWPGf3dGRG7QqepASMghyvafyh3Qqi4h
kjHlEuDBFpAL3ZYZUtafOY1g1itVE9KJGKXR2U3Pud6wcnyorA/UsTAJAyV4Isybze3stLMqWEZk
+uXQd+kXeTQZlVWroia/D0JZdVgNSfSCA+uRZQHiVH3Dk9gQOR935cN4GeLeniPiC3a3Si6GkSf7
0agU1WIn2HV9j5chB1MYxgzB80cF3lXWvKdZvNtZE9IEIt6V3spAS5GTbcZd2Tr4RvNWcyhfAhA1
ozX7U4WQf8qkdDSz4A+RdZ+qO1mSC9OYd6w/MKp1lCZhMJ6nfP2nzkfMTO/LV+o3fZQeiqSdsUiV
2Suisje6obdKh3tVN3QCcYdafHcE+MmUmdvjE1hhE2mp4K8IRQSv2yNV6n2vmTs2xjrWm2G/+nJ+
rhwlaSVDPKu0wkhTu3/XLX8OV9zPYqK7+7VvOxCe+mC5t6h0kRs6QkPQ/8PWdE9c2lykLRlFcVoa
aa1HfP2/7zXDUuP1XUmZ3lZi7bTQcPa5xqnF9wQ3fcWJBe58FtUxfVnt0hG9mZWFbc0W162MadMF
yxlguylM3WXS+ct+/AtNps8PuBondHkuMZjGVKQ5rzpbDgCVU5ikURnrJUjZrWme3KhC/w1HrOJn
yPwNUW2mLzfRJZwWWnVCJG5HRpDDsCEUSX6cVj5Eejw6oJgHb7CU1XtKCaLyQZTF0mkQCbz7Lqp6
aNrS9IVlbCkiGy8OAW/3N7vlO5r8OmH/AsJBSiHqhzI3kQqpEwa/qJ/N6E3uA2YWmD314h9M4giG
WlJ8e54OdTRiFyE2YePE6kcLapEBVRhrEcdz6zUAN9fym0BFCJT6PAtREOFYp88GX2sS0CsURiBj
+YyVPFSfGwFMvoxrnCbHEjvg0P7TvL5gJgSPfo8LGwtcAm8DAiXJKK+AnhKsI1UbRwVmU0EaXjBR
56O0k+i2NBNYTz1dgUNtNuYgplxpz2KiXM0c8S42k3L79WkYipHG2mBYUUBSkDvnWBTvCM9rszyY
YxCsZMiLaz8Qcv4lEDR8+8w0JsKKIcG/b13vFset87a6lRBiqaiO5G7PTN/NZ+/WIEB3romDxBQh
85jt+PSKid7j57L32OXWAGARsjFqVscHgGIg8vblG8RsyDt+1PptXLzYH5LROKaMGg2Pfvze8Ugv
cUlVbtdGErTpyNj/rkUOma1zV+gytb0oAB1/ApN5+FiXXEPtY05CShlFpVUUWpimdzEg+fKj2dpT
xpEHLQmChHJXL/s0GUmzcwKnnenIoiMQxidEXt0EWod6h6ut2dpKey1PuUOJ1HRFRseoMcswaSjJ
AIY5uOjIF2LTGf+RhP/5uv9f4MlGemdzjBwHEY+Kzv3oQWOOIb8PKNXiDJBE+U9pp8Wj4VG29UMq
hHg7VbsOQyg4kFPlRld1aM915oEeCz33ssGHapu/QBADNU4kb1m6dC6hWB2qosaF8zxo6y1KdGK7
CJ+yi35mijpp2r0pVimHMBtA7wQXFaX9DYZ+WqHbrlnK+E3yooPLCkdbx7lANYa4tffnnGrJU9b6
y0kianWs2ErzGNmyoI/IxNU9jXLRBqNEh1vH+4jCOCIQZp5cLvf5A8+CWN4zRoFTrlB96tPps7z1
Oe4pC7SpitKl8D58qTEKt9jFXtGp9vB+uAssalRUn3jMum8JeuuV1SCx7tzW1TXzUb+6rhRVigl9
X7EFGxgwikEYPaj4Aw5i6BR65W9+/jJwWHmHAAJEuNOFWzZ7PBDZd3UXt75HTpMbNLAvezzEmnhe
cBEKK/1Wf/cr5a3YfLAhog1sQR/0wkx8tBsKubODbkXsqoCWGREa8IDaRqHyERXbD6oPmz4MyAF0
LpVEJfk3Y8uvwH74sT6mpkIeb4RhNZfC8XstOojW/eaO0C/LfHtn4ttA8sxYKpbr1jXULu5VN3ac
fyTDpNqTn8MmKUZUICUmWSUEFgoe7ckdzlcFlJPR7U1qdVnJaWua+jUIU1h8vtQ42ss02R5MoncN
aV38g5SblKuZSI/e6YzRICSDLNyDrapt+h2XGjbv7yQYdQFNv5q+szgXlxMH5N+lhdO8e+SWYASR
xbcg9rT4+LoEtJ1fW9UzD49i9dZ6KQJe1XeeQzwL2NS6F4B16jGe8P+xJlhERcTrweZw4T+LOwCl
yoCK3TDnzWq8RiAyaJwRdpXiI6qLuCvqaXwibwnkjaoMLNMbskpyRgy1uqcTdYq9sV5g6L1bV7mQ
b+/cmA3siPaDV5lkJN6o/u6PDB+GFE5ieSvc2534g9I0VXxuo8xAu/UHqe1Laob0XJO2Q+dMfKQm
CZeGDgG7dHTwPmmId6xi0GfID3Zvyu064p/ZEp8OQhUFJzpY/PuDe0qYcgs5MrZF/p43vMtqMz/P
CK0+VqNqpyAU90nLTkBHEWIYfRdgOpRLmLj3fNX3uZedyD0MIsBCFhFIVuDyYYw5rl9akcHXlpPZ
xibm8xZtMhfoyhh0Et2YcDB2axN1Q5BEucB2WB6xKH7zEp7pftkSF3w00kwos3Uz4iVunyK3PF8Y
F1LDXa4Nz16PFnUgAaFz6esUDHEX0USEKnnykVEZqUJsRyhd5v5QdFXNDG1+S1NdRGVvtF0zeCmI
/S+WvX9YQY8WrjIlLBwQNZ0mHZ0gXlHCWQBRmSbtcLij8oVrSIkEv0JMfnqP++dKtjgAW/9ogvRe
DE8R3Nm1X9oDciPSmbMbve5m2Kuc2XMeMI7ezBnIz+0lV+wvdOYVUFTZg8OP4grMEWTXvn0pRM0B
uSuXrT1oWLPtnwtfeBrP1ny06W3NbykrMp9IJsQ3aXTQGJ0gH+tTJu8KzgWljZ3yJ0BfDQg/cX34
S3pP0Y8Dbnf4YD4vnIkFGvypiExbBR7aBhLP0nQKwLKVVKL+DUszgh70u5L+Y9AHNcrMuz+4fAU0
ttYmI95uEEN9h8kjD9MxvmUzuTdXIrddzsWIZELmfELhEQjT6nEhALbDX0je0jIEQm7q4Ge/Ayc0
fjI9cwp/OnIWogg9u29lNw23S5+Gsbf7GAHLJfCySkoLA/uVCgQ5obUMVHgcDb6Gkh6Rftol4HxP
k6UwlmrmhMhKCitBPNloj4vfVGwxOGpS0Jnna2wWZRDi645wamg9Qlr7g92vxw+R3VsNVy+SIqM0
Y1txLjHK8I90g16rEQkanlsyshxlhIx4XdJhBZ3/SmA4NI4VGQZZnsBEsYCWEMvUyY+iqEpsum/8
wiZOiqrp+cbA8OqxIcXRbX7lVf1AEQyw46HO62Thg7Nha5K1vRhi30JnB+FNxZRBpvo/jAmjGT60
lfMo36uGkD+OED+QIro/sJUaRT8tNE7T8dJ+IgfpMd2mKu3B3uZ5bQyH45s4m62rvnQ7IUuJT0tl
iYlJYee6qwA1dniXtNcBnjMuPQqHLMZ0rA4ncJsKFxq/N+RtQ3ce0fNKMM27UPcV7+j6rLSnghIj
M3aM8N/0MfJaGmDCIs3HwQezMd0kdPa0/zkfWaxx70p2u16bagiu8TyCX+OsfHGfShPG1gU/o0y7
vmKBnuKa5eVfN1St2Z+zIWzqaBaJ2kutrwJjsm6XoGTkUyeYr08cfvho2qDYPAQWWkqlrcr67k8r
rgg+r5AOCOAZAaoOh7EfiDyPeL15qDHcZ+sqze8738Hxn3/YlxfjRFK6vjKUbbNPqGA1qD4FPrNW
vtD/8MA47lxxeWy+pSKAVr8Ir+eMTKN3y4RY12B0RNUbiXLAxrvjJZzS+wMHeBLZIyZKjscTgdb6
KTFMNrdyvcxV1e+U1k+lnHGJlUuOs8IV7p44d1QsuxADWAwLzU+gvA9gE4KHZG4V7M2E7jBgCmNl
NaT+iCYh4o/xRgYuoY6SCjeLpgy1j+1VWGM0qlagwjdBitA/jO2Vn9DExaWNjZ9872rslyUu3T/Y
out145eNHR7DbmeXxNrUzVmue3dZx4wpGd3KZqq4HyIhLKKueOqfBo5v4FI7CzmXFbO03CFW4gV7
etvdw2loKQ5F4DyyfGT590+rEygHV9Ghrurmy7Xb+jvyHpH88R+QoAxQo28P9XaMcXZspowO1uPx
4Rd2R8ZYON++AhPCNeOPwISjAtH0fetI80G1EWWS7ANBr8ngLqlR2E0CG0UrKQxN6S9ZQrmdK0Hm
eFfK8UUeg8ilXELkEbEeKxBu6kd/zFsD6WfSr4jpARSAvHNKVtFqZY2xHByA36Xy4M8ADmgwOPsA
zgD5np75fHvdSaiD4ItwP0wtEpYoyxzeOsI6w6QCmNAVAkAhNduGFFkI1Szl2BQFd87xV2ta1B6p
m/Ei1PKGnV7jjImsqtd+SP3rzDPM1+b5IZpqrwlw7cubetCqN6FIvy2l5r9f252atZhp2SH0lj/p
Aq4sGJSwVD9TyCTKTHOhynOhLqKoQ91BSRCMisp5Jf/v0z0n1Qk30TYc57A1TkAFbBHYCKqEw/ft
MYQ0x1f893V5s9CPujy8TWvkawt04zqz2SPHjiS+XEJFgrz+bAqPH4OXF0QSKeGz75v50Njrxnk2
+lPfdHELZYBCQ5NrSqU/7jE13ZH5aM0uFcoC4q2+nT70isTrWL0vwjSJs/Hqmvkgfg/kMsLS4XZ5
oBWLVTTf1h4zqL/08jl2ytAy0ozEHKfkPv0cveF651L/AP14lpLOUSusShzPIxR5K+EJCW+RLgL8
H13MrQ5e3gN6RkyoqgSI2LGh+sz4dGh9D7Gx/WVdupkQbJrqSGW99tmmfIux+4fDaLxCQ4pd/TeR
l+Z8hTMCrKgw6huNsiSsOsnimk+fZ9OikO4Q21c5EDGzYFT/l2rW+CmqwIWK7sOFGswFPNcGnCbc
lHyxwU14j8pZR4+bUCYktpmaH5W07KFR15oYn/kdLHPkcjqYJTnYewsFFPby6smDLbsiYhkhQ8vl
rjEF2HLnR2GKHYacThdUI0/a/jbOqfDNcaZl+kcMyVZFciIETA9douQsZlXNrDYP0FIxIut86dcZ
UODxxxtZKoc5RHVfsO2vg+Xczph/hxeGRPgj1iRGu3YqjZRuAAilQMXMiL8fdlLdXDoSX5YkGe1p
gtFizi3j0DPboGMcFb6y5SKv214MtxsmDdXmhAD0vEc2p6M3SI/bP5v4A7nZN6w7+3UwBPFjThRI
+uAbp/Ccd0CBiF1JDk9xuNvcWeA+K7FgqLPIOards4sWas7kilvydyaIiyU9JOEj1QYZn3JZ4egX
7A4jPZ1b/c3y896LtXlF73jXWxQ5RBrOU4AeKo5JrNDvcpbpdmrEOcYkoFQedOJzJy4sfQRbZRZI
Ll9LqE2td9+4kXPCEjuI6pDfbM8tmYlQo8uriEbxjn5bqZsyJzSRryuYBfUSKaGMeyJ4EkRvs6Wj
4xfEBPEHgHotdl1NvBJT4T4mBYFLm8SaGI2VipCyEjp5NUiCa3fxmi8v+f59EWYLhNWjuoBWo01o
KOS4ghGh341+e2V6zrx/LzELVjBZoak/Niky9bSoHVk0EO4TGu34nHGGp+pLxpO5OCi4dPuSroRX
gSgFu2JUXTapVIA7V8PGHFeaA/KsNje4GtlwesWaA6liY4VGogxW/xQtb7zyAmYGAeCA7GcnNZ8c
j+Dv9M+E9eE9v1UeiEh7U78JQ+WPpioEa82SfpNKUSjtkbl40sQBbRuqgx14XfEUzqvaxRrxHWOZ
XuP2a6gjWemarjZf3PWRCo5PBIlAlWaIrTMjSfzzbrlBGahwMUAw4W6w0YqIgj72eE8BnKGdZrGF
AZ5yWPMfDTvFFpJnDd+PPB6XjbtwR/JZ8JAngJx6reh+99N6qxOHok0HVAnh9GWOnLrQHEPTSx8b
7rj/nRz7MQf23Aogc+mHli/fOrFr96SK5pNUO8YYJePblmP4e+QAFbNI9vWp29dkq8tZaXmW5HgK
eRF6kyw5jZBD40cEs6qSPOYH+BmKCwcZ7kFRfkqzqeTLV6jUmvdZluZwxu2CEYr4g3XBGqbo36oB
xu+MKVRXZ3GbIK2EP1LP1cEuwoUunz4rQ2ydkXrT/ENCgo4N4Vbl9zx8VMPa/ntBOBl9ahieyzvy
+5s5F1XdRxwlLrZwYuUZ9G0yj0MoWauJJCCGNoUJITsnP8DAR5AXffRmebkY+j518EcCc+hgOb7w
cu8Tdsc/LijRT2J9QeH+9hbpYTzTz+9ThkwClSd4kBCT8UKveT4GsNY/It876jZZ8hq0cmmaijKR
gGXklPmm/s+LLfWztqtFxR3YQP4cRYtsh6W7W81gmbsg98NnAjEOyy3E2RI/Q1h5gvp6t7uNp/Yw
vW1AcNCCrXKF+ztKDkEP/N5132vpetaUCBkXOOtfPLY4D2oDLwW7AKz9qM0a3O71FgMYG+q6LSlL
RlWvFCIJ58fwIXJUwHq6pxNrhqJEWG37gOK6k8z6+6rzZ8CeCEs1RoeG8dyFOXLh/TVUgV+qFawK
Y5k5Y+w2qL0bO057enLL1Bvgi0J3VSYOPm+50MsYBvaCW9jw0NipTRb+k+Grj/Vi7vhMtZGwGO7n
EA6U+jvBVwwuOSviv6i+w5sdkUQFhbAjBTD0IhPFvOIzrLRDEsIVa2Tq2PRoKlNJuV+DQIvN6uB1
3j2dC2XazQmcax7nBbZORlP6CiCOO+2eaI+sRKneGJ+2yKvJCc0PcuBPZaKchBHk0w6qkxcZADi8
PmPvlR2LJ97OEGN9v8mUzK7RTWPhPyIhnUNjUMRJ4gEgY1xz6sCbeZg/Gx+EAm09WQs+9vISnH7U
J26ZDcM90m0sHUvjwOPBsMeDHX+8tfp+CQNT2F+hzYUxUAxvMYWvqAMgS5OQc9NfFtppqHwcAtae
/R+FGx35LMnEw4FN9GbQG2rkTakHUdOz617+kXRxQm9O5Kk6oszU1GpCnB0jlIkDgwjP+Ga+mmxb
ujJNiudl0Riko74Fj+ubF9jsUv6sfN21koErGLqfQcjHNyaIwYve8YO7CeSYK/NXMMSthLSkHm9T
JXXtQuBU2Xfan1MVFXJnQsrakCUFKEFv++OU0GcIV2vwGzQXAGbirJPfPGX6relkd1pDKX+BobE+
TznNCbcSZrY+pemO77MXNqYGz/C8x+Ccy0QZ5EuNW5x6B+2+rfQR4HsYdK4c1LOoxXRGngwhm0F2
sRWfuq6CpJNMuOhHaxOIG9yfatKki6lN8Wct6y2e01nxufwAh+lyGUEOTTOIeRjvJzQ5cGjZFbVt
pRMCHJ40XueeotYyq4FbFOY6l0Eks+MolQ8SRr1cFLU0Et4nkvQ3Eer7G16b9DijWGX9LZLCS/eh
edfb4EdNhvQ5GrrImpICA5WxyWkP6+XIfPeq+cxmLLKec3Y62si+KPyKEfIeZh39Y2SDKQGm4xuL
wlnnmH82fvQNf9qE/CYKk8k1YwsjoqB1JA0y2YjtgUtBO3mGnwQw1aDCksnWOLWtktoafA3TD62v
u7JSPoRwg7kKe7do+4WqzufsuFPcm0gnb8Z19ZeEMGx+fwVVy9FGyvtStAzI86bM/6YZFuPgb1+Z
KuEwcThwax+4cx3dkPglyJPIWU0fIq/33u/V1spaOnKJmCwlWk5xFZLCuVp3yeMHljl+qUgQ0nih
QifsbVDqInkskp9evHOzkacksvtXfK8QZyb/qYjPANw/L/piFgWWSII0SWZtKENWusZ5XiZpElWS
cL2wPTf/LfV1xByAuSCYrh9r4tdPXo/YjB3liQaHoUqj8XhQscVXikpAfIiL1Xmv60nnRxPoOzGH
YOOEsj/9ZGzlJIlUEcvtX2BVPHbNGjAPSisgerjHS+OYaoT9/0U1WyeuXbK46/QK6wKxQw7iMGZL
vVHhPrweFfI/gkWJYfcEhep7tU+ubnRUah7Yde0wypqK4SzjH1DQ+65oG+oBdy3AoCYDAUUTpEF7
nzmBmA4xiiu+xvJK0vmEvQP4T7bAFeGGvav3SHowwmNcEQrU/tHC06BugRmEkYZQafLsD4b6XhkL
NBGUsPTySD9MDijoHa15DL8COCr7kBB7Z2tvn0qoIhqhHjG2vLFpzub7TAo4l1CcdMW9UuGJHpp8
yO79W5ZPfAGpPdoX0GkQZlyqaRR8wv0VN1cJTmvtY6bXkO1vmHBEO0ZNOSRH5Gmgh6bLjLolxr6u
G7TG29S6hQqhot08d3FInaFP9r9ppuTMj8mgFQjKodpGiE3XysrFuO0JI7z+3/+A107l7/a17dLX
pKpPTiXIoa9GJzr/Ho5EdWWLgqc1bQl7z26jX0yEOffV7tPi/9JAvMRRqjVMskFKnNNSzWRBpufv
vdA7jqZXJxGRwQoWe2kqjbJrkom2RXCsrABw1L40GVZ3U4v8+VJLffEH/ulV/ny5+djhlF48o6p4
82hKkrOn/QFnWBZuPyK+5/Ymup27PKvNRNcs/aMom6qSxsaNtFLJ0Oy3T5Gc8iLb+5Wj3qJuDnZa
I7OuSJtrgXDKygwJw12BuQ+dCKASVjTo4CjLgaa56CoZHYjmsSyjRHdWM02sluSq8gZ1+HkLcx6v
+2AXRSk3oRjJKvPmKQOXmXVh7y6UUICUnlYscZOTOlQMVxahf/ukZoW5at89kdwUOXLTpuS5HyDH
GYvPr9IDx4j0aFyiwkR25do+obrSdJs2nHOv3ksbu/fxKwXnY7i+NVytrPFWFmifjaYlyVwy38NU
p1FeCbDdYGTL21pW7J9t2YDZv/NHODfORpfu8LK/hplvcnvoFto17Lsr39PYldp9AayW0wjA+qZm
xcpawk1NkyJwKOd3MJIp6hEK3b3r7zBMC1ptbAM/lXNayuIpd1MOMnrk5oUWR/AEYW73EvTNteki
zCrlS8Rr3DmsnW4R7lYQiL0l2UL12kk/yaXVGedp12Uf95RH0cqOO2qb5ZIvsoZQlsAH9ESWpl8l
DoZUHZkvyXmCeION2h1MKgPl91iE2v3AN/+X75stGbk0JosB55CszJ4iwaUDxWYkH2h/WPrqdIDp
8vmbWhMLTtfdYy5PuFx83hWcvvDsS62vSgjMFpT6rnD+gzKP1aEbJ8IlxuutGq3Lm6MvTE7biLBZ
8l2BvHOzBmK7sl60hD7hPRjZmhna5Nj0GE9w2S9CO5lWKRF4C6Lv/gy/YbmLZNfhRK1637horRmO
7LX5SMmhKc1ClGp0iluGJQ0hKjc70IX8f3GTfvf0uz53oZLaBgARI/xAh/pjIl0K4O5sMo8IPXoh
tbLpwGBvrC/I7i1FqXnXgCBwo/RCkz+rElQVS2CGP99v95+Cows07q/+cIQHB8MsBI03eD7l/jA4
4My5xw+ZvwzVZhJUCwzWrthPnq60F6nwm3LS1PvgV4C+Elns71eLpNiiWd8siWT5r0ZCvfKI1lJr
M44GcHPhm8I3K0OOFWuYDk5+h97wx51M15quLdH5IWFCmJ4Hzq40V2CumZYpI8izL9VSY9G1IXwY
uBveC+5uHLS8ZD9zqgKjBNduGrrPrSk7LYLr5C1udV9TtOYdPX82IMleigTCYr3kmkTrMU3VeZ46
fLVDgZnrejNpBReXqXJyD1g0PuTAVDz4nRu8TDZuX7nMf6IXuCes3f6DO8EwUl0AH7HbH7jg6rBt
fSktwS/hgDTWePjxn1ScHm1G4HyZ2vNv2+C7tIRr0fr3RFRnJkJyfFB/3xM8ClkK+/0JJSRm8McF
iCxzAkIn260YfhtCZvbqSs1M0nIgnMvXMwBoXWmnRyyHdGTPGC4tDMd/GhIrbIjN7xEGfIhApkoS
7Bbt6Y6kWdI666USzJ8H2lYRvmW47lof2QrIhLBYghz+fEVSLxaV0g1pVRYzSoHBsNqP5lpzdlkK
mMCh7q7deT/VDXPJvOoBzTG/gVYcDHYkJaTZjICqtQvrEjETLOY2bBPkMprYgIVxKlml35YE/E5Q
wfV96srHo8Dj1CGsE8HTdzkBXUtereK07ubMOTrmCveb6a70nYaAgOMl4meM2Ful2WxKfJh+7ThV
QtzPNxKt95e/bnF05W71EvWO9db8+Wg0E1glub4M08akDCYFy3z5pbhTI74KzFyyFXGSM9+XE4mj
AV/efF36n4Jfz/UR49lUJq+L5yBmp4/gc51DY7v9QQgUSbnTMYXD/HDhXW63jfo+wdamP0TAkbuW
5ylBPNHlSn0N1Sm5tr01i9NXZdNBXIvaMGK/WbkGkS8EHsThvmKoPyzMW3OTr2hGSyVmTYysgJEM
ET7zoVzNEFTFJ8axUBVGy3BR+adXMBjEkUq3rFeLipSQAUeJSOtU7s0aRAoeDRwU7VX8g4J3W5k2
PS9ZyaOajI0Q+OkbjZZV1URLAoxhtWs25WHbsi2V71LCVvj/yxGuBktAgPvQRdzyKo0PSw3pHjim
MsiCDvqvM1nkV+9pRYx9ND28O4gn38exdUBpq8QGR9OKvxEnNd6Y4FYQaQ7TwDzAsxGtj5rFaAv+
INRX8q3LzIeQu794L5suKInkSBZJOJMjKxfob/FPVEmff7v/71GHxXd5PH76lihGNlk9QWeQeT4X
E4lkyMruFdADpwvYlUA//SHc53b6QGJrPFdiExdoIVrGzchmaWN4cxVvc8Wca/ainPz+Lf3xCIpd
YxiSW4WlttTGkXLhR+n31P+syPryXt6a0Cza2Hgzb71kjuoJ5xF/hhzd0T28CDBAJmUoSP1bQYz5
BTULOEnlEJslNTifDWIoI9k7ONjusbTv4OJJ/14xQR7XHOwNh2m8m/rcSMgEKFmt+Nf88vbRuCOE
CHcEX5ohwTvE+vsxzZxuCF9jfS2LSmqr3Td0ac+MkHIMhNBcanzAAsW6lUVyclNOwwnwwEqAbGWQ
DQoNVpcCf8ZgpvSUc8fDXyWiFMyaljQSOOuUmYdoOMcekuhTwajcH1qYHUZrfja1WgHDH/ohupZF
zbOCvKoSLEbuJhUqUjxG3oCHXcIO2CTyEslZ2fpAVv7lfUa3P8g8L2gG6+HkwHsCO7vVPHBXvESW
F1qDVg3EobLSUmwAlQWakQ5ha34Twd/NLSOngart38fM4pa1i7c6gqgnG7SO+56hErdDfKSQWkxh
bkliWUHF/vvL0JzpFyTBzGiCb70h7ME+JJ7VA2CaB55N8gKg6QxihiCPWEwpsCRfIQ6AaN7k5yFD
NnHUJnFxAt1FQrbES7iQgkxdarTq2dGhCvuRyJzufQJzAoRGUlNMwdzXeuCMKofggvChSQPzNWi8
Oi3UtboWjVEwIavz4cAh1+geThhK60L5bflCL+10FtK6rx+55vIUjBLqSYaB+9cVgThxuuuSEw+A
1TKjciOeXuc3j2FGf7ichFVabjh4yrzjUIIjWxERYMFm1t3DfTjVQtbyZfmiPjpxkEAFtaib1pMz
AluMafASZZ5BT7QOwF+kuYdOoDuVAEEqcm6/vRgxDpUXIkSlYKwtkQrWoIbp72Rf/zdwrhVuaXKx
eNXqeV26JgwYhL1SqSRhbDHHbuxoyB2KbAP0KRszJje7owBS8CePArQa7iC/VvZukYnUGmWPIrCG
rziw3gvJZtkVzLO9qAHmk1KY3EqLSfQhGOxnaYxMb/QuISA5HuDCUkptUaIurwuGFQV7+2BKYo/4
ikbTx5wmGmVUWQKIsxuLqqoyszVfV2ZVSY34j/Qx5MnUlouHfONpSUaBEFXcKNcKDQOXESD0FJPs
wxXm+NwKdgmQLwf7Kxrz3fJU+FoHsFLjLw3ko/ZbpNZWkNfboawPBq7K3V6INYkDiEmNF3xFCCPw
teR+z2ch88TS+2szdCWECFLUdv2d8RW67TD/VRq57DrBp1n0wQpzy7DV6fwR/bHz/o6sImfhWWQN
u7KjVGgmg/NvTUFrSCSjkJ2c0oSsJsaVX0kJN5L3bSbI7t8qgBXRUC2Dm6BSGRycrTvlelMfwH9T
Yic1tJvFJbJI9G2M+sZLSQh3pPL7b4mTq6Y64xmQOpu3wjPHN9+58TckwGkmLqjEUw1WZ8iS5rdV
Q9X1he8Dti7pPBqt2M/HRi0l4Jg3vxntWA/CPAE7vryKgoKXFIy9HwcnDHDt2RshImV8fK+hNbP5
/0tN5jOoJECr2d1Ml96agcPbw1Ejc+/XaLGfK+gaOFKMRJWzyDx+5rfdud/F9rbS6pla0O6tgPwn
Nz8KoIZgwddRncY4tTgR7CyDwVVM7O31I0D8ed3DfOCDl8iROrj8v6qttsP5Ftl7qRa5w0JQ4oEH
3Tq5zZdFxn7mUcMMSDk+df3dEBNXlOmQpwqYEmMhw1QEgQaInSo5euwOPQoRHBbr0432o1xC6pQo
+PVUXEjgrTua1YCq1KnZM3WfLeFLCezcwF5YudRMHBEqXdMBLcc8Qq8QcXtCgzOE1o53qrBXYFXP
zr+1ZA56TP1myFf9/x/R0auhigx/SqZCfWRbnRtVAgJeSXetq6Fyi//ZwSHo47NN8CtoFxyn2HuR
o+P+4M9iYkjzxFC2aM4366X6RiNWr6jN2iPDyV/3FLeOV5/fNOI5stVBBCHg5xy666+at6V7T7rW
UpCpiI0X93i84aAlk22cwd7hc3JvhJ26LQgLwKranQASKk9ohBnVSHeHnUz3z3uYx8MBxBQzwKUg
Jdjj4Mia0V5T0ZiBE6Yn6FeQ3aOnSqb0PF4DMjLj24zpR0gIAVskDea71O9TaDbilHzIyYCvxoTe
bSHbTU1DqUir2wLSsD3oOJSAwK/GdLNkhWAfl4r/PXlb+q+A5P8FRtc/0rSrFUGaJyFyOPUdXKk1
lcQ1j5xb8pNDcuKROPcWPdLdGd5zCS449E4et3yFAXZm0SnN8t8jUabzYSW952YqE6cMY4aJf6By
JwNVeN0hwBHelGN0da+P511jfySk/28WYz1FR1okec+uZnFQwwdqrOkqTUSAu36WkCbvHxKS6qkU
pzTkiqud2kpsCCNEh6nctu26uT30qNOfcOx8BMSoueog64pV6aroFuChQ0kDIGqLcBN8qJ1Izcbw
0d+r/jPqQkPnSvrCZKCXNAqlCtZTRpDiO7zFEscZFbs4JtluP6mA+LneqFVcv6Fs4tET7IvxxOsE
LCz19FbV5mJLcMcG6z8ifpcK+ZO3W00X32syWiEwLu3xweVBJ0tMKf4UCJmuAoogZyrXdMrJTZY1
EOKL3Jz6o+wUkcUDnRwOnOXv/mzrIb8CazVAAM6qRfhec88jjQf42jyCaYyf7VfoAlnUKpaIoDxx
Xb7Zyrj6jSwRBMuutd6SB2a6PhgkQYc/puIwW8NSEvqr2WZg3dJ8DPYa7xsLVXz7TiWVVD6eZiW1
SxOz55huJzzJ+jcis7uVM3k75tIGI90eETgELcgMDf2UVRmgkzMaIvMkvX6ycS1/VJ6CcoEWWS7j
4iFDPCbdFZLagCeziq0HDGNCQE/Xd8xkX82DM0BO9DmuMrS06gNe/jIJZcaMFXiaT1wjzpVcHDgY
bp+9goGY45d/E7BPfRYKedieMLN7tzFXiUXnh1Z73nA17KTU0/ppw54OXx2Br0ZY7j4OQmVfoJrY
+WlQXy6Lx+pzl7QTI42pOA8lZQiBzDIRz8CNKCs2O3C93TDYIrph7Dv05AzWx9misYZnXpqpj4wQ
wv80h5joDuDVf35bO248XKGIGpWkl2YwUvSR8hfCC/wo0/nofbw7sUd4FoCXxRgeUGi1lGcGKdRj
rzCbn2328zFX+StOZsk2HDXy0SImYu01RY+fmRK8m1X7bMKEstiyqwqwg6Q1uCUqbck/TowTGfsw
ZuRjSR+hvPkm8M5ig0JugNXkBCY4iA5Y//8yqAcl8zMNQP6BGzLZlenyIrNO3G5vAt+rAv0QcqDD
o48B/CSGZqsWfpy5jCNLgE3aQFflYqkZAWbX57qjYT95xJumZ7ipYMmunkGB/DXXSskYb62l+t24
ItpN52Qh7bIlWJQqLFmOc/Tp3xtgFdDgZtvNCz7mGg5qD6/jB+6yZKFS7KpjSgs07geCUq3/VgKl
4P05beIktHSPPc1Rookx8X0M4taeTkOmKGaOPwyQjFWQlT4wR+tWynrU/ojVMBhR1+AB/vnps5i3
J4HAwhPWyGaY5r/+R2nj+7OZEy27M6GHakP+gJaJBtRpP1bZkMD1BwINRjqw4e70Jtg5DLKIqau5
p5986FynDHpgGu+t5O/qci4SVyv0p28ZWZUa4Z5Kvkj+se4gdrt/f8o8q7qh2DZG57089qDhNLCp
6d22NEHEo0quaj86xGcjDSac5Y9chlJdH2QCKBW3t8pgPApbv6MpdzT0RqLp4kudsMesDaQMy5It
SXfIs/uFAG1c/ssM13HYs6HPFNWNf5udMUDsdpF44CPaTBrNKUy+inPw/Ul6OMaeCG3j9NHufvQG
2PDImOGnb93WJ9H9D5PSL7LyKTPlcfq7a8uHw6t9yARH/e1CetTFNzpkY98KRRxPMJXr0QybtVEN
KM7guQWBskt2a/xSaJtp7jn7h//tPj9EJXEscKkidzMzHH8w9Si+Pm6sSM+5XmCRw///8i/BfyB9
z7KCEeT45A5poZ4/6jpPjYm14eDI+BDSEOkoVb4wwIxpZ5z+HjSAmT6DkYIlw84eKzPxOhlHct3A
TYljoKywVPRmvG6gFZKhFAvbMAT2BtgvkqbNxaqyH41VSIysShFoMnTYCQCSMqqmN5ITfN3DaxmU
9SEkuQXtE3X6DEj1YBO3quVPUfWoI4KuCIQQyndt3cuqwB60LqTxBPjbEbcptIsBaSL1Fvkhhqhv
gYSA6RRjZlVGp+epHpCPpyHbWNszswSqngCwCwtcs8gGZxp1H4mDY5mdqIYTqXTQzSd7Fi3DkfoH
G8RhAkTpgS7pT/O88868K35oM75E0EMKEj2hqbA2JsF3b8cd5+F7yjrRs44XAWGilg74l9XDUB0R
RwID7+1BGEAr3Bt/1oFb5/XuZat/oL00jhhmKpwhgtf+xIO/c+vVXV0bkm94L1MzgCMQxNR3/r8T
xYAtB5nZlgsny6h0YcIqyWbRIJF8NU115A3xVacYxFXqCvLEc4nbOb9eL2iT5cq+o6Y4rfzNEjqs
hz8zzHs9N70uuxT/Jx9vzWtJ7/WgcJUPH+ibKdgfWh6EsSi4SJ5RueZu/a7Aeerecu4hxgHLfde6
NiE4AyCMBGAPIPBqGvm36oJFYW+QbTyZ1FpR/KfAYWFFNmmpb24suiulaFdRK5cwiNlQCx6c7N3b
fv0lnXFrA5V2v+7/9ltb+7RmB7rz5bMhGFq8c4ieY/NfHRirg8RVVib6Gykyp19EeYyCviyglmEL
XdRUko+RDHu2Lupp0J2EjvL1QDHG7ZAWtBdWUu6BI4acAvvEpT7cRyma7yB5DLq2Bcy1Q4EeG4O2
BYK6Jv0hGVDZzUh/dY8d7ZKwXY/Ivwp+LR6gjcHnPCla2nXtQ8p1JCdmeG0609kU0mOlA9DrcQ2s
Ib59AGpEoXEtH3YiOAEmGnLOE65nwvCJcw0W8Sui67qOBjGu2XgNuH6/0RXTLIiHuJrv0Oc1E9/g
S7TtfoHEpeosCjM8TsvfN8GL5NwPPJgV4qRUoaJCX7GrnlShYaVmTWMepBDjC9u0lXfPdVcduJuA
MxZkulNn3tFMsizJELbLmlWURHEN7DpA5++JidfQFhazd9kqXpccuoDawEZAhzmEoFHdX0i5H/ts
JNJLbhLSlNUPlQp3wpadQXWYswKaTdv26bqPizykKD0JC42nsnn0RraDHxvVByeXmIYgzWbYB4Mb
7HFhXpg1i5RuWMdsg+jmDjB8Ykm2k4L7pe8Q+Jo/8q2tVpYdziAY6MyjBpN3RjR5zsvlUpQuM6JX
r9FMXOo0yyznajoGj5hnGGv5nqgqYOwwKfTDFLZpTAl5VARRez/KimvwmeQsy9GDqneAvqB7SBbO
7lQ/D6UCNmnC7qOYU4o0K8zb2UHwI4ZQ5WWUhm8kpF+OalDwwHUws1RL/XRbwIkCS5L0t1Zk0/iL
R9P3xvFyq8JtMlfUixSgsgLCVp6kzWRtTAYBQNFbhEq9U1ga98dqMW/9ybgrhKJH+M0q4tFP4J1K
m4pPZ+BLgfDvO+WWEnkar4k7jwogSPT1aC77hqrQpxUE5gRkZGWzR5mlzAvbeNBCMtirZvfCD9/B
KgjjFpa/IDivS9RSmbObHATna1/d7I+XMpymqBTgKMhSUtaD6ZXDVlbtaBZczlmzb8VcdBbgajdO
pQGFV6Pxqq6LmCw93VadDkRC2wMLsJV2kfk1uNIja9yV9c09De4BetH1vKXOs/xrML+wX6yQO/lT
XVA1JFBDagNBnZxkdNu/mZItB7nFaVS3I/ttIgfdnvny+F5KhmIUXiDKs70deW7p/XtJDVvO6fiS
KKEp6YWil+4HpQ0Q3rwMJdR0KwCx31ILBT8FHmyQ8gyd2sNu+BXLKIfzmBi0C40xMUKF4E6MHUsi
CQ92dGMpGyhje77gojHT2ys/4m5xmdGfb/N1ASpiUVzRvI9TQZhEvoBEQoPryn8F8wwJFbN56uwk
zs20OGlIFQVzmWP1XIvzaedoAVoVWFpvSKMk/rDyAXn6uWpADLqCL9NfHiRQxaPkqRbP3/Oxi9eT
zZ5z4l8od+p24Np6BxT7USsh52MIvP0dNtAbP2QTHkKMz8RVBt6SLKYyEH9FggIGKvXi5Ua27llR
5U9XfGSAVgfeCmi5YV0mIuTXNPt7ggYhcHc1Nrc2ePR6bdJIHoTYwA+Yr6tX2YqaFNgBErPRD7U7
4ShBu/REfyVHqcbtsev3YDYYn9T3RsSXDOsnj98grbiT0tuUr2XI598dXnkLDEvREefJY42bRvNH
x+Gnixyw6zznmQECt9MxqXAYhB9blnw0Lw/yM0MNGR3Po0ysyxqU6IZs/V5MYyxJ7WvtKebHv2S2
IrRBpG3wDpywyHZrt2wTJTy37lO4P3i8YdvucUMbLgY2wLHW7DbecEqSgpykn0zTAQeBOZrVATsC
dJiL+77qyBHa69F/4RRUmH2Oxs5Nt943ZBfO/0rt6atOgtfVgGbRYItxYjtHfXfUY0oAJ8+soX4y
nHC0AcJEoklOJ/eUCPWQ6OBuJJ/kpTAGiRo4mDcwUhTjBwMClgmfpqkDcbqzjFT3GKQvFyjj1R5N
VUQFNFzlzbywrLQp0I/Dx4ALuLT/gyv6TxdHy7Y94l0mC7BuBoWPl7xbFMs2dVS43ezqFUe61CLG
w4B3A8hPiHiOTf3cms8is9HbS61QQZImkc9xB5EePBpUwj0JgqXYw4o1WffAjvvOoKNsF4Z9SyFD
ZojYMkRbSXgPAvS02x+1pkNPzPflX/G5/DwstUmd1mnAkAxMK1+25PxOC+4OgOyrGaklcoP4jehA
fFSz7Hh8dOlKffRtuzVwn5sYY0c4cfR0+cl/IVhs4BOATUCOBnAYGtZRGV74UeVk1S/RkWpSA48M
4hCTjA6RwIxkLrMs7aqlTCw0CArDJo/HYDt2oB5bCm/UmYZtG9BIZvXVQTls7PELvZsfBLso8Moy
xzAhXK3QKn4jiyRgYHf/Ydcu7XhDuz6fDn28/D5+FE1WAqnaP6fRu7+Jb2+pU4W6ZImwPLIEhUgX
4ARaIRJfDY3SseEz8U/xkdLfidLqLxQ2mg/FcK4AFHdXlPnxZbhf9FMTEPPBb4KdmCowSmGW2FQ4
5bCIfXdBWvBkLT24PLiZ4q1zMlx4fgxzxvujWhcPkE2sFKtk6KJyZOE7wcHWLWnAPNk+Wdz7t57o
TzP9EnMGIkyxCTTLtAbrMFOjFmHdqfa9N7kE8dHumv6JNI39WglsrGVjJXQt45IDagJq5l1qCXQE
jRoxrtvUSxCgbMlK5NC8rcEUyUrAPUM+hIugxBRhJFPTqHivqntO2b98QAr3KvB/TwkY4fkhGKLm
/uk5JEhMm98lKRK+ip+/6VeFqqlCfYsjhJ4GgaNbFIWvt0S1YsvWvgeZ8Nv2n84PfNgRZ0cwn3QB
tHjIy8lr1cdkFulby/R2WrcaCzjvdei2ckDF7NcZT7DbHuFKnNzKXW1S+K2sxIvBBbNi7jALxbcJ
ip230D3dUSCZ1s1sf0Cg4KPjkXMZ7fYwVnduEwZArJGla5LHkESTuUQ0Qb185YyHlp6BWCfdYkcl
DMscoM01AEcgDRhxgTVdSHKQe8elixpAvbEU2AeawmaRYNWgZm6w/xd0OQlQLC1o2O4MLfTKgY5+
oH7wAItFr+2DhpQqwixAj8ZGNC5IgeO5K5yBDi4g39dqeF2ZLCarCGcKsAaNRjFepkE2AxJfzwNK
FHzSkJOxPw33GaRL0ZstqxFg/X8J3FrRkERwHhhDteMNSCJqB6wpphVsgvXP7XNZXIQVTQ43/u9O
83Ap6I8oRTtUM6A2Y5OLhk48sl7pObJwGdDK07SvB+1n289pvhHh+GMJxRJUDYLYB4HK4sq+pPPu
e3b331w7DZgpLIcKRrd48yfjDlUY1QMASIHNh8fU2WfkWK9aTcthQDr689rdWVMC6rCb9dMF8/X0
tZWnGOLxk66+8QRZZ7QPYWYTtXKa24lVv3jvZ/7kcBH9LWWwsf8d7d4BmEt72CLaOmzrVulUpGhF
Ey7xZqz03IrKO2Ra/zZAcdt69wPo6MCjIBD2aPOp0sHUPG3/iDihLZO60wGHsj7bA9dd6io8XdXS
75xW0sMdfeW9qFjTka7DxNOv5u3a1AVclo/tGvzLusGYWQuUgGamap1dyqJgTvgYYYhelHSzf9GR
LNSeIA8iZ3wUzj4Hna+Pb9JYgCV86Mgk+cTuGKxO95piYaPUOZrMoWXHyw7otISB8AomsZ8Q95PA
KHQSVUr8eT833aCmnaSPc05O8Faeg5ZjwVMexQVho8BApBugfeaCdLWT7BVLizs0tnrloqqcadfv
yUhaRjwVNpWBg8hJWp0tFHQ8gr/fWXqpHMMuEpUUyevLW+VmAvQxXm3E6jmCOzXhJu9nagI3hYwy
kpyl8cREQhwdUlvQlTfcFars2XToUINGF0i89TeWmV7PAnH+ug8IZf2iH+UKl3D9QifG3LWvtFy1
5+LlW+q6fFWa7wajpbxLBsFyLX52KrI+24lO/7CG5Rv5gzX8z4CSLAtNLltSui6sOCfatPvVutHi
hUCGcdRTHEs0y3X5Lkge1togmnEIuYp/byRuJScjal3cPCLboXBXgC7H56NTpvXe04yz6GBFW0Om
9kGpK9k4TRcrOlLicnpTmTGwEiAcpuY65+JaFIT3xyLSJdzt4XVQJaLMJVxENHRlwC9lZTN3K/V1
cr+vl1WlFhZLi8G9SmLY7Jv7bPO8Av0UnaI0i0Af3Osvr7uekBB5DTx+WJR5bZ0pA3HxUUtN5m6U
jNKfvJVmRNdZpVKPSpzNBXd8bbQFEao1m+zoFcR3W3+efjUFbQ2YklJuIK/hFKuSEVtmx821xe6C
I/XoZlck6LbIJuglHLS69lx7QC98C397zCgXToWtrwxXjzZjCTm6/SH3o8eHnMdKs/XUpwmW2JFQ
yh2e5jIQnWYHLDkVZUZd+VF1znsQuyTjFYm+QfyWC00GHxrDrq0cg7HxDLKjUrDMMYOrIDvJKTsx
GxgnQPYL17ApnS3auW+yv790WRmf1gbR8sApAlj1/BMq904sE6/A7qhmkQ6yuLjDXqnplYlP1wDk
kN8D/WA1GV8LrpVT0IzITRVzU+tOhVRjhXGl2ZjlpdC9bf551ZCPnYTKYrtdpAelD6PZ5OXAkg1A
0d7iKhROB4xhVDXsWVw0/7f4IIc3klBVI6lLlqtH3IuENDf6FFkgKbgSCnEbR7rxktmadEpdb4N4
NB9X+ppEO0Etjcw1sHhqoDULNTnPAfnVfo0R4VEbH0xE9HN5WrJDk/Ae+kSg0Mp/De5+ty/kMNaf
If49lFjEJL/VC2jYOR+wzdDoLstyrbTk231VN9bxuZO8powHPEZ1Fpoq1cEJjII/K3gJrUNi8qal
oEAG3uaN34qoPM13kinvgar0tYFYzdqXBP0+RLt8bsbCXdQmrI6oGPOvxJSDSy2/xgZBN6deA9V8
Mv+l2l1kGaeiUa79xvmH2TG9RZHQgQPV42ITAtI/d0WbZjtlgl1qmkZYGkKV5nlRPLBE1bofTvJV
BD8aNH1rrmNMOx/pNxYOFRrEMQYR15N3OVvAgSqRtjhJulSjprkabYXI5NU0HrEcMi5jnDB37zeK
gzKGiYV6bHYK6VGRxICF8caRgpThN5N62mdM2nmmY8ZEoD9iAbBSaTsS/zSoe2vKPT2lWbJ5mrt5
SEmyxfb3joxpFa5uL/df38DiwGzGMo8ZM0l7oVnFM2A6tz4RbMaSYw0ZTyi2+n7TaY5bcyld8woe
NRxvq8V+1V5PJaWHknks4y2Dn+iiMpvCSXXgvKB9nVvZGpwvxZVBIHRcJkD5eUG8FLQ2L2BXzeTA
YLqMkk2bKWhpud11a+50etsvMoRv/gv0o9QJsUf2iDXMan6bCLIMbDieD9LqpzBwmXLrfppiLFhF
aKGv6AHkSEVfCddFH6AR4YWZLDeAcfvJkQ/jVhLKSIUXbbdGBrzHR8ZO8wwHLM4ljBrJvMlGFmy/
TOT3sCyrliODErFNcf5tN91muLVW+j/oyD+HPvA72i7D1j9yLaXQILCuaXdXmjKeIuUYAEBw9Uat
S4v9+EaA6JMTCZg8TTLh+WE7AwGN22H0k1jrr4A6H3lyUAmRaZKka3LLPcTfenVPokam4VEs+CjZ
8dlFVOKFzJcWFvcylw/isph61RSJyELW6p/sngWePtDgd9izeByaaeZXVBo5QkDkAjIwGzsqibHC
QiEMVWD7Abrfyqj4u720vcvObzvsT48Jt0oeHkbMJFAdBfY1z54DpTAds+Ngo/ei6m68u5AIBjI3
s9J/h1agr7aIhp0k4B7N3WiWWELPGxFlDCVUy/TPI1q3wsZwKPU90FWm8pIjrpBLBfNHRxzCafWp
1K/WMtCEH9eMMJR67Bg+c3LrfqvqhPB8FtujCX+nbOa1pfpwTW7ILRxc2J9yW0ZmLCDI+hFo/+bV
1lCdpNxDyLe5AyP8jvbyGLmeeOInRsQU50GTYMhWU58hGbNgp6TQRhgv+25ZGFhBwEhS1DhTRJEY
5ZZ+4ei6yWWHP96rUQKeYtU6I8dU5h8cBFzWJFuxfiobieQFSBH1Kr5lVkLV6BtKXYKnWib6CgrZ
Us/OxXOu76yRaph3l9OcaXChL/G0cwEBbx8+3YQO2j6ahk6ktDz1/dllKWqoic3v2FCbVBlegK/c
v1Bsu+56xVl7hJaRkoJj9WzC9Osa912rH1abhIkBS2v/oTGnpkglBmloBm6/YtBwjdrHmvWESG2S
AUASFHqbvPpBjjZYMY/D9U9/SCHUy9COt+P+XN0ePhrHGJcMYHCbq8gOPaQgPhwlc7ec+yTuvIEK
1aSdqDU5Yhry4i65ghTFC66ATfacFiIHEg5ozI5S2wmthSnYXsKHHXwzQFeQnJvnuj5tvoZ8zIKX
ArH0zxc8q4KgkzvjT03QM5GiRr0OHB8TwPXWFhmmR276VNZplTCBi2/B/FSPzorwDl/9A1x+MSfK
EBBzYXs0xXb2WbVdbrzPjXzaD2sI7iH35w7u/TzZjC7YWyhNx8k9dTM5+NNmkSn04CXnbvgQPVR3
kSXwX59Z/AoGtJBxVwF3n42bidxwK4DvxgwLsAx2maeUMO3Jk6FwO4/357ELtsX/J7lQIZptTePz
JTYFcFi35ttIVAu0CvSb2QGItRVjdxOd5Rh8zNOuyl47MNUFhZBvHVgj5omgDsUMfxx381U1yWMr
fOfwTlU62xuVlFPXgsV+edMnaiZ2YJ/8bkPkjE+AlH+eQLlzr766wIFWHo+FSuoDl/kS3bXfun/L
zqEWxJJRpEKUxMyXkBpMjBfJSNshRW6MIy4H66xG/Wbpcb1aN78S76k3c75GlFRwLimLHXcUT5oM
bVeeUlwAi8VwS1oIpqc7wnpRyVHGBWUOBnMPPmXhliqcor2/qm0zBXHHsg5qKfL8q1bD5uAnDTmw
t0Nbk7OlqBEw+9f8xrmXoYA8FqFaO4d3pTQQMnVpTDZFAJMIVS9enqWr14sA6yqSCU4ATyUi8NGn
EQ8jZ1I7HqcyYxWMt3IWjjus/rdXrv8mjXZWTtL8Kim+xKUObSXAH+6pWXb02u4UPyG7wQretoML
s5nyZFIR7xLyvHquzu7R09Nf+qrpTtSr/iCGBS2RqS1qlgTTZWW4Chd+qIfLzp17LJe78HWSkZPJ
SO+dTM/n97DrS5wKAPT7uk5lyjpuu47CzZ0LMPyBhugkBkOhVmjCROzIlcVb/vPNdGahieF6Hkdm
1VgnO4Lcs9UOAUH0LuuCdWSnvK3wKd964966ruM7POyiq/rAlWDAUC8kf8TyD0GCjKHxiWFtu4UD
h9sxB9RB0k7CM9qls2rleU+TcqqcvlUmSUXaG59L2TGCc5HjMj35aDaDr2SfEj+R64JL+NcL/awQ
KZzhbooo9qipVDXWCj5RpVHw06Fpa0azx8l7hXJWIwfCFn/k2MM0/Wu6Yk8l+xOzgtzLmbWgWIEc
zOdXZY9RsVIzoox6ByG5N5RNtC/Geg6DETsY8DRP6h0AUBXDDeaBoLExxm8DQtJTLo2fHiLpwahA
PXf1LA7x7GbiFAf6hJ74kmc/xRz60Wirk+cvlxKfStQISgkUbqUuRsQ+kvTwXBuOz73/dGwKqLRh
ixeNQyY0ag2WbxySBNivDFjBO7hEuTZs1wgTpkOjtIMxgwEiV4g5b5vDqLoLbF2o5XASRcuzTCz2
tSR/o3js7pqdQOlx8e42vPtuCRX9wxgC/a9neG307R6TqTM3PHZ/XWRnFZDXg7uXC1pcuq+u//PX
RfnAbNaCmLYm/levVMM36hTYZztaaOMwOb1BpIqZv7kUOPepDeKnlyiF5ZhmxknSKpJMdSCFjoVr
iukBj9cuky8o0Gpn6CKud4I2bdb31SG9Dp+hrOwNNVb+nfmjyfhqxEIMzmg/B9zk6H1CnF5rtq7D
FIw1GjN0nnvqIfX0MK92HwZUpsiDrUUr1BlEul5wF0sFUY/1mo6wQFmkvxODwh0dxXhbpDGlwQvR
HuMFsq5W5giGijR4ITVeqQBUJrgj4VWeTJSP9d483Y14pqPHvDAEceTEBdECOGnEbkl98HIU1V1z
/2LDdZJ9EB1I4rarpO3Bq0K4smZck34YxrRajHjhuHBJRtydmrpf5k7GRPsdUleZnjbvKujH/FMW
OAk5RNFUzj6fhaE633hS/zNksBTqnCSFeo1MNZ+Q/KDQIr/ypmgNQV4plo2G2CXUUMLlXs8i6jKW
EKvhmJffm5eNXHOoQTDOiRMhdm0FUd1s/NbJlsgjqib1CDgQ8uBNee9cqJpo0SNKVLp8KCVnzAUg
2RiF/g+N8S6C19ysOnN6JTZHpSFFh0Mapyw6aN/JioJ81fclJS4gIHI5A2iVzGZ68oEK/5XUgzGf
uQJVFr7zDgcRKwl8VGQHPyG8ccszlpcqedhSLp/JbCmR/HQFfJKYWs7ilXZNhLu10ug8EScYTVKF
iCpRQ0HE/dCN7jTqKCfTWtsJXePhIh0Wdk8GYpvfriKm2BVFTV2Sd82lYkG2n139LLUKVQqPgnP7
c+kA0umtfWtq4k1x6KKXsqCluWDgMJW8fLOFQre067l6Yh0V7AR5RnnSed42RzymmgyMaLlnsdbL
c7yOB9uroH+gfj7uUmnETkBR8EBTl34FDorR9y1Cxm1S3SMMSVPiS0lG3CTLN28WwZmJ7K+nMnAI
+vyCKHYE2coOOWHyVPs6VsrCHE7tsR+SbfYMppTPsCj/TXITkheGEC+vbwz9bc+wyr8WSu5yFQ5Z
8whpJppNTKxzEYlOVY6nvK4F53WMpuGSMnrv59oz1auy1nd1dfHoqlEO5Ip+gIVBLGNZhrUt/803
RXIx29Jyw070xc2wzIQmDwR2Eptbb2DdfJWMMAWH9Rdi9cOz1xo+67PxS3nG836JB4mESEYNwuiJ
sMdD2DsGSZCdCRmGmMrbjQCE0DWTu8MMJMaMd5v5H1R+LGq+TLwx4tbT9e7WztD5nkDQj8Sh90Be
Okg8wRD1q3B9lE/OZ7dvgO17LXk66y3lMBjrI0/4yIE9SsVEdVf2W/hAxH+kg0VXfn0Wfy7VzANC
hP7VRd3DNZzO0JlStQn3GyHcgdfY/yf/WNNYuaFksfiEq3lmD64/hdp80GQKQSQJYGhzeVwc6Z0I
713kdrhMsMWcaBZ+YX8WXEiJhkKjT4q+jRAhbx42kE37iNzOz3xqfWbd4K5fMpzrk9KuQ9otGOSt
ArC2EAeZ+7Z+b5gogSgm8/ws6rXZGOE0Lpz1zfsua1RES0iHLHb88JL6mEJGnH05huxachFnmAs3
pdJoJ7kcrkeZpm0nTD3scjb8UvyjXx1R+1GlvqOrd7hkC8Zp85x25YrciCnlmzyJKAG7sShM8O2Q
OJNsAqWCeRNKqfcx9t6oNolKexPjfWnYUteRUPByAf8oyQTUk4aTOmjXAEIwG+61BqrQnN2Ciwxv
wJtdgCRgWMzVD/FIJxJG/dsRLLsvq1NhOqDpAWLfxJYTZNo1hh7hPIWRMau10BK89hHmbiWAm6BK
Hc31Y9Xp9Ej11boL7X/+n/Tf9BbMdVyOQXHknnGNTsTrBD2L3A+AkoLry4SqQQqWCfYqT7MpYFlR
0BcAxuRO+Vp2PMGkCrvpC6kZ5U2XoBSoMxsIsKuIx81ByKwtflPp/lZQYHO0Op0DaWnjE58en7nF
swi/54cJQayXsNpo0VnzkKuO7YQC4lFbUlMn1cMgAwNyfDJrSPXOPSBpc8YAnbeEXBg4KUZgT9ho
7hImjT2KK/NuubOmXkSdEtmq3HM+U8NO06vVthdNP5BiwKRFqF8j3GLfuTaAi1PjawyrqYNFVzkE
Kp1pgwKocQ1qVXIjnHSyuqDJvQ3xyeJwmShCjRZuR4ogRRyY9/mNULeh8FztbOihQZwYIKUUqxmv
fUNB0IvRi/ULd/eKflg6WjHF2uaFu9NhsS8WaCOlZmkw2Hkor57Nw9UAUyOnc+rlcCBUocDOInWg
Jp5r/LuXBg6co0rg/tX3PZU/4IRCVeMaWaAi4gedIiGe/Qz1K2HhP1/8ELyixOcYXaN6vfSFM7Kb
KjCT+9urC1GVZnh9D/TztZ0QNX+pp4lKbtU55IkZkYeL8/Sj/PnpNBSjTMKz9bpNqRI/zMY1ae3u
sF5QV6nFyzTGfmRN+Fey0+p7dtSEEINefPq3e/BeSvbGrjpCPsBNEFcMrDvFb2MVJW7p26ahf8XL
ftMeW/2eb4lkhVWcizJXYOtxWjwGRex5qVXMn2CuVKNBusdBcM4gqkDeTfRwLpi7wtJGKcKyM1W4
Cq6QWF7FzgCt1mtanpwy1xDuga7Bjy4W56tdlCrjTwztcDaBtPfdJl+cYQIl56llMarasoz4ju9s
VottYE7eK91oMIxwA2m8zwOTP6n0eX1BNS/f7vthEHSq0p3gCRNeZFa4Xem7/RQYH/7in1gdSRwc
rK05DaeU7JpgI1Kh2/mXx5jSorrj5Okrl07sY0cHL7W+hDagQQ4pJbTwIafSc67wB7YqQVT3WDaS
4Rk8vgNkJcKaEtX2lMBtDxGS2yRkNrghffjxdZRjwbXLBpBBxXPOnO2lErLACQOIfkZr1vSl8YrX
r4S/91tk/V39L4eN+VzBmZohdro5U0JGcRhSjpV9B6PyXNVNuR2bsoLCKronXGvjqPEdRu0vsMYm
z9z9C+5L8vfV7KbFusTUpdsYCWW4szT+yMB6jBRzoOo544bDNHQ3DqvYCbz0Tt/zMiYY3dXIO+OC
gYkBHloMtgI7R05LzNydRDZsngebVpEWztt52Y5u7QqOxb/eYdQNmGaWOfTKTE1I/ZIjYjBFsDv1
IGlQ9z3i8RkhIgIJ3N+anel+9FemQERcHfj8CZJKYfNiA0h/WB8wuN5amLnRCwV/F8L4wi7CFshL
Z/9afiCaMAATk5OTwcbyAGwnsgoAJ2hj4Ed+sO116bMo96OII5OO4Alr/1p1/ixZiYfpn46S++3F
TcUsBkhg5+tnyvz4mBaubI8mUUWb7YdTvEkqnvNY54tLGlOs4peWtOuWeiY8Ir1kIuatDeJcfINA
bEgQxbF+zYVz/P6duVgqg5saAROfyLFGy19TSK1ELAuJAsQtnz1pnzjdnclGEr1WpkpiykZgEAB7
UdzSRZAuQSiZ3ARmutm5fW7immYnuo7sfxsv6bHj1W6GepmqzQ9ua+v987ad8xXuFSmTwRnwtXRX
8kKbvvflNDx4gYZ5++BQgJtUJwehsZWdxQ5ZE/F06o3qQSghlWDa0QALuuz02FFQGTlsuOn9QdmU
Tq6O9hhAV/hyQbG84Gf+N39jljMp4VwVrSX+Pv6KvyF1EzKcjOEw9ifoy0/38artdpK3mKEZtIax
1+eEHP7NPGHJuhB2Ivz4QqDi7+LX0bT6pHqAYgTfZ8AR+FfijQ/1LO2TFgkplbNf/mFOkmIgCrbK
JbuNt80Fzr4Fl6I1XNtnxdB1rnNcb09ED9/d42lhVwm2dcUghDf2wTXgrvTfUHyXbSegTMomfuAv
VSY7n7feoOYNVvlAXDzuTLlmwzEYIFIiDoCAG4PxYvluFG66MdPvjg7+M3nJvwTcGWnYVTSIE9DO
kUlaxG3mbctLoZooNGQzBGqMLFs0/2fSmioK1W/AN1qTCbMUaaIx+Wte+GtKh/Y90lAS5XRei8JC
juNZ0Sd/l8gC0W6fAYmPLaGi2WcoYqIGK3YIWuQYxKEGu0HoGig/PIBtlu603P/Uz4+Ktv0tlXLA
+RI9Z/qBzpsZDLSQ6Epy8iNA7pDTOEyu2GeHEt12hCw0v6ll9TLw8NH2x9rOcCV5Pfjnna/PFeSS
JED6SypSdWyaZ5vAQhXcGLEB9GFfVofqlR2OHyV2gwTou81+jPw9BC6BiLaSpVNse+HMSMIOXBsl
J4oEgdV9+AtYyX7qZYLEruiNZQBJLsQN34wiWYhB6QZlWPR58k+voTjBuE8QYVDhuIN8kc5QwRDr
e4MUHT+iiBkDVtBLrPDeU1GoqMnqhZRa17EO6sF4/mkjpguHYh32slhzV1ELIvgWlk5FNFZuMtHO
ptRMYai9pR11GsIGw7qXS6lra3A+WiWgQB7Vfe5xYrp4WHBcrxHJymi/+vMN068G0uzTmTj3fO75
hSGYt/7UNSXYRuheXZeP+TTf8RCQYdtCR3BNt0VLIuLcpuW+iuI0RtrtZj6mDIZbR6wQkCX+rQCP
fIMuHJsewpcxBqc0AUWrNjXJqIfV7ndanVZGk+iQhFoCynIX48GisNkSZ4WCIS7OminiOAwGCJNV
cNGzee3+3NC4b4/7rIdI3NRE9GHV24C+I9pjeuLyyfg2gNW9aTWV+H7jpSVhl3U6MiRtz2yTyD6g
n5kBoLeUv2iXgu6wlkx/yJ6jub6Sn9zNiTkvMuYhuWyJLioO5RKhTP5lWkgjKSA0yVCGoPLD7E/U
cDrLefBFpYolXtkO85PcC8GvIrpYMYqVs8uTLnx/0FNJjPOP9mCqX4Dt0an3PGuTVzFxodv+DdXt
b5dpI9AMrk2cPLYB9hS+wBnbqfA/tqYqh6lBD7hwadFZslZu/1eqcMjtpw/aBtRvhNjup9QuYKgf
HWLT0fQoN2Z+BXQhdVb/q/iDygGUQAAHeYl05Ofc5fkB056NLLLGVnKnkniMlyO+nVPHVpajUCo1
3w3thjZSmwA4DcX4gidzDhtF0c8oM50DLrNCGr8hTDTpXc5jNcVa17en42ezqCHJmAFZW6xnURU2
s89y9AQ8qki+lxc4HQhGI52ObEo/o9dHZ221ldgQX2SkWNokiMkSizfaUKbSePYgwhvJQkp7rH/o
R3IFoTH2adwfbIWmhpCiyaq4+s4MzFutSry0Nzu0a8lrFenCXVFWy4SDRbDqZj2c6z3LoSfg0MHv
IdH8RqQlUg9Cyp4fkCrq/nVAq2Daa83UaRui203PIDJtZmY8MssUzeAX9IUkFReKkinXEkaShsDq
DQg2fzrrHo8EafZuw9L528RQEcNvJMyBWAwMU8Vp1zW6Jn01aNKFQ1+ZqM+1idPeC5nmOuu/L5/d
9+pbMOmHSrngmjmXm0Ke41UCqhgppVLSv1ghZHpQQ7Mu7pD4x8snfHCzMDUXoBWkZhXu/mDMYD9l
jyaCoj+WDoB/3CngFqTcSutYa7EkBbMwhUoUF9L72tG7gnsQmW0xuJEgXqIf7FVnL+AAAm79jUfv
tw040czJKxh3XstfpEqsvrLqLizJmtkhCcnsvCSzsqaGIjPbkbfnhHK2+xi13L6d8kY9cN9uTcKN
Js+etf5YwzCxrx28d8T+rmqNavlYmJMnztWSSG/Pzo0BlIf87mI7H/yDNBnI7DCyX3FQUcEPUYf1
0RGjur9YjcGbqYju9HCkfbLcHde8HuCXk3Uw4ISk000cS8tFqeus6LEO3nT65cyAsaG2Vo7oZ/Y3
DDK3ZtH2XtOixQC4NUidTajJhVYLbscNfYjTHJAhfUa3tHFx/5O+2iUiUFE34DQWPHULM2jWuduR
GG6s5d7Mt+GEv9vLXBNgTWAsVHKtitlJMRngdPDj+sENifDg3xhgQvdJtKtoTDHkRYzwgcyRdeOV
hzOtlR9BFqFNF8Zphq/CDSnOuVsS+0c8oBMxSOUMXEvRa+d2cqQ2EEB72l6gGN/fx3QLOxMoS3R7
jVtLBpNhVTqNe6LZo3JTtupYR7WOWDHAD3rOSvZI8/okAq267tgnVHotJSDB7lth4x7hmkvusUSP
Sps+q35SKlm+sqQtMgUDFXU0xeDBWWxeW9jnnCRqYrMDy2xQNZtDmHuP0dMC/YvEnvuHbufbNIzu
5zPnMp9xUgCVsMOHFnDYgHzvM8rGKcx801LWTAHwMnh76/Uhb1I0Zf+Dp/uOhk7CLBHj/1/h3ap1
dkZhn9U0TcnazbOTE0kcTW1gJHtplAljTAt8ScOxBnGtZCE5nYnw8WlViera+tNv4mYmpJ+yeebk
5BGZd+TELHSG0ULXb57L3UJR2kA6g0uN6oS1wuoxkPAABCLuMhQozJj/bAYVUjAAlIJLnDAa11ZU
3Gdpk8iQF10GNssjlrdv6J5vWr2OEmd9ie5y9KMA+R2q1cif+8Jw5XkYluiJ+Md1fB+084mlr9oI
skmJrFNcrERObdoqj7El2c8/0Kq3dNuz3QoVe3lIzk6GkT2iqdBJSIF94b9WhJTnXgqdrkaI7zdE
cBtCj2v1aayGtb0+Yp7epuREID8pCVPdUuG1kAbA3GzdLhgikFSq2e/NRMOsgF/EILEVnCHg1zru
6WdVnVM1F05g/57+7ozjrrCOrOVPgJYehC0Bf7AFL2Cr8MVA7GNfoXFHQ0KE2Fd3IlehlCy0oWiy
JrgI+4/SjulcEDd1T0rAv53W63AgTPK/9zbRDZRh+RnJ9YwCnKLpvnR3iN8e+qEji182qJ1DWvc5
cfz1s/oUOzGXJxSpCd6oU/QhRb91yZ4RUQ/O/XhfVF3oQdULVKy1WDA0yEU03ajZL/+BxcrDoZ4v
nLze9/yxwmRuUl+mPPo5wAdQzalhEjMafSHmeV4Fsp/KIROw+0JmJYJ9/QHQy0dGIhxDXjqXV32X
rLq+eNgFI4wvPjtmCI+toRRNsPdz+cD6BVGzDzeGYfgtoNaFGnw/KYbm5wrf6+D0tjSoXKpR/77f
hRB+pCecrMJ4ZbdQKF3wWUz/4yE15TiqsIgWaEIaUMj+u3cvWA8o5X3hKQ/7atl5GdiOnIXIx34d
EHxfKPG6frvYQOiYKasz4BUNGVkPpdHsFolEonhL39geLY1pCUC9p8vKyN+/ciVbQWWH9N8F3fXQ
/CcuroPSc1nVYNBQl30Ac5OSiS5Mw1lsSD/XWNxqdZ9r01ywdx4g+IXxJ0NuQ0LcJOeYt1fGZEcQ
4tXuTfeHRzIqtNjaccMN0dI2Y0iMejdvWcurnPWPn1ARvvrRgOh3iS0YZ2PX6fjW0CwilRmfeK/n
1izQXhGc2eRb53TFfQ5+fonBIllQ0+mR8h50SeR6DrhiO43acntSo2cTuvKoWfMZIq4wndT2QUnP
SOIz0GwgEu+PvbUGvLy+pVt65MlN7D2voJUl0vt3kkxfDe9vAUeIBBZPiuQNCZ8Lms2L3u90gEEn
oFH/FQj82xzz4CgdP/Yu2PdwUMJCp9FVsPqJCN8UvW1sJEl9P0qxiU7PsUV4z7GFVAwenqGyYGHd
5iHTOdKTPQ6/YpqvTNLcCvnoI284cCI4hXVWeaj/nulReftCokvc5wE7G4DRYrtzIaA1s72cQki9
Wvgqtf1Pm6bBjX7Pvvb+TNwiEpK7qLJtuQouz9mYCFpsz93BffkGptT7AK0LUGBGqBUgXZWDH+Nu
XdvAhlIzLz3F0A61jl2PS/bwI9cHmgLaZllFEnVcLwophP7+2gPoloK7DguD8xS5TlimFKMRKBpe
U5bwpzTXxnRWzMnAOMZIxe2DL9Czp22Dpt0B1lusT8f8to2IWTOQOFjxYfY9MX91qGdI8qQ0WGaG
f8Z3bvMC60H6XIiTO8v9fLeg8PLpPFV02FJ5TEQ6X5VLhcn2D6/dMlB1ebzgqQxyYzlZVDCdvAOF
tMVwZzoQNF7Eut7+c5J5/FNcSA5oUUzVNK8g4USSYNljLDXsLSWbs0+L87IqDnkfNN5zdWIjtbgP
XIyCEczPIMERZC9RNrtYSh5nVRWS1DAkpmbii+lHGn441WZIqlR0ALCyXelLTz0KQmHpzrCv8Ovr
WPU5VybzaZXGbZQc2hJ54tY/Ppn2/pP+5gkfyXzfSg74Q3YDCml0EC1wYeUZSzonYrA6BDFrnZZB
OJ6qy1G98m4OIXSA8zDsqK/8+ClAWa+lI+ICH8bkJRoP5hJEkqRHVBh/xqhM4s7pclE06eMEIp8m
rehoG+VSxgC7tXMZot4tkpwH+9SqVMTZDFHdLHrx5ELFi+ByLWJK62WEYQuQxBH5Y/4rPM4WKGCU
AUyDG77gRvTgaFDskM4RJJcMWacXCeJ82wTBtLGAy9TRDhwaZOF9L9sayfzSg5MefiBxoQvQqN71
WAS9xac9Sty8Tq9/pIA2ONbaxoJUsyZXCgxckkSSJnLjQuH8MI37i0zpX6VQOZ+F8hOdEigJHagN
iz4D+jmxQPzrQ9eLh7/0qHTohli6Ar5RXicqUAKjnyU6OzW4jQ1K2aiG8TmL3IUb7nc1UiA2nGL3
Uw6xZ2BUHWlo45XF8WaXGL3yV5fk8alci9oSYB6nV7bsHwAPSKUa5G5lsIh52wV1RUcXD7o8Cuc0
h5W9Bdahsaeuc10I7ahSYTjR5g57OO0oZzerZoNfLftGUnpAokzfg7CQ1AGndRWz+lIyS7ERzy9q
VAviVfuYN6q2QuC5/I1it42SEg/pL3TLS8kEpJMjdpTMG7AY0Pen0xcL+P7JtJo1qVJfM4JpD6Fk
z1LMy3iVekJFLVJfwe7zxLlwRAqE3pdp2joQw4FwzSVXWzoj8jCaMMMBl0Uk2lGb22xRo4/boF/a
prvVSjZroooKay4iwV32JPKVVkbeNRz1qYj+DML/b1zsrYCxysBnLyTfWpOBm8nR7HzHDs3lJRHJ
wcghln3adKXYNMJmUxMbW5BHjFnQgJJJ4V5Emmpgj0UnSFenABNi+y8UW/7cC73+oclCgxqpSjUj
lKWam5K+JOHMI1mQBCpmojxD2FMZdYhZFHUz4ZbJWHYloRXwV+64Ay8fAjXibBo/OOBDT/2NYeAv
9CxOG33O/u9+un+P24/gyZ+U9DtlqS0sEa8JJwn6GJm1D4M453HnjxxhYfBgdisnD/W4yOvIA7KD
I4bIboCma4sJOXxoT2mRwik523jnP6UlazvBFGO+xQnF9ZoUUi8NsAw2Z6gxU7fKU1HyeFxTzz4b
JFQy1QNG8W1rdpr8hbSYqSRSMkTEfvzmv3Wfr96jtK+0rUW7Uhjzp4a6TuWiGaoQ6d+9vFZaRPD/
QHBCTGQcVJjEE/xiKT4XZZKzCDPG3yIAJvfDG1HOzPvsQRlWhzflFLFyLr3zxcpIQaCFuT6JrHBm
neDCxbiJJwV6shCVZn9+KYemxF24Yd+oVuJvZD5whwtniMTcaFIQ/swWjnk7Rn7oLBszMHXUe5UC
sEt5xKKFyjy3UZuHycA/owJBTvvzl5QtUjNMv0EkJbtFkMpDyDSjb/C4RNmsuvkTow5h3hWHV0Vs
UnfhaCNlZhW3hACAB6+SggpWLXByicbRIOqLDVA2OApaxlpBVOATEwQfhHSNe80dHYi2OKHaNy6z
6JL8ribeyTFkdCpH2JPqN98BdW4/vWNDEG1b9UC8+jshhGHfHr45fbr+lGPAglZZsE27zmEhitff
aapoBxCmugSxI4iUlL8pxVTogleau7dLupwXj0KrholxPOzezv5Rfxr6qVvCUL6zVPStE3idYjzg
IkPJgnKrr9L8JJBkXQD0PCaPpraXHmcPeDMsAExHNoDKFC0rkAYTUKCV9X+PKN04cRuvXgtYA9ov
sdO43+4qgz8c/vqn8q9yVjlGaUqSNdsld4+qJU7wgyCBN0IbC+afHIrdKsmF7ZGJ6ysEZuQqVeA8
inO9TtVh7f5LFj7Ymo3np83Uzl7g99l0/fhbFLruGDIF8dUgFnok0igbyQcb5cdMhpRgCwNxt6g3
0+c2X0XPO1EZQptYJiL54M8pbT/S9qNwmWYUAYW69YShtBGgnSgdQHMIoNw0DVptjrSM62YmRlV4
XCr9QYkDMdnjXaFpOAIPgZcdWw3iiMKk6ForZ4bFuUJkiRJJpoTQZDF4k4dGWqkcc4Zmq/hfpSHj
lw3v8JE3RY7qqyOXlR4qYlyC6N0W+wKvgo7MpZAl+gSPTaR8Lmj67B3wzPapdqvfl8ZsRxswWp6m
ZtwGSBiBQf/EaMjyTn4U2UMHnf8HB1le7mqhxB7KNr2k5AqL91Bvg8yG9J9syUPaEqXhbiBeNK/j
IhxOfvfjtmtVZ2Hk9buvWmCgGb4UibOy4KZMjSpKE4Hb6CMaL07BSht5DxbRtO+Se8p/p7+RjZT5
vg++1BUM0boWMieIXkUvr6DHGjMMRoExQZPQ/vu2NZPofC5hXgznoNbT/zVhs76E9f1EtnTzh75R
YIcL7UUjSQsekrfJ58ZBTJZfeyMPxP0MFF+bNy9TRsekQe/1GoyW7M0R0VXa23yEa+T+/ZGlBbXL
b21g8A0NxzwOZArIx/XgJs4MjtxkBeRlorK0li19yNgI5f2zzd7Y+mGhuCuSql064960tkVqOml6
dSeScy5a39om4R683YhRrc7F0l/1cyckH79PVY/OWdSdBEDLF1T5MJkkqYUHuCbaiIyQxDI6FzPD
ovAKaYWMp1fTgG/vM8HHrRF1w8itQpcF9HY8GFygLE6O58f/HxmE/9iqmJ+TD2VO9DUDlX7S91li
+oa9YS/AdM9zJ3TOpXe90GgU4XUAHT1/Il1TZRYGQUixRcLY+k/Gw5G40fq7iFiFs3044Nh8YCQM
ymXSpGuIUNjFlC/MiR3uX+iGXLfUwjRcxyl7wpBJ1tEVbN5m4YnPjty/jwRUZ2QqHaHE3/AR/pnd
i+O5z6Z5ED1p3uP3yXKuDJ7zdOb83cAXpRyO873LHsOs+24p9ZAGLe/nsQBRSTToE+ujulzwT+vh
QI2Fjp3P/iQyj3Q7FdSxH4GmVlFyEZvgS/lSF9pnYKHkcaaF0cLlvMuLr8qV28C0En/iiIqEkgZV
D8z23ed3w6XrbLN8YK+XU+MGbfjZhyUaBDcFqSna1kuYrojt1EzgjtQlwyZ8cWTR4AfJV/SNhcLl
J/G0f6pVjrrKhF8iZkThS7dJ1qoryf9aYvWG+FBEA5Gi4VIFpSQ2wKZvrpLtDSe+BJgUouSIUPxl
dEG7rLRUbXlzMFDOD23GUAQ3WLdnpLdFuH/XBiks4VLY0ubB+9H61Tirsovy9PDjtnn4aszOGWCX
rDnVhyomATowmdJYo+wO2fhkSrl5U4ljYJGSPPllUWAEHDiGhPBrCZEsc2Axcip+u3l5S74gn+Jd
cq6XMJDdc7jVoJ3YSb5rdkffLCcdxxv0Z0EAtfI5jJx/Radhw2zursWeM6xhw8VMhkgQlzd3EN1H
3SGhb68pxQrdSBxbADICIs/vhCRFk0uZVCU2wbz+E9hT9dIW9driDaQPDQPghI1SW0XFjAO3xc1E
zWiFLGm2N27n43mD1bOpewjAa0ArMa7jzt/QHdsQkRvnuxfyq7gNTpJ/Wn/W+xRPu6HJ4ukFZgKt
RSQC7evaqWT4d0MRRmsIKAxdZblkSlC2ECvGQyL4IzHgE1bXRThb/WPmIzmBv6YK4FecnAkea1uR
l0klBgqjpF1XUD8wsG/BzvSQH9udJer8AdOaR7kpCAZkCicsko7fC7UiSSK56NhzyCliyPFu7duO
tHB28q6gHJMNdQoWEh4PUwvxPmbBkLwYxx6qvpytBdgD2soxrOeRDAKPEhYX9d2JrCedo9JBcD5U
OmDzl8mtln2WW1XzofVhTcDk2MWnRK/pUn/6GMn92gTa19vVjWxN8ijbr5ICX4tKwOykCY2zPAJx
rLOQDm9av/1Q2tt04/hIRiYrTfQmeONLW/fpUzPRdxUR6sXq1X6XOjwFskak7nSVy67Yvr99LUhJ
VDjiMizMadLfe8sbonBMifEDRC7TXlwG2rWmw3sCaD+tUOMt7gMy1DeTJJSkH4Dvtz/5GehYgICw
x1afvqL+WIuu9OctjCWZbwXF+7SGDms+M4iq9leMNvH4HGTrRRsoxJQuBRAdD7exI1Kf5YiiKu0x
s76wFKqWLPfRSNYwrDFgb6ACpsLPibzUoOhqle+6IuokuaV1mhFQyUORxEuMnlPZHrk5vo/R2FrZ
heGyeWaBBc282TerBX/aMvFDJYb8gLpJ2BtHI8Z2uKlDGJ9x0fcS7BwcUKKG2y+t29pyl+T5ioBC
ZqIPd9fSPAHTBUZde6uBBiv2oL8a9SKP6nWvc+Uwlpq8l2cjD4ulY/Y+pdduCDwvPhFo0eUvufkN
6NJyue3f/iR/KR4Z65Tv9duJLddvt7HJnBV8anGYx+ciPeOFIrAL+74M9xHv4dKhXK/BZlDUU2g4
KPShaa7ceEekgHImlxEsdY7D5jYzGLLhRWW3ZH/KjoNmehWGXzDXeHEfi1d/mdg3ZIS4niND3tvp
HYbnFb9JUHFNuCv4IJbTGvNpgnY64KoRx8a9gcWdWn8hm8WUfPH+vnxDZeG/s/62Jl7kZb/Lp2qa
sK0S4vyhJlBnDJz+QYoVRbuHK4kMZ8oh9KuzOOFTYQouJ/45mEJZwLZ5cX2okNwTU/XYH+7bCkra
8Vl9RqW/yWtNG3GaWp8a/azSPMQJgAgPy7SDE5CERW2JnRe75XdM8vjnqpp1fNqyyJNWnN5S2UBj
k9Lfg0/owXXYRM13rQPRFHkJvPg+h7r/UATCd6Q0/X/bUswQYa2s571w+pMVbdTzuHCnadd11bkO
DIWyvx8JLiaEZQggAJebPqE0+RhwskPSrBfOzUvLuDa9X9OGKYNtkecXMcmmzq0Kvamto7jp+2uQ
F+v4pKqqBxdCkk4RySNyQ49WU501ZPJSgYn+h4QakDlgcTNy1rlhSofWwsVrEcA+GZT6H0dvrrCM
tMHFszq9blIfSV6vEjL7nkuAgSyvoFs9/8eAI2xyZFi/LqkwDBGYNQuLz0Xvh9IWVZAKppbASqaC
8zfYm9LobBZUY9yb9HXWelcTvApn5x1BAsC6YDffri1mvWJlChyuV67lTgkOUWQ0RkY3XaxxXPF3
tXxMwaFpePNLc5hlfABclBQWLidO08I3mg1tapBTxzqNYvZt38HaZW/yDfqmolsNtQcUy0bI/qKI
uvDiU8nQuYmiMe8Ycz5O92jMpO98nf6cfmMMgndlfnYHpZ0aMgQWPxkn8c3nsO3bmG2ovv6YRy2J
eBNLpaR+ETnFselaUqxMoXaLVlnVGxgFH9MNVT85R92l5wtEHnHoo3uyFq+muVvgVgMPJu1ZF+um
kQ61MFxD2MYxinDqA5I+2+YeKPzZ4q5Nc6sMFNT1RXGidOwdaA1VB881Yrsq8UO0Lh7nlg+l+Vj1
DZQnS1vxfoP1f8z3ZXGKw3Xm4LXWd47Q9pEvFmJWFQb7++KaYKOZ801bXXl1zU4PvIjFB1fRgTOo
mXy6DdBHpSxLHVLB1zJLBAfR0mK0NOQ5WFSPGjYuGlW+kzcqTpJ2gQNHDSFVmZWY5jESk7phrcbF
hcyXoqFEBtiulTa7hCrFxJzjUEyTSVH50dZP3vV97v3LvPlWfRYso/ts6nj6kpVOqyMlmkEgD+Pc
V0vNcdZ+jnwB0pGztOVZT/yxMuBtnfEIgir9hQKndSW7igbYKarupmavaCo/jm2tBr8YUuEQ2bKi
lDSw6RpapyCAbX6dRPvlzT5aPPMnX3ia+dvl9rzxgkvfMF2a254eGx+Wt6UaXhzZHiu1Rvq9xH6g
o0PRBZCpq0HWScmVFpGHEEmacUWQdk+GI8VfHE9DxKQ5nDHkCDrWTvVsseV25Yf6nkiTr8EzS/jA
5T8aZyfs87ZCE/l2S5D/x9jczFAncTGseS8MYlEl2RQVz4XIvbTWTnmFfjuk86XC3HTmM4eSiKFG
AePkIo7KlaTOFRyMgcblbmK4v0rzF8y2kKsK4S+Vs+0zoNODb8il+p31BANUyPD/LQH+fuyTgsWo
qs6fYrWjtr2IaVCyAQCMJYdnCOcpCw8wuouolbHNeJGT1b97B8MDnlrZqr+8/fQg3/Uk18+3fjOe
bRBwU9wl48TeoAQN0q4Irc5GnpBfPamcoacVtJCE6ZUP5D/qe4nsFAb8lQB2U/5K7bOUA1HXa+d3
9z8mC2bMilbQqrwPW5hcCdoOt2mu/mFY31mrnV+DyKpmWOWfY5GOPiSpZZrDF7dpySR1sIvivUk6
pfb/7iSXgT9jPt8POcz8Jc6xzLS7aDCpcFCA+Z45i6LQjFPa3fIwVtU9JDDInqYqqtlifn14bVpl
AM/sfFEudAaW9gj7/izSL42xn8M/7WkHglXpDbrQU0xGjMGcavLNiQSuh35dqj8AbZpZsUT4Y16s
UZ+kUkfj3Hfet+BqzoCg29H4qcDKaLyTR18zVVh25JSrcbMpUxq8voP7DnXQv/nflqtTYwe/Mqzn
FjqaemdVVtTqpKwUJ8EcKBZbzhpAASdHvDj1CGbTK3UN7vrlW7uoJoiq6nQUPBODvHxnWRT0cSa8
DTQUjgEONWto7ZolBvnb2XzqGN4Y8ILZasgxJlPgQWGUaFJ7xUU6CD9257uHP/rwhCuO56PUX8T8
hXCbVNrZLNmjveZoi9+56cLzzGkz2tNS9LfkGlVWYAOIqu8iYorTnx8WJTpT4tfk5fETUTWvknBs
+wWmZXVi1PEZ3/+dMAJ7ze1OPH1/Pdnj5Gly9SgeS0gHEq5hVfbR1cWQzPwVfTHTm4H31wvTEKjO
fUn3yVkceM2JLuqYtCzWkgFeNkwSKGnoXHqClfQZZlkfp/mRpyTOGKiY5r0d+jruBDFpYsNoL2rH
tWChVTfaSVQBpMOnEr2SqB2ue8irY7TkKt3MWxrXdaHEUk1N45Kso/aPQJtkQjlAyg1jU3o2xDMm
APYqYX/ow1pqtyR1ntS52oVFvhpCpuNVJUYNA9Tc2TeUbU+ADZqXxakg2EKa/JhEPSa9dARkJtQ3
wH+nUDPxU2DNQc5E1xHvURKqOxlI8FE7yIOns28omyF4NARq2EBDcfEI4IiOku+htipleUVfHOxY
PQgCwtDc8qswWz33vQOxoN0FYGGsYo/4i0gY89WavnIfX7Ge17S4JEp9KtyZ7sh8+npJ6b0kUJfW
yzizXr5UgKjTZPscfO7gsfIssGV489WIhVR1e0jiMRrw3hdbTmCWoabNxboHEp2ghK6MESPbJOek
lQV/8T2awiFLg8Fhjpbm/u/weeB4xz7zWv79jArxZ96BrwGq5dxuSCpU+JzvhtWz7Qb1lHD7SF0h
c3Ch6d1f8kap83mJU8cFuZ38NV+kUezul6mvPgAfgly2CpbOMSelLG2E52rrdWRfIqH2CZ1ULAUn
7+Bm1bTNUYImqrgps0ZvafB0OZ909jqvUoOd/wpMQ8MTpT6nCTrX34V/OrL0RokoZkQCZzaWzPe9
4751F4OFpimQ/NwotQZ4/7yP/Kxi2IwKhvfiDETejWWB6VTNQh2Rc3tZbhq+wIkWwvCDwFHwnBcY
KD0mZpM3u2/h0nk0X3gaPuN4QFazg6orYVbCT8YGGCH9qvLeKhDP11YrhBEfUAbO9/+Mw6hs34wk
fdcBwcl+cB1DgjfmqyGbyRIwTEYFKd7y4tCea8AkAGU1U2E37ETKw6T+ZDEHbRvqjd4oHmM/Ptvq
BUcmti7a/r30by86NjIy7LaC26jWoROw9VD+gVFjfOs9KUXzE8UCagn0qbXgPcAmWmihUGr/vuNK
0P7aTGzCVn2JtdCwBRaIj8QjuQHbAd98oCWdKEGXXDBdM0zyt7mGgxStoKPV0ihjlSG7+/r+a37r
6g3cTXjyrI2e0IG61fRWtcrCHvXpQNAClCAsVKYBJB2iEErNUisPKkyRVThMH5P3h+xUJcmQiFuy
tgUxas4nwJXgFlgxjf4LQNedcghZsh1s9G5uIyzOnW/IW50exMHi3ifuafQ8UFwvoRrJHCDEf1f8
NXew218djAnaLvwdt+/Y5tubUPx1yekb/VNMBcJQv1JCKFmHepd9pHYDALTXiLvfJ2UaR/jQ70Sq
rc4BGAFF444RlXpO3qXWF3I0kZ6sYgy32SdiRN5bPov9S/Ro5Gu0M4q8C8onOzsVZggxFieKLkqe
bqhQQxUkbDBWdk/JjwfjO2L8bJj9/gImJXML4UDROFt1BGMTmUPVKZ+bmiIcnj/4k8GWBxjNAodu
Gjm2Wqd7ZHE7yXnyr6SNpW2lKA1W9RbaqTEKh9N0asIxu6q3mIQFJIHIqkfqknTPkq7Q7iSHyd5I
iQCTjPqiUWqUjfAcMD1cer8LflFG3ZglicQ0AAKUuDALKIvOu9TifOeCylISAU0w8Rup9K4hl8PK
n2YBvtygmwzYM2sTjU1JxjaDCTYJmMNeKz4LwpCZnYIz8nzz5mg2n/arDBnugueQmdlmQy0yvrnQ
t/xouyJoy2Fqf3HGY8U+y0trsngw4rk10+9bkYPloLsXIlTuOYdmpQx0+ZWIVgn1ciA+iek7ITgR
/q2A0X7wnAAV4jFzuU9QYj3KdfSkOASeQrGOeZxbeS4c0rwx1WtW9B88PDrbzz7THCoLeJUBS+9J
M7epNcu/apCed1OB/r9BGEcEc/NPZRwf2z62y1p88qRGxXao+LgYIYFmC7D378gA3oiIiYs7aeSE
ZtTEmrbm4giLjDw8I29XSZCDe/cXADPM2D3g2gtFQw+k4KBwAlB3LXOcTOOUio3o3BI0pV7ah3hq
2erkFUhMemaJ1PNXBj/AwV6ZiEGZXxyV8RgrR32lRuFW3HI5l+9rSxTM1KEV2p2eqW6/DckW2ykC
Wil0Vts2Zywuqh2hAaVZ2yKWbetTj4U243XHYZ3YKfZ2DRq+J6nAcOgJHKqTcJLDIunL87o3B5dC
jzt3bw7ybJez7p8khrgTk7ARubzRRvlAJg5bXLkYSqhORumFHx1RVG9umQ/xD5343O6g4XoFrqJx
cgEw7+4BDBLPc43lHv+uWa4fxOkgSqNj9StdGa9VY9YuL11X1qvkeJ64Q4TJ76kzGrC1UDQbh/R+
lx0I37F9pY7D47Bhi59gVpOcsyvvQzCdJmlJVbDnLSKpXApBAD6myencJBoBx0zkospH+Ka0GQQM
dJ1heFNfzGKYDpfhb8ichfjGKyBzix8cQvXDNJeSK+2ZrEGiDp7jf1/QlZbLzqjcsfVsm1YP5MTO
pfNJTtbUn2KBDbgWyx/RD+OBRl8NTGYHqUROntHJCnC0N0rJd1X9LBeT26c9o9JLLQ2sUTxp47HC
vyIXvdi3JP13oLMvyE8JgtUaJKuCFTUsxWHeCgV4VYzVV7Txa/Uy2mejxdd91bB2OU/BB1F5LSb3
o4W1tT75kkitNvPlZJ5CVZoWn2vkNyN83Mt75YnOPee8S6rwHE4X6e5fIerbsJt2Ovp7KiXUzO/F
XFVHIDzJcAbT7Gf3vi4Rod0U3IETvmC0F+DW2o2j8vEKB90yhl8kq5/b7jTKXLfbyCGnZvTJKxwS
4jJxr6d5gwOUknBgeFWsZDFUGSyw+MJKMYo6BmfussVpWHrYqCRloUg21LYNPW3QJPG4dlVuXRa3
5vj5RbiyHl6J8ljxxHbgprAj50l3IcZHqI/00c52SzUBxPpkOGUTAIFZOCMvV4iRcfTktUZfmF7D
rOljgzR9LFYv+odioOz4XVQPPlwH67ck/6ibKQbsEVazpuufELZw6ndHuiMdtCPUXhcDLkAr94Ze
GOUNsvBdY8DLE77JxHLzUCgPuFEumRO0pRo9q639TCsUTDAu9zqcJZ0Xiggsg4L9SbrczXxc44pw
DTRdZ5oK/i9aUPqDedQ0Df1O4y22b7hmp1RbrZkzzBWQ8pESM6AEo7ET+TzAhYDMNlylYWk9roYo
iCOeDMkzZ2FFGbwgHgBJfO6mLAN+H8c6ISwJyHvbjTqWPS/9dkeTOuPJMYxFfTJWAttiMfvmnTnE
GEs1qRgH6d3BX+RH97oMeGEZn+mhLA0H+VBe1NaQjh7zebWnOlNVFMqCIh671bq9L8x6r19afFZD
ZdXyCDeBWnQiBNz8bJSMMah9JuLuZMdFVztrOwVhtEWT0FyLiPwrtOZys8xeoMWn1lQE2EasKiap
LdQGoB3duv1jiOs08hxt5pGBBx5e/5KJG9DDukAJHccUj5m7H/iWeiiZpqotuVKnvby87alJxIBC
UfpZFEyG8GIEQ5uZEibjTiGKowxgcAEUzLZZBIsQXXV4wLZKiS3q8DCTZkuXSDn56rwvjnZomLKK
HQAMzakre07SQx4ESCmaXwMEy/Q9tWhQgN3WzAMlkPGKswbfOrvE36WNxTGgtdg0EJ2g0UI5Zb6Q
j3OBsQRIXd3MnZHAlqoTKcy3wWCGlc0DlMN3FEt7znkU23hag1aARshpn1lL3tXQaPCIAo2Zx9/K
FI52DGp37c92pETB0R1ATRGCnGolgbjW9x+/zrj+qEUOMq2QSFRT3ACpqVYLPqCmzOhpgV+WpQK5
n+RFvDDmMsBtoQE9n6sxSjDATbqjvTE6ULEcudlIM/e0K0GrPwwi+CCaminnKNDia5k46P2mSSUa
4ynZZVN3YY36VKKwTTCSPMJ5rBShx2d9SULYWHRYWiT0K3RzzmQq+hQAoXZmV5/FVGv4FzKDP2HD
xxX8j/DN+ZeMvsOAhMiFnux07upvWIJ75KhmiyXYgCRTg5qhuZoTEKz2XzqYP3+ug1vFl7WDkiV5
KAfbrlaSxfFrAAoS4jxpbtJIE2njjTkU1BVF6zVc3mRBv4Kv7WdeIwuyVBbpLorC3j1Ssvb3RD6X
KrRR/55usSmvHTKCPszK07yY713rN/K0Ah2GZzCLvTkIVrOQ73TrhDok4bv+bPjS1HYhMAw1NyDa
zVD1tOI6gL1GDaYPKv3SAkskpMoRaIRISsw06WrhkeuBqYnVul1HVO6OuDIDuCYNbco9sVpbw3dt
OQ2omWjEF0w1HJxbEkeTYHOG9AWd2KJT+LCUaLrV6+UTGwXTTA6IeHrzpIcsM73gtSzUWsJaz9Jl
TydNcIWI4upWTPRUMyUDsB6hzz1rb/TWNsVdIT+6dlaiUyB/24tFCDEb1lAwS5nBjs4cN42edq0w
UkDnZ9WH3x/5mwW4wB22+REhhaRlZ6dD+b6bFVHDsji7RaPX6KJ6YutHWsnGsKrGdn4QSTu4slKS
40794Wdilc0jkkLmKwJbdlmMHmChmc0O/SfdY7f7dHn2jOKU7FD6x5NZO7oxJuIkbaxhUlnCncc2
HtT3Bg8GPXmJ0nZc5mixOkWv6Wu98TgSuLfh/SctGrgmhhjEFjQYwZOTnvBtnNb4/cS8n9pQHJk0
W27pykYsw6Q6I7x0qXvQJqZ/ujg5BorwJMP3TsF7xoLijLqhaFtiYzOQxvmiZQpWUP5o/+mxihU5
E06/93g5++NN+vlMXpUlvcrNv0BN9bT94gnMlJAqOOdT0uw/i4jRLob72hzX8qFlyoFB3CuGeBMN
2j0hBB69IRWl23ZG+vXMUFcP5j+tFphtF4tqYL5UrfxkaK55G96+Y8+Qbbu7wLfTjvNsm3opfDC2
vo4ufj3llCKLiaMXgFVbYPkzq/PDLIcfjWN/0iUfKHgJPjxXCBS3yc5oeE1BbsviQ6L4dbqh69nt
2gfuovvh0egOZmCeHUxJrouPNW0NbpgoRWbOq61wGEqTb71dna39wdM7siFBMZ6ygPe21ZdUp3U8
lEFkx9RSDjDjKkaVSbr6Lxt/6rTCnZbEyABjpnbzug63kRBp5b5KxWK+z98PfKybhjfevu37iis6
LCa6MOwzJoNcG9OA3cpxOb5cbyzg2WTcxduzPTrv89+sFx23G0BPGvetoCxJEfVieWuOMvQ3XCg5
vfrYHnDgTghDq/yBWFxBAM1a0c4PpcLfyPYV2v3iyGVEiEJzDhWIsrJ6PPp1ZTRO1lslM1qHXtpx
rKBbR6tq+csOjJiSxR49buXrwRuT20Qa1rJXZbTjtJzW/f6ymoxHCBYwnLVjb+WN7jmldqdr6Mqn
iqQac4MCmCYSTgZTTiTNzpl1Ckiciwjnpq5u9dRHs/M9B3QtFpdKBmUksfowfgxmjgQ8oxTza8Nn
gYaLwa/H1hH+qY5fGoEPkq/mwa7j1vDSa1YnuOrV+ZMrTxw/mtQdx9+JOfw61odyD5sCX/jdE0JE
aw74yyJFDCskers3lUz9an+u+42XaudEx3alA/oY/9I1u2qMJRICNP9yXslUJ3Nt1SwgS3/u8Gdp
gD/sfqtwicF2tHdRt2haXn1b4pYOGnt9J78RNoFYPTwKaVQ5R2Z2xMvxpSPEFddqG57fYR21yezT
8N+rRJdZ2KrRqrccloFTyzuaDmMdnhr5HnfrLVVWFavAdebb6/NXu6ZX3XUHQQLNrO67J3CXmCyX
Xf9Oifqb0PDOUkSiBKXWPwqNKiWJWN7EmuG7RvTUDXBZdbpvnJLUFZDMWAPs1tdjbIe4BG3rFjby
Oaf4q2DLhv6QNsiEF7TyI+hus+kRdIdWEKQ++1UrAbCOFiJlZQh3L4CssdiZkE4B9Bc4SSa+1gcU
s5n1eHmSJZqKFPK2WVMtaG2/FWBxbQo6JZzM/t5WiIOFEbm5gvRHg3njLseKM8EHVo0BDQ95pKP7
VciqzxFbufT1M/Pp/Le1LStpbhnj9Yoptto0dEcfcsEPiIof8TtfGcyom/33ha88R1we9CvYN16e
4As7GNSUwG8L7eY2bD0tzq7nMzvaGIGbq2uSRZeJ57dMXabyPzlgyxGF8Pk1o3T1ryGppXXQf3qU
2ttdjVQ5xpoaafvFYZo0Cqc4Jwcocr3mV5y2IslOsD5l026Oc92lK3DSaq4o5RbHA5p3s0JUG2SB
2FrrY8FA8zQIoMoqZ8N0FtC1jsJUoCZ+TXEqPam9nDedae7Aj0zlj6s9XR8RVkzOZtAW/S5k3xKb
fGC/nMponeYVT2OPqgR29n62aP5yZXR0pvCW2Tn0Aiz+VutFnlM+66szTM8bb3+E7Jhwa6oDQoeo
GeHqVdmXo75qDKWsGL/zloXAxxOrj4ge2a/WEYvUwZR//Vzq268K5NFyLrzJWLWC6ZCa31ikmKMB
rPN05MeMxTpjgOo5znAZkA8/gUSGqlyDWoa/fZlE+e6wYH/YLNzlWr0NbWdO6uclDEV+STgGWeE7
pDWQIolu4Dcc1lUbU3a/Vj7GJV74AP2ECjI/52vF2leRkRyBTCOh9qDO67Z8GRdFZyiYvZaVAaXL
OdWfgQyfILyhhKAh4+UWcC3VRbJUaKVndAHDq68UVlWS0vehAE25hjmXqmI0qUcgLAb9PR+rsMu2
tj42nXyfatQKCwuMdRpUvMus4w2CDO4FfF6qHg8qp6GOUKIgvK5qp93cuJZpM3gNuFvd/wWv6OND
s0i5K7x2ZG355v7wDaao2AVCGSv28xszGeFQNGrkPRw2LAb1FeVvO0HoJ0GF/eBnJWugS9oYc6Xx
Qj538IqOz/RxXSy16cJNd3T5Jv8zu16E7Wzo04QBujvVqqcRMfM7mehk8YgZA86Py6ayXNgghxlM
oGsIh0xU+5OSlsXArbtehd8B0r6QmnH2SSjIxna+6GH1QK1OmKBPIhYvbi1C3LJisTJd8yCY+aix
xkULp0zNnmo1Gr/PuVnfQqKJ83MOO0slyas69fEdngDs6RDbqZxgiBiNzkg3yWmhq2ReMAt9ThBz
LO2n1QuwYoE/X1MwuOJ6To5QyD0VmTESsUZNZ4TgyHpNUij0wVBwi4FDPjlzmaUowQ0zrDCxSy6A
tLozKerxBl2LH3agBwtYIMKGVEWy8T6zQ3R24yGxWBZ9mbwlhjvK/qIhp6wXVoyZQAKGfhaSfOFq
i7fCsN4N/M2cHWp8oyoDa7+nNpFFglh19ADj6e9XfFU3LT5r1n6l3VwDWCI8vcHTVqoVrxWzKqdy
2klR9/I4A/VD7v6jenYgIfB6+UNBbSDUsl4eE1L8/EA+7GgHc0p7bb0yATnC17/LamDyYUBIK0oT
BxD7cJXMU3kkzJ7BOx9Wxy/kW3iKACkIivKqaNSO6f47jq75uMAZzJ6PdrkPsaGKZIkgO85BU2Cf
D1+GNSzb6CsXe5lJz1bOFmrG4oKCVTWP36wBRrxeMbxoc6dutue/pMmQ+nwgaVv4tzGg/z0aiuZb
bNNXgZT8r2FGhLDVYnLsFEod7hjBY8pWhAuvgFtf9P/qgkG9JzvgB/10BzJRpXxGolNB4UlLEaOG
KFCd0z0Czebzh1BohwOot+/1v76HuMmTBcq0lZ2wdp8dtB1N8vvl8bXVu6vw9OQXjZnbBaWJspR8
ApM5viirwhamBDQO9gQtimWCXJEKIvxaO1NTTlrBtJQ+Cy82tOQQOa6JS8qTHmA7t1d71PZWr1S1
KodddJBxpfRxCX9Htlw9dn37W2Mf8eD3XBwOY6/TWMrhHTffgD2NSutEjMZhNxqHSlg3WsVok9wa
Iu/JxMCYlqrjlPlDcFKcGHpdkgwoHFPDIQNHmybqgu6dmDTj5u8voX8lpWL7yqiOhH8GPolXUR6G
jKbGgmFqUkQjqn7LVOAy2UAaGX5At+XUfvpkmOc/Cv5LJtQ8U872BBcBPQWjMswqFeuJ0FpngX5s
1o8tyBvpAVGWAYmi40Bo3QN3pVVWKokspuLefXEkxmZXFQLGlzyQXmfS6km+LAZmr8THyS1bvMSH
tF6X0C/Ea5qAUFxYWrQeYvC/QKxl3ropTvK7oiI0eUGOwGiEu3LPQt2QPS62wtwzxNUi77Hc+rF7
KPr4WcSuBIz0ryAkhwiKOiNbT3h9SzxDSpCFkQab3GAL9ppDimqroq1lkoLEmwP23Y4bIviLti59
3Nh7Sl3I8nf5kGm8ccrMsWpdrD/uuBOtVgrmOfOEi49+RQ1V592gUYG5vsBGNBKvqS22Ir6B/66E
Z8g/Lp0v/zI04PruBasc2ZflEIrOKSYm1JBeM8nLIKJVB5ipWEgv+Yq+YmiIhQuW6lqmt0LrOpuf
jvWDMnoX5SsSX5eWtywn/4K42wjxE2+Jeg8SPiqExrqWv+2CRbs6zLIfDoYwWzZ9IVYf9gcB7dcx
pkw2ojgMhQzu4z6RVAr3n9yA4lpuuDx6RkfPjLylXPP/ApTwU9Cz0oIC4NOEJGLt7BkSzzPwvISP
IAXjmmJPSyxL4Khlyced/w+zgQKg2WdNzhCtHBGSzcEiN6Fkd5Y9JNQEkun/RNUBM0/Y5MyTZdN5
vxCZJy7gwrdVBfu2p4lwEtITzLJFAr19K+jf558dQ83cZziCfvs8keZnH2XeiWdgL9vfJeuRrkT8
BxKJRHqDGrYNNEzTk7gZ5jdn/BeFN0zHI35INp6ztEQRTbRYKzCOZ+nofQcJnMoN8LMBN1PTkOeP
FlBsl8P5wmFhF0iXukehafcvqovUbM5z/YOKXOkfQfbHgCZ5dKAZ4AKEgBjl4u4g3PEMOlpzXJbi
zn+AYHqEpfXUWKu/XuBO1KMDmbqSPd+D7Twni/DwHqvhsJ4sxqAXY9APhO2aeI3HepjSzDA1Ivfn
iNjMJgXNhC+ctu9tOJchTaGfT15eBWxc1NkmLo0uxOVOiI7Ekn7jnnpTWC3x70wUexuNKB0JM3Yt
EUvUOAcznRiutHWj5lNiZ9y+G+XUltfTNfC72uG2pKICtRsq3O6z49MnuI3Pnns6nZWmONXLkxrB
Xq/Wf9EqjWOfttN0l4UoYGNrfcQjfTMPMy+Sb2LItql43+/w8K3YlMp6E6ZaNSTwRfqFNoqwpSJ1
GlucNdVzhtvpAb/L8Se+4KOeVUyKIPYlR+mHg8UhZ3u3FRL9tMfvskt6UWSkLfMipo2TacMXTExd
j6RGb26JgqobD4+Rh907M0DdHc2GWYOW7O2dzcWFwAJxvmUeeW1B112v50rYRQZi30G2bUUDkGqK
LwI1J9nvCRL9g/iMO0ThIj/lH1titVjChA2PQzNM+bKH9E88m/Z6W6ymrJi6g2XBRgCsZWxEBu4r
wXhC1x7swv2YANk0rLIFbQJG4VA7TX+0U9W8Y+IXgbgTEvc/I2Pg5489qd6lXj/iRtAwRO5aSgS7
+AOEBpQjaAnyBA6MnZWvgNoWrjGmBCuk99gOMsbWcuJil8dwSLGnvhxDFvg0WhgJJeaLicSYF5r7
HOYU+OnHWwPfVxLetFzshBHSLhFCw4h9JpR4b6SeZIIDRfPfKRaKLiXbTjbaFmg8wDjlmCKLvWoN
EMSHav8ctHwO08ISIpfMqTzLAHlc2O+6bxhDSyledhwsy1sFqVHAf2g4nKz8buvgTn45rNIVtcZV
EBoY0LoSIWSeCItK0pWEhoCgkysCMuXHajfTkh5l2nqnqzimwwuhSsv59EKd4O3qNXiFT/fqXvVz
Bhd+A4t/2HkAx8cfm/1vAcib5IW60R9QYi1olg69wLqijorXV1WhSYC8YLh0dDgU1mls7PZOMxki
MxKfwU+ssZJhPO5Hn8YYf7FnOyzxOmAtpu0rU6J+z8IKLZTrJ9AYrT4XpflQ1eZbC9LHDn24zhi4
zUnceJ/XysMi6PkOoRNUYAs65fhalTG433cYyhutIhsom5N+6RvzlrNP/lGb/XTVAE1dDXbGpI6S
0EtUHtSqrmdF7GrkNApXbIt82DCnl0RneQJWhHseY40Hnfj2JpCOYONARk2xo1uRTvRzuk4WcKCI
dG8PYXSd2Yt7WxcebwlIDV82jKc0h9IFRZ3lByGHc9510YG61OSOgA80CW1BI9ctfBTe8ND+x+5Z
OqO37XP9xlToyLf+SSJwi1bOQ7T7idGL/g7DSoQzlr1An1rbLwh4C4ibO0m9M/auzbk/pvMj7Lfj
hJldlVxj4jmtnDlLwXtX8sw0f/rtyaCYkptKPTOILzo4dYeA+p4XsJE5FoN1OBFm0exMR2mCnHTQ
KJ1iP45DZQA/N5vTrxEq7mnGG8cJztp1w+WRrWGnqQ1SjAgiTucU6euVpIR5y9RNBVWpUezwTneD
RXJcU9zfd/F9dif+UTSgIgqD7lHqLplg5bgksV38gbll+trFD/mrX7Tcqo4PQZo9qhY/jYBj4uIQ
12GV0ZJjazdo3wNHiZINm5h2NmcjukxQD9cOObVirPhFiSODneH5J9GRrWmdOTQEjHPrq4IvApEP
ldyksdEa5oO78coO/G9RziSJc3DVbMhI4ytqSm9eaJxFZJpc4NfLXkTLuN9Js5Q+FfwH7H8IZL0i
yG5PmAZBikOBKS7jG1yNw7N9+1QPJssMgQ3XvkdUUxmLIj+eFrVUeE7j9NQ2kOLw3jYEblQZidWd
Frvn7ZQzf3iPMwfug1ugJnXJkRC+AxOlDMKiLxUyXHZWrLuqlwCPBOI8atxF00L8gH0vNtedUsgG
ODpUMYrGTvr7DF8/vCgANMdKYR9FB0/lCTeFK9ocyXCWGseJAzLs7MDk0O3sq2KbnVG6AE6py3im
0MZku39U0tM3Iyqc2Z5Pf7152XorKgTsvwGJFtL0RoBFRWfgMVcWLdN3FqWoXWL5acMV8QZvCcpL
OFQRzTTlIJbUWZQnh0F2ZOMLJa1Ww9KXJ6kq3VZhjuGAHTOHadymktkyDbYhdL2XjEf7FhLkWYVg
Oy2e4FNH5pPRRM7LXCfsrLwCEyYzS7LdPBCQSivcps35k7+GutJZ1+mCHuIXojWDI6mXHQrDdPF5
f0AjUGX8FjeyLtNrVas+wrtkrM5hUHI7Qn2w03X3ATTZp7Dn2lZwhpL/ago7IQgb53MMyNAlSvVV
3OrQ5d7/jK5oRbjVDV+C3/9GNhEe5wmYIAAqvBnGqYEAF2XUc3U2SAH8r8hfZw/YNtpyjLXa4lbN
p3s8MAsFhGirSTaHOkAORJIBi+An/9NV7DyupkuEeFR6mMBf/PK1sYSNu41UH1j9dTcoB53g35nK
huYYoCIfCaBb0yMRNKJk1Th+BpbRKVuMuLoJl2uufRq/Qzq353v6SxYKZgYPHoOd6lfnLpHutXt/
S4CvPy9N2qHAouGdMTdJ6wvpT1oOAzItl7dARQGgX1dNOI1yuWF/9hZO8kyv02+JZKSLs6hK9WGU
08OrP6IpJbHzKpY8gyKcSaWE+Rklr38T4bYQq0FsZgTEnMfONp+GQN6IEDNUj174HueP9FNzogHJ
R3mjhBagtstyEAZqwR46pXXuMMA30Me1fPycF1ezNp5OGDWKoIjbuSwg83hPws9Mwfi2G7Q6c0wc
46Gl5+4XI3FVKnmWUgaU7FuAlMg/W8hGimpJCX3VKe1DuZOWIrQgTZ9tmzvsaOxjKDReh9qOTuWB
jah5sSsCa8RBQnd4NaCPmFXAcgm3F6v3KJjSYiKrnZdzjqI6v7TAax5CfKAJODFNeLrseQ5Y/ZZh
irUiO3fOY5XFTFngiNNlbCPYbbxFDIDpecxpZrMwL1AoTb1T0Jwc03zGPUkrQiXdEApzWBR9qA5U
onw40M+TbsRJ/fTgdCR0BcmTsdnnHqsGZ4Jasaw/TmDL7cQ1X0wnV5+71OF26QKq0QIM9Z7k7tpJ
/DITF/dUBrhhW1aYX9webUOmslfs5wn+d9anDKP5aOTFI/HX4iWjFKYvjKJPg3S4eK8R0qtv1yQ0
hFfeAQkkQrXsgS8CeVMvq1rInVCzHnIgkUAsQOW1XAbwzrM6owQmfeSWS9EmG1B9uvQvI/8BlM7D
4s9EFVL9dA+c4sCGarVaCiqnkU2z9Z/BwSuZDh/ySz2nmL4Y1iOblyua5ALApmAXPBGEh3ZskKUg
yhGUYVG96TOw+kVfrz/m1V9XoZ1xH81l1+bEQ0b8S5rtfgokteCSgDfaegjGxCbMzYQysj5SeTDa
l7NM8TVUjXJ7QjBGwBPl8yW04mms9shqE1juXEhDfb8sKPElzfCjdXdB0oLtQjzpxsNMsn02sU/4
sUtopuoyDmE4XHCjbPXvEDqHuzGtEBQo3ICi99eNLH31qHhIrZB9sDPHFtadyR+Zr2j23C3XpQ6H
7z2JkOpzU3mr3r6KdwKxAgtc1YhcVBCIjlm0b+/sSEdAvGectewVxrWukKggHEIwEfOrkZA31B+p
Rvzwr1xp7W1lzvEmU3hOLNY7n7OEAqkAm9L9UdFIjOD+PD5MESOrER3PRSDX8MFP4rS19YpbQnhV
EkeWiyOMT4wFOB1aKffVrVGc+nLop5D3pRlrNz7LODevF1W9uJUkVai6DoHFF6AHmVJNI5zu8VB2
vvJ7tSEABuE7/wQVNwSybSPTiyTb92TvdIS7XdVPuWH2+8oQ6yOYxajQG4J3yhJTBQ03II5Sjwcc
HRA6RU2JVcX/CkaINnlRaRo7lBPEgYLZC7E4tzrkyM4szFRGB5GGYcKjf82wScCqGk27SegqRK6U
6/4tVaULv2FduPRhiVqhi1/qXrtsmhvCrLVtJkqbsfJxKSt/Uzq+kTzHfLCEJan4M/1JEgDabBRq
Ip6/x5OjenYxLaP2B3bjDAm31xRIjczaxXNiZod6oFavQroM3Kv2y2hIZIVu9p2pFusm44ft2vXJ
8+j0FZhrpai3TecGy80uvAikIntoKdgnQUz7BQAXB/f8Wg6hVurOmnB6MY8NbstqrdICjN1tBhvY
MCR6DDGBgpQATXUYK4Z5+4tsezAauiknYkvNYwXjCIcE1s9be3l7nZjtDLBwbWlOF5Rz8LTGWNNs
tPn1Q43JD1iQz28zxHnWONQrwd/+GIhMm942aaO3AgzPjPKuUMWB7sEcZFOgttuUiJ1QidWl7cLv
3XQ5VW4TUuJYFSBRJxTj8Ifv2AMmtCJq4fJ1N1PEPQ6Wd/WitHOilXwXH98Zr8BprEzpcuVQe4Gy
KGwGxSL9uNWe5FXj5ESOGTmT4NY5rrqerblxpWKs2oAo+ngG1UixO3oQS0gZupoup/3RXt34j/YV
T+WDYWO9gYGMWxrGJY7U2LuvDwHF1qCGk3pUeIIQ99XYxv1NaZM/8VemF/xhIrBV0BkD2hH0wRVB
bllNULiaiKEg0HWRImjI1fQzwiJN5feZ6dlMZxICy46HQ6cizq9DHBlJuYC/oCWaFsuhcn6LncHK
Ga5Tp1XMoYNlBfQQK+WLC1AUxqVxvnq+SQASJh4qyUz44KBf3rIdDwqR7aLjg4B5MeSvsTS/U0W7
ovJSithsXItdBChCmDhL8aRmdOyX2tXl9loe9bYq5JYjcYQ1iwcWRVV6SZ6wkrvy+JsRDGQr64CS
P4c3vIDWZ86Byyh3tRRJ/tB9yxRIDbmECIespavmYGLoILhzW+8l/tcYDZbtDl74gjQYbpNoTygF
WEF+BXwcMWpfe2iIQBhgWaKt9BPVgG2Auahmn26usRPi5lVvDnXspIkXsCyG9Mpm2DF13PMt8cgI
PpRYhZANsqtK9vbaoBR41zr8gvm+esf6F2IO87r7p1d+9uJ4JXi4Rsdp1f4J2z3PTkJ/3Ue/B47B
H9vrtC9xluOlJQc4IP21qFVnSKtIQVZbWxncNEnWDJTLYXr39aLLqmjKHn2vqhMt2Y8gTOmwNRAb
UWC7SsGtSUxsHIxLdb8roagwaUNg30F8bz8NUxO42uuYfSMwKpTQ4l8bIuqX+yQ+2pNFvkpIfvWN
XN8qQzVUzwPjldLAGmeYhf4dOAYlLwmUwiaI/j+PSm1vdXB6HfjGR/tYG9VqT+c5PepWBdzp0Eo9
4g0X/RW92ZETd+OhWIFHPt2FZgNrpFj+YcodLyqAU6wRkAP8yLhdNqGcYKkkLPPzU+wctfe9GeV3
6g3yGPUvyBTV+XIU1ZT/SUkjOGr4ldh6yzwxYU66K1cxglNZQHVGuOaoJaW0g3ZhU2UVv6Q5e7U5
5HwpFSn+R4UiIm0cUzPMkxDnifnFBR71IlZIcWwldYZlHeOvEybvm+h3SiHJ2tQu6p5DDeFt2DX3
sbD7ADWZoFvqeAJVZmkB3FWXDUd3Tks22h6L7kx9UUpN9hgXpI0mM2YjNTDL+SW7QEFTsx3wtEWm
xTKCnsst97OXEbnzS9FSIR6ma2qWoPII9GY3Mp7ThEnPCckJeqfaELg3nte25CeSwAPtzeP5pIH1
U5GZP/MDt2aQOPUmnl+MpUTNKi7TDAJInLGEdvtbGvM3kYpEvPsvEgS+IlURW502REPTutUZUxih
z006bysBkTeK5ul+f2OyerWoViiF0DDL+0HG8/cJmwtdIhSO0LkkBR4p3rlLt3TNSrHEcyiuaNdd
ssfcISgq5+eluDCFrMElpwVTdQiqU8netkGuHhzeZdQjc7utN+kWPIS2mSkh1zNTILs3xOH2EAR8
DsTV8L5mUFHKunN6ruRd4Tmh4btA0heJrW2K/veYdftLQZfBbFLccJyYHujY7CME4+4epqjzF47V
lQd9pkkTFSpY2du44/kwo3VFaz2UySA7h1hByz4dbHBhMkY0OZhPXCqU8YkVC02+yHa50K4n5DVl
jN7OsukzmhZy1mpBlg2iCbIt7pR4jpYw5yRWyfrBq77PmyhINibw6751vCjF65PbLJgD4yCj8kE4
DYeYuvsGJv/joI7aOSAEekb55kV4oPavf3SJ8SclIK8xCgf8imTPyVsankSozDg5kzXYhj4xiZl9
OthfwY19cGdu2vBA3ortvrRhSNslLEJvJOvqF/F+AgpEj4bwficU4M7ShZxEHg2Mwa9BnFtFsRZf
dU1mo4hy6TZ3SgE8M63dHvfZBTG7y+EQ8dum3mKDuqS7TtxxCR4aQFOyFy+yFfMUPJ6vLiCilapy
vWzTaQGi5mz1JEptM3UisnLy/HFa4Kps5xWtdo3KdfGGmfzUj3AmOpqYaiCGN7noLZ3uyjEQJNu7
yp0mrI5v22eRYNH0A9wzS0uCb2S/VRLUTuuqgcPS8Z8c5BgmxXCI3GcSHnU2axio1Q77HdABi5bq
AmyM9NCUjHlJ2lST3NqnYcrZrUYc9f0FAlExElT4QXpJ42ly+B05JYVyrIKOsIpSykLR0T8o9nGI
EYtluHNhUOn3ddvpuM1+2OaNo3fp8CAy3ev+pAAgmUCLxN8iJbAAvuh7MBIbjgGkR09weDgK2tQB
pBj3okzCY8DHbHTZLOFu0DkhYQ9uFcOBff3Huwg+K1B8tCmOU2f4pcEs09uUB7lLIKTNL4jJ7gpj
Dnkf5MGUnR7UOF/LZhaJrGxpJpq0ugxC1zrfnd510Tlg5VE+ojQ6UC0cl7clV+KRfWkaZcM1TJD3
NF2UnfvmomNQ1sMfoGkqi1gYPBOliIZjcubXk03VN54tYTcKid+Zt/N4HNlNoUp2nPV7IViHTKav
SjisSwDK8a+PidOjYG0B+1NVkgKwuPrAwq1So+2/Wzx1C9UnKcW8qtw/x9rOK0tyeKYkO9ATUfdP
9FsoBTl9V+Z5qsRXB3eFfk5zcJLWQsrYOVCD9b1+MWjAv3GKQg5unIdLKKqMgBLOeNPbHWKo9Hp8
irEGcV+frIwE3ECda6SJxEmHZlZ0X3zd2vIZX4ty88r7OJ5fdL8ahWF7WQzU0HV0Kn9RkFO2lfXO
ZkuArZjmaMsuKs7c+qZAxlVVD3QdSta0W8RrYDLC5jcpHN2OhYQI+B5ia+ClBpZkEXMS56u+ckdF
ofLaJj4VQJL+5ImQ8Yz7ckgrrBS/zy9h3G3y/ceA99yXCZY2Fs4B62FnvRkw38sqi872iVZIUUu7
Lru/+0W6oNWoYioy+rP18vvpCUVygs08OZtldEOsn9h2rTnfe4Z2J9bKB8fMN8GMBUmfn8mTC2EK
mRqsFIv7A/UumhjCiZ+XY4YSW1Je/V+rzh7T8E2/F9xGzcUeO4bKrkpqkO7ubJScJiywlKYSdatS
AH4c8C83P1lplknb55j7AIKV+5ur0bUE1WbccqkAUNXm0NSWHMFl13aikBs6QQzdMWBqbPHCQa15
wvsR/Pg5eEpWquZVhQF/y+M0ySyjA75I6cPD6hJVfCkF68ERqUzFTbYXSg+paGtV4/kCprhPSokP
dkn+5PUPaV7b1JF13v16LyOh2LB0hP4QUqoJeQs6GD+5wm5O3O3EosG+L/FxXHRYni+UaJX9ll8l
0PbiKcVs5wTESm9oL9N3VDsjO7XPKhOqWjDb6Yzlt592eznVcpuYXjYNpeMpDny1U0lUbbpUEyHn
3CWApI7YKlT/byBHH7pWds/1X+6+gIkBeHs93l5ohU+7dkkaly0UPKI5gc/L/l8IeXAQA33SrVyr
WhcIs19cjVa5kMKJ1UhffcqUDTXKdvKmlg2/NQ3eR4jN2WyeMeHcH4rfsVzZEku2gJufJIRxYJfv
iR1MyJuJrijh/gZMsomp0SsCvLPhz0pAbg9Aezb1B8blRec2QuMET5LrhuIVvnEGgWAJZxOzMcrB
HqOgmJiCMDiF5o0elnjeiWQKXNX/5VCXP3WFQc/ghDYCng4NbTmyN5PjuKDwGes1Arb5P4851zzg
rpNHoLBYAZhA8zotNeOzI8D3S5hjA2KSIfvbaXN8df+cHyOHYZmdCjeTKf2g++Osvhj+zZ8oR7XC
sZbP1dwW7cuDz/aU+W74a/osmTocuRERlgo6u9baoUgbYVJtuEssP18kQrnuMkiord7NG8GgUtL1
e34OdVwfH6AI5uxY9vALudmr453PKHC5IDqECh1YmYGYtPka3IeQKNWVhHTktQcYZs0F5BGF8/4T
shrJgPazUCJcq49Ltyx9AyW+MPeitLo4Zvfo1Z+dsaAYNnYzP56Vt60XzDVmhgNQeUexlf90fdE3
WtMsVXdnVuqxrHrdvSSy/VHMu5M1eeUQJ6LFVOC4HFQKEQkYAA3sfzNaFVpo1w8DeNpZwS+LRn+0
oLDpWottSgcmhEygq2XZ/C6dxhAFp7QoqhEA/H7hLsvwoTke2ih1bH/QNyz9p79u3rXk+uuT+w7F
Rhb+LxzJe8GdVgDNJCPj61p7UKKV0I4ADf5bBgFp5f62aDQEJf2eEI8LhJgfvz66tMu8UH1akWuf
ESPrIsZms28evCA7xTv9xx/VYwi19t7UzIZCwURoxDHFq7RM1gUYq33NErRlkO5ilrn5lEeh5hGQ
dASQoGvRyaFTQOhGP61jvljrX+RqMW3UEzCXc+8CNsKD1dqpC4gHbtQod3090t+Dd1fOAjKZsLLw
me/kwxLkcvJXqpySg8xThEEaq2J8BVeJ8Ne96DRc3Xr6BVqnLEM5uqrvrR/N8wKpP9Ye+6VeWGd5
SaA3Wcq2R63G7vNMBTgF7Px4kOfc7QLHg/yGvTXLF7ZqSEjEqhX8odVgSyEnkqhf240+LjusmP5W
obsqIHjZAzvQK5dnJfOZPkT5ABcYozmz0PjNzsAFPB+WAzMlCMBWUpj5+oxLtKk80uXp1jiGScBU
A5uTvyRm77bwWGMPxTE1TnoYKQPeJGO8EWzsAsPvF18cAXvb6uDnUz/n+xkx7jTqxmVta9pBBQ76
II/RgrWC1ldppggApEiujcjR2Daak+TouBf5aNCn1sfHhoen3Mh7uP9uz7fujFHoGl9nxAvUo/Ma
DK2hco22ryJDVheQsqdnHcjytKEcYuQhkdijSboEldONAZ1rrN2Fx8N+1kCPPq8gBjYPSU2qSEDf
lEJKjDJzmUFQ3luZZQsw3iHx1DuF7GAKbrlJK55rP5HJXg5j4/SPCa5bMzitxA4YyFs/Cd1RvTuL
zHmO/u+DZYZEaFATe2ptqckL/OuxJDRlTkrudpAaKrgamkGFnfxoX2n0V1GoA9kT6CdIG/7eFLh7
JJ14o2Gm4RxVjzX62sur2zkzMZEaKpQ68eV3z6q9pk8afvy0QBwFLuAVU5kg3ElEFmC8/b+a4tSF
JrPM0W7w6NL/pzXHCPfZgFKgDR49+CFRT4tMxazIgdBTKb9W+qQERIQXyiQIw7JxyJPZwJsb6GTm
HRqoiNOcM6ZaLctggkf7VoM9YH9lfR3livd5oI2D45qxZZYkeG62ZQa4TVvGC3m7yQxGB3fzsHZq
skdNTjk/iu9HxGd/ABtj/xAQ7T/rF+7SrbwTvK5a52Pcljno923EMd46/2zluRdVBhDpr+n6M3BZ
iv9gyvIHVVBxgLmJGY3rqHjJRyHJLmU8pi0o7UXeAPLd4WU0L1652rPMO3FR29I/RmKgFkYdAhr8
SHhOCBdmP4CPACEACPjSnPO3LM/XAwRMrmUQx3K0ImQ5hfcCE6J0TGNOje6x1ssdhps/ziGxjKBD
dVaEMdX1ItzXdUUtBqg73vs+cLd2StDY5wjbTJ6t8qhtLGKxqHeKQA6Ue5xwnm+fp869gvhB7r8H
MDBW3ecXd5G6h3kjAEr3VTmHVI8VVfaUqgO3VeocSXkCVchgSV8Cz8vS3mgbFZdExlTQUvfGPCM3
VYejlYMSt1U8DbuOeeAmMzy44vO/FOCtlMcWnPjADPwap0QP5Kd6KUzTGGGqrpERqN6yES1F3Ic/
OsxEJ4QyKXYA3Hr+GpPMV1J/h90vqxeinUWYNTXBZ/t078ctfhcBweJcFHhDRgvkotLdW705KXYO
ZV5rkDM1g2I33znB8ZUaL/j/E/EWIV+Ocm3z0xV8tgxGnChIc2nfGUnf/GBGjft+dzfZFeYW7idB
9Wu8EIlVcM3SE54cvnwAvxBbbfd9N2ePDd4BbtwdNFSuEIdFMLJL/5KnUS1CIvtvjvP0oNiUkbVN
tefBfbkm9JSHdUVfPRUI/uCdOETXd/WYOZaVLnKc6ATo8T/9iQDINlksTdvjJ8Vvmgfn+LeY/xOb
xaBGSFxrJOj6KfN4/o6TsGwGE69w0+g5I25r3u17A2Y3yymVZlD+Zxpbyls3SA3Fe9sn0iypsL+X
VAp/ZCBXaLIS1l3ANqPm6pfdIdSKPGtP+VFR0nPnboLUtgogtV3LX6TJXk648c8PAhEH3RCn/NKm
uxsIWvCcfxqNYlQ5sSQoi/L5caNbANce6XysqtbIp/M+bvUCDup88xTpqowxG5CiR5rELlaDERas
17J+nI7xKgrmrSb/FWP/3/zcK5QQebZhePeQ3ZVTNd/ZZf2fDSnlIyrW1vCs+0snPSfKzfPdJO18
WbOnfiIhLFSDfqGyZ5MouQEVL5AJEgySCdVZrLU3Q6sAtz5wfs30wLMXR7xJw23xwrFAIHy5VwLH
9C/DSonwvNu3XkjN5A6IcjJPCI7I1EwfZvvioPSYx76fGrmf27U9kEX9IIgb3/IWSQBkGw8KVq1M
teC921gKjHr/D7Ot8t3VIfqzF/xfbKxwZmOdMktEci37SFiPDPVD+BUMm+77/0Qqxa8g6Te/Bk2m
or2dwTz0rNMuaNhv59a6cXmOUQYmlC1wiA4jZY0XNPLbhqKL5lPDRD/FvWcflwK6Am1LTzSmL3gM
w3XaG/RimRj44uIh7bHfF2yf8b0vZKLoBJVrDUmrzN7KzOIFVBmSkJ6epqXbDoj5xnC6k0R31B/X
y54gvRjIdJ51Uw7J559k4VuSXAdinyhrOoiiFbtaKRdMuHsuahffCpKGbnWuRVMTXncRJ7MNVFHt
ej1fuq7pCNbfOkxxrsbCl5iMuFqSkUK8WwVibXPYL9kAACrKA2TShYqGkdhlLDHdP9cX/KQ7h4rW
1XwnFmEmusRHSTSSuAcr0Gmzy/yNSl4HydwhC3bGUHfHtmIHj9r3uw6Rhjf4y9XHQTVK7xaGgqgG
6vFrKapXlNaAlqis8vVJGnJKRO6ho6yrJ5HUKJO5DeKnb9WlfPgGRepy4ThE+VTeMYJJkNwz2KRB
mFCIf4kPZyn1g0seyOADgCn6eTVitgwTEcOs6D8RhYTqyL5v5zg5o6T71KR2pdleMY65lkiI4JyF
kadGB/yZ7TXa5miUGqPprWa+YRMOpPGXYdehE+5J4ecbcT8HuohJtAt1Henu/alimalnn9qKqkoN
wSAjwjRgyQVpqwiF6Q3OBnIJhOgP8Fcm2twWkjRivVOSdBAYsStAlBeWwlOL8aGYEo66VUhLuAdz
IAPIkWrpiGm2Zt/G/QkymYzLGJstk1tUnx+OcYK6FE+/NE/6Jn34Nfeb4v06aw8qNFHXmOq7Edgt
IKcNTZpJ2JTcE/cTMBWAUICSSPIkhfXs6arSUS8659vQIpPnu2q7FEG8x9RlI0bXvFA3mEh9oH8N
tv1zo8up9oD8llWMerweqipXTuzrcas+g2WAqryBSRZZmL1H/i/4WQuqA979Yxwm/zp3KiMBhKyC
l58/orQoWX3K592iBLV7dAqcawnQdMJffAPG4J+p8tAeL7nsKBJ2y+fMC1rI2sWyku4M/AnBHIzh
T4yGgd/Xdji/c5wgKliMQ9ssdvXJ7QRk8Dxc+zbHMXGHRuPRamU9KWPnSfe027TdlrB072E4MTji
sVxyKw1fCNcBFMVK+TCGS9KUWg1ZR8PxYE8PqEdG6kcLmBo7aSbCCF/ynKf7um4dg7FpnV6K5Ncq
d4oHS8cC1D8jDXmmFY6vOUcqLLjPtlQwbFzKRKzvcPZ16E562Qoc5Ixg4QRJPlOl5rFqJLCTlxLW
FgpyfQ8rY/sT8hduWEWBl73pbSWfGjXbkfWJxUMdiP6ZsbmMAF8tLt8EpaDsdPtWcxzXE+5yl5ds
lblGQqkranleLh6KnV26CSLZ7QCd7Gt5XXIeUfb76gDFsfSURrmrRIKD2PY3Dobg/yy4n402fat5
AYWXN0q5VmUwRzjctw7SefcaidzE7S78L5uohGIRCMQSJucwAsyW2AS7f0WOoaRXAFQvkqOpuk7F
Sa0JKsHhZIblmXxfNuLV/lMwsK0R26nx+MQsT6WT9xVyXvV2W0JQCFMYK9gWJDGdqDuEAvunZ9NT
0jE37Nru3IAsoP9sO0AQkr1ccCzhSxTRuXOPj8NCvcPWnIxfHLCk/60mr7wPWkjt8bllxqwL4CZ+
D/3YgfZ1l5Z5LHkUSoGvukf1DsLNFkXcTOKWsdqdZPWETb3sXeCuawr8yJIZ4TJPbm58bsR1wkbg
T7HR3DrsLRO+PCOvxBG2rUUPe9kG8BNMKVVQLAXkQ6AKBPcdCh4OvZgs6qfwK9xXhwlYmb38QmnR
+/mdMheGNl4TAHr+aItmH6Ler99lAyG3KKGyJsvxD5Y/r9iKzhYjzVyHKlg+H3kqraHh0uQJlK1k
ZqTTQbJDu0/Vn1T8F1l/j0gwi1emW8owUy4oi+9vypIhuei/Rl5Fuyuv/3CfBgAJC2K+nhLH5Z2b
oH1MPFov63Hl+QdTZuPWY+SN0DgMvGc/Bpy18tBj8vvIKBPtEX+JlcY2z/FCLL7rprzdmJcHyGSe
ngDnsrzfiZadbxnEYuvn3HdFCwZoUKwsD9wi/j28eOkBqggBjFQG1/6kWx4cRiFURLWivoyEa5j6
ltSGD4po4Z6+1WFZ2PrsKoWyo+KfAJ4PeDwKPTtu+U0L+GTWS11aJte7cQE8pgR4Zi7/14U3JavU
rHhxw3wUXZld+GRzzvMsMWdzPj9epz/r54qSnvKgkRWCg8/Fklk0NhR5I7RpdbFra7s2fiTIdsMW
7G7rYN1ylWdaHjEwvoaQAZ/6diM0LrqIKNYkcdV2LYFKXKqTwAtjOukS1oYNz4PK61XaKhznBqA1
LcsOqYU5fGy0H561fE/Oj3Sfhn8HIkuIFoCtFG2rzHcXyvNByXYazyAdQ7dEK5xTtK65ZZ5KWvPZ
qZgZdLhdsQpcXasAEl9VuFweWazFaQ2y/PNndaOsyMKhVsF3nZAWNAJxzplqATiuKG13lsqx/ezo
ehmkQLYzKpjjcz71abxpu5y9ccsjUc2n1baMoabi0QMfoRvepfoaT810dJPbx963MZMK+o6OPAd4
gspSOPo5+pkjWMBPrtzZgDAnhKG76TD8nCVil7N2gNVWq/bLn0ECXgEqkUbWysZKfjRof0RsWICX
Bt04Ed405pHJxFwxdUTnfvqF6hRBPPNSRHrKHanCm9B3fbdN+BbztbR6m8hg6lFR9N+KKJhyCbKc
4RQtooZiSpyI5YbFLAZwH4RyebbRXKhJ0IzJduH11IIgte87/BKUiCgzKfQss+2tw/S8Y8m0GR/4
vW7iqu+cTGJ/XZpz3VHQxrMe0QFKQgPXQIFwy4or1oCxzhcD/79+JHNI9wvQRqesTWMCsJsHlBxw
A1DGZ0/y083D/HQdrbR9ar1vIjzKrI2i9e4aIMg04u/SLBCD9ZhfDk98qbKxnEO3Wee8gvmoOn6w
8T1TJAkNLkXi7dxMrLYSnG8KUampJ6ihblMRsG2eiz/Q7yZuofMLdfOfnW4fVY63KhB9OUD+OjgX
+TOGoTRkJ7ClnVU0A6Ga0Vfo/kyvkB3NLOXTKHHHHHGrMsICPsrVB1QPieusTW1gjVnQZLZeEGCz
iM6NMSN25qMiRIpEBPOT05ME+U3mpGgmO4SK8VGaBDPrVp/irlEGPhG8UFULpISPD1DESxZVniSf
MCImHdDu8at5fzlC+u+GAzbvPLTlIoa3brPMUPOYCwKVVELXyrBqmiTUMY6YI49bk97xpNu4a8KR
9Nf1shg2zuK7SHGbvHV0ljPtb/49hwG2e2Rznz5vARuQm7bogBVloAUaaRXVHvlGVrwY3vVWlpeW
n7g6ybuB020UCoqBgk0ry9qVxYLxWAMUP289n1BLkuG/VGXyWGhbzKm//0NF++xJWMHqTP4nGJ08
9qC/Su7gYftKbB1RbsWEfev+NCTqA4+3h7CrLqRpJJL1A+Te+lx/i00UoDRVys7q8NifxzJ3RO40
P89HDnLq9uET70AxdvKqK0TOHF9YQ8Q3k1cq3Q1rUpNRjfdd4iD53AiUO0P46u0/VDr4hJDtWvyP
SVugfBhAfu7wrX3o3fEvnWm5NXOvIIV0uyJQ26vv9rwwiBBHxIsutvi3g2TbKVzISuECKM7qCCoN
FB+CQC1zkA2h9ap0RgajkS2fLFoqsFQ1Ad19Ket81scBGUX70ekWKEukuqCMOhojXouJQYs6eY7k
hUL/JthVvtHOxC6xVI4YTEEKunEpwW0bO599uWaFaGfc5NuNYS7btVM+BidvlqJZ6sa2Fe7frhhk
OsuS/J15T5/Qf6AQRu+uAHFGgoERkXD1I3ewSisCfly3KEOgumuZc/4teCjdN0F9myZgVX8jvGq2
DZRFkHVb8lZEGVh/iI3AnNmMkLTxfJcseQ3wzILeUmnvYcrllmqMmTaWCDnU7CodLUBz+zPPwqlb
LjMJAY44Nhq5JG1VFn4LEuIQ5aMM6KAtsIk5IXnNMH2s/SfCATQAm/eEuKseAIMuB5j/doQo10lD
wtQ8RbS9OTh3nsa0QvuMTsutr1HhFKWgeA6ZFr8rb2Q3td18KhVgX+/AeqpJ+sTYv5gP6xBCjeJy
jkvxi9r7ZXa+2OrEB8UBqznKZoWpJ3bAlUwRpjISlHgNTAB0NDK7FGV9Abt7XtoDKa/VOPApRgf6
saLt7RbFc3oYDEOA6NR9nGdZIFCjdfXg8n+F+JB0DTIX4RWD3Vku6E0uwbPPon+HVOWV/HbRguUC
CidlKu4TkuOvrzH56DTKVBh7YZjlsiRem2yp42ty3Hra6bIWHIyVQGqADQ8d0jlqxp+jTF+WbMjd
XR0WR8T9fwdqta7frnjkon80O7uJKrYG04dLxe606FMLgayrLddHxF1HqzwXiK81GmrBOOTNHlHC
Q2lbq075mCC0mcX+HyBcNsc6mcwfGQqv5bAttnPsNAJ6/kQkCNi2H2FLDbAFaTxfaKTljPPzwBrH
p/pnUk2DMWDnUUz1EKlxfbpj8IVzxQCMBH15prseONoDEi8VZP0bn0ctsDhzOoWUt5XhnYTLDAsa
RQYoM6F8aRVuCEMV/25tugHyXu+h+lb3sOqhYn/bfrORWNJgKvfdbNB3/6TmoeTr0UKuazwoYr5V
056ibiCeTf881gDcOHr0OFBAD6AVDBEoiuo5k7xAVKeXPjrmEyrJcshKUFC1OKTQzealpK+EoYxj
1xnjo/0EjyB4NCTLMWNaZroM85+SmZdqwm04/MT57iNPh9Pvt3ON5671lBOk7lWxu24VU7nLI8iI
cpsI98sDR9NtgVp5vA6ik7FEG1CDIUYc1Mr12zsCLhYFwHPutB4ZngWnByAiziLrTide2pZD/v/i
tW5syTb29nSjmqQFnCzWLYniP42zvIpOpBVfSqzO+2yJKjZYEA+jP4xe8MH7m/JHXSLLTjJpxvB+
kQugVKDjlQ3OJbQQPbS2am8zbEK8xlCmKzJwYgn9vb/d/xJPcd78B63rUI2UN+MTjewdft/LpptN
kELMK35JcFYg9C3coslkZdztyNTVNnaeiU8iqLSR4+yLN8HUd5b36x7nQmRpGNAYGt4wF9LPQfz3
wQ5hmvwNaTnbDXUbGwUk5/tinqvuMkMSwTcQerPG2A6yBqnskeOgtDDLrApTz8n7zzN5u7TaEU92
zMhjZbOkCfwEfgGW6iJRKzECxcbXn2i4o8eFeI7Pck+6VQ2cNMLZhUsm83u0TrMyyBa+mlUDI308
oQNJ3ELqPTEY5KjrunORFEbS0CZYIvLf0groiPuKVrTeZvXZgTsDqPP6Dcb0UrD5Oy5nljdpkiGC
LvKYWNxZ0CSy5KV1kk9bQaEsB70YnAxUx7icW+MiMJ083ISM6eQ63tOccOWo0ZKMQupJQUW45+3V
aQt7wgxotRjgH70tJ1ac5jTWFGPrOqRUwHEQ/KIPnuw/rDFeRhHCzP5H0aYO9CW/SkKNdUQVNfcE
0jEJRApxFnqn4AwnJVN48RUHsMXeQs08nUaUafzgQZFpHcIYujNc9SBKW6Pnn2gi1a47K1UBdEus
vb88J0VIJn+DV5PKv5c+JOknQohIKJ3VlchSFww9x8+OPoFGaXgdFl5/Ahfdr83ZeD8YYbzWuBSK
ltXHKrNn6PxbBp/4yIsVCqNVVfhGvSwyajN5G1fCLy8hSJdONMJO6n9qjPwXDnKajm15Nxe+EUuw
3egBDWP4QoMESB60pU1AnI4UpBnjUfNtlgRB7BKM0bXkVURALcwkXYq2Uv6PF0wNRM1nikOCNUhL
3zbLIDtXe4Pi4mpTXLJWQZ/sXieCZsy1mNYcK/WZmohVko/5hzJu5+IY0vl/uQwYlPoPeUcri0rp
1L7ZdwNI6Ff4PXr9An/dHu0XHsqzpTLhy/cwv+c88uzaH94j91wXOQ20FrAfoSbyuSd5+jghGHw7
LtgzfTlbAi4N/5Dasj5oJELWYTsrI0Li0vp0MLbQuwZnjFcAqGNSpEgB+DQx/p1gqnGtWB9B5JPv
zu/l1bRoOu0nsqLQSG0D7g+6yWDA7kCqEeahVHJqApWddrNUksQlhW7pklOeDCTzgG/UkMFEXEGj
QoMsAb8ArY1pDneZN6rAJMwafgpdzSCtCaeC71zQzeRRMUTutyguUBXpbUfEi6vsbtMrj2KPFC06
ACCi+WVyLHwQWkpEWpzX3B4mEf3D7ensMVdw8Vg7avElWRnKHycEg6tnuBtPVXJ2vn0PTCR8PNSc
k9bT+7LO5BI0d+fzTV2VDCm/VLYu5zVgNnb1RL3wJb9gl7pwqRagcxAPBJyCxKa6pPMJs8Gn9yOb
DAIv696mcxUOjMJ6pPHYtbHdAvDZa6XXSyIzmqmZXysXykIfcHlLm5JMeu/BjaLRxBsOVnTEW3kl
tbsVzyWI6Zoz5WUyMeZ6U98WTcBn2+tGwATPRoBsGnpC1yJB0aILekhZYaXAC3osaE5trzh5mrB5
tHLfTb4a3KoiebO0vxuounXJcE0H1HsbmlECqedsAVn9KJeld1CJtlVte9UPQL0EMoaJorw2jPp2
C5Kv79PNwb+Rt+g+m+JKgSkqKohEK4b8Wy1Hfh7zk/1CE1QssAHujF0P20680YY9neQMYWMIzDuR
GQ75GAYVn/qF87rp1LTcsV858mX83xUX9GF0SLwbaQw2xWQx8s0908QtSCrLHdKP8uR3lGZaF4MN
195Dn9DwonQxtyJ05Xbm1gHrFrcZrscsmpXWA4yjbz2SYurcCJq3qnQq4rDmk3CutpahPCA18uNz
YgIgZFO6hSBWJwNvSkv/eO9n2Nx5c+KK2sfP4BhH5nEI4KFpEVsXlCB6O8eRg70Dy6GbadyqsE5q
+BNTOdMgB+4zJ5960b0b/wNCfqmaCFIB3hwqDQ+HybFlqMwKfZSX1Q/cMRxvmK3usUPilm3HWzu4
LxjpNCzcshHWUrCQa20cib3yu5XuY/5AkMWLH5jWNEEJtBUKUK4NxDu8g4OKDGPcou/tb4zu9WqA
0pqixEJHqkAafh6SeoLf6PrAo/8W7C2LPOf0bu3ng7eD3DmbzmSxgUUGmUfQDQO3YFwDKOQIWAIt
XBHmLRGGX8Wj6xMOtC4Nn/azDw3kJoI3nLjVtbIS888EOgZV6m1ziC9xB2zqoij/y5J2ZHureGtw
9C7pzfJbBYtZqk20znCtK22R3TPMVtbtruBTlvpb++Ph0d/qN67IOKX9OIoIPLNzmCcOWha8/QEG
iGY2oSXPQTQevvoti+tD4KhUtVkhh1GkZhvfGhOi8RDw9tg4Sr1xLoHnFtD1QEXa0oiYG58M5i7G
bs41G5N55PTjJdVyd5kDfnVtPyD6r/KD1AbR1OCZB7skV6kyJOXEU+P+7ZQjhEcWAzcwST3HnefF
kHczue4XOT6fG4EIRr77FTIH+M+uJeJuHMGTgqAfmsNNZ0p6BwfNsmDQ/kGcUa8TJRKPyFUuBIMH
5EMmQmm2xknvljRI0JSeMxpCDL8Brxn/P6pdxS/+Fnd3B6PQkhTRhZkW56/TebNnXYehO+eSSMxa
/DJS5iNiS6rYDQY9D3gTbsUHb1mdh/u1xt2d/CU1+k1fDfmx6K+GZiJxzX2qMRqnomx/AZy7EDHI
kuniLAfJG+n6Quv/3QT/wKU5FKoq13+0Xs2Aztus1tPMqLPT1YL0VKAdocyf5SOsga3+xbbbmUfn
kKrDOUpncMxscQhUfi4uo3Sx89ObZviDnMYHZ+XoQ1kSVkkES5tnYSU2Wylsfsrb6mtvOVWK55zg
vAT+cnItPj1jxskZPibYzDqg12+b4kBD07s7tcKANRidqlodTQ7dghjpbab7JViujdsXsvz0zQkg
Nl9KlLGoBa8KY2j1Gcs3c+Biu9nxwbrrIB860Blj85WIYxj4RFXA+VtjbgFI3unIirkGdyxZAr3L
zwqp4hkZDYNb1hTzW+aac8Zf5NTWQi2h39z5xfBxf5UmsCpzPUVvFbm2daDeAo90Fq7TbGn1l1k/
kNscBMasbYH14KicinCXRS9NyrjXj5OpKAntv6s8H+q1/XQJK1VweMj4QbSXBIVmRI6+rnXyKDiQ
aspc5VN9R105Q4xWHXw+EJkhHadqQd81I3AwUWkzpN/3++F/XQKHi2krJESeMRi5SdT+CjxHabFq
C/R5a1IBkPqkIOeHuaquKQAwOTnjky28VbAy2ryyUa/3HY/PTcVvAwcBo4+V6WfD8P3yGlAv9Lg7
xPEUJ0+n8TxX4FQSWfmSmvzvH1f4CFMhqzDhLHf2sGjH2W1kp5QOy0C9bO5eH0GrRRZvm/OJPot1
uoGYSM/yPAznyL7Ytfc1OpY8HlFezz/ct6g9WWrY/FqC8iQtmV5h2g0MeEgTIu6zdnRZNmj9E9HX
NCMKJ6LNyKIyIaeOH4TrJhl/f/+G/8p1Kmnrq4MThWdkX2pH5/b2ZtAPwuLLdUIR5f8NlFP0unjp
0AVqsKQdi+6ibnxaZsVIwdtCDHKez5NRINSILoH3LiLTx4HaTupc7EPse3a7KO7YRy80K0wt7P8L
1Y8MQQswV6EhedGBpUzm8uA//4QpjOr7tbwgES6l0StYpZMXXop1RKBpSfaSGrUeZqg6rzZ4doWU
8DpovUuWefwupamr3PoHJaMFG9vsOjssRWIJ5AiNsBFqrpOKGIEIhDOBjKFXk+Dvj1dKeP0eIAj9
fpFfYHS8gk+7qGcOTANG9KXdVrZNaAzLpRJZNI4Wl0KVZ4dHS1F9zBQWSS1anRC7W3Au7mk/xw5h
UklhlKvb/+NGqqu7JMXe5VjZy6xNOI8RL/Q3mf5lHHb/+XeQC8Hn2Pt/pE8kUg25BhbiJl2KQnS4
UfgFkyaVsJ2VxGLAhG9RyCENsO+exG+/Vwxe3axKxfmoXL/qnaOSBKsiTkiEhmTp8DTCoPzkcj9i
CshoKBn42ivbw4EB1dowN4LV1AwtOhsIeZ+hzJNnVQsOl86Fpvas7QbEAfYSRZ5RLkY0ilz7kgaS
4EI6pxyLto2WZuWI8uV/OrzLbTE9J3asVm5xbTgqQJvaJoruhMcyjdoAKcukdio3H11OQLHIXE3w
PAah5AdDmwrMBNZo1yJsWQtLc4XvsHZUzoyU1ieqt0W+/4O3QORt5gbOkZWQOVUhpU/CPL6Q9HJu
JcXWEgbciI4cRcdFeCdnrgl6abObMyb5I9JoI6BitnMitHF0ffs/RjOBc9ARZj/K4zMyt8hHDAV1
r+ns+lMkneJtLMmkVa0ugwRiq+qQfELHA/TBkIGqU9oAS4V93mx2kcDg6uCVxa/sjw7ttNVZavAV
zX9wh0cOd+kObwLSjfTw9i3zgdL6jTTHqLFQqoV570i5v1uKyzZ1hZ/aqgHr8M/vujjAegz9rT+R
jb+j1H2emxEobUbop7PcBnXj+1mGY8hfEFpQSsU3oe3JxMrJ/lRvLwPoY3uIrW6nnUcdi0Qzdvvt
VpgLsryMdo/A/ydvDCUqbOiyK20cCkc0K83Lbi+ufc7/Xt/1YDjz/vENVkn2AKXjuY33CR/MK22L
Qkgfi1fS5AOseYSQ49kr0u89+mEWaM5vIE/TGU9908flBK9RO835w176RspGKN8TGcX4rY8/qJ3q
fpLKxUrRqQL9/6kTLlxc7BLPeuuaqHK4TuDRkr8VtklToQtzeL6SYEVDUhZvzB/4unOWfk9UH1T6
p0ZCldOV6IS3/P6i9mz37RUAb4T4Jf3yZ/VvgjZLHVUUw6xlfiszozVV4lSdC84fXHwiVwgeyZEt
a/w7XVuHJyKya8AchpehNuaLWMlrU4uGkyjobGVChRRKb2Ur0qxpdrl2EyxUnZfASFFjR3kxW6mS
jMTXQinQhfNkCBQuzxM4u6cBML/MlrkrRDrlDjlDvCcLMrRCrVLn20T6Y8riEBFZTrVyW8JebWhG
qd3BBVfymcZJg88CuA/yTUtUvAuPtrBl0o2D2XCRF1nuttsHzkDvRATeyBRr+uTVX2ef/vaH4YDr
KHjff+DWMT9b/2Y2YPbuFiuqb+5+NR6vqhciir+iqlmTF4lx5IHV+71k0WSHP5qLGZrWg4xFVR1r
Z0MqNu8oBmeVoxGB9lpx33YgDZjXgHCmHZgxKw4E6BGNJ4VEHaXRgXZn2z46MS31YTsSo+htdiiM
WNShC68cW+Pke20H4jCAyt3eyBh31kvQ4xJrMUQdYM7KbtEdmTUISq7StyuIB7XdcbGOo6JcGW4q
VvC5h+oRyJ2Ky85aMR4wH+JC7PIzMlSmbk1RLnAmd8fu9Gz05OrBaWo96WWOqNBDAg4L+5oAxKO8
nMKWLu32CNm8VsCR9UcLy1V/Axu/Gl1+dQdjNT827lXrBqYux/iTeqcVZFJ3dWuWMHKvoQ69ipXr
09BYVm4dRAAGFs4Qq3kcmedSnCJ4jbYtUVO1gh1hPJ1nnccQgieW38m5G7xp7KOBKTmDp6WASnKQ
q0HN0Wy3iLUvEL4R08THdVmgNWewBW2ZGy9if7Z9HxA6msX0wL1RPZDwolnEyb1rnWRAh6R44qBa
OOpsQn0oaxVwOR+VXe35TEdmRD2y+9O/xlU/Jh5yFiUxp9nwtNdjpMjrFijJDCyS0pQYEW0Cv6O7
Tw9ucEe6X2KUaVHyQnY+o/RPKoc/eK4jHXlE3MxEWNa6mRIICNAU1rkfGUfUBK+EwC1tokwqM7KI
K54F2SMbDHDEGNtDo+GlzaEG8FG7GLBag6q0TgoXnHyolJktKn/L/S6jbYY3j3oFcAY14zUWMHdk
fP/cCRc66rRcsXf4P+kxqZqKo4p1i+RX1+87dCy8UtaVPsOCa7/PqyEXIjWW29hi67f/BSFZ9Uzl
tUjZp+O4ZLUNwLZuzNwakcwr9x+lmNYjgtSJEsjl55SVz96M5DG8oSRNRU7e7xwiBnJKcw1zXwVm
xD3TzG+CWTh11Orv92KSQyUDLyVABi4Wddo4xWTDhm2EUBt/TBSJe0OMPWumXftzxvYaBKvgdb6g
3suX1AI3nzfWEGaJArv66H6rvYLomnozKR6DvNZYLeN/KjpiVcnjyhNd+joa+am7ARBITTTyTt8n
Ma0w+UnMptVO3nBOwRzK6z/t7g0XsYnVPj6Ru3Bi0WnKcYOxG6m6STbHpnneQgARbmbzETSZ68h/
0LzmPVxDcRpwU0kVamTikoXrEbZ/oujepoouaUqV8XcwV09VglKCp9TPxhz/TfasRS5Bgekss0fb
b/aKiqtGLKA7R4mGw0Ix5789bN8uR4U2JKNK1s1tBokF9larFhIhVp6JysSTt6gGQ6TF5ng7aw4T
vg7PLeHmJOUWdpGi8UyO+9XGIyQ0yJzsu0lLcW3icAL1d60lpYwmUjW3IVMjbMaF+WwWEJhGAqUp
Ybp1M3q1+CNjNFa8UFoug/fPvHyrJNfnnE+/XgH8gqhUdcH9/TA/nPTCBytPoQtyp8DXmiI52ytc
lr3fQk9qxP5taF34OOXzA4l1zKhnDA40MEGtPZoNMCOjKdmJEOqptH+EVg1He7Ce1S9IDi8S6Rvf
ayT31n7SwJpzL4EmTQGEA3l9iOaAbBGepg2eGK3O5QQ+e1oQVdQlrEe/uh3V6DPG/hrbJiBLH8+9
cF4Swf4Y0jrQ5Yiktf87U3Vvz6o51zTdgCvQJ6YxsRfOQcYFCiDgBFhzTT74V8msgZP+l5NfpjeW
cdEIhnJIT8GAkxcbMRMeNPAenLuzTpWtkCElkn275XCOgbaBnkkbSDB8v0NfFKqHfGm7Jjw4S6r9
H4qc0c/kq5zY/Wt2ur6UwXlXnOFS2jSV54FAGs48CTFUcVB/PI4efEC5sX1GSB3KoZQLpfFeUHpt
iJGTnc1wUdm24Bc2ZcAE06ikjRrj/IIkbRGidi20sSDAbM3UzDnitmYhwaPyhO7/3D7wgRS8g4yo
X4wafstAfTOYi5oYbXYcPbzWYHoj6P+Mo6cevFYV5xXfdILv/zAky9hbyF5UOsPlLPHAwsYKS3/a
xh+O+2gE+aZRy6SSwmAhuHhPdGVUplzHSFNWfuuh1+F6YV0Xcs1TV3QAjhwjsYsw7/liFJaBFaLX
R4/eQHMAGCc8Ed1DiW3OtTFTuQJTn4LAPbHaYIql1uEUvZMa0uyrfIuZxU0rqCxOameO7ulVEjFQ
X7V9hbpdSGTqHFE2BD6eFVxurCbtklSV7qFJrooWIIOQcE5foeg9C/0XF6RTdmOynPLCISKwWrkn
ysyGVHB8RoqG4b7Ugoyg4YyJbUAbhXLQeSMSgm1R8XsliB71SJx1BN91c9H7oavN63LgSIWyF2xm
PV+e5RgtWc0Aq0YGWq3Bm4nb8bmTOf2LhcuI/8f2t5DvU9RJlTD12HN9U9lOmHttrRQndluTEcJo
8N5H4XxBg+6GI/dIi7b8AhvgzSOw9IUpZpdbhCtMK2o2nU0LU5gjmWxz4FKUNKQonWtQDoluIA5I
ACKYunpecdJoSWgFKC7OEoNskH+hZwiUTHUA2YlOk/6EdXYjOzy2AUi/a0YonfkEXI7XK83NlZ2z
sIDWgU1bP/DTDgI2KKxriic0X+KEQym5Swj66PlaMsd0FtGiP22Zaqa1wObIcqr7O47DsHjJgUKM
TbVb82W6/npH9s/jWnYS76pRcX7256kJYwxZSvNRxP32Pc9WvXRhNe8AzgvPHdFKX2z6EQMx/Gq+
wds5/vEmPNup2ESTSvwE/iJjmy0BiDYSs95RMGF2Xook04ob4CMwY5xeqz76+aLDngoIa5FMsEbU
RBH+vBCdcbVWaEMFS5Dt9ioabiau5wXbSAyvpkh54Xle2PbpmmdGzu8B7WFEoRjCRua33mbdKphF
XU7xVda7PmOYtlX9hSzg7xdCCV9yuSIHPhPx9JA7EXWX2YMDzbyWSqSkFS/PdeTQFGcPDF6af310
/kvKZTUtl2EF5BKxpEw9x/L6EbMhb7yZJcOPbJ1bO/CoW4KkWvUBYCgBJ5XDWR0e7oWQ9wPhqRVJ
sB14tSRjMKhRoZ7sDRBPzRjPIvmoBIDXlHTFdvBCIf5HPWv8OAL4hldjUk/Fc3/3xFRhz9A1G4dO
LRgMdSdOTQlc7w1HIBDf5M4fQ29gHPVoFX/lpBmIiLz8UGXFmgfAMzCqTSBVJo8a3LC5SbhkGGH2
XYyAaUJ2j3gPTBHMIjZbr7fibFVsxxO/5bIVGG57mNiONXsUWpegJI4OwUaalq9GTyKfK1DynNqp
1Hkh5omK30EHoq1m+cjSj7jZREl85w0hOwR1OfAAw3SRbuBcrT1rCESRQOvVILFiqNIUGxfWs2CZ
zMR0TRdf2TgHwAn9tb67L3vlp4kR+Mk2/ahBtI/EhWe2OyGoXsDZHXBKb1YAi3qZGzhflXLF9V3Z
86P4SBM9k6o3vwJWsNSthoR/PpGCPR3iF13ubwlDMMNMtl7A8OGga6089VTa32PCfFyXH2sK8q1B
awTOj3nen+pIFQBajYCrzIJ7IWbISK2C1oADcfx4E4KJR1V2s0RhisW0cUw8EeZeCBiC58CWnlRF
b/kKGKm35mJZtl1HK857YN+MWBLguywD1++Vdqve2vHifj6UoO8Pem6QsPxvlFyel5hX58Tmadp5
ojiSUCaC1ULPnwOJ1hG38kHhPOqtFWfU/LjsYjpiUoz0nZxIvcQbM4PjzZldziM54K9zwC+fzS1n
HHELgqILx1IZe3G21hNYa/42yikiRsp+wXQP0xW0wLMDbehnu1C8104HjjnWjQbjHMgHv7x+IKb3
VhnS6W+R6OX72NFBMeCPf1f0k4THnVLjG+SHObVZxEf7ByfI7+Al55HnvjKVnoiSaj6oqZHLkHJu
2NkZ/KwUsM3QVcMc/06mFI+y0x3FJ8pbx/VqxwoSiaf3YQRWAqgK7fZ+EjRwH3l/SwKsNMHnIaR0
sBlTCBDdg5pVUaUgqbsveIN+sIySTgobAajDiO8IBrp9XuBAa4VzfANQ13aveHQSzxT70+nHqVrb
h006QENM1CYLKQGoByHy6ub30h8CQgsnphBpCnTs92Z/VlwHOjZCC2kD1u10/2Pgt4bIpwCpn2Kl
Rmto5CHkTBKacNN/4JnSDKOIsBLyhJhH8PemUbvKGn/yhN4vdNb1qEuhr7Sm8Glb26TQWIlA+ply
w6rLzf7htJnkYyfDDRjI8Zs+foxgEszt155NvM0HP9DLs0MAapV7eJ2ofXhuoYePamWvYa8jUdMf
I1UMPJU+dBjgmrqUtQTmEAIvTf4Ca7EaCBD1lnfoV2VizcqmDYeFvsZdlgmZRg93d+ttkzk93/IW
ZWRn5opCRQa4COgvSW1PQh12ta2E2TwL0jOuQCGsKBytLNeJ5i921s6raoCl+s1/GwdJnsvrMqMQ
oHfejrwyENHHOh0zfltH65qytjTKgFX+eNH4KvJuAt3qsDVfCg3QBsD2Q+qC5Aa98OSK9LLSNTv0
BCoev9OF9FNBFjuDl/TWKa6kdJHakWiWgVMlbpoJjYlLMlFQ4ALz/0bgz0gV4FeY5xtDNi6IU6br
enV/Tqx6PHBQsxEgJPeTBqjJ07pSJIYbrySdcQoNp/1ZcBrSNjWVX88JdLH86MQNMKNbmcB2tlau
6GiBVE5nkYkNDHdnK5f4sctFbP2vtxEaP1yrAe2Ejwoy21bzQp1Q6+8WOgksRIgwCt8XEA2xCNSM
LoXTTAUt3vmKuakUFJQA0WSBv6+N2DvPxfLUAnfmsH2FNGJidaDDKYmBB3Vwnnmg+/Ebq5f7FDP2
RWzw3gkvXkadQLTorbxE2ZJ/v+pLSwBeuHckc/Byxp3QOsaOdaNizuCIjEHe2PY8S39I2DgB8SUL
BVPy3s4IB34ESfJyaF0cg5rg6xumQN+QGagld56gBGmGM08u8illPXsH124GzPgVMiMUKbI2Ky+Y
c4OvZ/MjcMTynqgPr1HgA6ZVrJawXL7B4+O44eSJuzFBTOq4b8ypKu9uffRZv/ckekKqqghG+Z6D
Wa2lmBxrNq0XALYXcIo5y9aG8a0X/AXIxEsX3edvvH0v4fH4g1pzbs8POE7k3tH6HmwCwyMyROw7
OXngFOSQUt+maMjhwJzS+qtUGYPrxMtldsrmpnDQkEjsY4qpXF38vfzHtbvvtVs+H2QFoenbfbB9
74pDEdG0M5TutBADzacPkHcJr8XTk4w26vHU8WCSgMtyRGLWkP1r1m0lnLSRAGzbVyYhfSISKt0l
wCuYhzxzSluJMEQNAuCn8SPC4VcbsZunoPM2uSkYnY+pF6xQ3YKmFFz9kDFv/pumrOBbmrXQhAHR
6Qh6wbjOiwcDItyS8AHrNr5NvzaQm22Z+H832EstUnMpVw5Luzwq/XRfqVIvq8OyJqusqZyufciz
Pc8tfZlBgCJJpBIWd0Edqawkim7QQDhiLoaYYthVOk5gaEnpS84o9mDxJ+1xktwkAAya+c1AFp1w
OMNFJMBkLe4dlFx/I0W87HN8Yv1vV7uxthRdcXlxNquDeKlje+EWHIn4XJSkOvIOtWdQPJjS7yc6
eIPsxwmv88z4pyrIYwnqAEtG2bl0mPmRzHwFBdtPVfiY2m+98kdZaCq/IuUMi16yb6+0ZeRA5X8l
Fh9JQeiJV6u3o7rDU1UDhjy34COr4dh8oYWEVGiDOxKTBEcZBNluro3Lhuj1GujHcIwfdwXMB0Al
JsBc3iNMAptL1RHEDZX7KeeETv3GI0KJf4O+DEkAc3M+RNXNhljr5kpUyZWSWgOKnkyUASFBO4hz
GzUd1VHj/k5D8R0bsbL0xEribOaNaCmlbpodYI9Uh0IPwRocPYu+1auhYH1WOy8PF4i2kTBDYPvj
oW/7RlwJv+w6LIFP1nTAtNzL16CUTQjT1i89aNKxXxEOOun17jMe8ewXzrMf6lOW5tfbxJepEen/
nrLZCfEtpDyRXXrpqUypMpWtYhKWDtPvaIoKSQ/VCa81wJd+u6unKWBFm9wy36WS7HSSLNvvjClN
miJLu7GHW2zbw2Ixhua5dsruUrmvIrZsCbgubpUyv98oDu//PunpEppeXEibbeFacyTbMqK7CZpr
jdfXp+4Q7t0pw8j12/Nq8oMlQrRfkjyS8vb6l6esGA51QSvo2kolERmMAe0qe49mPuuOPUVXJYWt
OB7qw2FHAhgTFR4XMneLrqQcvV25qIy3lmlwvEwnaWxWLGM5Ux2EsxXcm2qFrHbQgt0SFwVLSCHw
A/ZouYqP2r17rWhyu6tgttjNqQ1pMItRLIvsfY51ebNMfmrxuvMjcE+MiDbjhbBLJFrMIpUgFgJu
weleh6TXx4JX7DufUvzbdRXNA6mNFA8p5BTPjtT5BXn6HACAMqaA7zSxZGqmWvFhmgWOLzFcnKBR
Stug7uKkIb4F/bSlfkOKGu6IPYb/xOYZ6TF2cSpEs99A/QYuaK2rw7gt176jVlmUedFvI4BuNqb0
IhAc+RVaQWHbtQiXiQPthTBdWuuK2fO2IYuDUNAHtJnvlvNZOcgLZt0qS+oYqANEybFY+TigiV4I
oT4wdI4QyqdNRK18moQH6lvpYcMc3x/YGWfkAyvK7xHtr4u7Ap9JJc2kDpSosv1+/RHtdZ63Qu4P
ks3fWiAMsTssiMOSNGxOEFcQUIEZcNE1D3DsGRWHpbe6hbEt/Lai/glqdLcc21SAJ14PZ5WGKpbu
RoSO342jnlo/WcHxDv7T+XKjmAuDd0xCHZJXciNAep71odBNB+bIo/B/cgvo3tD27Fi9JT8k6YMW
CNi5vQSrbYYNv4ppeWUFzQKsEPqgslAOrkmfesSe2lkRvrjVvo/FFOhRp8rghcKDk7oq5tFvb220
jod7CnciQBIaXdMhQc+AcejBz2Dwin9h6v8u6wTq9DzB6GNL8C88xqmgvrtk94W2LjiKwMtmO48J
627T9fkAb1L/VEIYBxz+XQiqkkGCmx8/BU/nPbcYxqNEWsaWAFMS8ND1qEYMELBfgIFY29Pd4W19
ytFoTk6sWGT6Kdg0vKO7TumZYgGG+p4JhvV0Za/axgowDYuZ5G2PBey4ax1kKjrmhTOfo0XA0tb/
O765P7QXiURWDN2gZvcfse58YUkpQuT2TfLBJ2g81ojKhcjzZzG+Sa6VYZr2Z1D11jrxuE6XmHO2
DENiEFCpHeidPMkqDrF3Q31YmGQknqd5FcN53nM2M7yRF83++qaylTAUhV3agZHBJggErzI4rr6M
vxLlOYosOaysrMtYDjeEF1FRitjWtBbsRpBoF00IGmhLGj1D+stVUPnbZ28Sgg6MI1kkda/jStnB
/IXYpr10kuc02oXtZauBT3arWCnjWKJ5fTeZVyQBLgfyxlW+bggeAXr/ZM/+5A9MLAd+IGQa9A+n
2p0/g90xMOYm/aZXJxhcC8a0ngBNSYgSouMwmTTTDR603+c0+9bXEVqT/b1CWiOWDeoXt7vWZArS
cBv8bp17SzDxzXtmB2ndyWrrsS0/Bb1loT49KhqtHSndLybeCVM3xFvGvKy7y83MiRrSzaWlnyay
W4jsUd3Y+0WqSB1+9hCrg+OSA+hNk1or1ekNalNEMWr+EgNty2J0aGrewP1EmJZ/ibMLpYNDXcD0
wq5PqVAUdqDIn2k24i4b/Ov82E5s2/cf4yP2MJzhFpHuw91qxKMGEVb1+EekshdZGi4ap3cPDj0L
Z7ZjDY8iYcaokoar65pAoopbTgsA0N397sfDHWJX1nY7ixcpNtCrRI+yEuBaCg3Ybvo8iOX8HjQr
SlKyvgz3Dqo4QhOSYEplpQXPOjB2QPv9EGWCYu5giM4Ikq8jI4tg20FzF/yv3+SwO9wJJ8ZhwK3e
Jt3DrMR5R3M2npSLArarY+hlvbWTvTjAkOOkoewPlKF2/vRYnOutwmt3ATi2hy2v3AeqrXdBxjkT
7yFNA2UDttns8354sF/1x213FNCSadnludoFWDdCbxYNgYcflgvixhEHV8cEjetle8pB4GzsFKAS
MK8F63yxg0eONPt7/Xpo+7lauCxIh1p7zDcGWm/wsxT8wA/eZgu144b3eXiemi9LX2uO1PhY7j5U
rem/SRgqjQYR8QoRLmnoqdhqR5LT7ZMu8bK7tR6w0GH+/RjcaeRbaHu099TL1nxXTsDd4mvTNReu
v9VK3lcHfimZnXLZn9EEFYOZouqZH0ZaujT8V+BOqZuJCqX56o205UOwX9vYPjvt2+kE7k2fbdpP
dIJNyajV1cZcjkAvr9f8Q8cHvCWgIM0CT+Had47Sfb+YlSv2Y0Z1sdbnaNMASbLrOolMcI4wp4q1
RASVOVa1DTShKC7nkEvRnG7zJWSc5u0a4VOqrHDjhdko5fWaD9XREbldQbXKsaT3chU7onD0Hjtb
Ew7vaw7OP63ATzY/6HoboPVr6aEkiPGrlx//HbOkR9/kzw4k4It/hA9/lxaxiisfRbqPrJIy1rCY
Tf+VApRAyiaplQSpw+OGiHLVzGaVgUh6sdNSuHQCz5MLKKBiJOOWYn6mppeDcT1UkGCrCxVsAKui
G0ixgrtmru07gHlGKeBy0yKxHSo/hsiWQ4zSZ2dBZ69TYD3yGFHq8E002j/R9XKIn7+4pTe59Vjh
iB3Pouo/iwteUr64YrTGmDobehFcPR5hpt5qsq/UV15fabSXkcPrQTsuWKwxBq+33OK1TqYU7b9y
uMDMUHNXOebfFw8PTy6cCcdZR9neuv9HJA9AynjCES00rsTJUEsB/mRguevaqxe084xB0itHiBZg
DwyS0LO0NPnFpJqUEaPGPjCebC7RfLNxopRe+++7lDphZzz/Bdw5AMYVJzDANKjUjQH/X4B/QoDR
kSn/T7XHK6tKO8I3snbVEjk9ELOHwoO3tf3UmIfZyoK3yoAtrQf97IxZRYGtiW/s3ggAdSKaHmJl
gmZkNgkZxIf6YQ88wytEItkSu/gawNrBEfhbvyvynD8wItQFG1M+euClYQPlOzhdMy/CVUAqLtsL
g5oxHzRrIa2M0T6XsefKwuyRPQArfk8xdb5YAn83QJyhpDJMRPi/zhQELDjq/q/nMfIhs20Rmk4h
uPZQKyIClshfa1+kzgVhDoUfowiD4J5FBN+NyRKTcBkAd2iRSOoze8W4xjoAzXJQSJo8WlHV6LKw
JWv+xxsAshI2QE8NjY9hd6OCCqSxdDmWFjLN43anEjaM+udCcp81ZdKbMuY0/Q+BFAPXJfkVJFD0
k1wY1yXNncynpt7PkvPDwcgL2aMpMqVBDnjlaf3FsQeck3P1H10suwxOokfIyKG1rLlvR9le+A77
cDldCNkkQKVCUcjlZp1T5lRlXCzx9Fok2NOqRUGgtg3/ei2zYCXtVQpg01PRwJVmQWBfCbbXGqm1
6v5zrbkVFZwX82OomJmbkyvDuhp2kOt7+i8EHx4iJtPrEDGk9eGLvjLnxFcpPFgvQkwK9kU2bvm5
BqYsr7SUtELxly8fQ1MaJpR2/W41Lz5csNON/aGA58prc272hONK90q7C2LtwDTXOG3F+IzNh9Ne
Ay5wxCfxEULYqHvgP3MB9h/BR7L/64AjKCfNKn7zxTEp/6jtatczIfy3hydQeMaoDpSy3qIrAyPL
N1Rflbv8N+JG4htfz8y5VX+cBfunJfF4gtBrdO87YMoVt8UBPpKvPRiTTfGX7ZqcT8ZmFLN4EP9t
RAXx4e+7rBrLpoijikS63UB6NTKDuc0I5qIM3jrY+oM6xZSUxifCcDGqWFutXkV4CsSgSE+/rMuw
LgDWj24/3eIoLVJG9HfFZWxupPdYDT94ELajJXUccY38AFcgL3AiBhTUZBdxiYcljhO6tSiwAEVi
54vtqLIlEC9xYVgI1wzP+VMHJhUwBdJe9+2QNoj4h33TPfDdE7YmLUR9ESYkWwRVcQH58mYBdMD4
EFidarTS/uk20RtywhXDTREzwrX8Yc/sW/5f9z9QJl+vnrivUYqezUMr5Hdb6IhCHv/HszRWX6S6
hMpopm7MayNqR4sZRa+CfFLbkbY5SKcOHZ3c4LXitnxpDx1tjOwDyoJBVgdOEKIFccHtEURqspRk
i6B3bebERs9FZlUyWUej41aiOpmGdqVewo86HTTkyDX+t3a7c9ml3tzd5y0AJ8v+11Fc2GRdYxU5
25qMheE+7TPmZm3PJNxpxBTmfBFMM+LPcnyDH2/GAR7MyDUoqacjDysamH9H+DY98gR+hUXb9Zsb
A+ssY8QFwqYzsc7QNxsKl/icous366UvPx/flL81Pz8lAqwbvB3I3xrjiWE3rPshFdSSVN/+1NKH
PBeiJKVlEPxx1TIKQwtYKrCoEL9Y5y9BGtX18hyIdI2p5jdN82LBvom54XOLNbZLiz8bEORkYDGQ
4Q5UKVn43W8elgFKv9f4LjLMyT7M9O/fI6qF40E4zhKCOLJePKcJ9kjGQw3Dv9YJdgzf1c02eg0N
HmnHOpvulh9XVpH66FOdRe7J/i3vF0FuyY0+FbZX3zKoV4jxsVYXNJ7o/hXtuDbWhTGvGZ0icCvo
Z8z+g6FRy62MG6N1U1bQY0SxAWJI9x2QQgKis5u151+KIa+nueMhjtZpTWDMWdOUX+dlmr3L7Q5h
Yb1hfR2GO0Jt2Ex9x346LAru+gR9OBVnyeYuSk2jKn0DQwrTWnbVNanLlfIiMNhBhadmWN5ZmiwT
AUnAXUiSVC8QDh1i5BPnAqqM2akp/8VQyBKVnNxCmRYo3XiUajWkdRDYZ7O1sHUO881DsZbYVHw2
2UzuJ6wZwHMps5hZ2/DvOg8JNlBscNwyF64V6NGGevd9l7rIHpDDBcC49XRSB3MquzuM2cEmAFk2
8rBPws2l8b5V4M3EqUTNGVEfgWcJnVUCHhqBouyhXy5jH8oq7ydphsBsmiQayWE5hpO0bUHr4GGc
1QyfU3F9EWZkWmrbtG0vgwwVE3yWAH9IfyJLdXZc1U4QFHpar/31l2hOmEBt8v3rFBlCfn2KOu5x
1CkuO8mCJXqQrSH+E+KvaZp3WJIKt6vBWoff/3ZDyiWnc6bDBkArINhxPHN/AMXDr43no8eABrd8
h0RcCUoFTYteebzbMVXbzYV4sf0dzB6yQ11TeuSu8H9hQQ/2tDk12yJiTHQkdtDZLzvGN3zkxd5c
1lu+zCkdOFAN6r4GZHWIJyIC5NoVDOxAn9E4KghwbJMpJV34So+uytQfYcwpk4WT4ePhlhXEcTut
rWd5dFWJ9jyhpXeZYFGghnjLw4Cd1ow/Fnj3KM0o4FOE50cRvkrI92v0sWzPdkvFSCG09Scnatuv
411KvY8uc4UTIbUwEBKThNppr8nBQkz9tkXwldSi6aTkP2ZK7wcx5v8gE/Kcc7nXqpTsSfjgTx//
K4q9eM6Zmg/9DSttukVpqj07fsbg5HuBJaB5ZkvWu7HY946wcCeKIKzp2jfKyQLgD3RnU6uH8US0
4Czs8EK/TQ8aWAnihow+X2LkZqN9POacI9kdR64UAfRcuxenQEhtvZQVwixcKoemyY82eaf3o4vA
Do9ETkEQnfruWl4oPxmgXdsMBDVEP368odvVtwVt9VwlfHGmEHI4LZManylGQ7fAa0yyzz88ZDCF
1CmOupil6SUJiBgKpi3DKnS3/X8nQUqzMuM5Y2Zrpfr9a6IZOMRjNS4w6F7pWbb16goGCFwu8RiM
LEq8cQeTlzY8AMsbD+yBLPDknh+sITOmgsBUpQaNrjgAKJnGOqTiNFD+Reh+qKiuW9uAx0c0yj8w
/gFkWV+BINTzouDexm6zLpqLZPWPgAZmdJp2e01aA4+0wNiiJQ49EVaIuz8F01GL9N0EqN+SlV3Q
lE8MGQpdJjoftJy19SLEtBtTaISFemMnrCl8Eb99lIIMLr6no78DUsHAhBHfRf3r5+19URTbvbN4
l+QtIDMsQ8lEhKrz4RPo+qcFLLGWxUDYzL5OSf4o8MGVvZyTlgfhMV7v2KGQyX7F7vVNWJC7KWTW
hNQ8mR71RaQa/UJBzr9ul9jPR5XFjbh4vt5P5RZnQPmgG+c77GPH3ncKVNaoG9SMBE+/HVxrEA/h
gt/SM1DvNDrnkLIYlNvPwc1RK8tAw/dnmozwJXhMDfqwiqyQ1R0DgjWansoh2YDPmMVWcIvYOSFl
Jp7kcfkaxFaWFf/V11qVAAybmgXwKj6Ur8LpIRFWScOWFLs8YUjou0XtCxt4DteCEPTTceCQi6YS
zUQl1LZ1FITI1UOYYEqIAh5ZHspGCtGADbZWhj1YO0jFMF1R3SEQITa90RLn1r/AIaMKfJx1Rafl
ZNJYdzRYXk4GijzJ/lScU+sBkqcaTX+I7SiZ0bgI7/pEsgehDEOCLqm6wu8itwlnKDSBcLdEU+Yr
nvY5gk3qCykubLG+XTvV5gzyLEE+jhzHUvB73o+4tNmloTHEbFDRX9kWAeaPV+Doknpfb6CErGWn
OLxHZdmC/aau6ck0h0NSuTccK6Lvhf+UG7TCHGfhc6uCwF2C+/S2CtmZGorYiePeszRpxoa4q1M0
x6Bd4sZWFjQXgYzJOj7v89/iyebBBIVs2vHRi0nJ5w2J8wJNXQF8cf9vD+vkESRDeQRZwM/Um+h1
OK6xIqozUtaGA2SjSxK+vpiNuKbWfDl9A0WIc9pl1EeA7KbkB+H6dnqVB2+bCyjerrxlzviv4WYg
zMitvSkzO+MjmYAoRtkDxX91yXzs6XKf5N6JQj+0TvjN+4Yf4bhMPxosGo9yjzTvFxiASJspZ6Kx
D/DYFjhEWDbBHiNdCWSTtB7sYxs4nox52VQiFDcQFdNo/KtiIqrrLZyXhDDZf5XdGiPTxirea4nq
sbU9895kGBoz/lcgTPEDnmyaA282gUVYAD1quUN4iL374y0CBJo+xX6oVnrEB8W1s1d3nWjPRJre
AHBxzZ+sVfEvv9+mX+8UyFkYhm+gLJQwahB5cGRBUEKzme5Vhc8TfNut0vIEvX+KQVMaJu4aIjKf
JF/aQt99l2NJ6B/SSeLw8q9wL7yACONl4JFr+IWHR2nOvPmvIgoaLh7l3C1jlYaFsKjjnG51+FhR
mJNrDZN5wm7WtZsNtmAdd+2XqreGx1RFs1ndV/n8VIBv2HNLKqGj31fKb9bKSyXTEmS+vveCsT+E
XRUUDaic0k4UZLsFO2j5UqWo9to6sWYdaK3y2/15zrLC2U1T7XUlOC79F2mD3mn/8kK7rQX/FU57
0HUrusw9WHP3wik9GJCss0dVpUGJ3YNxwNKozVWufaBhF0IyExLMB5rjozrgJiBY5Ai1IncBsv7z
pRWOUCaPXA81TqLbD3/zDHGq068xlHTl/z34YTFVV8PXPZnWGpIol2URPDiHKoNDNkGDSmQ/sVtb
qeUZ4QMcPh9l5y1jkQxfcxmah0Kak594GeIuI2IkSfzPFPkcpftA62ao7HwoI5LMvqEaXDXlvcWs
8ZaVIHnKuC8Xczj+LFSL/1ac5n7T3U1Kxc9nYukWXaQ0oL9NR+2mZJi6f6nAb8fXT19V75f6tNAK
oAs1mzbX0YgcBjgWtfjxM8XdNkreH4qRgfCOxZ44zlN6anjLJUo15+x+/tpb40EJBdJDjjrtQD9a
wxucPKSYIWEEP+UO8AvJUBbd8hj3DA/EaNExY13ZGqpDYMXiAWA07rORvuQg6WwC5pz5EFSljL/H
/DVcpDCo44BUDJ202ig/Ea5PRJZAT0WH2RZ0pKIx7Tf4IiO4kj6JV+jZ0j/KSIJ+k+dzIWhJOqf8
v/CQv+30jqxDbpzwA5TF8fb/zPKRaJlsZDG+FGNNNPYdfuE1wW2Z8TX0dayXqD6sA47ymkHy8bJS
sCOgCh9x4Wc9JfGzIitCkElfNWFO9Z7kDxZyfEc9rfQptpje02/GCrBHueOPQs4LuCnWdgx04SXl
0gkqFu4Y752Pq/UOH84QWvvszEgCOt7jjT40kQOPMeSNZGHDtvpdJFGzwvUCjG0VPcEPzzNyeeiN
zvxqbKCagCnGxXpRtcT/Fj2g6YEmkEO7z1fqWvxocpl04JtqTgkTbt6ADmMnij/11kTMThXcW94b
UmPRLELyWIvjeaxaP2wvSHk4H/8Xk06wavmy9NOVb7nb4uBMGW9Si/xVA91oP6xFL2S3iKBOOvhC
llFNW914g54Ea2iY4ohR508wWelB+QJNgpDyFLWwYqPRgKA4stlFvrMNbmKweh9Bo02J800tI4oK
h2Sl7dqRNdLiiVlrb2mtB86Uik6vqkKXMbHsx//rRVeCR9oOCjmH79Xu0gajvtiAcEHbxbJdq63c
gIyyWg5El/oS7ImDLRm1DPHUCKKKxoGsyA97jhWbSN36ltvnxxi0uxwlvc7DlEcMdTc+zkMSZ2Rx
KNIQMAuZhC99o63aXBdfk/RvzM1T4Em52FJKqdm5WzgUKbuQ3nVXJDLaPka63HAQz2/V0fO0QYU7
XM1YolNyhDBobl9Dkd6Lb+V78ARpzhKF+Bnz6pN2yPYtUWlK1iAezVTQxI/jNBUZ61ADymjHm1gD
ewrNzOkRIE1GXfxHzRJ8UGXd4PzBFv9zqMqK3R5nuELdxePZFXpheYU0CKFgWauczGuBSGkWuLKU
kXy5Tc6L1UiK+P4bcayS6BQZQ+7iObujtCJTihVDL32qIck4M+FSwQ46t1h3CB+1MuMwtOXg0j0V
ykwmnjz1buOHvAXlxRUjknZrqitYbuebKpcO55SyU8ZEUFFU00e3Xo6yN2CDZ0lAjef6MG9l/2Wt
Q0pqQD69V2snKKy+bWEUSdyfP+vy4TcalD+hrIj4Eum1EpMzigDieBUnPC4zUXnZ+KgnGw+dyZYB
mw4XVq1kM+GVp1g4QJ0atHhULjUsyXwgTUICXzMWXmeGy7+mw3h1cQ7oePr/cejkPOlozBh5g3vC
ZbhVjjsSg6Aof+MgJoPaged99AGR1D+RZZ4klMJrPgSqZHhj08YUJ1XtctvWFEi+40XlkSknl996
nLZJiB+yGpB4apvxBUIq0j9nTN/DhKN71tXAoBjbZG5zboTYo9C51qf+HlBxfHrC5XF7c3A2oe4N
ECczVEPYiGTvpWfPo+PbGm2EUa+8uadrInBXqBcUX+fB8iKGe6OGElPjPd/j7qSeGMJnUVapqqeL
btHEfhqm4lvGvJclPc46Znw3klDLewn3sNeCGK4btgPyfLZj3z3yHDcRwD9ag9SbMK6ug6/P2njc
IHuZfKCDh/CyHvCq3OvN4wjMyiiNmOYsvtRlb37nrAgD+wtoeoqhfHajvcKESL/pKOknGwOSXdne
luA5V6RRGhQZhgU9B9hk+reLh4p5A8EofNKd9Td3mTA2wikp+g+KJk5fj7XMkV5nUU/N9s0MI3QE
2lffyKyvYF2K/04AODlJ1vYvKZqVmt1ukszsknhIzwCCvIkQEI+0yE1UblHkDQ+lpSMxwkDgMa/L
CXn1lh8Pqc/KnXSWWr9l7d8zY+WDbLm4FrpKpZzNhjuujddctxZSTXtajI+fh4lx5/c/hoqFmwMr
jG41ArkjNZpDkIcUMT7Eq3M9GnutbysKzwW/POyamVW5GzioCGYNqmEhgICUphPTa04/8O9tQALg
3VrOulNtuzStiuf4ni7w/DjwvXI+qEu5fIUeKFTQnHAjfJskwLHupNVD5lLOBPJEfWeRLwZggTdF
DHa7tD12KYTWdbmUV8abv3Tw+8WNxN9g6MSObDBksHddMMcBx2Gk6UMiOutSwkUCV6/PqpVyvcg5
ooWz3mMf4Nlqe6y5ykHWhOGy5hYGyiA2ZuVk3RHKX0LDClqe9u1OhZvQW1DwrMhFLguZCB/o9qks
PHI69az4ufIRhb/7AuTcaBR6jw5K1DAlOussytmWXWHadWheuP5XEO3uAGhZQj2/OYb0U6RWPfEf
OHgKfPGjnr7ClGKTYaFDFrF/1oFspzD5OkpvVsEo1o5kKhW2TFrtZfB5NGBFXtMSNYE4MsnMrYl1
Mwx08d+VvQUWDnBJtEcuvkEzADqZZTMh9trAn6+XdbLmJmnQ6Ti4WTucCJ333z3vhqJTnq0mCVeD
C3FBTaNpB+cupXs8zHTviNXIk68W0z/TS25zo1lUbH9iPPgVd1bqj+rxP6/umK6PxGcswu8ojLNM
2qBD3+lvA+35S5+U6EBBHvKHsb8CHBbuJzH/6qvf0K/zRt5RtF12GYX8+f4MmmTlFaNo4nbzwmUp
gmmI/6JneaBIxFYw7kBuBet6VYPIST2Mg3WsJ0IROwuiyq/ZG68ZDBdRwTY/n6k/QdvnXfmIgp8v
tVJhMyt5ofQn4IKQKad+skh2YVcZWZtWsTgAkl9H1w4DVOPLrzfkQ5TM00JHxsAZxqtkmZBsLnpi
7dNiUXzC2NaxI2Xo3VP52LdYmuqyuPigiGXZNXIL++mXz5LIpsytDjU05+7je7AmN6tWDn9u36cf
O90xDxat008RCsR7ahgMq0pe6ukH5lG8RzKEeiJfJDj7Sor6WI7tzN1e2WrOF5sjZEyVX0pheQOj
GvmMsOUI0bq2sF2d++i099cyQ89Ux8dBCL5yQTIN1Zh8/YC50M+hnrkRPaH93zONGcot+CgtDRRR
OF7vCTPNR4yNiKgasWAfX8T7XRUN80i0MJWy16B0ioY7qt4CrKDQZ60CygQuE6bOGrFx+ffKsIfs
2Ht6svvs8gzaBm509vbHKVTwmQFgVPlAaHVHFQgWAV6ZAxr31w+PVeBybhLDlcR9LPbMXJz2z8QL
2H6Mi7DlKSD1ch3hBApmvLql3vt8463xXZtsVas4MgxQp0EGMSHIDkBb69rWsI0qG4e9hNUF4j+z
6En0QOElc8GeFYSq9o4Toqq69VhO1YqtfaQuXM1NE2b7ZK75ve2IamNQL90VK6/G6NP3zwWUNMNQ
8Kc3wUgHBTdZcZjw7F3ZOW9FthVNuYBN0LMt86ma1IQ7hDbEtPJLAkHah1AjkB7aKjaCjdGy4b4P
L2HCGC4zpBxpYQVxvJMLvSViQAfJVjKOZZPhZXHOnekyoOEhlkZoSyHA7ZPBXdoiUOLClNZ+tGdi
X0+zYiykP91Ootl6VPnT8T8/Z/mjb5lGGkAcIwvmM7nYtDwZogDlbMDQqfZa8JywSmwRCOEHhCdC
vB99CAL34cXBOtO/mD8mmvOM9+KaZMzXF+tllyDfvdnDREh8y/q9TVuDxk1ku3CXl9hP0nISzq2C
JjZiApHfvS0gv61+TyZSGoUE05sel41qbW7rbJQZgsN5OHyQyf/6qVLb5t++Oy2ilIPmKcy1DPUR
IEDFPlekm7GCE6jy3FdK/3tQvz9anYGdEcYNp3eQayvdUN/53GevXrhvd/mJv/NH3erK8Y3RKQV+
MF3KX3vlAB6W0ZAH8InuRbI2HD1AWY5+xpZS4jdAN0aC8VeAsayCXpBL5gCzmhGMDl/mnlgjcFGH
DhULqsj7g0LtEhkLBqaUpeprMZcRFtc4mks009kurYsf7F4aNnmidpy7jNMX45hAWQTh6zE0VuLE
eEL/f7/MH76HSLAulyIVz6RERDAZKyVF2dq4ykYoy1gWgswq2fwFcCPzUaIBaCwVe6MBbyHjf7yX
hls5ihgck8UxeG3vhReGEQEWuPo4p8waMcFoB4T35fzWdYpO67Y0h9yWwWC1EI3ujDb05RHmtY1a
2epQYqaIqHdCM55LB9XG3efz1SitZ9IfOwPQ1tUF6wpi5mLMjUJP6pggMheKZE//gghB1W8ZKjjl
6c476/A7uBNNKIZe63UKvm4Qdn+vQNkMaCvhSIdZL7OXDKNG0L8zdG7nwm+f69EQOF15HW++9Kul
1/H+Acbuzu2rrM+jaIkLe6Uj2Eb4ianAuqgaRN/ONEz3n5JxaBJN6T94hPFqcFdNf8Vq1Ex1wP0s
m4fcGIzsB8L4ySOGAPl8zCQcHeFCdXAjboBGq8lW4SgcqU++83zHT70QgX8ySiSOOnptdVnGmqBf
/b6kXjpSGI7FETnA4X+hf394QPDBMvG6RTr1ioYofevMrDlnRf2hamKjtR16KsZ6JYLzzlAXtKxf
0mDBpkRi/5umMRYaDsa4LQ0N/kG5Bb75LfGrdrxBgP7CvPajHzyHbAJPShMs7rSz/w8AX4rIOumt
MfKgFo71f/Zz+vpVmG5c8hml5I4Tg8M7YsQFnuNWaXtUWrPs2lBSjg3B2/weONm71giK8k8SGxhv
yLaa7vtH1OBX8P8qQDGqwDxeKouEAkSru19hEoHl0niTUXcuIbet7/fR5/ZrHy+h8j6+1J2ALLhZ
uXKigESb+Iw4fJ7wB+7KKetW3B37rs5UiwGh/VMsxclP6h26ThX2dWFvUDeFBKVfOxHWg/eK1zXC
QW3YSU4+z+8rtFXB0QdqH1qvwFjL4wvvJ7TbmS5txMU1bvURty+XW7z36r1y9/SMkQoa92dwiAcJ
VGdt6rAcOGGvY4WNIp92wkNwztGQ7X6am5NGA2cOBiKWbgazDrbPF1ZT1VjpxAjILjAFlal9hDn5
2G4z9VCohibfO3vqsW1jO6JAt+CXv/QGADdKlR1fKNd/lmS2w//l2Rg7ocqa+avkMCaQ0S8QSXvp
IzSOaj+oXqlj3cWPe1ou76jc3R5cj86faN60llgXsvB4rNCQ1JY/5QUXRQklnqOUF1KTAizD+/dL
6yPulBDz5f8fFlAd3zNGTsRZMDLn/NGxJ7K/WBJV4+bovVJHuU3rPqraJ3cxjcYfVQ0i85H0n3Ie
/4AQldNlBl1sbaW8qolbN5EZCvMveqV7eDXRAhEInZgdXj+r6BwsB3Fsd+wUhMZRrlu0uMXOLwF+
AmIBjgOfOy+p0gKG1xwN6TpXGjhTVjalQ0MMU0Wb2Apz0pl2HGtiM/BIkoqxpLvLwxIDVAHNL4Jl
QxJ21mXZltHYDniAwDrRiYJ2RI0h1wM0F9VQe3ws0FUoW7IMkcdOCEvKpzNo61vryKhRDN9DTyLf
GdE8de0+Mo7sJ6yKDgUZD3UIoIps69HTWuNJy9pQaGekEmvTUtYnvcZ0Jz6ec+ffAprSrtUeC9Z1
tsfeB3Tt7qmPAorsEfB4zV8166fC8eGxX3A30h4f999P2fINttAxI4oZln0TFPx9kSj53kawK5xe
I1SRQUwUzD2P1vc8OegM261sP7QIXphcew7mHwja0oEzW4Xtp1lA1hL01bmhRFHsmrEDBLAJc1ej
ozljgRSxxIJybxAh7P6VkRXC9tDnBlG3XESOt5wSrzOvTJ3rQhbl2il5jb/0libKwef+GoQtrB0l
g1YaseT+G/D+kMkZIQ3UnL8bAht5hdfe62lJn7S8cQZzjbLsYE8jWtShuV/uJefA93J7zLhZXvMe
U+/6A+oQahXgLkRa1lxwAXnzIRG5Vr1JVJlupxbTjgCpFL/Y5SB49ZXU45fZvNJGhdE8ytLt8vCx
iQix8WsdHvGjS9RofB4cffvtu87UFxwbYubgW0e4Cz/3RWBnAeLyrePBWym7GmpVidbE999rEvyg
x8CWOEZAptyVKaYm/DDuBNu7ZsNHHNZVvOU4B2P0ReJcoc5FyqMyPSbCp7r7aY5T1vH/99JvsXMX
j5+mGafcqzkV5p2vK139dwN8DZdhXxBQvMkqRN55HqJFRtQzsbiSkeZyvZoMMIxg2UABliXyVkje
wAVzmyFBO7soKGADzKdlfcIvThk+LQMT5uODpqSic3+DCgfpZCYvFEbcEHrvswda0STt5bfx7t3A
b99IfENSk6tGNs0x0QGHIoCmQPubYnoHZ2gIee7pkjg8CfP8W3hGst0tdBzocTZCoXY5rfAIQYic
xgeUlHrqo+OOU49/VCtSUBRZt6bzKu+wjM4yjirxHkoQvSGgZlKIO6aKLqdAPexOr2E3R3c0mOlY
r+lX/udlaNEWBFKILdyy2We5iMCWRrAtnJ848LlnnpXMI6jW8r+s3iGZJVvMOf2w2O3ZStldU68W
nNimiSXg+b2k/+HuSP4F0XTOnqq2WPab/HxnQR+pWq+y19HZYbb9G12SHWI5x6XR0s/uTahCxVFV
5p4zQToksf2JyUZWppyw0R1cYc2RlOkiJcag0w4zW18OLKerziBENcEBABaQc2TYlJ/qworEgckA
TDZKA0bNVMhz5fCgxQRLJMQlOBYPyc47uoAU/u4xOYyB0/UrPx8SV8ZnBExKWeslNFIMCjGVROZb
ClCch2z6plLGF4HtLcuq/uEWUuijRylENn2p9MT0GOO3GMv5/xEIxoGgtz+4WegdWjeFsdadcWPP
ydmTXFJcgiPowsu3DTrXeCCrE1f9F24aPyKbR6Bcpmuwo60bBat36l8cD2iYeXbUkR3RxzkNNb2r
zUSjNXnffxxtbz/two50StT2gYPKgEuE6kX81hO/Jk/WcZmqdL6CRmQzTytmrU6iyWtZ/4f2FqFA
Gg23YNaaCXAUX+8lAv1UwnLv69smkbBrPLODHuQeLVL0CIfX7b631THawI3upYMQ5QV/hya1QukU
OXjF02XZ+Nx54kdRNuCV41SEuRaHPF4GZvlGvmv9MzcYNW46ZyoVusR38drcwETiWHCKCc/DRitf
6zs6rnnYvybj0GA6cADkyfOX5Zuaif/+0RtI4XYwCSwswCECWKmRNowOWb5nx05Jt5234zcoihX9
94sfFLUh3fncWP8PABXRgjvsJgVwfLfUTZSLNfzclR/QTEwkTIGe7TRscTxAepZcXWorS41yC+iD
EJx19D2B8Uq9kPvzk/1KgeZ9JFk2gARmH3uiEtBDK27FlT565VPQRU/cuEnOPfjTCdF4mhhGoNN1
MMa4lV6mcfYvCf0A4t7Hrm2zA7AE8JHmCPVqyyTIRSOlVFFwfXJM3FA1Xb6xbkRR8HTeH2VMpfDb
7F6rFbn79NXO70cQe3CxOAQFW6rFJHYZU4MzQGm+9KU8WEp1YfTncP/qrtA07BdodbX8TZ7/fMI5
ZytmokPaAkQb50wNSTRoXVnPYkjmvFSgbekKK7oGOBv0NBKbzhwoMZmoGuqsP/307wuGmX7laYK0
g7mKguZV7TLlShnTNuRQdSwGY7btb8BUSD7vdH44nu/uYklePeickroKfXwE5dWLVDwtnVrJAQT5
nLyFv99NwoTcd1270TESmTbBh7S6J5b6PgnmXYYvoyRJmYI/Uzz6Dq9x8uH1nebDlxNw3ZwafHA7
d1fgX7y0U6VsY9MQAXaWyiX0J1PxvdAV63u023bBSvwqqM4YPXXfVgkpkjG7qqkkT9ADq9IWARhm
K09lx+EJiaN99SAKbb78xr8DYqxZyEYolaF5vNMVkhpX1KmtEYjUXYMXG17XlSCM3SP0nndtcDCN
kktLeNdhw9Bq1OUpzVAv23v3W7a3+Z72jqLaKVQDRu8WAiEHVp3T3HWln2oTJxq1WMBUz/JuMY7p
9YC7qeA/qoZCqF1V5f/au4hdKmCYX8Qk4nmfgCteotXqbd3DSVO3Y3UfZlJ2+inTq0f+InbjnC6K
YMAMe8aKzADpYraMHCQh0qiMZ0OCx7a/xXxBi5RQKcUUdmq6nwUU+OE1wYDotZo7TH5m0gWgJ5WV
4wAuIddFF1GBjKvceETO+8/0SXT+r3wUOKOMQFsJC4y5NMAW2ck4f5kUYX4BEQ5eh3D8sJ83ocQW
fqpbocEZD62Nr8JZ3nGFeOkhh7wYrF/LHjyaZl1pnBXnCkrlRUDI7azzWk21qoXyvaaQLh1nMUTq
ybsV1fTwCZIgGCzN6lTSejn3dmMLCbSFROnQwK7pn3BvbNIZ7gTIZqT5Oa2y3fsTNSOTPIFi0QuH
aSGWeroms6HSM3lNfEzSd0jGPiThvO+4sOUvhjNS3KR8hf7ttmsAaClKzuDLyyqz3649ydWqhMTL
LgOe/w9OOk8QGcYwaTbIc3RG9CM03PsQTsD/yB5rKiYRugOhbOe5J0aT2Tv4TCKkNSs6IYM1JCDF
HrcBmdySwoBMAZzK8EwEyXduP9n7B2w736pUS3gW2o5Q2ZNKtykwzyJ4hQrUNSUwsiihFnF7eKBq
im92X0mp58KdSRO96gdL28q+TG6ZbHzytn2dAXn3U7Bhmnur0Fs7O36BjLD8oXORSYse+Zs++Pcg
XCyntJv789aeNLhbNn9a3IKcQHswD/fDPVJDp+ZEK6xilKaS8MLPuoyQNu21aM8wrYwzqjIOrZxR
33NNBd9bcf8ZUc3tMI7KQ5DusktGgg7BpuGTEr7I9gBrjczsGxwTD9M3U5Pb1EyU0axSZX2uqr9t
FUZXuIa4vajmwttsZmJzmnzHlDYWkz5gWqUTXqkDDZiXcXQySXCSsV13vFqLK+VFRnjPbrKJiiJf
YLgl9xzNSV3C4uRbF6uOinV7zgrS+/cV40Znz38nSpJ9wg1izsa2OiMECotmhwrXbL9Rh//OBzCQ
L4yDGifiTveaW0E2h4swqpuGD6+7jtO1OyZpBXdGnfiHBZDwbM9GJZcOG+q19uUorCfleXjfKvd5
W1SC5tDD+txyQ7zBJCUC9bvLQWAkufATEiCG+MDsa9OzbEjZwLYcBDqShAbC3P2CmDgm+Ib3FLcI
3wLzhn/fvnhfnxSJF7OT/5/Jpu6KWjW2fZ1W506+wHQwaW6Q2lTeOHTAl5eWrYKGIvyE4dkvPaqM
mAqiP/FHiuNZAEO/LfOnJE5zO4TnIMSDLGJm1yp+I3AFmHEwJ7gNAmsz6CGlOmhPXJUUoD8pWJb6
zOfsdGpiFgHVPP2B4039Q0u167kQHMNeFwCYfZkIuS+QpndaJKNbrYG12Xb05j5lygnA7Ivp0QY2
uOKQCUR/cRpwCpSdSrOu8jrw2g1rnASI1iIHdg8LDRs2akjQdX/7GniptOBB0BggIlxFjvOYoSDY
GWVHqRfYtTYM3/2Vugwg/VOQYFinwve/K4zrKhWuwcxvH4di/pbH3pA2WvJfAzdG3AqE3RDqlgZx
YC1p8LH/1u/7ByKBeXpIPrtAstNEirMao7o6PsVgMq3WTbeWian+dbi33KZusBXrnq7cXYJWLgW1
MCxOifWA8VhH1OGqrouUXt6/+mrk6gDWfAjt6yqpa2HAA4o/R2J+F11mLce6zJpTS3AhoL1IQYWw
UZhfHXFObVX9cJ7jTjAskIB9GalIz9Y616OqAvAIu5yLJHsa6n/uzKslFZBIcsCPNOtRHfYx5wdP
T23lx1pj39RJbdKvVZD5STvissgSffW6QXyGR+aH8w7aarLNrUiSfZgCJWRA6Czr1VPSttC6ROZu
KY36nZ2EL4rdLl4b6agpma2pvecVUmPNq4wjvnmjYUmwSJFvrVLncB/iCtNzxg7QVU6UD7r1KB+K
TCACBvVgrW2PXdZKmUgjBhaodbBGiObgRhS6CdS7L3qoT6yTxrK4w6PaAlGkb6cUoEFFJxbpM2by
GjfNl8RrqmJr/lIzQYNEANL6dW5wlFcfMkk/rBraad9txnkggTxxxATa0gFiTVBzPw0QMf9gWHd3
FBVWxy86m5Q5BZnUvtFHqCaxV0IxsNt+VIhryqv6ojRk20yMeZ17KLIlxT8bf/9g6zvM5xSEM07B
St4X5o9iFQM2PQl1KHxL1VBTVLK3fiQS9/vog3CtPoovSrqUUOoOWOZ0TKo3oQxC9y5qUOaf/Guu
qdgv6ufoxInJmiSFMnV2u6urFg1PMZjmuOliHxuP0dWBn7ci6/eOJcvbRPU2JCAoIQZVDPl7gnU/
U7UqjDwxPopOemINlvs++baaoLxWz8ynbTpwQSV3NqQE71aytsexGpirMzmK3b2f0TBqi7Ro3VH7
HX3b4bDR90Eq25l2MSE+5QYccJVeOwe8RNAL/pVt3tRGaOYNVsBXdGhTe8PIjp8nZld4JPDXSCDh
XlMQpUZDJvqE8WoQv6QPm/D+hwkbdqdY2kGECUBmjUZgKvXNMndz5RNrq8LZCkza8df2pwNhTZ8N
AlpgKTUyM4qPZqlk8x6dPWnLQp2qd4aK0Hga4UHpLM/kUpxs9Ih16RdmcSRyqjzxpZphqe5mO3mk
WltD9b/odQfEcNAIW7MD7GvGqemgyp3IgyNUAzW2HGsFiz1f2ooNNWSAwqIxKNu4WNjuHFIovguj
N3UQPvE7lDIGZgLHCB1gaQI4uQNwWrlI/ODHwYQ5x7WLPblCCrlFH9hElTqy5EiI9zvMKbSvlGEs
6m/eWCDeL12QJeaKWjkxmOFGwDawITQ7rbNIx0vYjXG3t3/xIiPWw1mDeBkI0jruIy01zMBaR5aO
tW+mceHpkX6YzsNswNUKUq/NtdKKx3aKJNaftNF88ri5oziNXG1Gj8gp/6taQZChP70xkPQrjq4W
8jJsAZwiyov+xXldhX4D8ghq0I51AEPJ6Y3g8ltPaigL29Iy3ap+Xs/s9RXGGb76i+eqeoirW9T/
PL/fapoz8bwetRcVVtuyicKIlrrLkay20tM12sLV2RKyc1sre5+UnJcXXZHCVq/OXPh63NWRSQ7M
Gy3fua2egnIcoh3S5eyOkpaJJsRqpKAMcViCytqNyqKd7YXBzi/kLSJmbprenAMe79LBZgNd5z6/
/oK9kBiUlMmVyNjMa7qPdvgMvzDYBZ4GXRwQzoHB0VpIdmCDiyw0hMwOGEu1+1nVyJ0YpPtL/jhv
wPFXWn64aPmgbragkLtKJ4vAr0O8tN3zjzWCxg/EZfOCAj9rIkKXZhTDYZK9fWl+d+zqa8By+Or6
2Ex3ydxmLxSaeXO1LuEbyWF8aMke7KYIzvQ0FebFd51p+Ww1XKGA47gv3siUSSLUjfFKWar+rpfB
TxoD0W7LmatetbeiAdlBVKOcNSTDBOs5nEJ52DUc5+F45tsvl4OCK0Q2YIWaUzXiJ6izfRvy8EyG
cvMJjf3l4mP5wIbtumSHXSUqsulHts6U7k/vX20SIZFEzcprsYh8IXdSaF493wYC8ZvSs2hIVgdO
GsngBSfsQqTTQnK6SQ3LnJSfObnUELQwFvD0Q+O+lrR9gBREs9p92i3OiSyupAa3zEHF8cvrNQJ7
dpl6Cvsy8rVdof32aYGQ8beDJ7ZDb35RHTiwjM8in+UKa2n9NG7UYUz9gOYt/cP68ml0c61XS1S/
ruWkyu81gxaQt6NTEDHQCXX3AoaZi85mzwm1ReEItcmXjjlVemqxSC1CGpj4e9MPQWzWxKiehKze
aSIsHw8c/ecbZaCaz0qPKMaYo2/eKeIR+J5ZFCcROFkRlK0zJs5yhWr0IIiJfIAzpNGREF+vdqNg
P72MbhUpH8xh7v5cYKUNE9xYYXytCUB/OjuHS7QTcFfMuLeRVZTU28ka4XKq1dm+MMiCDTEzQ4/Z
zd/amWe5l1YWOBR00i7fL/6ZdBZ/FuhO9WrsuZD5yIH98Gnaz49McgI4CQ0LGMTvMmehTan3CxWY
2XZBGF5lYzGPxCOuwWEyqYBIg8RObY7VLeRRmJp43KF/eE5wqnYxYUUGGOBOK4trrwtIvy9u9RI6
Mxj1i9UKjntp/khLNQf5Klc6qFFVGKfUgCoUqTAIt2PMdhL1hcE1tTWPAD/W3O539cCsZV1lxfBK
QqXwu75ugY13i7UqJeTXe4kMxmLMWLm3y0Ri9kmkh+BNSVtIFljIkCQV6/Bfe8ZEBlM6dlUMj97+
Ocr6MCm/VbRdiqituUpOZFBo2/wwFTDqrHolEy4OiliHQsqouwZpnBrZ+O7NML9nZL2RdzoZ/ioT
ATaR+4qoS9Wsi2tehUAvo170kNZOxE/oAp61eA7iuTj3AdGK5ITHXV7qprg2JlUoi/Tx/AYfSW5C
uxmnwLDoWoBmN5MiTeHSTXH3xAJnMm6JoofD2GWwtyzjUDpvDTLXUTM5lz/jLg+GQrbxuqs3ZdDv
LZS9rLt5XvoqPUtfeuwcNKLefTtjRF095dS7tBUeBfcFB3oN2yL713UHzbM15vdRNKywb6mpVD52
zgKrIPyorZxlcTjcNvpUm4/UvQtHnRvhwseBReGGtlMBk1UBinWyU97Y5CGykiajh+2TMBXb4XYe
tu4IM//ri9ZYduljF7UPh0HoFMxycRYhiJrGEXukPeMqO1MyFF4h/JhtJL1MqebEv2ltkphErVkU
DW4MVVBV/F8EvvFYHt7CsgIL9U7EtB5yXFIoDdJ/Wc57+/cKLeLrAJvX1OswJX6QqWALswx3ZNuo
7dC1eFkVKk0z2f7eulKJglj0DV+xDNGFrI906l2S5/FCjUMi7Lel3HenJjbIFUKV0A5HF6r20J4b
3M/VD5ExOGncfGP74mdJ2zXCPP9Rwxk3Fl7hdqgvAQzPjNoj9x1X3K8N6JN2bzW39ePueEJmR2Pt
pVUeoZ/k9Ya9JwKw11OfPK58bYNHoDSRfk1g5VU38Se/iBI7DuidmuuyUUn9Z/+kzsB3v+fQGo0M
vVSs3VB+o77yB0gp8aDBsLUQvVnkjjSemKABEAgn7r+SVBdKCPazR77DlrfUSpgjTSQtKZmc03EV
CAvA5FZCDGg1sMMhr7X5KJIqLlqxmR6c2VsHOIsdRvhgq2VhGWRAQNmD6HloD0mORxrCXJ493ecz
ujjNCm0eW0QnL2XhEAwJHZRqRyxkez6bU7/vYZA5DBkznv5tPIMVP50LKBta49C3SDxlNFaMQjL7
CTjHeny68egZW7/K5bO/OdxYAHYixwwHit0hKGb4z1ylxyH5aEuyzdWGO27fuUpCxBWIbU2jbtkM
GGQ+pPZg+bj/DXhradIX5upOsH/mz1HX72j3zKDCHrDMhoR9DPdBg9+5PD9fiNhSfaKRfKvNDuwS
nr/PveIlpckzvoOS29bpPCCSD1GQqrZG8HzCzIKKGVRPjWGCIXCUdMFxxbGkLHFNW5P+06oPGrQw
+5O/oC8K0mMaWUL7CVH8rmD/kxuN5s+oFeFZ1mX6ncWfd3JjXWEsE9n1dfsoacq60rlmR7rqX8vY
47vXBdrNoCz7k8F9nqCJxPrG+oLlXT9TGplhI0JlvXKq1eEmuuFvsBhJNPeaNV5IPf6u/FS50eoT
3Cs3dw0XaGAaSrn42OH66/sdSlbRfjmpcbPvRRCKO0BxMUkk0V+pZrWuQmXdlsNF+q19ojiMKi+K
Y/NMQ2OozCLPP5z+kCxxyjm8xZJ8SpSxFnfXMER4bPLPLcP57ccI4gWWXdK6bUtJ/K5KV+d0BYGM
h6Z5kJwoQ0VbidJjOtWYAlZy9SDNyB3zWLf3atw979+DTBrvr9xkZAAoQUh86TFXXRRIWSV/iOZB
FrWe8I0FIHf5sGLiFCKXKSt4OygWwRGkf8tcY4woal1Qbz2q4EpOxQ1GqRoCKbV9wTPjLHTTaXal
3ixxVkxc6jJ6YfRoc6i1CypPagupDYAmgk0XWreiZvggiSZ+raojMj46KtPi2C8TvEf+YKvTtFbS
jlbof4EHPWasUec50YPmS0wff7hONLp28BggcBp2hdM1qfgOIVq2536jbpiX6O5K3Hic69Z9aw38
TN+o8SsbGAlwic2dprWDgwCrgrgXeEqMsNndrB+f+2+KzcyKotItksXHAzAk+PrUzT69LL4CxkIu
N6g1mvHMe7oDi6NvATu1jfvyANa93BTfWPBpc0zWIvXjqYTPn1kSSJ/1qEFLeuyfcZPvZjWOIgY/
rDK9KAUCfl0SOdyhF9aLHoFu3No58LLxu0iT7vMo11YP+B3JbfAC6vuq7Gd9iW51TgqjALoI4U9q
5AtvXdyL9Uaa3xoRPIe4alyL/3+RAeZUabjW48DPU+Jl6iNG0QxaUnxXIKwaNrEL8q9Br+Bw04qE
M+6TJLjlsdrigktGRaqJT53sQQpyCozC/JFRCDC29Bcm46uQbS96nI028OUFcynMV1MxW/XdkHTB
aWMHcwjjtvAR5jCjoJ4xcZ1XkgO49uS+vdlgEJr7kqZoyq7UHeFpVh+EODHLp3NxlV0ghuPaeA8O
ekgmHE3AOFy+6TvidYIuVX8en4rXQ1ctNqWmDWEF3qycH0eHoinZF6C9yEFTVpKn9AnMst5WorWG
dBxdt3nYITRhfAPzhKi4ZOyqbZfyDfPfw0pOPoiQ9tjVhn+bA6EZoe+KtGZ2QJhaxJ5T7DiTmcGs
gDrdFbuYKvrEI++USbbUxEXAjNB6hEqv1y9+HbydhLMTIrZ+rUL4dqOl6b3qPP9UWILvnE8GRl7U
uhnZ3TSkR6AIeRKz3DO+8dJ8ingP9Q/vsM29h3BYoTOIfSKaFlNhv7smmVVyNDMQzcU0sVbUfVQa
b3AbVR282zTrMKB3ewPhJzp393krRfnRNui62Zp8JMbd8/RmM/JdsJrLML04mywmgwd+Qv0dLS5+
Fxk3E2NneEiA86qcOQBtX/7U+2SAneVhKDLA376lUya2pXjXJOmSFZL3q7SMSp55psi4s0ZAH9NX
+5KnzVMTXisFlIUUYiaDjM5xjTfhYJpodXdI54RHH10E8fQjrHCqB8kqiaukb2yVhrDD+0otr1ve
cCEyB/4ML7jlwYgGQ44R5EVXIXHtqEODSeWQoGn7JdMD5E19mSvcYCkpYzhBxJKrSEJMJX8/0+Ny
fKBDcmreJAcftyVVvNaIUx6lTKFxdrvLvirgR0mso2i94LlmDqiY2mtYhb6+POWpv7Ylqp0aO8qY
MkLjgh2KX14GSO9pVL6aVUuLSVDClwYBehgE7AXr2TFwJNa9a55q1R4xMjt+inQnRWFmW56rrcrX
sLB1UGJP48s740BAqDutr6d+mLfGIYistMmmo7gvbIFn6Eo6I7pAMq40oxA1W258kz/KNugRlAWX
KpVKfQiJB+wBwWsDh6k6FP9i4imYubZP+hkrY9byEMt9ZzrIvqNUgcQqSHmcxWgpfpTO874zs1gi
0Y0kQKeZHxX9Qfv+LUC3CQkIoYIMCpX9sJqRJof3I3eQRQIHBm5IpPxRFnre6EFsOKdtHhRZfjj+
NKd9kiTJ+EjNN3VwJcyJwg3xsO7eRlzOKfvK4lK8D+0Bk0s09fgsh7UG4xrUBie5uc3EvYEz4LlX
m0o3lT0xAMiv6/JYikrM8pPYvd1H6lxWVK3Xppd+Oh+RpcAcQAqHOI0NooIKzNT6zCaQbHgVf4DX
q1INfupZOc3I5RsyYDIHeBCqMOs/oUmdeFMnYRHNUEZsU+6VPOx6ZpUpBh87KBroXR+NwZdQeGTK
5+UJ+QL+6JPQX5wjX5ktEtIgtJ2CbRWAVYMUS9ggIgbNSRL+YGqdf8Jz2v5VLqEwWZEDoegD1Cgu
/Kp/otLldiZ8aMylVwUNm4ihqfjx6F78VkNDjzdPV9CDBM2qCmJRmCb/odGChRZPba0D/FWTQOP6
KtWyrIb+7EuXBdWtH9YCZdeHQrf2lacDpGjb2uKKMnaYrvSuM/dqNK75oScc76Llllz5LlB5ufum
0rIdiULwl1RCivGKtuk83qanST4bzpQUx+niKdKxdVphWzhul9Uf5auL3D5T+EclGMVPOYqdS2i8
p5U0eJjD5sdUnSfHDgFwq+RzBqZMzF+hKTkqNoDpIrCbxbZuHEL0FTJqQwcV3Jb0F4KdVT5xEDi2
rxtLPz7dYzTmyiF6LWuBlpQNO9rKHvnkjGvMHWZEyngJ2s8NBqB1T8plUoFlTwnnRm6MC16ZFEWk
B3OQrJy3JXI0sfNPaHE2RrQzDVAorTOBJxcjfvSlJ3IG0ztFdnhXOSeLIogdJ8vBbFpxBmeg/88N
Lixbj58NuksFgW8+j4y2IAM/laG+qqx2xktBKDdvtvRnzAf2aDW86BoL384cmFGQxxw4TSJF1/SL
1/nCVj5d3xJ3dxF9RfLHkUQkqRlbLkY18g2U2cpDPdyoRV0rlb25FScyPFOhSzTiL1SUXpFEi+UF
VzNzaYO9s6rRgrXQPMoAN5BnC9imHE63Rvm1rLIfi9fR5zrlX80dqqRaVyZJSCMOsT0fos62vHGn
qr7FgRyPPr0wt6UbWiqCgWiWGWKCxH7Pp78MpnMxKFdsVmYRgjKKhFijYBlkxEdM9piKvda/e368
OqepxmUlvyZK8/hK59pmy8o1WepK6uLukRRbNSiOISIUdMpYT8OqPl5B/G45ixKqu6exnMFDFRoz
1xvMcjsP1+HzZjoj41R4vhDZsyiTMWRNaxRWth4PwFOainjsmeVWd2s+Nv4Ru73TV23lwROoqtB0
7je/2+keY5cMYyrmn8BrbIdbAXo0AcJJCC4Yzo6scJzsY8Pj8gMLLGiTBfEXEwRpUL+BodMcn7u4
7zzXj5vq6I8QT5TGZSqQuBe8W306r/TdK4PMX/g89QDUL1jWIFT/u+CpEjXnK61Mi8Ep8xtM8uLU
mxIyimmQ7+z8kkmuCPsPQm+bZ7Tb4LZuV10tQJ8N6VNEwlx7Ki0VuM+J1YZw7nqxX0zY6DUcVu2d
ehP24b8I3NY6q3F5YVA3ZaEynnvhidH2y3VjsYQgk3gCXAmI0KZPmPow8m9NX0478EwSoSj3EBUj
Si/6gL0kXbPnRRNl0+Tcd5BSHKjOb1oMSXns3l78kcdvwcXrBetbAMJFkUHIgbG85J6b5H++LjHu
KSjbf+a2FDyMoICiAJ0veXFtbVUBVz0JuPqeuBFC67vF22f4VutCBwqfuar9YeX3+mUbBRu82jwq
rybzz6qPiF2UAE2Cnytk/rLphif6z/me/ipAMN0SIpgu41uc1q/pNXkDfdVQ/vV7/s/eVIX0ND4P
H0cTY+4QBKWDl6bwxVP21vxfVDzL+77h8P6kT9KHkpBPul9hBllGdl9suzsutZT0YIL7Ouz/3B9d
aW541DwbvRNGWvieV8NU0tTQi/hVkuYTLsoR1Z/AutIOwFjqfbCxYqFNqda/hV/dlsldALC+2+Me
EYnRZEdq7xOApNaV3Pm16lhXXk/6xvHig1wrddqVy5zlI3Xbi7LmVy/kJcI7PvWCSvoGystv0FY6
btzmUqu4V82y0G4V4e7AZ+DOMJayyX1TArR6qeKCZp7fFlZqLTQ16fGG6RgiQ28i2tVrMTTr4Ysh
cjiW015/CakqT6zBvIJqyewv/dh4SdsnwclAwe8leGlvgRZMGA2AG0+j/3DkFGpEOqlm6wgbOt8i
5uND5zC8tNgQsu2frUgf9Rzt8VtakjNhhE6Xacnt/EFEag+Fc55Fo3eLf2JRBMds+8qtxuZ3tgRL
H8+A0HQm3mp7K2vyBDLpjuKGs0lSKJXUALzlKcQMBEFIjbc6DYzqUhQUcn/DX19/GWqBFeNihT/A
Hb7c+a3+6a5kMs9Q8j5+IK/KFYTHeaHz+PigFtL25x5ZlXjy1Bng3yCFb8YtiSNhK/dFL/JpNxnr
qhtx8RIzJNwLr5ekeZS15UsATBpSyU/r5/dRpwMVEqiZ553KNTLKXHO7y0ZICMjRuzBPzp/SJ7lT
/BX+oP5EPk6TeNYuRC4jijDz3lCXp8CaTuWA5Sa2g6kzW7PEsOlyUCX8xd0Uai3URFiAJk4sxuDO
zY724GlPv6iwala1ghwCPS6tS0ps5Z3jjwqK0RJzLDu9d8fyH7VHoCjYPxPhuuN9dv9ttomUmwyV
S2PwKnHJKPZG2J0R7dAxak0k3MsFbw1gZbFE1bkmy6qgbKg4fXSO2ogzGYmX0gGer3utp6ep2t/5
/RmC6NG2Y11dt0DlrxZuLcBCCsJEphRcZNr11LYQ6Zzdo4reYPmR5SoT/JW28HsU9yf+adVNBfiG
HhzyRc5E/gnKrGLpEqo7Eo3lGVUhPaGzVCmJ4LETpkS7BTAlerZgzJD8Frf8KdR9pgj4sAWKSVFa
IwgGdO/Izm96FiMh14Rx5tpG4GfmiQ0cKq19w8CGY9LEZpDQBa6wbJNgwjgy2csE5StDiFy+0J5v
QZ8twpxboZPdzTl/sF82MhsA8rMELY0P68lzYdDMS7iVGnLl39D3ZNDFWJPQe+pfNE9l7mk5Aqin
xQcoZR16B1ZLYQVGR2Oe+5NDbfKNMRwJsWN+QdETDdzB4vcbnVoDhdscJE1tR+x/H2n829xAvb4D
GEiEpBYPDRf8ct61PopKHiw37fJFuyjIryZcU8XPCA0Vt9bghZ8x1SbbnMLAvEmWKzqmCYOudY6s
XL97QUkRhZQlVr8H1oCFnJDUgsHr9BU/CZiy/IxfMjPwhpFFk4aVRKJvvwgfRHpRZflJY4w/fCLX
f0LGvG3iZHo+IWD7CXxs++40JYnKhEK+psMq7cYb5KuIoEJiNQuWlCCCt0Szu1x6GWTcTpZOFdRg
zSJ7iBIPOxKEUlLiVM1+XwWS4Mqn5p5EqAI37hwRkNTbucd+oFBmSL1dPYPu7JqpPCxtLq5eb6WV
G0M3VpEOEVYhvgElamZAxY/NI+XCnGqOIxDhOXzYUUM/dPs5sRDJ2OeiB3bVD9OrUNWra34eT+Kn
leyvwowsVg+jZumR41Gq1r6a2VNjZtlvDWMT+h6dr8fnc4K5fed9Cq35pWWvRsqMxT7fMqlatLyD
sIOvolfImlyZjFXm6h5//RyADzyfx3Zo4JAwp6S0eha/BmrblShIPVNcXZU2i/89wviXoex32A74
Y8RHPfeETKMBbEBFZycojiVBzBrgT1e03Los2D7Xbwgnql/f2N4/2ecbxHdXB26sjbPMs/HiL6/g
IUnnaXrGpdvbhb6MWTq90AQHQUmv4Xkl1ANDFkLXO8MyiMOWnN7IsOia3bMURLT3xGkw3hTIHYnX
rqubiuQoP3UEsdpAAOFBdnGZCz8be0Oeth47KsJIEIg1ObeJjHmfgbWtfCaNZ105/3SLCci0LUjF
7l2ZCwPy6ywScQ1lZlG2l6tSuOsal3Zpo4zizinAwR7qDoB790WUWNu7LY9uZUUyg+h2YU+fZvB5
4hzV7ld0BhIX6Q6/B8DgJR+3QuMJOAbWi3nVKQtPVtbzstHfZAuG3WjKu20pZShzN/PLgxLlpXKz
AZnRJt1oqEaTFMbriN6ViB34K272RCreyq13zg1j/hIqTUHnZW15zlzF77DilwFXIjuoWFkrjY4B
gMBfAbqMCtxRMHwQUgr1szthTFNUqBnLI8efXOhfljy39z9eqp0okfee1c1PIhrKlkeo7JuB2LAO
xEY83VBdzpO9BSONz7aeGtwN4y8WS4H4JCPsg3X1Tf158Q2Y2kBVp2Qy8eIv1gzH0ttHmCOF1b9O
QwV5VMQALHYdf/vcck9TSQqyOzV2sQUFPEK5hzofMQov1Oaphifr171oFMbOvMUEQtFBNZw1+e5I
d+07//JyOK7PXHMMje1P67QpCTEbujfF+IQBWO2Z5HEnnsaiCeKVI/tAEJoqzmRuctLuNuTsu3n8
yZS50lpvwd6uJt2jUBIM4JFMQVEY0NJ8q+dFDWtEedrV58Z0XanJUvwY7OrHqxI6h/MWDXaXYOKz
lvPQWP4DrXB+1KlzGjsa83HykEQHFAk3H6BEhqeT9M334V1R2JdErrsfhdIpYEE5LEmiXEyvt3mO
oIoAPNXSISQvwleKmVCICEQBvZS8pLG/cr83N/a3w9FyBpuI6gi6pJohVhy1cJj0oplBHgE5cM7R
4m99DznyrS108FG56fl1Qp2bzs20CGXjy2QCx4Tka/fnqP/lCgdqsY6ciuqIi2VJYINaFALuuOZp
Ujnfi6pCNbnIBnrrsdclOUj6Ba3htvNlk4ydTNrYQ2oOPu626/1ZKL19POnY3T9K713LWa0c85ms
jlU2HMsgo+jvgcosvRMROPbTPhnqhK5+zy/BI1JBde0YFOxzR+ECTZhftNxX3A/fXKJWsa6U6Q/K
DYINxRKmtTCxb6Ok85ahELHiM3QBFmLXilBqQwR6bcvu87lUBnUzOOuwCLQcsbM/79gChPsGQ5j0
jB3UuOBlXiV7+vXYV32+TdimYVnQPsvdPinlpe+AT2KhZpo6E56gb7GppcmrYtL1S54H8rnyeM0Q
LlVH5Erl9dxuE47rtMwNq+vrrPd6A6fnDXpb6MUrClyh/c2hZsbLyycIScRMBlT/L3HTzFzeA30/
VbRa58dWtUMQMSXrfag4Zo0fRMDGHJBoq77+/pnWa2NgoIljPLy8apf+3xVLXNOH7oa8CpublHPx
dMMEbM04omo8wKtfhxeHTVexFbgv4Xxj6y8NrjhjBEwX/OpoYHAtPJ1SmoKOVkntF0/CgpDfMI3s
p/DVc6eyyr6ln9IldY2GHWSfheRYgipv7IkjlZeLKccNQJvb1uZB9/51Ox5/do89ahZNbuD7G1dy
pGeoLpDz/JUAPuusKQPn5GH1aJqSWE6tEmcDK4o1PPW8zHnTvjnmGV9YcDuEUlvAaAcMhhhb9nju
1LUqpHASgr1p1z/aU2mSyoVt065+X6Fb4rvqDcn1VCwoGXs2NnIbS6G9r4tXJI4Ie4sbPKv89HoG
6iWNsHHdif3AduU2sfImYEVcjLXNehtOcEQdSel1dFbx548gNmwnEQRIads3wT6ohan/Bznf7Z/I
XT5tCcGjtDRlqMfZwpG6MRSF+yq3+MSu3HXHcPm0OwF43LUk3cZzTH35xVzUdizwWvOkZMwfyHTV
31yESCodTfSa6BSup9Qi2sYrArQuhCG3kvk+0NXwR9ZcBRxnbzs+G1s1L8qashth4aE/TEiGju5u
seLa646/PEhXvouJxU1jqRvupXvPefCYrCSgS9wMlA9k2iYTwYQH8ZRM4DzjjnMq+Zy24QWGp0WT
ngZgAwghVBWFYABRAOHB5EcNfE7CgVWr8OwBN9SZA5RhJXn86iTUXxu6ORIyMQZrclNdExklxk2o
O7ErmEiJd+hhPsWTGk2jNcW4LFbLOo69aIB2eRpJDkjKnwS870ACOtcjVWWemBbDzizqs5+509Ne
+YuXGLXPDeAv0BlEiV99KY6qKBdhIF5pnwbV8ZZPyWPzRhppcsGZ1Vi4Q8JDLZ9DzUl035kdQdij
ce0QFXGM5IaVL3NtqH0uSq7swmYcJi5v37t6w6WEKLLBUmzmZ93Y60pWNx3TrwtaiYCPJ252kJjs
lQEnBhUI5K/BElmnRu/QykPK6mY/CAfJ9uUM/Vj6GJu68Xmf8zhx39I8dxEW8PtriY8zWxtcGiv+
CPo2cI+dz1nSrADJ6/YeUjJEpAW0HzkQeZvZJcM3nb3PJQJKK2wadNPt9cwI5dSvvas6UA0RpieJ
DstG1C2vHvHjZl7yfV+68em2MjqRvxLJ9d+df72243JS4+nkqukYu5e1ZxhMQp08c+JPLnj4+Rul
4ObfD9jdIaJDBlwpvanIOSVB7G1iRNTs5hYh7pEP4AIg5fCpyuUJ3LXCdTK7DoCUm+XfhGrOIAcC
2EEmDQ7RkBmG7ALEhSM1XGZHcPRGviPZOTIkMg8qevZx9n1yRiornka2Vk+paYh5eLJ04nwLSh9+
Ch+kaK13Wk3N6aHLCq8e+PiRVqyi4mYQPbqsMlAQ3RZXLar6Fb7mac7SHqdKd2hf3Wyx3hWK3eNr
kyDhlVRKEc/opTNl1HdfuB5OgVoNWxzhisJpSIzKwhNpJ+tn/9fbaja4ED36xg/meishUPAR31Gf
JVYDpeseqO6XYrcrnyvfDyjR3llQ5bBAr1pgEDRHwlBuIzicu1VqIe+Isfgg6vSy74JWBAHfweNc
RtZBsqWZMXEtf6f5EZTmxEJ0fqX5DhKbS/Mx+BLZYDHfc1duUtbqheBZ0vi1ZWM+r5+ontg8Mw/j
ODIOY4ejXITBLrudLg2FIpUNLtkeGdmfNAZF1dWkiQND7Q/jwSncc3JI3IRcVr68bSR7uxfzhEcq
THxtPTsaGT/6L2YsfLUR5F3NL4rsGGsK3Z9AZBRtC1Mh6fnv5VXO3YhZFM0CuE+qCKWmwAV8xz2o
qJFscHzT7pOEthZKV+Z/Xzu/Nc+uDklo8YDs9FKuhHL5AMcRVMFMERwpUc6qYSraXQSuVhX74qbb
8W0zqfTotwqICDw5tEkdukmsx2T+EeCnSKnl1PcHVpigZ7Ta2f2JFex+O1BwZo9KUiltnSeqvIld
Phhdwki6zpUKT0m3LIjh3HJNgLW6Yr7IFjNSY9eb8tSw5HY09zZfIyqQtLe2RNarqZQAlJBqW55y
R5lxjc7vsYoA1nzul7LNvpLq1mi43FTMA5eeKrKAswIXlFjXA8i0E5x4NgrJLilg5OMiDxF2hQC8
aQnyNDZziyE4mp6zwf8VkztX5E+2IaRaNYrsUhHdP0XdN8Ije8gAIuzFgoCzFEUK3AMigFAXWMk3
n5aWfqu+IPpjAbu3tIzBWSP68ay/k0O5nrVoQnoV3LSKclpT5Vt9uknUQqB8Z89IotH0TWYPfoEv
2mzsHt/nZc4TuDXKIndb7zTOONgbcZ5Q9GpDeBIqaL15ilNqXdnIUTg38UO5PIUJTCg4pdxTyUQx
HXXV1z4ESlfPU5iTcLbaYai8EBK9ZuUMSMN7hhGwhPKEKcUxSyZMDlb+DGH9/fM0eCGG15AiEuGJ
4wtfU2kT6+VvuwGEfSI4RQESYhlKyO/uh0Up0ray1sBYWolw5UMvBpuQ9+RgbAffpTrltnMrKQvp
pdK/9C4wYHKCVzQqU/n4eU5s9UQFgDjA+v0D/eTmMpA65QXEJGPDTb4FIufINBGlT6l+itQ9h6aY
0+O6szHMxSVCqNpF/m/+F8qHDrDVYAKh0xMRMk++t9OZW4X8b6FKgTufEUjEXnP/kZ/raOafOzFT
wMSd7HTzamHi3NFXI2w2RBdxkL+OFWrHscvCY23jiV+JxTtjawnAQ2n3muyyhmOFq84+8Yh6nfdH
WM9y2C7sthDGfClIEMClMy4WwwlCDskhXy4HSGMoI2vPr9dcPk6hHtXK7Zz+Kvhe1kPcc9HkfhsX
c+hMOLevyRkYaTHHLGSU8fLdvYp1ZrsImwXU9fyBXRC7UNgAHbcd57YAfJcGwdjH/IlKVCrW31A0
VSVkPJ+W1virk1vZNgFW4rYnw2s6fV6/fal94KEGNHaFgD+3l5Q3rsyQHAF0MEFWg6i+QM0hT4dV
CAGQK4g7Lacu2kOng6M7tPedKzOW0A1b2oBKkdT8DCoR5DvXb2rJkqFtCBqRiqBdCceawJn176m1
PAHvrk4GUDyO1JjKszswbha7UQBOdfesMYOW0YGlc6JZIIQ6nT8gV4h9IzK6WJqyBkF7Ql9LFY0z
Dzt9Nf+37ZIHWAMYP82Fi3lMbEIl4KyYN4bKjO9D22CavrXljwwHw7G+VYbkXuHMT/JXPdW9KBJ/
qorCFN83iJqjdjqMlaS+i00Ps3r1iAGU9UeGJJJ6ZpNp2r4mCbvZk5dHOg6AaFBBDWd2SA4aHdff
ct6LAEnuCANS82TDUhLfiOm3JmOWn8WQ1PUB05TtCctioX6SFyJhQNYM/c3FVHf7tVPHc3DrpI4W
wZnLObvqKaZ9FlPVIZ0W4JKk0icMZf7Ekgs7IBK7ALMtDP2MwmkrAbl+i2Yk4tlMwMVF95Pi+X/v
CxMnqzqV1C0JRy/xOxImywWefHcdlmgqmqT0KB4n/dJb6xWExQFBvvxO0zAY1TEo9u/Zj63WAa23
P6tn8ZCUa3ZGUkFaxPt+WS3uLhq+BUdE5E0kFThqAlA+QvwLONGo+RS8msu1h06S6KOpGmdayvjQ
ud1Ob4mUQT5Ce+loqFDPHuApBYkXKKSzVEoMFoKa3Hyj+1dL/qaXrfEX+JnkC7UXIHE2t/GXVpRw
c28KeyijHdhvaDGvq5p2e3c3MhP2VUaJwJsYflk9CxkJxR+b+9OSL/oDNmtrNtLHfVV9JttP9vog
e/6EZvmB5ri+kFMetiJbMGNNNxIupgD6HI7SakhZnL+2FjbM9Yk8NlbVTxf8WKMUQHzjdOQHSBk8
ABZFz7PLBto63ncZXlvnoIlzqOU7N8UZgq7hc6WF+u/a5aJuGovD6izJXYlPeQiv2mpXB2ZwXw42
dJXxA48jlgWwhvFDrW8yAyKb2dcP3ADDY2BWxc3ao41M4jtZK2iHm58MBNB0JYsL6EoXjndrqP/I
ARukprVPmz9CS2Zi0IwFyjE6yL1J82CFlsWgvcMO7kqr2PrDiMp/atDakS93NGADJQmqzVUbd5bu
K+qX5Jc0T5UsfIZHT1Rhy9hGmoFbr0LwczqvomZhE6lmid02wAbYiwYu+ovbfJhWZwAf3Vny1SSL
r0O4wBrHeWC2h9VaI4Vptq6tYF2ic0hDHmhwXGjweeh2AK1B1/0tMiF0+dBsKQnUY7wLUJx+MGsq
Kg7V09I7XZDVZDvJGyOyXWEJkbYrMwBaSUSCF9PKLe753h/fwzYEoTXXaEiD0gEFJZOBdGn3T58G
P8egQwtGtDClsnI+gNl/FYI7akLucxz7RmGxVCfDvYxd36V8JV3CRVkxPhVz1kxOqp96lZhlY4KV
rZ04mcRVTfqQwdUCCTpU33AP3VCfPR2If9s4nu4E5XCxirfIcTwbY7h6L3Ohnmh/D1GfUHflDhw1
3YGpUA6GxEn0oNYocZ8j5HnVJQrgRoZFWHNdVxHFSzfBW8I4ZpQGdzOBlh5W6y0ptjgDQBq4tujP
Ideu8L9viZoc3d49JZOZpneEFpabPuLnKoz9YujeZSB9pYpmh+FtbaCC4B3qosI+yXLhhbVHtTFl
nk8FOpZ9Y5Y2fQpceaOc7Y8n9uJUNE1g+TZGxdIngp1HQ8rli+g3Mi/9WCy9/ch/4aiMLxVCXzG4
aJajfKKuK3L8NIo2JbQIyp3GCFrS5NWgsWJZHkNW5dy+a7ABi23D3ILJ1qkeEgK5JrhxhFF3/xcU
9qVJ+YwKT9o/irfW4rbP/bLicEhlHViSL3cEQOROFNV8iFAfU/GixtWHgqUsujLkoPBxWsxdYHcc
Pwap8ErOCRm76A0b9axHGxfpFUf45VJ/C3I60HbtcwRIOCcSeFxqDLV2pLlWGkMeGB2uo6aGx1Im
4kB40UdQj8uLrGrXma8ohDhmdiqRsNWDnbqCDhnrHt/X8yqDH/DxZvUXFqLO3DOiU4rvXbKH40fc
5q9u5jj2XTbxIk7QGqnIcX/q0qYTeS3oHRjeF7LDSXGQGuuPELXKHPPKkHSHrw/5WYUwU4P++pWZ
+kbC7tAQezAkLrr1Nigdk5SaIyAZHaqvk/LsY1WIwd0+oqcl/z/34Af4gQx3H3vS3LhlJTyrSYLb
dKlNHH3vpoeB/1hnL1nS2K+dF1ZWaxjuAhvcrU5LlHH1BrjHtCUs1grJ0hLjueGyk+5A7o94Az+8
b+hI0RWtqkMkQuQFwDoNysT8YdZ7DpBzY4qEqxjAHY3ywON0pV+h92yjI92od8FQdpLUPh/DPxjy
Q8MWtb3UAEvoxUOX/Ko/LpX8lyVIHQq8Lka9SAVY/AqtsP23GfFPQvyWT4V1lfDZOaUyNNeeuJW0
P27wFR430MmwLUfv0TYHy+3Ak9Uz2j0LROqskWHyHYNOWguaLnhHSw/1PRt+4C6y0dgHfIpXFgYC
JSdTUqCKJLt1AMeh2kM0A7safAcHuec1VWz69/SLIPBRa1nZCJhDGUxy0AdE4x5C/6pLt+Wsiqtf
k6KvkjMNh0piCJFvfAVxey0a4PsmHqYSwM9psJBqPk9knuPBK5bhr2S0zSXrHH/R796NGiaEd0eM
y3CYXajramEdbHd9FNrJb9TwWELn2nnw2MFbGCqX26QO3+6LOC+h4Zd05GL3ZcX1RYQW2Wp4i0fR
DpTCzuMP63bBy6xmXwN/0vifXh36HiS8AFBCBDGf8pghZ64VzF5+vGPhp7qnuzU28TzzuK64zVHh
lK4MFGODRRhmvg5aujxBmAWIaN4T3bD5ZrgIGoAomNRA+HH9Plf7fYwKs6K3U7CY/ukSiVvNQDmc
i8fl9e1oDNtGoVPbXUGVXyfJnEGO+htXheOA05pFEn6v2PXOCvkb0PzA7Tk3sTQxrYMdslGliTIP
mRTvHJ/37Hg28g8cxTzeJ0q2m5uU+8y8zlInv11VFtrPZxp7tIQuS6tqg7GEdcS+CuezdaaL09Ps
VjjNtI92r1o0K5X2GTjlzL3bwS+fgll2Ik1B2MG6Rh58ukm/HVZY9BL0ofJncL31RcwPOZrfQv/b
6V54QAibjkCV9/KzDPs7KtY8MpvEUdRoM4YNH5tgC35BROgllY63bUBbON6DdR6C33qwSqfm+WeL
7qgCG5C7QpVvE6/dIt2Q+iwuJAGWpHwh8F2vAmwTukT4UegWGUtHO31X8maB9tkcYYF1sTw1UYdV
cfwyhPnw6H2pFIs4/9k+sJ7yV3G6MfaWPOw0k9VtQIWnmU4dPMV6a5eS/+QJTA9N++IPeu+mem/6
aUd217eAhXI7RJszcGYjxL5eVYnPVcrEbU9owg7XLAIW1fo/2eNKRN8xbG17uuNaOyB6H+OCpNi7
g1ze2gAe4KFSlXj7sKgWfY3PfSnPMnoi0e/SytYo7ZmvuyE/ZTK0DxFj/lHLd0z/A93g79USiTo8
sh+7Q8exvU1fetoIfRaLzrQ3yioGl0IyBOl7EOvRyZPy8uu0+zPkKZaDnhoxBs/NQOd+87NTAfTE
uXtNQDd7q8f1+X0+I01jnO89ABaaSVqCMcvRqj2wXp6Nj8Clu+Ee4JTwx8IblqlvC/omT92nYits
UdnHkNLyZz8ghFhA7gVyYCCdtuvyWH3yfBou+8tX5c3Tl+GVhIEb3MFFxhUAjru66mfq8NvJKH5B
yyQyc23yZ4JISm5RuuIrqlh++CLXbmcMlZA/Ps3ktt01yvOHn156a5fBxY/R98y2X9IWXWLJZYag
ettjIcK8ndQxk/J226ihd+3RtgWpq52AtWm22Ir/jzQtFInZ4enoAM0yEX274CGpoQdIk7Ds/Tcg
nmkq+adjM/FhJi+oCK50w9WWIBD8qmeFgd3OazDcQALey7rn46OZIkxcOWb4i38Aity+HgXNHGwn
sS1wH1lYQH8uLD6XSzKfvDN3jtaCEbustFqNzNg8We+2OCJJCITG5nxqi8xbNSYJ4wGiMRS00KOH
O1KbRVg3f0fePn/HGYdf5R054yuJzZCTytWMzRRLKOcfs9n20JWvHn4wUCgkkWXG7/hdiqFudwVX
FACtHZoPXpgae7htCgIagq0c/IJKxYaMZPXRTveAWS5xc2MJq5EdOM5m2+7osrAaH+wUDZXr11QH
vzfBJlMIQige+3h7/SD6EGREaWpxNRElXTcs1mXTcC9Hn5//QGtBmOewoHVWKgMtXgpOPdhmQcFH
hP87mTVQp4qRnenaJX7j3Z0TvKUC/T2+ZJtVfL9fWAbGvIcRQqtwHedcA9eZQ7cvJn3LJ477oscv
iigaRJc57SCxPSjdcCINA5i8bKisHKTF0JROPyFKP0VXKsZ/a0uwjVWT0StEtFMagHXaE8nhzz4k
/tr7QA==
`protect end_protected

