

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R+TTV2BAhe9Ek8IveLCAIK+vyB2qa4TorazWyGCbrxCKkVhTBvAD6RqPeP/JqtRuh2zDPzraR9rT
gUyNSWD83A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XM2mYTm+gCT0AhW4S5p7IlzH34WHm/fa2tLSENK5xQp44huwLBqk+dBcYbe4GM+6wqA3pzoUNE9T
SluI3P6DpsOt14ispiaJSciB+VdlU+Q0e63sKyfq++TGO3CTW5OhLIxojUbYrTbdY4WbGkk4yG0Y
qGwauBBx1uBueCA2GC4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M9U+BjMD5E96pT2zTDB1OSiHn8IS+G+aDNa3MIF/jeClLSPAOJwufjuzRcyAtwx0354Pb7AaFOwR
6CcoWPQM1dcUC6avyG/0PRrtZP/KpXS3/9PiWsaFHPYVLfqBMCUDoraXwfpfMxmOy8hD0iI6TtWc
j1xJUXVsbv+kqOeTUloYmwdRx/8cs46FvZfnFpiZXMFMsTsT9zvmCyNxiZefgFKT064BWsCkg2fa
W2IXperFJQzpE9mXVwGSjl6xDUp55esPyEPcDI4xy0T+q2KtBQj2Qn2DJRZ8DKAvjXNQmo/tbweh
l+RGgbFge035kxDZ/t5pFweR/SYowAMdG2yOwA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
absLoVdCG0/WeiZ9M4NtAUjz+XnLze4vahkoVw40DL65GHoB/ikdBh+LyLQ7V3LckxaJp7Ihe1ow
2yXZZfuygvynBc+n/CI1EDwjo64cUTgVLg6gqySahs3D5Xkp8kFBBxARQmdoErJqqhefej6SXrxx
13OxNfq4vRGx7YG4l2M61gUhVtUX9poQdq5dxitmrLXD1kpdnUsj/YIpVBaLv/TBn9G44WiyRNIK
ojx9q2JyYKiWBfcBh+fpJV9PudrBUPMu8kvWsRizFr+r8Ya09D3o9iJUZ6FWOBiFsidvZNgmp1u/
nv56cp+qpaTesLtwmKiZbrhQtq6YXQvzPpDQXQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
t2oJ825g01R4DfbjT3g+VDPmL9PAyVC2t8Ozl94Xb2xucD77bNiPcvutyZFkA0lqWfRMp8Z3kkTE
OOo/FpGS3c1SP04/jMKLZD9E7DL6iVBRfxa3itPHxsSD0RAP4yPHw3yCiIsmB0q25x8+so3h/QOv
DKZh98m5ku9UnG+pY6c=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
koDeaCPE+GNu9rMKu+nnX8UvNKbOa7mKCRwRUXCmZNo0yL7JuxnKQiStr89+6Ws9bOIbY8P6XKLC
WoSokcQl2MIZuh7gUJ+LQSPTB9HIkHPuGGPibAaiYY3e/6TBvv0+QG5gTvuf18Nz0UQyxRzNBFY7
2e0fNw+zoh4XJubbVaqqBBqTNyIM/naqx2G+DBhvJF/RlcpsJUe2eVt+uttis5ukRD1ndenp7rvA
+Ub6MDtoxunfFJsXEQ8QZkuZiT5XfcmJdkquGywSafJqKksYNJZpGleQnak/ePqKq8cYIbfpqOo1
MlqTFX2khe/WU/cqsW+5jXmRAgWueTOvg5hW2A==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wZaMVki09KtetQFaQKbOEpc8bkgxHSc8zyuzh+dwZ44uN2hbx3K7ITnC8dDkn3EMZGwk7C0u4eBt
eru14n5jQ1LfuUg4cKuwRNAgFxc7GaymqPYSRK9OQZHWZ+w6Alh4X9YWb6UVcsv4sCJA8YT9QeZ2
8PJYA3L+OY2t8Dcx3JcdLeVgMWDrP/zfpXyfMdPpwgBSSCqJHFsYdlG06onoQq2DDJ/SpC0W2oHU
JJAOTss7Cf3giWx2XTrorU5k4KbClTaEv4QAsogatkMf+oa9OfJQg5b7OUNbNqSzTV2IvRXtKIBC
N3mFkAtau93JXZzbow8bF+Y708RmUyIR5AX9og==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gidhQdKtgCKZpycO58SKONz/x64JxoYiDvm7CY7FhAgR8N3zqVR49qh/d9ImLGjAjXhz9ISSvhiE
1TpzIsqbVIoSEHhHCsw8fW3eNfjSKG9+5c0qMghoZBwnf9txWcso6wczPV8wSYfFgOnId+/H4w2u
MtSdrp2j2HeGCN7hmduXDeRIcLF+ekxNNZVk0wscD3yxYdFDWscebLgM1N+Cx8uwWvloVVe1fNSl
IBecuxue/tBnCdqw10D1fC8gGorhdNUhO2bTYqZL/+voIIAXkux7Z0BGx6B2uSJYuZ0j2LS23yyk
r0QDrL3YOpbEPBbFhTy9LQz59rkITBRhVeBqVg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lv7TtlI9EkMH+4ifu40NSGcF5VLP+fQr0uBXzvHjgpvggoEPEBlbTyXFtewlIbLNuHO4GjqSxFa3
oGjcKGgjJ4JKEHh9NZ/42sDCCnN1TS1zrfhPhpg3aJ3aGsOq5GxB6oAuNGvsTC7HgKk9lvgZfAiC
9ubfhd8fCUCrbS2jYuGLkpNxtwRxEbxLfMa6l2yusSJt8g6sfH0aGGBJWZjKnUZ1SyA1DmzZW3ox
o1AE17uwesEX5+JGPaqlsN+jLpbHhpv24GF4NS806LjJrXOO9qXbZScc78Z/R2xMBhLYAC0AHR8o
o8hlz9kYq3NSGSCdEMOcxNjVxDMYBrdZ+Lc+ag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296400)
`protect data_block
Wz29/u0PWPYi8wFwXeBrJu9tlDebMGVFejp6UJFlBFcnMsap2a8Y9qROJVSrdhe5Yagr/HaoNxPB
4sbk5Ebidfns3Na//tAFu8XVI7DgD+K0X6GqXsTdIqo9Qa21nYtWNi/mt3neTlBuvP7naC036Bw6
Vs6xN1sfTkprWy0i5usy/kQZPekOtksLDlo2tsLe6DaahNb/WgCkdoS/DYeozfANJ/a8sowwFXAV
LGwkBTN1fhRjC3NXxzGBitwz7niwivGdGAQA9x/gWjY9lrxg+NPQ3mTmfVOtuKqoi1u3cdxllX7J
jeVyaEpPr5lBF0CHs2q/5nzzp1A8lgBRZ5qZ4YIxAWHtK7Ky9LXl1SdL1zCKvODhy0/9AHKo36hZ
mb1wq/j5z/9eAqcjMzStgt67yyxFtfxWCGxRaK7F/cRidlXK4/qaLkIi8hWb1urRi4ecx16cJzUZ
7Swg21ImWziaWX2BefPvjyhB5VraxpWamqpsH5c+gCly72PujRq1lqxuu9x2WS/KI9Nhl7sBzv4y
2skEK/67sQspn7MWtRm/x+7Qjneqk9CBo25mGXg9ceETCRuG23o/ccSH6Uh2ua+PrAI7bzxXGEAD
Tbe7TjXAW4iID2wnIW/Llk9UNmhUEsUoy1Oe/qUIsBF5bmLgHvU0b4M7V1cIX6wI/oBDC5ksJaD9
01uBn6Kg9AN6VKnnfKH6RyTHrImlVuQl+00iHyaarKF3A4dHYx3CwK8aAV0p60jJQfIvcF7wUA+V
md+eHZ535p0/Z9TtHyDGOuWSwM1fqkbg3YGu7ahJkuDVYOQwv6TfAQqncJH/1eJxg7uPpUMN/477
SwyjSGs3A1jOqs957U+uqZNWNLZYLIytVNkjlXnRqQcBWRcKA8fRBI/DcRLJWz1tg6JFm5BQhat8
H/zF2z1v6n342RIQS1TdNjdSi2+0c/0l0DKOtDG7FMhJpJLgI1JOoVtrEEh0RbeY5M178WOMBWn9
mwTyTNZbOxwhP6hvNMgJx3QWOysw+S4d6y8k7P8EJMGQCkfp7bU2NLRr3p8lqTqLeTHkZnfX9SR2
ivsBxXDAfmjpeSPNO0RE2xJaPjJf8wjyEWloZtXGCqfD3iND9P5SLYdYwUfxMQGU0DueImhZ6z4z
CTHG7fFfdK96LB4FmfN08sPPLqfbpZxj0bVP22d12+6HyKowkrJ/j4D6H5h9dq9yZRrv+ZulnCer
MOyFbjffcsUZDfcUB6bMzAHB/XKrPxT2HPEhtB2YpY/T+HmOeetUs9s/4OF3pCujjM2BfsozxfVR
8XJAs/BH8FMlFgIqMGDyFG9tqytBgKPk2rS2Apn+usbpO5sA/CbGe+WNZ0BdQBeA7rB3y/ykU7jI
x7xue4NCEoV7j+tq4YcxmjbKl7MuZH/6/jc+jGfV15nlen9S8ar8oX3LlZQ9iW0Qob07oaTef4n6
3R+ZuRF2/X/SbgSElFPvHxO9xZTBZOfhpUrCw2GyKxySQoFN0qosqx3a2ykoFQ7BSq58XOq4h/4C
u+4LL12JL/cJspBR7I0z4UoYG0Jd1zQy2K3d0vy3cTu4AM4xePtNean/xW1JSa6SlqM5J6JejIp3
0/kAg4DE0Ok7s5K4K9uLZkTqTP3GZYZ0N4rH3GQ5xMqU1bg0+lmzPp/CqzioV+FG5oTJL0XOJU9Q
Fm+RZId/y8bVWmirN41GKWFDglEXA5P1svp/+z3d9s9V1AT6xoPS/CfGxYFjyUZYmf/ILNMMA+i6
ORQen/4q9bncitzQlggngYA9e3q1JEi7Rk+rL4Umo72qZA7kmZ6YnwifX7RHTB5/+5rh4T2YiLJw
gcuQeRa4ALS8yStjY7xS903ZZobvy5o+4I6qK+ZhrzScoVugcNkETkANgMbqI5Q7sHtmrRwuQ6W8
MX/hxuEhVeoeLibBIf3mELfVgE/Z8GwYqNABHIx1L7aawaoS8z31tsYGt82z+91kjCZ3d44MWdug
esmwN475LBKWSNN8zlC2yW27dWne3fpPeO7u28/IYLet7MM+n/mkhi6kPP5yLSQB2ZgMxAU81Kt2
3Gm+bC/vIYvuJGTMvyrfGoRTy5SZZ3lUPxT7oG14MohXnV8Y4Fz+3lDp2k8SIxyaYrHhEbkjZhWM
UOja/7ZJFn1hWAz58lh8gY9JOJa8TZvaq9sv0kkmumh5gnSKOOobXhFc5wkAztYZAbXWKUrpyKXi
prlK9z4PSi8lFrYXmmTwtR1+HbzMLjs4FvJSvsnWSCL1hqf8gu5pLOPzReO1n0YXVVEMmoB6yDli
0KhxHB8Jtv5B8xnuLxsT+rklJvQvu0VzqQz9l3y8THhAjdHMQZcJs8enaak9PmRNj+84qAWqi3bc
zRA1HmD792QwAfQtBB4aAT295v84lmmkHZWV4x9XLR+hPLhpqjzg2a5pGuFw9PhtNuGdevWkUJH3
euBJLCOf5IiebHO5xTzLJvBqiUmBJGgHDwIXaWnPlggsU3DaAYoBHjteP4ByZU2L6zYjl96jcgwy
jFIUIhWB8x1k/qrKblWxM5brqNZxeXw0Nn38ZU8eqL+OJYrVuS/83qUtL0Rxu2atN/ZYNfHRmcdB
KLCzXAT+iUyslYkCkv7h2P3vnUIs/Pvk4shwjuVcNg0xdYfXjQvtNmLKD9IQmWmoQQCLrF2H7iet
VNeWYyXEV3KLxC9j+cWA6e1MbcdM8qQghKaGltdAjgmXpNpn27X7TLYAFR9RreHX1o2cmlt/29rE
lE6WCyI0uQdlCn0oUbxFh0qPO1LLon1diK9CeHNSMkqOa/y3pBQrjVLzr8x/TcYqRlnOti9SGCuP
4hXeaWA2fai4F2q5hFLteNMskOHlJDpWXdhCiZ/YNNxdmzc5rXyr7o9++pwPO6iqozrRy8jF7fXd
QiEB74vQwDfCgTHkF/iEeJtXWz3ADH8Npv0kvNOzH/f+LklNp7G8Rgcm90cBboxcLgnjK/HABBQL
Dkd3eEcQWSLBcWPd1v2ZDN6O2vFqvMGup0SCx53lxdH/ypSIz6FQ2c0j7Vw4mdncme5SFLg3wR1O
7dXB9tv2LTC1AggQg3DcGRy9zPZdiXfiKX41WBONzExGPh0SbX/PZM1UhlonF0Vezz2//cFPnVbx
iIbVExEjscGVGo5Yv/WaPX8vLvCi1eo/JoW9n2F99P9CFE3L8kz+MCzJT6OsAUUb9JZT5enIhy6s
VB6KZ+fwi2rSSoHVcOFYANSGRniCheiBf1C/1dYvSFOjYlGBQBbseSZGo8B/dOtviJT+xXAerA/t
HZe9HF0xGXdm6n7dIgYmE1Ia1Ry6JoK2LCvHlMX7qRXRQSRzoJIIFeT8Zc+cyQFWaAKvuPYRK8b/
bVGa+xxkrpvyyt791eM1MXDijzShmk+5mv4KRx+khesWC6frHotwJohwTYTmwHKTwRphQrN9haMs
2SOW+YodI4zgSuvZcpOgI8AdLzeXPfmLzjg2RSH4ia/3GD0CR7BNh7G+QqE1cI2YT9HDBEb9MTR4
oVmM8PhCTN5iu0rJ6yNxUd+u9CxFSleJRWe5cfP6CRF20dMifYAb3xgCFVEqJz2zOYGfm6HP/+a/
dX0DEEhhpDoKo7/Q6Fgn8wFoJu8cLhiJZGJXPLRtFZ5MHDRm9sYuHbpITNAmodnL8qw1MbiJUe0Z
dAfQUnZOTIh2P8enmE1fJZC6VhNCDIA7aO9ety93skdakbz1ePoQi1vYju/v21bd3IWP/ogAKDvU
b1EeFZSyGKmNZzfZrvPtT7DWk8v4DPloB5+xM00iWw1ABf9jBMPcJkW0Yplwqa4MemM25VWWf0iP
HpuMU4QLGNLQo5s0akFLEQrZx99cy4xKS1AbmwjvmddWtQyx7Ve7IlRsnjOyZ9gF+uxbYa1aX05J
4axq3HYUFMiOSE+SaBSjPpSuOBJQrCV00x0AOh8VgCykEtGcz52IRAIJvW+enQlUk6HuMFN+svMp
BApT8dlxeTSfrFgB4p8tecjAenXLpglpU/ADt+q8kwY+wjYhjCi7GdWebhaAsqHtiLUKp66Vadx7
fTFPOA3hkJiZYqJmRiIgEG7XF7b4WDSw8Ycrywx/3AvY9dWnfLRWkpyhDQ5hFYSDamIHoIPgAV/c
xz+uEEX5etTua/SGFa6CeCvggXAAvlF0rCWCd1ZVT2ZibXqZ5x+8YMmLGkfn7+IvGxqWefFVecIX
Px99Pi+t7uUtoD2WMA9Keat18KoUiSiP8K8o9Lo3hVaB4KuYOUoYAbEp8kM5281Tch05a9rJyM89
meIy2FMkNUgyyC78Fe+v1FRFim+UTLUzJd0PdOY9HAJeqJKpAChbg2vTQaVL6rTExZM+d7HBC5K7
bhZAWPi7GKAFivyAkmuj2DaSWA8BcoRmQjUs95m/IMa1c5jFCI0Sope3pbMpZKqq9pu+YCob1ub2
KH5ZrTWauICrAjyG5iMGMfu/HgQOg6yzOHu0vPaJrsqvU38V7TDJEJtohqC46YnZKPdhYHGktBpv
djZeZ9SIhir706Q50QWrSut/mMq1uxk6usW/Dsjbr0U8B8CaUQxQ/b2TWc+YQzfq7XR6qRqp7lzm
IWGOPAwWwTC/N7AhAy+yCI4txa3L9DVNSr8arsQVQpV2og2tRcSMUftuPaPl3nYhhDVBtxH31Bg6
8dvcKIOSnsWZcpfFm4iq8d2Lz0qLP7aQ+fJVkbuiOSITQ+joOTL82egytesra+Ce6zM9dXOL3oJ7
4eLEXsdd+mUapWPDc4kBqag8iyEY664nwXCk8IPXIXB2ZsyE2jgSX96hVb+0dvKnJI3KIF3ffAHC
SGeLjg3BsEyAN/27vxFixOrRXBGb6j9uNP86KkufKZ9SAt312+xLnpGtIv6k9BmDkITDNtVIMzDa
81E8IB9hts/au9EFOGyTjZxLMi9TGLLcFMHcAe2KKY6B9nvJYsZRAWWgSj9u9Y4fn7/nrphygwC/
xmmUEkKpCxN7dy4zYSrhU0CQSSZ7qFXVsKKHauTn18NsuZcw0iKgzN5/6lMEH/lQcAHhF/pPdAzQ
DQo35hULDPxghK1acZ9bBYk+LWWrTKL6fX82SfF6kdm5GYC4Ny4htgOpe68ARpdTsCr6I8yHTWEL
N027NhyE8XWk/NxDEzX28oG8cJptmUkDQTeu73VcPX9jXapf3KLvrS3vwkeHytw5mycjn95NFiJ+
5/rjoMdjrti2zwBnIR0I+oD2vMsSaMAKQDEN9KW5V+1RdUJsxgd78ZBG5ZemYY8Tr5ZquFyH+wcd
JnselxQ1ASgVpQ38TE9l+BskYP4sX3VhpAybYff0lBTDtaQslhxG2GxDi4tO+6bEhyP68pROeM/c
K7rQ11aoANG77gL6YNwqcQYENvE0+bD0eOkLAEzKO5Pqkdl6S70LIN3RB8jNQr//gIMFhguSVmAq
SYFb+HcXy58zIYenXa2xx9VdDmwAK6VgLwgdmtJyJsSSwJ7xiJlmp6prMLDqNTdb8/LQDvJflT0P
z7oBNzYCdvBU+C9waxPtVQrL0eUUbyIMEJ2+0ivYBJM/1/XsBGCu819wC1zdY7Idttbh9/VtuGP+
KthSZUVNgk+CQmuBVVfl1jDQNzKnKVhSubYsfyEb/+8filt/+YL2j/4AYUbSeyC8UkvhuydA3Zjw
iXj4fokZEU9pbI3hOD9H/m7VCq6yfuKxGU3o6/mObaOeKGze9Na9EpRazhqeoaXBRsmLVCRr63oE
5cKXliYwTwgZ1jnC0G/KY+idPgLysiOpIcOvDHbHxUCKOg4c/ma6JWf7Pq0G96dUhoJuKad1x0kA
08OYRrTfjYR2sTAhRO8oz15vYK28m0u+nf4GGq1Rhn62kpTcQUk14bGIZt5rDR2vOr81kFDLWtpm
4esOD4fKP39xzVvOkjXIlIiSBU/Q3ySV3jR/sT8/+HKMLIzshvFL6iCUQdejchBhJspW0Z0A1knF
iMIMBBK36UeEBqgRj/AJmil5YVdZkGH79LpTzEgFNgaOpYzOB37yLNlL8T4cscuw2B5EQqShOUQE
0Q3CTpQjLwl0DziA+FcVXB0PN4pIYlMR4dT/+9209b+WbFS1aF93RCoeX9Lx/Ak6qEV9aM+ipLGE
s8csNyEbGnfgrOgiw77djS7qpqUhcPVOyk80saeOGXr7xa/dsiGHswKogRMae17L6l3pAToQH5s/
we4W+UdNcXhDxJzR78w7xaiZjF5FBydR7NcBi6oI+2dfbVsh0YYak62ahUTMBOjmoYnPY5N7+dSo
PYJVYuoAtJ6bgu7hPNKNG3yo3ku/edoy/tCD7L+IQe3YsEF/o8UceRA/EnuKcbMZqJ9dsfJkhrNN
oWbcQajtdg5yP1/Ru656TjIC6y259QzDIPCrq7LokBvzV/tnoeDliHYu1408EpMZINfPTxt536aX
q5SX+CYVOc3Bz2ntPt/O2f8mpmDn34apKVkVvtDqyHX6IQCrC2xBL/BjdDRKNz9UsWa+qZraQa37
HqH1eMTLtDuHJnQGP1baovR5l+t21up9/SJm1tIFP/kYgBuSzgz4A7qt0UtCo+pwnrmCk8ys84MQ
RzpCEP6AzOhqNWkNKECbVuyHhWTEMoFxjCs8jN7BuIBg1qRVppjyjNPT0iUWpL5ICEh9S+UPvOEQ
tYjphv4Ke2nRfK6SXAgVaFi2oaPQbxRgB0mc4Z8AtGGLKDu5RqpTyFOqaZQ6BovywcUlmXLfQUlR
lvqLV7cw2Ph7fN0JN3cq8EqViftRVYiLHc/Tz4meU+Lt4UixV0Frolsyllpv3U3JIm9cJLmupedc
2whAd8bD2cfq4ZEgLrYykd027CS4QoDsnMz/N5y9O7q3wQKWyaYPdCU8/iUk0INl95a5kjGn2SPw
s/br7iWpo8lKDWS+UOCeC5uUjQ46q69Qti+valfvRQxlFdwRxKzgnaYxOn+4R1BVjtXhj6GioMDg
7nkzZQOlz7QxG2g4DcjmaRqNfG9KMIJ7KwafEEYcKSU6NowpSMCLooP3uwcH5pzGKcw82ejX9V5C
7iFT8AmmPQYa1qwXIIa0+kuNMBjnISHXszzm7BSfkc4CTTJFRF/AVYm4v0lkiwk6eE/99JVc9+cu
8tEPyng1SIgAn2Dblzn8XZRjuHgHJfwmlBx5EqYXRNwQHdFC6uXOSSX+JShKHSKjrdnbm4xhnbvI
FuRiq9hTsV4K0KTn6oPeRzPRuf3rpxYpaYsjn1Pi96245Nsx207y5gMSLEU2LzvBW1PpxLSLcdtB
yBuQuR+qr8lMf+4tvlM1sDa1BDH830dBk39fikLA2plIUbdwlM6t9rCPxqSl0XewZZHH0WPBolor
JT1Cx1mnvIj+KVN03hY3AX+Q1lM7juVhxS6/3oKr+vw/vCUDXjsZhS+vJI/eSJEy9Hx+konAXRCR
sa9fMme8GIUAgnY1bQAq2yDdbBq71xKjDRmUgXFI0sNfmh/R9o58I3hgk0CNXRco3UeBfeFb3Sbq
rvyTA6Rf/d59vlDWUP13PRsNaOKkcb3regh10dvNGASeZigi8iVAU6Wfyyq/vEjOJ+GKDX45kFkl
/H33ks5vGiT2A7CPGWbBErTzw1f75dRuS1p+CLmOXH1S+mR/JENGWb8e8iJbn20W32wUUpYh20CE
jtYEC6/l88UCeAyvC+zaZNqqupNOFS2xzrG9NzvWKp8VqA2Ly71YdOVgJe761dZwOtZkKeP44ChL
c+itSZfaBpO4LO8pjfbbl/+XFzEIBX6k3reHFg1oQUNscr4MCms8jMsygrHE+Ucb4EGioJdSNasH
HdlYFO++spH3hWUAz4vjAJx17KwMlIFJDWd1FF5GWtBe/3hjSOA+C7Ba5x6E5sVjG04vSrYkmDEt
yHj9qpKDdSrQZQ7/ATudK5Eiscl/Z+aJ13Xo3CXC2CM0VC7Gb1QsYxfnFh1oInkeqQ6bCg8wQoAJ
HF8pTaFqpXd46V1lGHTIdQKM237B3CobhwIG2EPZ6ZOLTA583xx5oTiXwsTxKdqmWtFET64o4329
k3o1BsfeZfKhfi8/hZnT4LU+8lvoF3vP8dGIafsHy0POz02tR/09SiXY9QcQkCTv9E3sTyHpvuna
CRV08vApByTJIuPtPWSHh+Dh7mhPUi00mYixwLBVxzmFTZniFiMI4cdIJm+9HDDeIURRjjFS5nYH
T6//hlBvdYYwNBIUE+yPbLGFlM0MHXbR3NtCqTnQAgaiIgl4M723ESNJ8M+CrzPbQaB1B17gcpWA
uwPcCI6ynUx6VyB88C4hMKwNcDvVY1w56NSIit2eNqcPDWyzDk3/LTzIwJup4PRjqqNjNkXFrV8F
qI6HmdkPROb63Oz/fEawMj5BPnPNjdheLYmwd5ewUr4ame/xZ6ZDP0Frk4SxORWZN0IDMd505cUA
zz4t5UwkOiNGzBqULRwuW7wMQOCUAesXnppAKreOL0pZOO9z6ayseRInCsAKDy28QvQ0HRQL945d
Yvq+VUOlUTXUc2rwb1pI0ANEUDNUPv5Kx83uSttF/+5FePqWC+CG7FQpsjW/zVhCYATj+WEdJUZf
vehEbM1YcnPK/BTu2tqdouU/WgoMLWmLTlCigJBkaEwpj2KFeLNgmuc2eGKtw1RcFs4x+9++GGH0
AADOylJjv5xZ4h7c4uNxj+OtqqkRJ6nIZvdNXZj67b844kTI934zqK2BnuB2Wr6Fz8v42o4yqKKM
g0SVs5UEVKclQBny0wCo3gEFHxuZ4Cw7mdSB5OZd45bUPmmI8gPx8NA+cwH5pXOnH55qwvNJNyfm
GMoLimNRGL+AufytJAUR8VS+Y44ASyHFkaP898Nfpps5v/lHWhy7osOBxrReFbhaYrWnsGlJnpZC
INBzvVEg3R3R9r7IoDXm47YgjdskP54/KXe896w8K8XgnPxGoFRBUkb+8HgaZmIx94UCF5usBjNm
XIuRv6OArgVfP0jtiyf8frDYZiFwwYdeTsS7kCNaU5rdyengF5T3G80ZjD662KZKtLca/wy3xzYJ
6vFIeDBufwPwQNEjMw48QXh2YOR912Igsobf24jl6QiDDOgCis9+/cLhTZ7ijGEq4HNx0oI2f7a9
1ncO6GLhkKgX2uO5TxHwxFWAaZITblDhmp3vAGsFc+6S9aKvMEj9HV1YH93w9BW194ep82VZtf48
SZDKyWt2Gj3G5amCmNt3hgLcVSQFyMOh9LGoSdHfsAwfqBze2xknjoQDRDIwsBrZ8bXPIi3OvQWc
nGo58RxfKIla+DklfW/DmpVDx+/bsMXAnaRDx1iQac8aA2qVmar1PP2Dv4mENcARs89ksOOE0/SC
i+onCHDrTULjQc4TblMVg3Mco0HDzJfVSxuVnG638++RLSVmsV+T1oGt6oHCK3/Ci3SNiCEB2j6T
1rvnuDdD/ZP/rfdmmSrk9Q9OMO37FolOuo9Brw5h0UxzHiFjd9aKBSEvZV8hVWJani4r6LsCuxk1
nu5QwZ+GxrEPy6G9ywtBlN4BHCVZan965tg+HGQjgHhPEvsQqHVxEej54QUIsDxJ7w23wlI/n6pI
uCvPcKwejUj5sQlYI7NrAsmwpcRg9uj2NrPXBR+lerInS5p9W+qhmXKgf3/YiYVVCn9AGEXeWWuG
JPz5NdmcDfxnFm9COq0BtwYLvtvyhOOuIIJHMWllyLFEulsZR1D9M3TbmZbQiaS5XAY1Zl+kkWQ7
EOplXWbSur2MtOSUO8fEqdnxvMG0eTTAJQ8PSqwJM5ZqVJiiA+UOIRkyr1sMdYLflm5tzNIHoTFP
kGMRTSMcpUOXEGkUZGq3IXMLgXKhkBGvIrE5td6+i8LPP4SAiycpFRrb5k+qpbSiEpUjMp58AwSC
XDftujO1FYZgiT/79NMO9Q8qhcKQX5NYOuG6zY33TpBS4q8vG4fUlFs4G4ApB53mLhEqf9KMmz6k
inMSmZNRNWgDxO+5uiRINhaVBrlS8EL/Sq5Fg61Mz40B8QGdafM3bAi0d0f5+4jouu20OaFil6td
s4HTcG3/DoIiBoIyjKinX5Xb3d94pXgjyfNh71jc4nPUNbgxU/f77JPP+HMMikh1g3qlre9LHnTe
0XTHtDrTrFIsbi/clF4XBV3igvjTDN2V3dKUVeHck0eN3TT2fNcN+Jc2uqiZO5/VT+XJsT8gTQK1
zxvi9AIx6wnPyAYtLQy/cBEF+mV8V5GSGK9s5q4ErFu9gXYeJc/7fUyc8UgES3G1nh3cvkxUlbDQ
ZgNGVEIAa0M4F9qosTbQTJ+nyjIWcTl0au35+5XcAV89Qte8pQ9O+wzpExL0EECi/RiMnE4p6x8s
DBk04xK8n3qrgQaUEEi20wyfhVVase/WGQ6M6nL6vSqqKqEpASdHxpU8T4/nRYgcQ6cetoK7DzkB
0RtN55Lac/1PifzHEKGKqPa95HbP2mhEtut36QEzw724i+C03xWZ242B8EyR3OeCa6107p7SkxL0
A0He++akDjoRe5BXfv8quxtBOpRGnOf3VooQvd4vuoLYIFomedtz00iVodcAx5wvt8VrbSMP/AJl
vkLJRKStCMik1POL2/NxLXjuWcn+XRZ+G+617tnoRoD9rhNG9tZMrB41cedUNsHYXJYnSZgwKvPh
JQs3VEds+FbYPRbH5X4OP99QY/3rXuF7HXGZ/yLXXaQ4RMTiD5Oj45omz+phFDlSxkWAT48eP/Iu
Jt/KQiCE6g5spzVVRZK6P/1dxzz9tgZBDdgErHaAml9PRDPTK4uirUaZRNxB3EIiCE9tHWNcg10o
CX86i8jjc2Tj8Rqz5raSeYCXl0lGeU5gIT7BRhvrbG3eMmWAkFdwblcZAQ9TTPGr7aEqAkaRpuPu
cK9qbqN8uaEJLWgtZ+TdbLRBsYb+2HxNZESaHnmHStlZnYr9ExehpQS7D3p14ludXLyxMG23T4vv
PzSfLF5bv1NzqtLr/I4E1Iij16rKqYkFCBjq0GcDVcJLoD7xxSM1o6ML/IzO0JQG8FP05vxt80dg
P/8nhnjwqsVv8z5VPMY6JwiNRuo6MoEgo6golPg4LhN8SVS436pqmoYO/y5I5fXunZcoBGUphThl
vIgPYIJVIiCo1wG4T/9cohABpqT8uEW13byo501b96FUgS446V1A2odnR+hxPOSDEl4pWt2VgXLh
NlfQqPvvxF86ws89U4/vLVnk18fxO3Wcyay23kdRuIM/rc/NWu+OcP5dXI611F6bsmSIvRW8R6Ni
QcOxBdUMe/QrpstTGduyKxTXS13B9ZNgjHc+2lvb7IhbSYrbcg9tYvL1w+Gzccrw7hhcdDuOupfC
OkEO4dfKXYHILCcZRsDx041bBSxSWSmpiO73S3Tkpi6wLQx/magAzjPTKGCVCAE3FNqwnO/lvd1e
oh5zK3/hqMvdY+dFcWDHg1lApM2OdDHhCqBboAfwVAWByhsR2iQousluj00DeU1uZPCxXwBzqO29
XkTSUlH/Pelb9kXppqjvFgA5VOItkY2GRDbudki+dZJvcpFLA2iOsB1jl52Ab2joBWThbSasp5rv
l8ij/vGfsruYNJy+kMIyAOoXpRi3cWseXIuJAtLb1VeAQycpNDthFmwSvjfz18UdyGUybSXwmP6t
Z6A4P15EEWwPeilRsVy4myOPBpl65qQatirvc/wqDglFYj+VpZFC7Ho/tbR2FZq4AezSy2y3Wng+
q7mCzPmykpu/YdIy1utfdZm/Pu1eKnkj8ffmHdG8EzjmKEZ3xmf6pXHBnm15/6REcCiWCM6NQHUQ
mS6TIowCRiV+OVej7LyXvH6Xa+cImxlIdsh83jsqdhibj0j+Ltig5QGz4LqT8Lm0KHfmlaVELTHZ
ujE1wbZd1zbtkCejVzqwXn5MOR6dLptdRTxU4XrYuHjylsfl5Wane90XF/ZVH1p4g8efaZmJrM7h
Cd5T4P8j3OQB1bzeqJzFKCMCAgsx11hKd/4UGKUuLqRL2gTwV1kIaCS244t6Y4iqESIKpZhxf4em
ewBcUCwVld/96lJdESpIw1SeT279N5UdDsVpZJok4eiBwRmNl8fQkUh1n0Mwke7l9WYDCsq5AOp0
bolonD6D+OKVNBL5VHUiu6LRIU70TjVR71vllUvngO2FtYIuEyf46UJDox9BjLMdvX3C6UPtf8pn
RYRbsdXLZIxFEvnwPN0ZuBlJBvqWLQORps8v5gBww7A9Gxocdrnk9iDhdydApbZlbsMUs+Kfn1NX
5GmODEt8R4Geted07my70/VW2qB1Wiub6mj8zSZB/dradhgVtoqeWoGM/Mmqed0lsb94upKAb6Un
5iA/flSluqOBi4XsX2WDgHbe9qpt7FoWe6k7aFhW7sYUq0ScbWpaw8y1wboFvBrtS3rSDp7RAh5o
qxHou2pFZLT4aTp7CfRxDAY2WQ8RViOre9tCHTA0dLiNy2sh/EWTEziWCAqRdF3J+b8oMPZqDsLK
FdTR76r327ev6/KE/lMEwC+pdwNOlfWWmj1N3hK0I1DPtNn9kyQno3Wi73tGdqc5BtHnukSYrrAX
KxmWCCmcHId1jV0lUE3n+ULWQZAgFWcsFDfMQndOVgyK14QiehrYxqIlhe+Wdzujl0SVWju9h9bW
eOoXDtvJiEz/LDF17v2sCBo07FBx9AnReaxtmOpoiV/14PoT7AbHu8YA40Ha4e8ZpJr7A1ICnMcc
tEIg/vIAhbzo6RejwHThGFq0i4EEqmlkhMoypbE4EGsgBZVpg8mNk4HCt/t6rCAk3SVSrgSyq9ns
aRx/RyW4yNR5nFjCUpSsxp5E273Yzoo6slfQDMLI3U/VPFK7Iz+OFGwtzNXn9/5FQK4PY2JEcnxV
eCy2lHu8agci0JFqVlhcwMhQiuFsWaDAhA67um259nrTNZCWthjKUqt+NDWlNlS38QE8+xHVdep5
eDeNxHqrD8AeE30Oc5fvR7j4i8Y8BrZ4owKW2jI/sdAZey+ulE4QY7njfGrHQvqJU/Y5z/+3URLH
dI6UpHDMUjYuzGLQCR/Fz99UJPSbI4XpzZCG3hclWjdT6bPVz/1MqHblbiPpzFncwJi1jV6PDDr5
2/6ZYQbicH8aJWrnoEZohPXS2lPoHU97rYItB/2MqGfQwAm3STVsYmyC5KLvgawrqAaoG1E/1IL7
tP4rv1RMWM8xzGl9eDxfq572jRFdkpgrheVb/JKpuvvxS73yGdqClucmn2n9AfH4yNELEq7mTDg0
jL9OLTougpHvd60uHpYQ52bDe6poBDPRNpe7Z0YieBb3+EbTbZMeBtZlZnEiUT6toIvXh8h72oEi
356YQRh7g8rCL3kbRZN6KBrOSJ8gdgtGoZ1NfvZ4T/yRUlSnKGzUAh8CPJLUGf++NBqDgzXwJHKy
v705G4l8LPATe7FMUWPk/plkDdR+vDfnR+VgRytQ70uzyN5q/YWT/VHCSiMznJdSEwHu0wZO34ij
Qq18FQCQ20Ef6OsR8eHrzsMdRDnZT3hcUs7ywnDb/Jc62ybVa3cpkHadLzEU+aBM98ch0uuyWGOM
4bAjZbePmgFgEW1kqeqwNgxaVO9dFy5rxD687FWwbHrPuiA7nvbTEmGZKqmh7ZGjNhK4qbe4rSTM
mU+vq9Q1pbfBpQc32eQGk7y81LFcgQj/n8Q3cDeEXuNH6rtRJ0YZtQl6jBbrR90LkJ9BpqYpLfQx
2nmWUO5rHVSkJ0vjNpnZen9U71ZO/I4168+X38/w2vsfXzoT8RKo8fGskch7IfZm4c5SvG9WqUNg
zxzUIpMeYQG5PRLwpB7swt6LRWQ5LhtgWPdE8fFDwEybDy93FWDHihkSKv/VBH9YCDpJKepOADPB
o1LlZ7Gjch+JbmNMhU1+Wr4STge1LJu4vT/lagexOob3vEZLgKAzg/rCWwRdTeshGK/ygUS//q/Y
0OUUWe7BdUHgDlDW0rx5xRkiXy9oyeoMxqaYBO3qX8bAy8oPwti6nXOsmSX27ZUd0pcu3e9x+LOt
ygvtuH9r168VuniqsLBSIiXzZ+h3mw+AfWDbSubxqZTmJUBe/JTMR0WK6RtHskFiRpVVMTQxy72e
pmYX9/JRK18PQMz3V/C++NGKworJrXgFXZKG5+pSvpvuJQ7eam+CH44IQ0MT/RS32FzoN/o2TY7C
ZmYz8qomQM5H1AdHB83r1PFZRv+yFiiuOMfvJtrvGnrTw3zawwVFsmCE195TEHLnwQnGKdYt93tN
Bwt2uzDGqY1mURLZRIrKQKTLue6oObb2EC82w69xEgB1jlIWehyAdQck4myMkOYO5bddGWILjd7x
qubZVg9yk4g0yszZBjwDk38IKcQBIMqOoBdVbc5a5HXxi+mb3rdMlB6D806XyGeR7a+yPSAvqt2X
ezAJKBsVZwuKuxajK5tZL45/dfIg+wDaGMV93Cl/iF2oxGuLukZzOwmq1UTV2tyMxzu2gMUKkwcD
imO7NrJ8+qfv9c+tU8swDdifsaRDiw02f7SUhbpaVZdiB2b/XZYLj2baKg1YWx3enBRQGOuo1h58
fmCJs/Wfx6m2ayqFH+GJSpf0lhqfoHjv2CH4Qe0jL8N32CSIf40PrUHtvldhVqXNDsJwXy2ZK2OK
LL8gRGRb3agEd50E0EbmpUYcOjYLCgxOIjKAXbQVzh67JY8v5XIvlIymx0IpdLayni1S/PrxDzhP
l53eOLlhHHHUBof+vNYCmhuwGlbIKEu2YiPo8lvMD/DrDX8GPceeo4BFbHPKnez8ApYpz4YjNgsf
IEtdPXs1A8Sv4jyV52E0nTZ21L7fr1qlqUPEW9DjEx0QAy6OLw2qW1uxDk6dOjcYK7OLpdJfczhD
SywTq2OMikBdM8Q6wc28CeXEZIpoxiKgErV6s3OpkrEz7sMU6K7+l4ez+udW00X88s+4hQYOxLpO
ahWLsfovpWJYWIOenedldoeU9YUQcGYTDuRJ54Fz6RajI8VvG0fmLYc2/avFxhANBYIwBnV2eyJu
vsEh0Q9BG/OYCQMUYEUzIwKacEgLY9+XyvIHkyeAogb4SOpBflm6qzrVXIpfwxEAN2pM2/gXtHNm
i18UpKhww70spBmxf5AmksRa5ib7RqFQUZ+pMQ3PuBEHI9xhx0d8DOkPZ4ml0jPCjT86Ap2cGH0Y
TgRh83HlWk4ymOHoiAifsWpOkiVKyNw0y3Z/B29PalTOQP0af4v7jdTnmiKFVqN1tH6doBlGDwTx
BiITh13Oft10V/43gbI28gV8/6tfCZDG5Y4+TiWQyIuzQbLGUJXvnF+P+QD0bEhgIXe7t27XYOwx
VhbeFmvG3OvRDe3J2ALm12z1r0XNt4jf2OGcBCaqT0w9M283Eq+Q8Jrh7Lg9JRlKyVNxBBpWVYkk
MEqPL5hFD5/7RRT1uZ+B+s2zO/Lzv/2BceZyKXvRhdNMwhJ6ClU06puOfmciIbpIdjtgyR05epIs
RbenGDJ5Nyi/VlvB4kzBgc08rkkbI7NnMdLNuerwGSOvp1pfzCnmLFJ//hEt8snmxK8oDuqSlNUU
Ucd/WbZpDpcryEjHWgN/RAOPQy2LoCpJWzuzPCGw4vBsJiXYB8eSi8PlHqyAjN3LJrerRpkIH4ea
KI/3WCzWKErrgR7GYrWdgQRvooejk0F00LLpsvIeqzzroJF+P62/ZYNyjoROcF54zlrleFx/2dnL
g0x8x9i87sPCwfWTiUiYLD2MFGfhxZ3nRoqicJ+KzOttdshUgHoyvz+UthRE7qeN6dyttuw/T9+d
6IWbU1wZvq2OTaFy0pp27jmgnTrNwYZO438r6e9/LliNmOofbqkY9E9DYMXawUYoZwvT8Rp+JeSS
YE4WuVjliIvbblML8pYdj3gZje/9pitviqGoZ7RYX/1D5yyk7b69E4Jb+LbS6h+hhdQoAPmfg0dI
1vyagMMJwZBFe6z53V3n/Yx4UpWOSAEB8mhwOHPgYvCJt0fu0puoKGsZelbWdi80lkc8F/AMbLSp
Qh0oZGp2V38rlkB97v3Om102jiBeL8QbYqgAc+IvP3Ih+yXrVLaPM9BCbv7Q28CB1HJJ5j2dlBMC
uTtyPbYXQnbbSKEU6QPvB34uucXq/HMjLUU2V6YHjKz/tPwMUL7nauc+D8LKwnQiFpJXW6s652X1
QSzCgsbuihpgXsojJyuDv9xmInttgcwm9XGG6ZqZfL/hpQJZl06yuygtviJt2hLXC+RSaF8bNdwB
eiSjrDEGEFPKYGlQeh3AQ06WSbRa1L2RcZ1dqmUgJp9JWuXInd5bd7+IkUlct1fw/QRH9v8ou+f8
ERbuU1u/PSNszSOlwcIKxZXGMBWAjAW2WU1qf8iEE0FK4ewihT/dsPkGKukXJbHRISDnFu+etj4c
qjuG06H9T1dT1gRgdGIzsOW2rtyigml7SxAwcGdCtFayHRT5OSodzOv/a9/YJGfqyNYR1E1nEGEK
Gsjp8tDmOMKLuxXwmeJjGJkZw6lFrAFEG35ZXNWJt0TE9dewNQe7KcqRVXK9+W1KMvXEV4gbEt3/
LFidz1TOWFljmqZ7wNS2kRsGNlqG1OtUn8InWI6GgXX8cZVwrO0aFbwnu10pJzMU8BL42ajAidub
hVdIlMyF7usbJ4Hnimr5zv4xpUUJw43X+SY3bACHzNLNKiqSXZhvjFbCjt9EBjv9UomXLLiFIF2M
YQ8gJNKGlbe1II/ygxB5WQKg4MiAeir5htM+kbL3Y/G20wKgM1pIu0Pt5Cct59dFMyqSebyDX4yG
R4oTkkQuS6EXFrxdVdcoaQfwpGuYWSpfJcciikP3sIQBpA6/ohQ+z3r4z96r/dsrNq4fsPoE/jjy
Zxy7EOrlLrLlnzzli8dUFgliNjI+Ky21FTvkv8m74DhLnox+7P3gdNtM6LKu9CcpW6Z/20yiEDbB
AGB4h9SevHAf7l8NQTYt3xuSR9yLURCpnKhScQtDGB56pFdwqeNOjEMbSebcPQdsowont11UwRnm
fPZXXRIj92DvYCg6Eh1FQ3ffMKpnFHllWP+Taw8NaXdcXAz3VrEB4PG5Oju4mUjcQ0JEZl9s7Bmk
1htQVPZwkBgXyI+sjaRuTJJmED/5Y+7280xjo8DSippW0tt8/mB425Am5h9SbTykFN07Pv5I9Qy8
4VJUBEO7Vgzly9PcmvQrwmVopBVwVFWBJItij1IOZT37AXTK95jv+0DviG5jbVa+k1yoATlyxKa1
PsmMniriFGFzE1yrwyOm6YGjBpZ/fehjZ+1J6i9KL9j3mnVrw1vKRnFBL8bGN13bn6jVHUX080Ys
yXLWdpRzI2duzQeLC6jAifW3so6koQnfU9pW3DHigKR/Mug+p6acDndw7Iv6pkRtL3NBp2/DLECq
g1F2LcBqLfdhgMQcTcKG9Rccpi4jZp/2i29WIpxvAphmRHMXQlSZVY+Toqbn5LBpRm667QFbYWci
PWuKWrNVz83CFk3/DqVeFaWI/W3t5RH+DFbBeIzFXKyvFEp5OeajiadM4TJSzOBJFQOQ3sEcfg0j
SWHGo/Gtc/rk3Vinorf7sG+73CvR4Ka7lyBd0IT2og74+2ftBhMBZm0u9m0pY6+JfZjMzcigtUlw
NxCMHOYJS47/50DK42pbcZM3WmpCNxTX9zR+Row0c+jo+JRioKT1uXKZR019L8X4WTc1wO3lqhIs
UoeYcuZ1wwNZfLXIyNwvDRM/bZeMp6r/W3+N9HX0tA2CeNkTyIOzXicODZaeBCFjQLjcoDGWXeye
YaayTf1J7J2Nxj1QOdRpo8TWu74SBI0R23fuM1JfrT3N79vS+9x34ZvQKhMYvBAM3VKPXfwPz30V
vFb1l9BGD6eAvgFnxa6Oy5o0yY3jXs9K/NHy2sRhNSF2S+iIsLrW/s3EODT3uLBXugWc3bNrsiiK
Pr9lXfF8fv/AP6WKSuqnAmZBJkHdtDjdtN/Swv1B0CbigRFXciVmOoBcxwTVITspQE4cU8qzA5Dg
m3JDaxRvPSesFKxmJ4ObCW86IV5zWjIwIrmx0tC4uOF0DQd9x4nUXK9E3F2px8G6MY+BZHyQo/xq
QEX3SVu+0JOtg1RuVXhc8loxB0+cEDZL2LwopTwAayW2odtbfCEQEq85JC1Xpe/i0oihWNWBlUpq
q3hVgn5dmLG6L6scnybQcjCxCTucm5RWwA/cPd/u+qTDlBGgZzG1q1HT2FtqFzUDYzCnQyAZmahd
4rZwOwdlQeyTyef+EmiRjSo3o9UC+ElregNsGMj5VnP5ivlQTu8hJMSiNLvH9GR9jkhVJ85CItom
kH8h5ND6PtGnaBoZdb6IDF912DjxHlbrZnNsw/7FYOARMdVPtAsYFuQ2HwTQ6xHLW1UuXwtPH5XC
yW+j9jg36rBP5JvTNnTDVpzL6dApFuxqciVyN3INqkC0d9dkWxvtgcRCQbtT777lYZkxyn156mT4
n4cKKj00NO9iD20We6UaAk94DVZoi0u4sw7YIin0j8EU1dz62uQktKBVYtw29Z6Bc+UW+QyaYnEe
5yXFVMKdwofdqacmnNX9JXJXHS2A7HiHDem/W6qQbrBbE2jt9BRt7pfwhP29n7/cDqFL7lanB24n
Eks7C89kmEjwDmI8LgKc6uHC2RU3/eozJYltyQcSMv450rOCCgCzoa9X60VWC83gYcCgC9ItxyRL
NbKXj+s0Tte5hqDlh3m8GXNmEbJvgEAkUTKF46GzGAzu6CxcZfoeGlJu2KoH6ig66J4ORkXux8a+
zpD4LebwPVRZkseYn2M8QR5A+r+u9uzQAKYQrP0pe9Mr2podeOHlGoE4Pg4G59hNQZdP4d5YFl8G
eRYtGuuZxsLtwV46cQzXWXWZXpJB9UfapU+UfbU95ol+Ws+oJ4pbCBxELcJS/QK5YKmb0aAAq4mf
pN1buQbgm3wltOcRwQn0gSUc7qGs+6xD6BZ9vhvl66IOddmGWRNhjmdUOUFi+s4SjBGntL283RJd
YNT9KTRCWZ1VGei1+6OM4v42RHOIr28uJi9eVNvZbS/MmJuhFnww44XnjQenqtPJLhVJa2czWYna
UrLqw82SR2I+V43qMhYAiC3hcakT0Y3naDIEc8gzxmUlgbUcRbtUrbBSP8rGUOnkUFYPJJ2aUttK
fAG7J06YzV606/wcz+WULAByC7iHE84UJ2P3+4TfJiB+kNoXcQrs/OVeKaGP896pTJ4rebYqp41q
GlDqrFiOkkXwGpXxBsTGRGBraaKPYZTcNECitirFoOOvbayMhLEvebj7x5+2CSMXWmqEtJplbNyf
gV7eGtHkK/UQ48Vx648rM742Pzrxruwe+Da2f2YaFaNOOu5WxM9fFXVt6CqyyaBfUe1OkuY0GPJL
jtvEv4Z5ruU7TsOfgtjLWaXsjIfu3WMTm7hNVXVrhirs78WNob+Hfb8VAGYpw/S1JqXdHib56ztO
sHnt/7LpTGM8lcQHPsQbm6YyD3QE/s6fQFcZuJJ0KWmPSJ3qnsZv3SMiF1PekF379ibWh0vqRPFF
bkSTJ9epOxhHnQMZPtqmTHhe6fRZPdonJ/PfnWgiN6KIRJUjPqZdupjDwbgzepPgFEbBgF+uMR9Z
w49jAYzZDPfcg2ZWoJS3kGjctWJIsGBSdIQb9BnLtLpCLneaq5ZFrWwYrsiu7l6m4TZbHYrjkDZi
Z3H/IhYe+tZCf3XLa7xkzpZX5/DcsQ4y+4QHxzP4ARQqSWyk4/zXRJkn8z3MOkhUj3ra4KIqz1nR
7BVftgKwGIOyQDaFkYNOoGJ/JDseEQ8MHa9U3d9XYREM76zUgXbrucpgFMnTmwdqn6YlMX9nka49
mezv6dwawHUzKQz3aU0IET4EI/JMEaD8vMEpmDlBsexwMwQQeJ2n64V1H0UWLVlGMVvKLYw8p6Mv
zMBxX/SbRQYSVpCqi/ET492E+iGIYArm2jaep+K93v++LEHuCgmSz5kZn0UtmrryN1BW9qyVaADV
jglFS0EBlqSYV58pMsH9QPxsyfCLhQeulbRsTQmKW2N06NP26xToUfztG8yxHR+qr7r2z74O+IeZ
v9RcO8Q7ZexSqhkeF+fBoUgHS8BB7LdknoIZD6BJu4lGBeY6f/PFbYm4LyrDCn28LTx9uxaxmb2P
fWRZoMIBQOqBYKIwtG/OySOwAacHMReqpCQuVtiNzRkJH1uQgvdmGuefJhsoaPM4K+K63yVQ8vF6
2cODlWQQV2z1FjozMJnDMWg4Nvv9p+9z7kWl8q/c9vdRcvuhvaox8Er4z8zUGmpKWOpX1WfMeXeN
WBYYdZgUVmLrpeizE5sWlT9f6TvXRpoiE3V4wIa/56Snmrd+lhx0YTYc354tDKQQp/9MgR2Aymiv
eFiEEwuqEcrVilY5sB3os2AB2Ci0IXNTYgSvtIjHSQSfuZ8arTGv/0lSWLHqYmwNleeHBiXbxTep
eJFiIonqqsL1Y6BSMtHkLnGuRorf9sEWy1FwyqkhZ5faiWRVqaukEax6dWDM7JT1fh2N85b4tsq8
fI3k2XUWSs3s6SoZtZnuBbZYx9eKVg6zwPqwURP6WJKpeaOsQmCCvNua3dNDyfn2+dpuFhBRgABd
3wxFdhyo5GP2oremNy22i09XZnWZ6DXJeiS0vxi9hCgdyguvyLDdJvewq8UWxrdxP0Uzox4xFS23
G3GM2WsSGIMQY6UbYCUWZr3SEV5sMT9A9yJa5nXIHwtlRMIwE+bg5Ofk2ivyMORdK7QZr4W1Q0Pg
kW3FmHCd8ysKCqsHrJkfPOHSRdlLCDgDwaRSEIAr+aTWe38J41aGW6xW4Afhbs6/nm/joU8hm+ES
8wrgFk+CD36c88GfUuaTVnkAo2+3q+o68if0vuE/H85FlQ0zNbT5HsvaYZIlKq9OReJ38ZnruYmX
Xx+GPvwFaatXJ+gYk8H5gHoNcd1YzUB19y0M4PSUER/pf2Cx0Ml6YxddqapVGCgGAFLgyMBW8QLl
Avtqy5MGcJ76OmTPUJFONVZXifDWEpLw7eBTf5p8CSK/ETiUMocW1mbonMd7qFsNoeg7XcfcmZea
oXx/GDktsEuMDnuRQZF9SWdKbameeFk4ubEod7cjkaFdie97hOsiILoIIY5BIcAeUYxjxQdPF8SJ
WEbGOYgVe/Aaye+JTlPaaHYwO7qz5Ik5+WG6/TkYKhB0Eoe9kAAixC2z30XJcsSq4wTdz6WYsHIF
rLedlQVeMets40dDs8fBHUQ+YOEXU6Bxcw9TKrCFsb70gJrfiTEwQV6zPzm0G203bKGHJtqqEzZd
ljKZ1HKnRksfNtdBqsxa5XpHPuoU3JqStfRyJHryWgteoOsO8u+igljiXRUhxqzkSPZv0AYfulcb
RpUEYeHv/n4tG2vAod6ouM6EWAHZmvwbY4xTL/XJfi0316nTxdUxMxP94FVQipxuXwtMSjzqquW0
bGNEoLKCEGTRZLd6XsCagNa+3bG7+2MvLp8smDNTQguktLoVx48E98vh3lIMmIPjJjHH9NbEldyb
PGzzaIFN5E93fG5s1y4w1JrZKmOi8OtRwkyOKgkbLIL4ajaN66UE+L8iNJemqJc76dRT8r9EDZxN
cythl4rDpMT7rKH8agimXQTQm2h7LqFfKzZcyA7ciisPuaEwPCcAABcWEbMJmN18dX3gotSN5yRE
+vl1QNYPfXbNU3TtA81ZCWPnBUg9f2OTSz/XuPPkB51zyYVS9cycD2YaFsmqwYczDMtKX0jq4nEr
MJZDxz62V+rhzyiXyqKtaSN8rsZhyxOFnEjZNMlPhrYUIAyetHuXbbOwD1VX6hoaEznsebYWjmQV
lbK7NwTGJJGRBsRpJNNU1KJwoB+osLA6AvJRUt9XEv8Mo3ki/YYRFawi4qnFkgvtWLT84H3XiU3k
1O6+sVi3GkkaTDCviuiK+i6Tvd+UC6JdoH/0fcaDPi8TD6HwlCplPIcCmh0f81g0zujVv0Ggb+MG
nR7R8qrwtenHKn0JzFZ6XCNrVvvco4/M1TTOc+gtJO6Y/3CNxXhFJn7j8TmDoqLs7u2WWajO8AuE
0p0eHeY7PEpRJfcQTgsZSzoE6YvaRTQQEfI/RES9jOsmsAx1VEIrEn9yG/vAIqzAodaLgvAHgOCH
5FA2cyUHfBOdPsEymUyJye/y1CMR+cr1GZzYpJJ4jOgjdZRMShuueTtWzbQBdEPu/yxjY1wsaVmb
VN/on3pMyNlPEbGyMitWzVQz8rpdoWXD5vaS88v4NAo5+2a2sgOL+NXGS3FZ821/fea8eSl1IZpC
BT58yk/7DCCkykoAJy4wNemzk0YXi2T3dphNoYkVXJ0K68bc4TQAJIdyRq+oGE/wqp08IIBONKaH
zbAYwCaXZrw2rIhb5QZ5jbz2Gmqmc9iwCKEK3SUChzedu82iQ3Af5MR6OxNGjGuCcFW6CB2gUoIC
MCxhbaV1R9eX02VLZtXsaizR32q28pUxHYkZ6KxwLWB4h2/Mok+w+TbA7hpJuN8I+thP+aHnch8M
5Kp5yHz27aQ2MRfX8qCSWZQBiCvR4rt1gdwMkOZb1LgC7mwUdKLjBfignqDtGNUs2KRO4Au8jYaj
qpP7nVGPXt7JR22I6yqR4eGyz+eQ/IchT8ySEih93roOg23YrLPPNy662v4HhdhCB+xnuUtfstkM
6zkzQYubfSgizK/iPcpKpCpKyy3xqQrglxlWaXqbHwEQRTarGZ1kyAkkYj2bTnij9DLoUw4royQ4
g6eEDObu8QzEW/YFpNfhUvgE/Qzom8Q35jfa3Wcn0DipIt5Vmj1gTSAQyZqKonebbOK6HtA9VIvh
oEbTSGB8Ag5rlDsV3n2vNzf52h71UOYQ6uC4yD0d+duNB8byxCr0be8mpFCy6fInUIz3EDmsMumS
Zv8AflrkkHyX5Uz1HvFQ6c55NLNTgm8FmrFHSU7ci5rMOF2g/5QuJZLUzv3oa9T9GhfR/gcrcyL9
i70ovK+icciR29xYY+Nz41pJQQr3Rj3lRuDNT+I2nq6N2JYwEWd6WKTXnPdoCJT3S0iYKKMtx8a1
aN9OSGAQO4812OWzLxxfrlxwaPCJw2WgSbnPzY/ZzMVMAbnk94RhqeyxFPnV/D0mWTcrD0gfQ+WC
wAhkSMffuJYh8wAltZ5RA8xGHlSGXP6n82jfjI7kv5wVewCp7ZnS/CEpm8d2U6vLAFWJGLbbQAZB
UImQpWe/6+MV+bXoeIiC11rZcEz3u6laf0+lDq+OPvtCIYnvZKH+DypfvJ1yBBvk3rOI+obi54SS
9N/wDSpqSXhqtr7pe8VYKZBl2lROH8/jeRIgY6GIVZqAGmiJu2JzylfsCe+U7ukiGphZqKxdF+Eo
+KHhCRoUtNtOCBuZmIjLOgF1iaMfQt8Dfyr5Y3GT93bE7rOmICIGE6KVrlpKPh0JtWNd7FBXQ36h
HmfZYcdt/s+1X2nht8FqB80Uhfg2b/3F6egJU340qYyHqpOq8y3VGU0GJBabYDpzHdXto2Z8Ibs9
/JcocqE1nebJJTp2erIie89O7HwonULQoHMUQ+mG4aI7G08cbB3UbTBvFlAPl+ClgOXtpUw3jVdD
xLKfAedo5EWFxXnHZiI0h6WIpuKD9yRSIVyLsDMgDachoKV4+YABSyiRHEJAYwC3vndKZvSZabsx
8rNKjK3Y1NZWXYGpIeRclmmGj5s1TEnbrbbsCEkHaiNdzXhI0DomDmXC82nwzZCHLr3ugkG+ualh
LIhVLK3V4aiSjngh2sBk5R9+DUGHQI6X+UZHFXqeEMRqPhp54Z20j13Nb0J0TkZYng8zbbausWnO
Z+81aspvFWIulLZrgrqyq3LYn9jM5x3US7MnG/YTsmhiAkFhWVKQrbYWu1/lg3KJ5IzAg1DFBFTb
XXKbft7JGXXr0NtD8DwO/XCI5lYfdyyJet/iRA4SU1qYG0/W3kqB6Ox8kxruYpBp6mTUYTYVCZcM
hslknTUbW38xhAMO3mqT9Qco3GoA6ejWV8EttJjy7clExz26L4UChfyDuN5PFUg8543KMUpg1gKj
eCRjZ5bjMGKDPYt1bMmPZ1zCtAMNtDbdCRpfIlE1VI6aTzWjYaQT6fH+EfvD3yOVt2ljaWdGE4F6
XTwHNwjKLqxVHnOMsD3JWmsYuKfuEnZoJVNXJkvvF+nbd9SDXJGrLxojcaZLfZ7TIQ9O3tdk6lhW
aFJJ3whFubDfqLYYyjZKI3nqPPaTl6altHKL7yWi46YS97wp3Gfv4XjbBEjW8MybBjsJYqoTGDSg
l/hEZOyXv81G7L0kLGkHr/8Oj2tt1RERtNJgpnY7FZJinPwhAFnRsxJjxnTUcYKK4m9bGkjBfjMd
ttvKrquh2lRj6t4rXPuxjS3OSJKu8KfR9EGsKl1rLq3ie1K9W73w6POXWC7NT7/8+5ckAhmeSat5
m/rZIB8ts/FVg4ZuukeMThnRDHy7hqqtIb8eUKwMZlZTD2DDskh1PXvzQPx1rF/+pfeLOsj8+/yf
+2YKRxrA36HU9Fcx3yV3FS6vEjOqcTiXi8a/OwlgfXaWQ6cR1vWlBxwgmWXHw2v9r9A1CVSfkRwE
qn2VdoAA+6RmjTSDMWx91OdxIebKqfc48E8FByU259iXCckJgJtpSh4IRuCOI7lKBq6FCiTEYI41
2wPsSKlgju9QwXYJoN3aIELe6D2AKSAEM0JlXeDci+T3LvqARx8KfH2TpZ9STydX5kTMDGhXurBw
ar4aNow4LhK1hbFeaP3OF/W9C+GrT+F2OeF/fa4Rj4lGktcYGI4Iq/OmcCr5cguChr8FaSIodNZv
MifECGB2vQpD93WfG2elkeu73HGLQBXiCqm9X/YY/s5Vr7BOV+B6MszablDPOdIssW2JoS3p4Cv+
cgjgea9ZM5nIOLwDI9c57Zc86Kb2Y0wvPwa0Mkw5AFuPLxkXm7NUJYutrpbi1frkCpt7QLINeUZA
52lqI0rrdERfMOCm/dYn5OM8/5EG7WWd0hlJCf1X4laqW+EaHckQMr8ByTWgtO10tuLqsT611HwQ
uwvHBXtXccFuuDfvRQ9IIIJ4i81Q2WeDTg66TH18TMr0pWmYbcNFS0EgvwIDKE5/zW5ncRX9+htb
dms4SmPPM/U2YdlV9QI7F6JYZaohlr+vuVQvaM7I/ohlcl5xWVMvUTfjAl5uoMdiDR6byc78jXmh
kZydYwnCO2ljjboJOYX/hesqAS3W5aUK6InBFzA5rwzKK/x30aMOAtF8E34qPzYV+cogMBpNSpFG
ifiJE8UdNI3+lvSlIw5zA9L8ipguk4JHXH9+SGJe3hqGv9tqqtKJurm88Avpa3V7VuHYtrSmEK4e
4gQgv15R3V8U++ff8/6iT3UJKC56z4XrtWByIUsoy69T1AEaQshFvon1iZzLg7k+yQxtgpqRS/va
1a077rRKASdtjGHoqwnj2yn+Z/0tZlCFQqyheYxDZE4+KqGXEtOWqbbOhMkxNVPabW7nmwcW59cN
PXpEb1CC6N+ulOxEBRoGjM87XZrlHZsgWLUvvWFsAPrV0l+e/Cavj87yORy5iY7wSRuR0Svq534b
5SSMHtWt7XtisT0Nd97Roz1hTuU/pTb0pSFqfrjFQoRpgq50Pf1/+HY9UIaib3lsc8gvmgKK2+F4
F+sXOmrwXnCnBfaKGhp/c2RQWbeZi7buUMRbGDHfFi2DwmGscJfNihzvQDl9+xwpJI9mCcEO+rnr
hSGND5brQlwb95V47jU6NoUMPuXOYlZUS9+vzG7HMNaF5j+PCvGO0DWYlGlozfBdGFgCpB5727uY
ijn3Aqbl2C13ulUBxiGVVbj+XSk3B2NX3XIvCDP66qb0RVvWlj/gET71TJfhGYR3hYddtVZ1ZJ04
5rRNNjFRCjEMvaTQgIBWQly5ZkwyuxW3yZFYNX0KMlMSgvM5XBUQ2ZQnO1jojKJFT9BYPljYWKAc
i8Q4N6Cc3zcPmGiFCs3tnPw7edX0yEu1Gvr7P6Nmjm1lGiD47rpPlkO4EcBBfhy31r2HKZ7Bea3i
bcDd/NZJ+VBNBu/hQPk/BD9qTatDHzdcVBlAmFWJqYfpURLrnfaZhXTDgt0DV9WFWpAPePm8Ps21
lxa7IZBAs998cIzTt/VwJdT+maQChdAFDlCyj+NvzPAzG6vqp8gI8cC5hMlJ2Lhy+ngOVpIgcMHD
TwwWRRe3IbD4izFPmdTKg1vcooHHlrNZfqgrzdMvP+K0BJnJlFhgaklT2OVYMzautZEZ4f8syX2N
FqQ1AT7MMiDOpVmUKgjz4nRkz0kPwECOPZ/LKlpv9C6WMiwiymB/tNaBu0G315M6FmiO1oOXo23E
dKIbHP/Eczfqds5cuq5sKT/9g4Pkpbn83bS/BJbaxCW9ezZujQ9BDbJZcCqk3pon3UWG8+62ua8X
OLuBKbTCSyf1YNyjUrusNbaY9OsAiLQeUkP0iPe+1qOyd2cBEbKrLhffJvb0ucHqASwp1AaDqkJ2
zRkThsSnFE9GZC15QkYfqxrqKxwT4Fxk53+zBYfeeZ0FrGsM1DEjho6jZrQCRbvCPbw5gdVc8QrQ
Lm8soQ1MpXtk3m5JFKPjqiO48p7D/7ue1oxP4Wnfez/zO6SV45YEifzoeftTnNYGWOA6JwEbkKQ6
GWh91qE9pUdC00InBAJ20v5MONKlfCXMmAjgEzua0bKLJ1YuKdVLlvP9IUZ82LenwHpV/aulSvjj
QH7UMB2qrUtV4hwLFWm7s/5BwZAeZtLJwgNM4d3goLpa4jRIZC94aRfULk+Tgq74RFbLDJDhYHMe
j7bj2HORrxHVjPB+jlVUOAsLTkM3Myhxl5IbBimDW5Oy684nbe4PCxWVButzkA02yL1s7TjnTDNk
fwPol1H93kC/Jp861cjUoTdeG81T8ai0ko74+GrycIwHfr0AcDbA2FzTT9+TwdqlIEtZoALjkgiA
0XBWGs3lZhZjUkL5lazW2oRnwbhGlRZIRqmU7KM7CfjHSMd2SaNk8CU8o1cKPQrCLCCnKALoDpFq
7QMINFyY3ywtkFlpHhlpnxEJ8qM4aQWiMqno8m//02nj2r12PGeUPuBDiaUBBR4QAJHXZ4pNM/4c
40bwHP6OmKF3H5GpTw92mCzNpDLYO1pOaD3DAWWBYMrpkRg/cBC1+oQbbpsEP6UV8x8dl2KgH4c4
4yUmzGycwjprBxHUGnRnyi543CyNr8yxsXIdXLz8gulTlVMS9WanSksaI3vpcg69NAvW63dMkEVy
01XPbwncCiAUC5DGKW1EF9yA86GaaySMuwu9p9THlSGxv2uIFx+Lc3XxoLBavuPjMyNx7irkxRhA
5cWzmRE4lk9qgIx9/uvntY+uEC/et8jw642ZnX3ga6wzFNwyExEDFCjiMvPq6qz7fD7+9cDkfv25
+JQoYFaVxsEBH3wQz0PX65PM792Vo6vfUPKwyUhUt1CCNRJjwOPoCS2QWEpHqmOFS261/8BeId4A
PBBv+ml0tMZ6sGMD25HB75LT3ERhDtHO7YVTHNxTTU4H4xfdTJIF9pPtxVq+ieAMvlAMAfKsz5eJ
fF5e+UnE8zPUfsuRS+CFAMa2HDYrX/tPHKqjM8XFsXYPjqzsJqxCDHq87R0Yvc3NSMpfvXbpMyLv
MZP7wYWFaj3L/kGKztw7H4YAvN5yC9kXaC+endQJtBr4lxJ++9wuWHNL39W0Jp6zWml/09argQf6
kNqPBozlI3bQzK884Zbqn5+gdkM6W9F7AHyEsUsz59pI3oZf+1Smzlkkfo0jxtoUYeIKrbgU7q2Q
NV3cDtVv4bXS4oqzSUCR58YPRarivclqIEKxHQMlQIR2XmIMiTHmYiueSNvrE9oQsSrcwW2J8PKW
GgqhLbDQQTSLtNEpisnEzM6Om+lGauweRiWoWUABdgm+aNQSNY/uOa57TyxxLcL43vOtaceJ/sTl
m5nXx5sKF6jJpcLMB/RO1dDlmr1W4KKPZNMdmihSzcjhKn31CVkOZo0LlO8yN2T21ihV+WDxII1E
k6r7yWdgavQXSBvMgGoc1fY5P+RvGn56N/JbH0+EiM4d48BPHMTFYBwO4IB3YfXKWnonpksy03CJ
Us228T2zpvkCQ3gKIgpuGPpLL929VFWHUMXgRuWEK+7+XWuh8sIy065boR1Hq73xRHjtrDrotVi3
hdoJ2MKyINP5udOnCOZtbh/qt3zeOTnIwexUjy/3qj4fsKr1dDNA7GEeKldiIiMB0YpygxIe5TlS
uHIohkDVEnL6bGxK1ibzla/9+nf2/eHKwNS7lPr02H2WvVF+izJzLoryu+zpEGhqnxp7xTHD+RJc
HyHE165vBqSDi4SNfxPnhjLq2MZ5+e88UBQrWpxcZVGMV4EaIUM2JcoOhvvbmwEAuMq4eszUJOA7
NtLCVoPNPbPGwZ/VUpZi8JyXcaHZM0S6sZu1NCKLkPAoAUbpNanPZzjfTRXzl/OhNWulT9DR+LEf
8Ava+ymo8j4+pxTd6u+RyrUSxo49lr+C5DecfvXqNccaFrAXurjnm2RC5stSw5598tBaO0SjnRsW
VE9E7Y68nfimES1xIZCOAsxf3uesfYOOlkoAF5ZHgiit9yz6OntKOFmwS/c/RpjlonJiujH/lLYW
Gg2nzQA3PKecJb5+OV3LpCFMTeB1ltcBlToajaGrqqeyqfXTQXeuhKBzK8+wOg+oASh1vLRplEM0
6Mft2VQZRPWx1aRFJCveVsG7QSgzzoq+CWvXE4fwiugq8RSKh6UceTS40cpsF/3dSHnHx7rJy2Qn
l95I1ZZUCqOgFyQJEqA+3LSdN2c/AkmDMu/BswQzgbzUpd5NYuzkakkiQbO13aNCLVdsa7MW67z0
uSPScF36t2LxRLhEr1ZZNAVdjH+EkMuq48PhBB0X7RGcx9lh5Cj5S0jkTQXz6elae1zt3NjiDchY
4BJZGkA7GhA9O9sicuJwtVSZfT4/rP7C+WN9uSShojgwMNVLrYKFdOEaOI7pSlVSfCObnPYQicaB
xB238NLPj4+2ljcln4kKV8ZiBtyy65zvYSO890cfC0W1+Gd47xIACA2fg7KJnM2kEknzBu2wf1uo
MHMIqJ5OM5zPXD2QQfZLc4Pp/UpYzaFpNSc3/Zx1NQFfRCn3tF9AbbZuPpzXyyj/p1m0OImFFTLP
+LGHAL2NHVaawKaifTkFTAV46LhRfMN81+afF5Qlilt0fsol7TuTQxNH5NOgkxr7RdxnsJuDPOiQ
Y/M6WDpdhLMltV3aJvtuDtSLLunbfmOrp5sm1S5FxWxAX6LH0u4jeTngspeDQo6qIxzagPOOo1o2
pAz6rjFsB/ANK6yQG54puCi41eVP2QUIup2tps5oswJADa+KWfEo30vpmkTkvqt9z+3K8odRH750
G/lMjIdUCg5QAvTiLp21x1mWbwjeEV/Jojo/VS2zx+r40zQsHDVEaKVZ8Ty8SGiFFQnUad4fRRnL
i2aCCfJg/x42MyDxQbKmq/ZnsVWAEyhWDahH1RIkLm2I53MEmOJTg2jTSqkxfkkPrdQARi3yaQTt
dk1EClTChLLGAy/wmsNjTZfp87gcoSjCiy0QnM3oR+TjE4VS4ACkaedbxmev6QTs0ZIMZA9HDtz+
SOdmCf59MCSwi5Ghptya/EWr7WsOihmRR+wxSlWHEP8gOsHOcPYvEXafGxEzuTWKK/U0ArF0i2X3
lm7C0ZECpJI7quzmuSDsTRB0grvOtt7gBtdNDJH0/gFEonkQKIxNeAgdXs3zam9mEtOllrVjHGY3
YhPDZtg1aNrs8B7BAL9Ofaglj6s20wrOF+eifQb7m80JegtyXbyXsAySEQkBfRVYcc+Xuw/stFty
9kFqWh+3w17F9Srw90HZby0HyPcOvBLt6J1B6AOqdM6bh4pPqBkmlDY9V5V0UjWXCXR782owb705
fUl1NiipyDXVSFsKFidHzS6pRUh21CJlfVs62QCLd1kN+5bV1n1lVgwKEZrA/ryFDavNeKE3x6QH
pc2nYV2husn3f1yiduR7+VyBXV6+IgOnZ6MTQTu6JlXaYVDhwk+Vy0fyWpzRUZ/S0dDRMIHFTSrK
4b2I4oHqQlvzVKL56EcE8jWvwvADyNUvaxQUPc8BCfkH2lzAZ+HFUfdA1VH9/QKsww+WgfX+HIkJ
/mBU97V1DpgxKQnM2KNt8Q/DKZX14VGraIhDqDs0Nd6AsLCBGdPlZivYhCu+PdgDyzR9ggi+/EOX
1+d0jEXI0B/SRmUwgviuVe3ZAyzb3T6HVq6gK5yGUczIQR1ThUVV15CI1Ppd/IhdL8eN/y4ZTTvw
fUPC0g7xbBrrwhqRryawitKbxd4j+bxOg54fG+W1jOWhvejooYqr8Tx2f3D4UfKcWp2dZIf+m8cr
5JgLjBXQAA0HbxrksYr9aAb4y/5jH37JFUChkB/qCxTGApMbDE4Beo21p9P9G9r+1iRw+5q81z+7
o3x2e0C8wTMSNWH21LZygkuyk9BBIe0C4zhxFyGoYEskQTmaVEoknPikZ3JBLDUH8xcul/FyRXD+
zsV4KDrzWhA3qwRIs9JQnTtuj5L19cn3omwQdDXUjZH/mGoYIMV6sDrb3mehKjkNsFJRHujWMx4B
sDSu+cSl4UzLns/uKqXVxuCJBMiTII1pfzj6AehG5z2mV+Y/W8hd4c24pvGka9u6EEDiIYhEdMhQ
RoVRA1f5AcFtjBTdtiHgChMW0SLtkfmn6Twh1pKtNilUAj03GSGMs4wz/okBK3fHzK4Qbp9iTxVT
fcfXKxSGUGJAldy8QiND02W7B+hKTrhdvbuBHH/znlP2DIUZobIOa606VX+vKF1sqZmpdG5uba7j
lgdSrCrCGLMRYDIJZ/nSK8gGksFTMsQd9zrAKizx1EUkr2QIRHy+aG62WkAHETZAcDR784HIM6yN
GBCH+Jbpf4RWs9L63CUlgu67S4luV/99H0p09Lw704N2Jud7qcywnZPlts6HxyaV+p+33ohQhusQ
BaBBRqM5FG2fkJx0pfYQo9YCyIjyLgnbDglzgKjd3dE7PfswppIbXBKBWdLpqJOA8ibtcoxlEzt2
Gx/hYwX1dncTHmWPWE0uurqKTU2qRlKSC/+IQS30wkchm1bamYrIZ2Mhj1ik67VeFobfltF+GdnY
x4jnSG1U/MjEFXrgJL7TV0CRYiRK2wb3M4FBsM/TNAex+p6dDBhjN2dPq4vuFXwLKPVWfJI/Y4Hr
nAy0RG3byczn0cKsSyor0dpuJIjZajUi9F8Dyzo25PKtryYmvk0iIEsJPPEb4CORzoAtZNWfAhvD
LprWrUg+Kl+AOGcL7n5fBxLclORm9FMNA/dIfDeQ+QYj/diGQb361bqmkxDt34KvoD0MKXP+sKY5
z0DPm1EuFRdl1CnF0sopbXkuW4GcokA1PR2M1rHri5e8b/o6SPaukYla7dQSk6zoBk1vItrvPC3g
OC4Kdx0Be/T6DDgBTp2z4VhFBuM8iGtwEpFj2WgqU09jC9m+3sH/9yjs7AMJBd8btc995ILwCCAt
rUO2IL+/iFFiGbJ80Ads3M1lU31p2p+d00KM9YD5ttuhvjtYAOoKJyIlDJ7CvYclm6oLMj++ponD
sp62VJIBrs10oFpXjGAJ/3yplUlCyRh/5aJiBBGffZD6jybn60JJjsOJu9hKaoKBteRJxwBXfs6Y
3nJDLjmGnwsrMpdxbNQNEXQ1vhDwdKOmeh5MRcLzmsukOzn9ly+45Bfb0sXASUKYcIIlc44sHO8f
xQxMpieXHd75yGdAYVSpZgG1M2rPGOUP1kkr9DsiJG0xrsBJWfYdGaqVXU4UCPK/K9nMUhdFKtgN
e4KxB7/Xyv+7ArE4xjwAvcCeH2+sJ1WXfCYAigTi7SJaqxg/rjwtL39grPIUnq9AXYBi3++gZUiV
cgkHHs2BvM0HRyVUEARMp1t/bN9SS7K+fbfRkcCss/bAOH+2IcJEQgcLo/kWUekRsWH8B/9WNfg8
ub4eEPj/ZGEPG/nWlM3s9VL9EuwxglA6F7ebo4q3DZTCbHFVGcyWVV8/mZ3k3ga1xwtTtBamVqRq
0nwZWBZFWZpNxjj9E7AuGb1GkP+VA5cedqCEYlJMHuSe3vQDN2W2MhYyNz3es2ycNZbN5HONZzgc
A1uwz/gkaGQdrsZxjbpzaqEXCQnwv4b7qZ3+1rXJ4FbmfLZLCiDtR4Nybs6wfzn3hmsxS7o8+SSh
pI3mZ1sR5ruwr5S/cG+1ZRE5q19uxADllLA0c0hcnhL9ykemuq6iV4gHmLvME3rgzJsZfOXnoorc
/X2lXCQh6ButxhExu4YfaBo+o3CnYcwDnja6nLotGaGjojFVqjHXRUVdGBlt7sjSdlcvl1dZy09N
42/at2ILREGv94fuGaU1x+MIlJZlCkBZOjM0mLk+FpGc65/+2oZQ5zrmX3PnVwa4hndEKodiqnTa
kiyrHpWIgPw8CdRUcqmmmW1VAHG3onj6VfSRPBUkLydrHs2r6iNnxlLlS/IY4P651dHlxlR1uli0
4QaXMgJD4FC7H5kGmH6PgihE62aTS4OkhlxsYEUtnGlvgaSq/vBkB9n6W7QCR2DhHddWmSZA8dgE
AfRJn1kVQGPawDFTxWFVtbaJd32GPvn9siwMiWldGpDwwKJT0/sWk9g6Mpkm5avzih3vQE/7cEMd
o3q1vOMhfETLZ3cIQExTmqBM6Xz2lEKwI2hgdOWtwf6A5HvkzXK83BTG9VEtzHzArYT85KZByG67
1IzmUZ3os5e2HzL9aBrHV8uOutSls+rlLyi5pUwG5lcR3Okn0Rh/1WKRJYfPV/gaSSX3eRaC0mxB
Kl6mkqJF8ffZmpnxZw2eqfQokJiRpN+ViSe3uqLusKB5PNoPPeljG6iDnB4nBLUplwm0jF1wH2wM
MwwuXTPK78FbkvTiEiONmqZbltJvEbPcoK9S4C3YVh7W90rd6HKjWMs0naqLj+j1PZRBy+VsNnC9
cekudTXRV833Vh2hacwJU2DRapAgS6WKeD1KUzT1YxSDWHLc7L3124d6enNr4Gn66uOR4d7gyOrB
hdMw6CgooV1njXPOcUHRO+WhymJP4u4Ci5NiRBBp41tmICFT3PGmM+tzPeHdedquxrLTtqBy68pr
ukHT3ppO0NdSVo0SqoiebN187pCpAEjTc+dqRxwMhOou2sjsqzzE7ZIaa4lFsF1Clan1aG0n4vp3
r8Jd2DghxiTt9FVSYWYMy/HH1lR4Es/s72yYIQKZAc6qfaM4NZwVhqTbDbuN58VkULOyCWgXE/Ce
AfaZcE/yJQNTR3AlI4gsZIxx6D3Fv3R1cMByKlvu2IM2rieflwJw50Lo37JD60jLY+akq3545v2N
K06BguHxL081dlCvNs32YDmd4pr0zcLIeDlpQL9j4qbJ6H8bUXXBF1nrHpJOaFve/X3fo9R77hPg
hBmM762kXvnY7yaSlepVhoQRRvy7zM2ifaWBm2WFvBNXBXQZpHQXmG02lFmvRV1i6M4XbRa4KCRe
wWe3fYrXKmLu7b9vjoUX60CFSG9yL39U8kav70LQtBnvKo73l5mkFJpljcMKJrFYaV6mtD3s5KAf
MicTjayGTu8CLRWV32xz41Ri0v+b2joVMMtyDrTMvAwN7spuILOiNEQBmV/0A2aWHEAAjLk0LdQ7
Fbr/i4Do+QV300Rgch/AtGbPwdVxBAs71OaObzPVzrLzVQRS1O1ZE1oPXqwU0sJmeA3iZvipYp/f
NTcWIMn2Cf7YL4Yn2N92hKK24QHhYevIGukzFrP3tb1XKuHU4Xl8LePawKVgPRFgHjBsEM9yGtu5
NKDfLGLFQ6bQ3XRSDcP8iC06Xj/a2QlL+Zd5B3B0GQauuLDiMBWEP4oZu5qNBTM1qhGd+ElHNu0u
yKXiHQ8lpWPj11uGo/JC4KUxCRIG0IlYRthwLl1tPfsrOTJqRYrCdiGWk2shG8Y3AG82bqu2FlmH
DAMylxR+B8VtRRPX/Fmg0V+zvnmfj9y6PiTGtd0GtqaHjBosW2HOnNclxsW0fC0tL7pOlxVxBlcR
zY3yp6mgr6Xadkn4TJ0I9r7EwMqgTBHky2Mc5moH6aEmXhhTYGbxR/ozsYuHQVEvhNWiox8n9ZGb
YtpK1H3QUNALZKBl07NCjzo+3vp0AGxFRgKMDC+oujlZHmtvuq/vWUVuo5egEjxhBCXwZs8hXbBo
etWGq2CyYXwSGmpcmvt2+eNuwYObJUwU6+yq7c0s0iHWZUGPPPAC1BUjdCOxh2Ub23o9IbTvEY0C
ohcykFvv1Q8oCMMIS7ChSESQAZS5aoiyAi05GaDf8F7HrKH8OakULHQobDmDsTzzfJbMiAf88Wyi
OWkSmTAMYQBEy4P8IXn7W//HYTrc49eUf75XQfS1MdMclUmua596QmkbV+g7XoyWWycy5zkqCxl5
aUzH1n5CoBefW8nEvWfBGSTtCowlM+UpqgKWuK3MgTKpRboPuoXQkcn7CLaYnBA99bvcLVLVi+nF
Y/Zb1suE/8LNzd0Tzz8Fu6bvLMKTYzBj5VQcNBSJZtL2Eg43jAhH1MX29XYGukF/JpDlhrVii3Mg
JUoK+fY2ZeVjRpfQ0ljC9uWDEbnADgndjGGYM6zQsaz9APZM/5EMzvBM9U/YDLLCyZXel5hfj3sh
vmrshRY3tJRa2KWSYOpie85EwonFfAzMVdOWCBcvgyzIc+CL2wSxev+vJWz047qdjvwXFF6UnrVT
3jwv8tSO62NxXqiy/GEBTjnsRuBwYFpP3T/YwPwRJloazeM+XmDPAr3Zv5fKw/GIbA0c+b2AHCvj
TM4SXrefIVxlki3yLE6QbdSxbP8XZY6Ks5zPcYA7kP4pArJooX/bCp0VgSmJIP+va913L9e66SDe
XuVYE5kNuFTJUWz4PreJ77vVaxIukdV/m5jKQPfusvitpOgMbIjcC428YstaKXnZvNMTaexJDn23
ROHBCgtYXouy72OhzzmPPIKFZ3pEsIp7iYQXwdCANUl+cwIjyN/B/A5L4F4h1Jr1fESsm5rtrsW/
3/sC91oZv90UmcWnzA/0Rf5HdVEdOiywQeiH7zYUGtAeIY4Q77e1H9+n8KZMLmkX9JghD/gE1nL/
hzQUcT+YgB1QOcYviZ6EHXvwUp0ch7KhULjOluyV5NFFh5PDyv91pY9/Fc8be6e70IiMsZdBFaVU
T7Ek+ajgP8SU1sutfCpDesfTTfQxK7M+NVkrqqARSm0XaN68Uc5RM65a/BthvJMPeCzysiPrDY2s
C8KVLKRmOqOqxaQpKTP+hEWcNqE4zESW+ujYuTHKDoRH2ckuIvrEK4UXMIMHoevEOHSruUIWG5aE
T/EqM69SPw6xFAtox0I2/7QziH+hUqN8aUXXVOwo3Hy/IcYdV6bziyhN+V213cRiiREK7jKt5z2W
Y/eR1UAAUXT4b0DJ8pAm/nzN+3IJlWCA3wtnvUBdYLQjeiWGxM1pbfTzIAeY9s6ZgS6hz8UTKEtK
c5BN1Y+sFTkDlfFz2af6/IvtUbONu6qOQgyeC6z94/QGvX1DXNzMbcOneRmaA9Tu5nhW0NFq8Eha
v7hgIfWSmlEtaYuBWKXF/W0o4iqDN0qOPnI4P1A+Clj31s0itPF0fwBmvkcUd594+Wi+v4wFrFaE
zcQ926Jo6WKCTq9Gun73WDmGE4G7XU3rzCqfRhm3aJgeB6SOIb7t6Cz+Y1fyPxWevlWTKcwGRocq
Rvo9BrzjoojDLdg4mho4WChyDH+FsEojcMEPqgZbs9lxgzbTLsQcL1mwFyVLYQL5eY5X6erH3ADz
DZG7tQ0bueqWo7qWzOyfVpWhSBc5++uBvzJwNy/5ACyQLVJ3vwSc36F24lVXbl/YqiDwMAirWHos
9DK80ELQO1t/VuCDh+nmXPaRrrWLc5Z3hbJYaXk2VtkfqIPgnKZkXz94zO+nbzC3YLXUDg6pu3pO
je1NmxWlvuisHnn3OVGs6ei0hvHNMBbB+QE2x/atEBDhT855JfEl65cpjdTi41K9ww7rKvIQYmp/
rb9F/d0pJc59+Pd+DLXYRkmJ5B9wUN4wxflq/NsFk90yBNMqRdxqt2hvtT83Q7Z6SrRTxm8RP9M0
D0As8uYkJYHsw2Dc7UflkSmTR4/Fcv1mt6xDAZ5a2QwGQKz1loodLPeVY2IePFMWL2mK7gfjmhdW
z3I5YMfVTgpTOdJEC1VpVClM1+5XSw8VoAZ5OlSZ+QeZmAu2brHshSiHewhI+qG6firU0AfIpAT0
ArSnYDEtB6sjir21nJhYqn2SfLiGYlX7rTfknP8cCAwRlqEsTPxqqpM3mZMpnG1+ywqfdap9DMmd
LkUkw/mGxDoBBjNGhOlwZ8ql/cEQOcGCeAxHCn6FejepqoRcoQK83hl4kupB5tfeHF3VVhiuJZKP
NEZ6GPRqyROEI4wsANbrYgmjR1Srid2Xlug8O8DC/AXdOjaG7dkuc4Y5Nud++C9I4LBxKqrvYUuv
thw3p6YwpT4lpcj1WqglqlbzxduwEjiawZAvxFR5WTmBxknrvgT+DBohZ4ni0EyjSf4IfWez0wJW
jBqCxgBKkMJRWsKIDH7ipcTgGa3iqRDESlYUn2ceSyGXEWh4/YoowFt/lDHFX62GKEh3UErYROtL
gGbVl+gpfSXV5Yd1Jto3VPKrWhV/L+ZGWcZId5Xgaj70xp/nKskvdWFDvl042lKvb5ruSOwh07/3
Dt21Z3L4gD7yIVg8akFhX7or5GvSGkeN28Un84K+1gT+vzIc0qKAqonXy3U2W4XL7aNlAGWrMj8Q
mYd/Yy+oCuLaklCAMluYtaYqOsnYfEhGgSgahlXBX196GTs3B2IubweZ7OFexO3HkMxs0ZI5vxAa
n7yaqaDEq3h7EQvOlAUcJjZAFAE+iWZCOEP619DPmdw6BSdrD1+QtkcrzlEEPcayUf/Ro1BGinwZ
RcAg2zC/BrHC8WhiUiPHQuEMDz19RWQWLMgRB9Wu325mkEqUUIhAxOSBlSwSBMEeTTlJD7aZwW0T
FIVE9p/trOCs4jzKCDCF7CRGNNuf4LcHubV7+MKQIM+atULAF/l7FV4gN7WOU/nLqtzsT/IBlENZ
WCxZuztwTe2jUgKGrnyqpmB6pJrLwuMtT9n0jeVXRnE/7C/1hnwnj0OK8wCJIsm5oiPG/vlwmPEw
TuXQ5R7oC4WpOuJgykmAYyUozsx+kKQtRuzHb49iurshzG7uXfT/9wA3tjBJiqCEgmFXce/NLSbh
fxzkHlrD8Ycmy9nxe153vCKRxWT6cT2v819Lg7Ql0geC1yaUdSsHqAnvtg8Vq8FD0/J2Yp9R4hRf
eKthLX+hEyHtqzNxLFEos1drIET9WroN2BYO8FWcLa3dz5VphdRAq2K7KPXdroJN50/e+AQbDwUA
JQ7RBBRXzVAJccuyic86ba4uEuWCCgMn7KQQlIJZV2IQILNO+x3vaJFBHdT/OyjD8gJAlCXaRsyI
enSZiPfBwjShrqoj9WGso5xQ3+qE/0H06r1fajf9nIWm6wiykr44/n5m0kZRSTR2x5s6VGtIobVv
3FtvtdQILalH/P1R+kELZoEpMwnywNeyCmduH6yj0BsF7Wqxq4HOn5Q9Z/PiVVA/oTfJT77S8PC6
SoJaQ5l+hy0BCoBLGaltlr3yIVI/N9BeJRxT6baTcXb/Ax++APLjaVk5XJ2BMrmj8HfQqwLpKx4x
smQ2hWBKRZjp1+LJHz+fxpc65vfti29q+s1iuIe0wR8RoTHhgkMA/NRCgyNe8dkMRjGkGFkI4OOt
nl//7QAZEHdvDV9mQwu/BoOvuNZbyBoMduRKoDd89vsjMDUQd3UJew8uDw5YsPqKI8CcqN5JgJmS
xihdtoPlqYrHLvdElHqixF00tBJr9vAXa7xRJiQqD1Nh36fzrtz0V27Zm0vQX4uXjz6LQz6dulO+
+mY7my+pWhchvDhtfCns1xzA0qPhBrmZ9iUx2HrEDmV86aShzPL5Io4aC5ROs0kDnhkMWKn16W9s
e0Nupm1biZFT1BLRkyAryX0QAAp2SfC2R81ZJ2X3OKa4unJMQ2wx75ayUo1jvGGyGtiDuLH2q1kV
P/WGMGoDkdZVLH1i5IuwLmM07C/oCkXUbm35uv6PXy8pyIFIJ7WT9zUqs1XMKWq5rEXk/d+mx7RB
iOeFddlYC+ZxUFDZR44wh0LB/aAW+zIsvOye9zD/XLo/tldilIyFB7xzDe5NRZ4JjDlxSuK0uSRg
qxInp0Pv39pmNk9U1RC5+pTdhqnYRjeTpCUr7fs5hxbCRh8LHl6Bm8xCdwnOvG5O8g5oDDuAszCS
GrU9oR2WrzSeXjtKuyinbG+1qmhfs/Wo+kh+ecHtKvl42T2WY81XtseQKjco4bJTylgDMOU6bwNw
X6nUtLSLJkRvWBuBFGVdcbkftyNNTKMR7Oq+xikizQsWmRxi0u7qyrYxpeGJSgOdrX374p92DS+j
IpVuGrgXVvDDXCjwqC9ljt9O1+dLycybqaxhFUDldtSmXokrsPTFm+bLmxUAfL3oHOTTQl48rRZN
kJhZAr+7nL4+7jOVJ2t4b/QmKqitZkldD3Z7bUWfBiSdQx+arCUOk5r9f2Mcu34+aWP9lvsgdJmg
ZbExlKipNJc3cpC/pQLIFiy6bZEO1ge2Uual36IUJ/D1TWtTWhcGHWOqur4hER5OeTZZdSo8zIpG
XVCgH9VdT4AllwVoIkDGJbp34H/k8OUo/+aeeQj7PaI7WEhtww8PuD7SueXaMvDTk/xRCeLKf8Me
/PIYckMrHtwH+roQehjT7Y0vJlSs6JmVUBJWEznpK4iEaU/jA/zYx63OEHJjZlTyzFFkipGLiCoP
L8hHaSkM2D+DqY+jT+fm7NrhH28eLrCVIwUx76xFEqlGM/E6m2b9i/EPo0tuzb1WMVbJrAGz5iCs
/XbQEGGFmtZPLX9lIxi6HwtChbS8lTD4elk/rOlCmaspoICxbSVp5hxIHrgGQoq1y3xPaJ2E3Osu
jOUgi0bvBFivWy6iG2l8gL/M8r7w+A2e/rC/84FSisZEJtrhJikRt0JsOlIbGlN4voJoyCPS+LQ9
lp7kYZYboOLRQXc/mEEMTV5GbKExfw9PM56PBjtm3xbEmC2jgA1HzhfO5cr7oU1P+DZ8zxoA+d26
3JkSyt81Mn+89tV9nZkT1GAENbRlYLaPfFBA7Xk9CsXpfJX/dFcqAgovQeEpEPEFevOwuPUh+em+
azB48inNBbR3ZHX8X7yF8sMCMuc9SHVgiLjIKT7RpvR86Nn1oDm6UQf1GF+G94b4tRgAVfXyY4A6
HwBYwYR+KJaRMhd0M+RfXbCkxNxmh97IrDPTXcuBt7HqqN9bfvHySqwAIHHqE/2CkiYG+E1jVRSS
0qZmwqfS0siaSIu9zoqXbZVrDK1a7Ic8PzFhQb0uWEPOR9nXgHEU2F1YaLBk99k/UH7TdCRqkGhD
xOX2DVi/gB6hKdnvayygtBNSOBnixRGNGqlazcSNRFAG103hgrw3dQKF0xCC67epQWCn/kv53ShQ
CROsNmvSdBcrvrVQTIzJNEp6VsXjytlV5I2ijq16HA5rNujMqATPMSD/XSZRzhXutzBFTRiKmTrg
U/ZRLFPp1X42yiQJXpOTuZfSrzYbG2iOUDXrdFFhGUrWJ/WlAt7e7sghwMRqXGVyuXpqln2FZpsy
/t7NPCJQTQRREIWbcrPib9N20kv5oGnkq1T9Y1YWdmJduiC0u4WqLMvuFTVzZtJcUvzaOIX64EyL
r7fyJRa4hggjq3XsySh25vsGw/gT44qOpPUokgZUNqq60k+aYm6ihylNckVlA5dBrpckADG2heiH
dVqknJOSZiX7jreQIRPITx9n20oImt3F4DqtVqlkkGeEGC+zmL1EHHTgFefAA81x8M2pkgkQyFxI
mB7mSQBovKzq60an6FHlHojRn/Xfpr9XubJETNjaBcgWTDkNYZkXnZMMi9DzWIK7Akup4KHo10SA
Y2ziNM7DF0O/gaaa8ht+D0/WenyEknILeWzKibWdFAItv3ZoSlzET45MtaEWzcTYMZm18VFzOwFf
AX170Zxd2VmdRdPDhVeM6UzgFXst8EN1qNy48OyvANaAy1b2ppxBILZ5IUsDrTDdhdH+5BStXTcD
LKDWOtVxh027WvJCosnxqbtSoEFxCSCsEYZqLdAONzf7UB86okH5LuuRcfiWVHhKdDRc39ud3qsD
vfNKjgkQj59srm3tOLYqYkt/5akYff6tnLycFus8QMjO6Mi67NsD2eafyGcHWhhgOS15xHtQxuFU
M1/WiZ+8dofRG4pq+z7fv28Un6QVG8bHT+xkI7uranq780RA3oaJXtFwHiP6/Wd7Js8den3PvBvN
4uGiV42WXic0EYhXqHXBLTO8izGp5LHtXUmtbzH79qSGhqIUqTv3B+YounjCN51uIq9Y8oqlszRR
M9CPo+OllSGmHQdRWQpdxaCWOcyZ/xN2BY/8aaX8m3J4COOuynZWngKMf1p1QrQt7EPm9LDxwdmm
RGCUrQTodmtl0Urw6DxTYL6VubdGp/nZvtHftQIysZ4QGiAQ15rH80qPTJfpXyaW4ZHaSB8YwnlF
HRycz68kiTRozftuXxsOBAa/HQ/ic6fptK/HX4yUrTxpXcAV3VBu8+x9ux0l74v4F/gqRjZuzMm7
9x6q0a7zG2fpWdlCjN4V88UG7L3jHuvR2s4YN68uFQbMUk0Cm4LJPAw92/ipzIOfMFQrDv3apq2E
LhV8TjLFqoqq9OHOfAD5DbKBfGnCz4G1IRHByuFrLbFhzhtqSavZ/ZXEqmdtexuKZYkTwR/ffcPu
3T/AvwhqYi3WRiuyYpo+CZxjU3+4uqfVHJsTTRt/A2Pb6tC/K9U8q50XzzBr1uPZVNbLUI+wcth6
cfqMpmQi5Hd+RqTCUcLeiLC3E+bO58mY8k5EBUfbZ1wCcQOoqbfWwW4IO2s7MYelAdCgwFDlIId+
HXs4KRb81BArmBeHqi9sJ+/qXTCufXkGghifgX5rBck+N6qU+uOgOFb6+Sxg4U3aVsX6x4d1NLMi
RdsIvSfK7akYmFOnmi54Phra/Hnmtvmhgn0oCSBneH8+mksP5onoiC+vDhMY5Is1Rxw/Yf4TMaPq
9dHv3AA5XP5Tpl+DcuZpv1rBYYoK3OSX/SyoAyboRMyyMKtQcBEyRgrMUj7NUAJPMqaBQOl6pBQg
Ii4qV7JHljQGo3bPu9dFuW+2XmjyWzMO4YaNySMsmpirJFebWzl9qHCDP8ikAowk2NvgmVSIP3lq
PfI9uie/kieqxBn6Z1ENxqxE7gxFNoofQIbOzgZuptwy/CEjE5tL/FQ4ybM0S+rWlyEYMzROAgOl
T/0P/when8GEAnzzGmZcdWNDlQMc4LdRMmTN46lmX701GN8i6do7M/oZU+/gKn8R9ypf5rNksExA
9SwFj/RUXKcfgSf6/ZBeJAEkj/HAShcZu0FVIZF/CZmzzCWdmOA17hejWFxW2hbupx7OaBujInuG
QUTbDwu9WhSQpJnu2qTNpeVv+INuPK29n/xiIWUtQRkAXXsOhZmQ3GfQmjvWHKsrqhdOjOtycs8W
yIApMVd2KzEW4iLp9+xeWQmsYxTUDPWx1zLUEif5oWblJZBH0A0XID8LZv0+Olxs0mWQMGO37aZa
m0F85UhDp3oIYXfaZ/TpG97xNlAvgPeKMw6XSc7jDlxN1eePwl+CYssg/Gq5Zv1Zin4ufMUIAJKp
HHMnlMMUntDAJYUR5kC5veIpwRVEjsOCBViT2PJcEeB1/4nYW5ryergqn3+pqqXiPoDU193iMuBF
1PKBprq/bnaMcucUBHsLpJTnsAYgnLNUdNYqqhedj13seEN4TsRvHRz1g8I1vRw2Bj1NmcCESs4B
pux9EcbbVtHvF0jsU+dzOQxBiXQJ4wnZWQIVI4HzJOzee4e9FHwgBLfusqjfbJ1uCtS9b+wDvZgH
MnEumWfC9OUJjnv/H+Bb0C77ovTMEygPxr6NzTDMfWOSx/s/5VCalR6P42gpCj7H517mqY9d3a6L
gQK/2zX1gSOP6jhnjJ2nhvvf/q5pIVrBlwmrzt+hO9l0smowHzUxtLS6LftHca0DlAWU+KOPQ6eG
Fb1cWHiPc4SXLsF14LYteqlgN30SiNPAGTtWXiXQPua3dAGebrhe0KA2tiY79X+XvM2c8JGL+9vc
H8dBStNEZzRqzdNohV+qaA5x8cjhqmWsN8iY1VuVXMU50/8X1k4ij1DKimwHL685UflA3ZkjwJlu
11BxNnSGLHLtPzxa5PRM2EhkzNBOZdF2PbvPbF7WBDlxPqyzfNNJ6kWCObEYXRdgcVOd/FPomtOS
b8+SWITco6AOqU8ONI8MmtHuMgl1NgpyQd0f6bRIsWD8UsmqnwiCqNuDBMNXF+EpkTcXTMOAa1uT
ph1t0OpzzXcKQiUdUEcOzftY0YGun5lEdV07zOzjwXBSRWatg7dJS3Li21tTUeAGjqc1cufADfE8
8hGGHyzEVRItmrgHXHvzdbd/vB4YjmBF9HGG72H11QMVqMmm/VDKGfTiLN9k0P+bItZzgcplUnZn
2654NBZZZnpubp099eND/Mz3j2cpU+FGV3YB7FAkLbdJGLXAl2QFdpUI/MkB4wX/6+nlkDkaP3uq
tK2QHnIA06w833P7ML3wchT6GdqvSD+TFHF3yetbQ9iJSlxVSm9/vuYBmlRSZk/5iZUNRxCpiobc
IrOKl4h9rM/HoXevyRc2Hcq6qOv1Wjqm5RTI8kokKRbfBCchfcn5nnV7glPzmtgV1p78EdcSBGkt
ssAPW3QYgzbFUpTMy/+MWXJEnOdA64GH0+4B21SOPBiGMOOhDnqhiPoTETcyTtdT3Rja26uZhi6g
E0phLxR3uXKYrkjxGbPf9PLnFOMnwKa5NMZKqvCAv7UCkzA/dRKBQszBJHK5c1rai8XEuJ5GDVP6
GtYsM3q5kCb/Lq2xhQqvlGl6UX6myBftHZALaQgnGPSeSG4VV3lVwpK6qz6VHwA9pIUXmWAkcGVp
XFkFkMYKNmp69Do8oMpHFFL3JyTQMHYA+8H+PrPN3CVYx12H90xL2IhWl38xVY1Zx33bokH1CnVD
BJ00/LXl0IPW7V+vrqQZh1U9ATVYPDwc/tUjkMcFXrP8CZ59HAwgGS68hjFDe9nrFbzrti2Wki5n
eCPNBVb9zlpiCA35ItYaVDrVaX1r1O3lKYZ07cqAlXpxQb5e00Qb8gJSv9eCys+WQpOg3EaVeYDd
5IoTg8NfXSOJpkRlPz2CM2Ke1+EwBMrdymoUy2cfAHzld469gzd0Y+f+fn018gY2ORPra77818d6
HMDDwHh2cJKgvnC0NK5it3hPhIMrDt9Am0CrzdF9vXwzE9wWIi3uAJs0VVJD74ElQ1IbcXpJdXAX
OdaKZkJ/Mf7vrRnRaMG9lAHoyxyp+WqBe+jVt4ltwGdmyTDrHJHeIitX3EMIUx9iPeY5sDWzaVdH
vFdaYgHtXd0dtLLV/F6sZX2Xzd48qGuV8OK5SnT77neFWHP3p8r0blORdne3mec00hIOfhaCyPwu
nlWkgi8F8I1PqTPyJCWlt552l7+sY85B35tE1lyvVWJ6LmM+1e84gReSBNBIKwGeME91kSZYAxE9
nu1PyxJmQB7X6+NzJmENeOzCAbkPg2Hm76AZL5SuTT039UKY7ie7oE4/uyv3RaTJBPRLR8Q+13b9
mdz6ByqnOiswSXf79dKbH9bMWRHCxKfKwlLVYaqxNIciP5JDJg0ONT0ZbMvz/1PmPNkqUEqinwhb
APDApgj7ggHLzfUITw8u9xfnLazAMGPvy9cqG8gbuObYtGO9d/vpgCb6i3UoDELpbG05ndr3XMQC
YqOHthM/wMafJcmfS2PtZvy1zmh40LNg4PB9SRURLibIElqlxsYYVwt2WbRHbFXWjihQopODIvIV
ni0STEvmtrjG2Oxyw0xcZ7MJaNrqc/w04p3c4MK339yihPkbznA5XiswaYRKF8gL7sdvQWu/R8bz
tEcYiI3dpkHTBL+seMo2rK7GVlC7puyEcGQ54P8KStxW0aiRUa3aEuicd7+vH9iN+ssgWLobFLoY
tSvCDLmS3c5Vy90fN6p5LyOyUrWR0cCW5/pnAPBmuUZoWAUT21vXDzOXijMHVVFPGBWQIXCG0Txk
Fow8hfA4UQgr1cWRavTi2+NJxsEBWqFubVHYu/aIEV/vMDSGz9a/D6TTrOGayUcACMK278B0kaDn
EDWYE5R5Rm83wAvINoWZVKl3nA+rbJNR6EodL47UfKtw6gENJR8ii4nxluW0z6JPhceG2DLdZuwh
bt92mpad+ffW14T3HBRE8kmqOBuKCL4Yo2htTHm7ceSLQRmUKxqfJ6SOOYDc0rUoPhpVVHxUEU3B
fYjuWHlfm94iwtX/cs4WXNYxyLbf0Mhh3juMR7J0a+AZNsXpFEfY16xI1juk2ZaXYpHoOIlaQJ5s
Pf/WikIlx3fe8TNtzxFZL9fbj1+o3TesmdML46RoMQk5/uoOJeqa9RkAy4JqgUEM6wcQYdVH81mG
ND7U2PH7qqNIvMsQkGP3W9hTdcRMP52taytdaLOz0QDZYUMBx4kW+dIVohYBkRac5dF+32rnMOFg
FD56ICUF9seLhK0HjhYOK8+zhnuKAOK0xyY4ysunuRS8kSgHFqF0hzVmSy2D5cn8hVPy+rju3pei
N8+gQ4Kx7mB62FPI2964gxnXdX4yJWywtOIWFDBDci6s6KFQAx06mYVSuDppQm3vgivygW1Z0y+I
JYRwW6frm52Ar9z0e+7blp/3UPCx0YDcwnlBH0Y6SneHt4wN4uLzkk+5emP4BsJ0iaNm+Q+7J/T+
WTKHJq58Vb9M5sbuTwvJ0QuNyyozYk+/wf7Hq+VQ+cGyGqrbWCA7AhUlgOpwJLU75oSBgLSiaiqd
RIF8eqqEobEBdGgTKJfN2iPxgF/WR++mP8fKr9LIQEcQNNcHdvtPYOEwzQU3HOGoZ9sPrnkn18N3
3xxSWEsMGPAc5mJM7MRYT7aatXdjqBYscau/pmA5dq2CMDuAUo089Xe6+kCH3mTv9oT2p1FKWH/I
7DbqzLmpUcgbnKo3auqVXz+eF5MJl1bsB9oeXlbdKmlofRNEP6t/zqQf55qdT4SbU8BB3hkJTL3H
qg5fx2LwPqLj1wzzdTTxVY8phts3NJUy8pGm18dyU9dTklixvttPVnYupJwCqQYn5fq3c1u3G9kl
mU0UesMUC3Uk++FbGNW/fAB1bvZ1h/ePxMv1edS5qYv5UUP3r9Np8LAsTfVt2fyEVPTohuOLmI0v
A5CxJPPE8htIP88KN61e6yhvgy2F+AXBppeLHQ1sCRwhnzUyi705/mJHIHWIR2L/S+lR3RWQTvMa
5DTcv5ku9d1Hq46R9sJUp/r2faIIXfl6QkIDWRje6J7qGlyQzaQPldf/GqcwWsBYc7YS+me/t0Fy
g2B+HFa4wAPbTUDUt22Tc8WD9s2Q3hPGneWlknbRnKhBCeRCPmcmT/ekhOiPb4w8u5hI9h4tHxi1
H5fjThblttziIDJtsGX2zLa/YZ1ccOC1Sr8IoWFuaBkC4bQhMt7icUsaCSlODg86uyuWPEAthFI7
5tb4hT5EVScGGIuOHHcArHCxqrms7DAoZQ3dPU3uAYgySubR7ROjqOgmLM546fYjkxSUbQScWmX8
y8jI51k6wb++YCg4+lq0DboUCt10MTsHjR04gWw81bSZOkkECscuzewUfzp4fHnPgX9rS41A16dw
0QajEf495YcYZsJFZxiFi12oELd6jgBiWevtl1pukna25FXCvvytEU2fxlPi1lbRVKZu2ST6qBLq
UlAv7XiUgxogJR0P9Gvt/AS3Uo0A8CWj870UJeKwdEYLsULsObYKtcISY/ATLmYrpjCKjN6ct/t4
G8J7BQn1vBkNSxLMGZzBDRgvYfrM/da2YcgFApjwxRHeMXEftv/RH40PmrN1elu7gewEEJLTMPB3
FJDxNVUJ4O6O/0J9vG8Br3JbvSPoaOR+KG7Z3gjxTfK9O3y8advCZMqHEyGNrlcrfijIlAc9uxEU
pL2/B1u9s1o86pWqAzarTDOk2K+PaQWoiBbC5eCwsQsJGxzOWo9rtTfC+inv/EtT9ivMMQm8oNrR
NdtFjpyhv9VM2L1umdw2Dz1yj2boqWFkD2YJ9NcrGv0ywyKPp0ZwTOyMM2UW1+WyHF3g2b0uWeYv
CraGheBZ1WBZfOoD5ir0aNxh2TN+eZ85MKKpTE8xk8zSGRlgsdukd7ayGfUHVIQMo8KBsZd+zgRc
iZrxzBMGNURDm0tV7cvJdfEfCvGKNMZ0OZOi5bHrJifAfbQ7g3Xq3ZgEztHdOT2A9x576Ikh/XR4
D+WVnJxpkHyV/u7cKssNvo6cjm+QvxQtFJblLUdF51jMXSweOFOipGpWHP3pbSb7v9vsnsg/zBkh
/R4055uFEv0l3iCM37v7KBCMfhsvEH2YZvasc8UlOewaXTz5vdXOcCLKuOryVpuRnkcITCFkkXjz
cvdtfDEZPEMMOL7UGj0ZkucAD9gRuO5BzcLUAW0gIxF80MaAfTUTmd3HNokEtDbuXJNioRnuuBSF
a1QdcDLiCUpdobY1FrDKqRUTkXHN7ygxoFpDu+UQ3AzF/TPI+FVeBEXyJOEQ1GBhSuq/L+q0XeEw
ahzBvPViHXdT5yNl/LRe9NZuic2gSECkU5aJzXtG13lD8TMFBrp2wmH3YPNuRAmK4dk7A474MB1N
ajS1sXBN4a4HxoQuQD2oaEjd+xb//wEwbP5iV0qnsuY5h8+xUm7lAf7Pb1bGgvlf1fSjquTYK7Wd
SIUeuvKoCbVCqHBSv/Ayqv6fhnk76mc6nS+pP/1J96cYD0/5HYGyyZRPHcbMjghaL0i2eq/TnMXC
NBP14TPyXGhThv2oUjB58Z4qes/YpaPIB1yOvh44AvTaUHz+4EOH8asFLkaX87D8i4R7UgrhbeQO
Qe63Ma38gV0cUaCslDSZtPoKh4U/lNXo2ig7CXepa6NP3kGeZFFM+kOZJUNsAaVtW2OfZA/ZJ5FY
vMZplgmtlWu0o/p0I6/Qy6tjWljUtxQ5XN1mzLWc9krKB3XS3TwKNHcDBFogsdiWP8tm6E3VtyQN
FRR02xJ2iktxPz2Rmo3uBXa7U/Uw1FV9Fst1+jKytzCREV3vmgBLImv9rNh5pY9NFw871rNGoYDt
meGK4rhv3wIizXmHJfTY4IuyV+U31J1An4xt5x1bHyveJePZSMqdNxEodias9hb6em9Cj+N63y2w
DR8KBOL+pcxlyglyaXOXY8dtji0uOuRoMlGGbcwiTKmhZmuFnziZlVTwcU9WEctlUp/0Y6X5ZIOy
+tgMnigGHSA9olvMJkFFlGmQNphf0ZBsh/9I/BoJ0LbZlsa+wnVluQ5+KhWzrZy7MyqGr9KF/6MK
/5rIx2Qn5g4fLRqpVoLffx4ppGoxN1Kd7YG7e4ZHRPcOoFVFotTUk//QUGTXV44XDa42kEyinS0J
scZHSgUi7W6Ft2LR+HPnaMZcrQrgZZpT3A9wNZ4mjiv4DrxahzWi9f6IprvccPKVLpOwciKB4TfU
33YFYW8kpKVxS0d5fGUBcviS+nN/mVf+w6djaSNFN4fNbrV6M2MwK3kKYIHS/Pwn1AjSAixGGrkA
AuO/fpdrO5UUyp+MZIReV5Qpjz5TBDkYvNOlsA2cwKozdrXxOxc05Gj+65kZJWWGqibDfAk4MkCY
6LSCbwMm1xg0Q4/f0/vUB0oHwbzRBlfypHNV1/3IEuGP6mXeM8DIb3ynXlzCebZCBhz0jzeD/Sb2
Lsl2zoR7vrDfIF7AW9y7EYVO2Nn/88Co9aOc3thtJ6dZ9rmSH5qRrEC9K7dxxmTjxhFcyxeO7pP5
neOcu0Ey/Rf9Kqh1sEPpBi2A25LVLRPvCjvyMpD2BKwW2EWJYNX/L0bzaaUVlzFxhe1PpIwjzdOp
DWZdsu8TtNCNl8DyiFr4PjXiqy/lMfNU5ncZxquFB4l7FmBB1oy/ZkqkGJzrmCqaLH1EFoz6r+Ic
++NgnoAl35tjqyRrx5CtmDxuo9uFt6gFNNke45xucBhSs2XDhPnrEhgrTC3KVwlbaKd/sHMppJWK
5sCpaVNbYbT+fjoUqXQMSrsY5VCiJ1iVpPD46CDpp/zwlgFATxY9jSC2alusWi2R6PWCnzBvz6jE
hw6hTjBkKfz2dN01/+ygox7ZWNEb3m1Zi3U3MUM7TbPchtdxzHLneYAa3trtu8ZPBRBYMSB4ysBc
7m7qhNWU/2pPnmJ4roZQlRaTqDYcVLBJ1QcS8Jy2b/E6D/oSSQlT7g6Dv1l79VznvW9QDKPn0eVT
XZyFaV2NwyLbgLUC3YDw8m/QNae86h8tdCah1bqIM4OeoBcckuChv80kl0H5MgMcUqd9jk8rTKII
TNA4xQH5kqSFMVWvqzc3XqW0ewFlZDTW+CVSd3oeCQ1fAPE6sEdoRgaZOZc9cggASHnJlU6pxoWt
ugs2NHlQZ8D9lVi50bIIvUPLPHKCR5G/sCawkXDo6KAKKUcogfPr5x2d0LS4lzr7ccaswS7Ulxbo
HRua8gkvHwJJLK7l0Fr1dLVjeRJeEWmD53Zcm6TJcKTR/q5ti4CPMxJldfZL6bTfzEw1/6IN6fCB
4soFdipD3B1+1dUbozu0PHzT10LXsshD2bUAgOkWWmA3GNUc4CAkWcHrZYIplyM8f4hbJ3AlMXUq
at4akQQsItZwy+1t4YECPU1rKnpBNdfa95B7a+rrbNjT7FshYuZg65pqyfv4CTW/2izyeTnPGSfL
LvH89B/rUsQ3fdA+dJbOqf/bBoaM+Bp/REiZfRlpKkZ881OovlAdNTI8g6ryRLHyTewUUnRDKmN4
9WgKvpEKC672b4ihgHJoBsN5qVI5RqPmDIFmAggbBJMOVfOi1tDGKgZ6gI8II25ooZlc7r72sGRl
nPaio5VsE7JXg+8+8tqH0Cjvb7HfitNC5xIb5JCgOKRC3OiogRs6FQkzwNyf9wjO4dtHutX/bkq4
fPmzbkLxTsM0ZnxqPkMehZpAYakOeCr+iFLXF7Ds/83I7H1OaSUGII9Gm2dMkoAOiwTfOxOhnYsv
rEzUqSFQa66y3YFbAZ9OpFODtGbU5XViNDku7+25l0OPfHv9KrFHnOZmEuuvRzSnxcQLUse6KtTy
d+fh13JlHe/oBPV+dR2ncKK4a05LLjYafF8/yZj5OZU1UAhBE7eeVQng7C9X7yKiFFZ+7N+VO7f/
b4Z2vlsFRPFC1Opgeev5jbyIaZiHbqlR4nJQQ3dQe174kH+UEEdMjshe5P2xWkWPxVSEuN30DLJP
aUbtxllBOeCdJtjE1un2DHSQvXDsyVPBMias6y6kcBAKHIHY03Ck8vJVW+yPP2JC1SUPHmep6mvr
VkhaIXGvnEaCivz7wAU84oStcHOus6m0m4TthnTsO2KuhQkcowY02NaIemD1NXXNGxkpRoFBTFa9
HzkyaWAd8S1WQ/LEPztRSTXMiczBaqgcQdY/YOofihZYCDcWU/j7CDDjOee9k2pBhQe+n2iNZOM8
thfXaeovtOX1eRZ0AXcebrudaNzWPCSQPf3Z0pPml8CsV+sOHzyyScWguLlZ4NM6DMyIsxCuK+4q
8Ihd0HVqWdDUPMhJC8Cue5IzV6w4CPDq9dGn7uCYflIphaI6GwMrZacDj4vLoUPl4KtrlusUjw01
TdFLoIH7Pt7E+zry73JBwFxQcMaalaDt9o8fvvO/4I3bt2RBkf4r2ClchahgNXl8DHEposzuOc7t
5T+hi6eWKMZh1myU9EShq9CctyfIIU/LwE+5h2jZ21KrfYCNO83G753pUau42vOXZ+/lITj8Uzrn
cZTiixiahae9xDgwjPNXSLCoPPxHZAAC5OmCBB2pG3bvvNQ+DMUsf1TtUkA20AMzkZy2YNuAz+VH
SlUkgGRxCaYxQWOmXSsW0rqbSO8UG5m4c/g3I/6w5yNljdnSNjeSFFTVqbGeDu0vr3qSaGJam+Wb
J6dwA99c9vO6EGWPWsXQ2bDIreZcuX/Y3nYln2DYjx1yRHpVQvhCvgQYA0QbT92LxUEm8ldlpn8t
pYspmYbGyU3Z92qzxXOho6d8mMPEDhz8KqxgXu6CA1PzX+9GjMiwadHGcLwhllHT2efm5owY4BLM
uV+Yr1ylV5uIuP+GI4A/j9L+S7TC8OpiRv0tBzl5cZPutgGOlVvH+Xtxiicv9A4Qp7k39nszOZRb
tww87hWeaGxtlCMJL/kI+31yntTp8q2WeVeRp4XRWgwzqT6/pvG70sbyojzOLF1fEUTaigW0aDmb
Wc/pyRlEGoH+4cUMevLNcfMdDpxRuAI3o3SANYT/Emq6yFVqhwpFZMKg7JZT9MMEso3RqPDLHrs8
qar7arS2gPGdm/u6yIk7Zo9OTeWaE3HiwS7hwELt31JNQvijnBHOXb1OhSfZscsSHu7hjKaSBFnk
n5NV8nGjBddRYJO53wXCnsHcg0kAIS9SmAAxwFtWd4cAi1d4tnxfelvmX7qIzAtPOK0TiCbcG5oC
zxeDqOdwUmUk2+eGdfsWF4Mh8XV5fXnUG2TppZ9kV8/+bGsoz/Z0w5a6YEA1I9rPlCROrLRX9bXQ
qDKYXh5U2vbmREFcwBrRsZQ5K5DJK3TZs5k6xMyVAdVHnyWDR1FOEsqNGU428Pb+XbUBPZyRbwkm
OSh8cEc/tWi1QwcjTpchXi9dlFx50Ys9JDoM1EEJGFDam84lACv2I2Vo4JMDmZUIYohfhwTBEwxH
mfRa1DiZCL2QTPS8Z/FCWwqdhx5xUxcl3JI88/XAkFtDHA0nh+DUs0sYCSFXjw1q4Q9nP1NuXLM0
8hY9E3TrDGWAhn/TNvrpul/f3sK16w1WxU7tXvkEE4c2Sa9FoHxVLJqZX9NoxDiHvtJpQU3H5HHB
fBqpDrkIcgxSNAd5Hh4lVqyhl3/VlLasBNMS9XWE2q633kanjegkIPTDZNCn99rhEbuOUifKQra9
ZI1Tw3FQi2RB5oUQZAQDVNvPqDUnIoecpP747csGOmO5WJ1GxDFSK8vIlJCDn1PEjDmWbMvBTvf4
GjQTyYYxw99kLukEtjWkU8nPveyYP2+AHvBENO7m+JzGGogAJMzSdoLz0q9c0531SJrEhiXrTld8
W3N5ZSwKs4XjHmk5bINu8XIuzn7Jf5HJHduku+OqB/aR/1LIl620aXc+3kpsaKU0LqPLXqiREUlL
Ng23XJiR5V3b98ZJV9Bj6fjQjLdhRG2nZK85xy/gWTMo3Qg0RdCrLXS5bmiv197Zc2I3YljjZG1g
W6u6kac3WcDTwXP5IYurs/iyPgBc1IYsORCH54RMLsR0fK7mjxLtYKXw+FEOWgCugXwaAqCoSTPI
UCFnLEAsYT6QsThrQ+L25kvLOkibkEi/e0I1dtJeyQG7MrjQffaEAj93ZEbwNnZboYT/uCAGrcub
XsKBr7drzzBOhLQVT/2QIe+ogel1Uca+sP+Hq2QXosSwx4U9M5N/XiLbx9vSdLfELsUeh9rxcuSb
c/KxfAMAF3zsYUNBP0zV54NkKJyiS7Qehn245mhpa7iL7DvTi4HKxW1Cke+69UdJRYSWwnGZiZHg
7GlKG3aThLUAUx2nu697B8kN/geB7/beccA+RyztOyjeHugZ1MG/kFwfRrVhKVi5qLdp9n12KGvk
omVxIOyHaMjovMyhSwM6xJU2pMxoGyCLDprSqjKvlWSzU4fahQ1zxwWab/jhReMa49W6CGbXYJ42
4zp9+s7/B/RDG68Tz2v0eTCbZqSPF+Ns6b60CCxiovS225JhhZ8a3XRdJmJWGSLuRCQ1X/+T1jgi
CWYs2Sj7gf3UCZO3e7PI6x6qq2INgOCV0Vkvo/rAVqXXYSV+Ml3pOb6G/P7krgZ6dcaBNSNcok28
nvmIvVmurci9bJSfitVTs6E1oXH32jmOjSv+zZaSpvYWiVlKQ2ZD0a4DxADLUAmIjK4438kLfZpB
qoCHmblsvyL7/260KYmoLPjecEY1wLzBqAyAUMFP3D3iWcSi3EWcTM4MvDOPaCx43hbyvKv3mDVh
a1PRD/jIUvO+ZuqzdMNS3Yi25sCkLtLo6J/pwdiIeHZacivz9g/Hik/Q9EurYZANPd7kQ8pTS9pw
qmYOkVIBpvplpbNeMR+FHyGosvIcjLFFM2C5iIxLEpIP9W2cb7uz6jNPPRjHt5xw0bWnkz3ACiTX
uJVRGgh9dn0Pasj5vptgKPB8xsKOvsTYcJhKKEu+hzEaCRxbXuSvqoIg1dHXziruA0+OVs1fO/82
FB4Jp4rKubAKlqDg6WRa6L8keZ4XaVqsTyPg+3L+YHfTyMRDVA1W02fhwi/474i9BMRhX/j2x2GJ
KsVGP5RSR0bOX1u3flhuC4KawdZ7ZKjyyTrYzGzKCki91r4A4veOTMGC7WT6HflCdqqiLCu784E/
sK6DEnaOhUjVrn4n69fZBRPNmShafhdvjDpa04BsTNhg1CoPhwtTnmacYCQOlXvE1UA7crH8cU/T
joYveeT9oolUVF1avloTnQjr639emtw4JmDYBdpfHR0NpqE5GFov9RXOPkeQtIYk5/N3zgOGu9d9
nTjX5YI0ntMjFXuBmK2p6GvGgcWrKRTkYn18nFYpzc1pbBlAZoNk41AkOxj3ThSR3owRPbmOVpeP
fw4QUfXNTM9UdkjPMVKSDflL+dRR2d0fedYB0b9ooKkrrZTDTM+YCjxfDayxARTH4J6BpJOM/5FY
IbEE3ajyRFOB8sPeOFJxpiFeVhyILm/AeNlLYU2LlEgu7XUg2xQPxurVkjmBmiW3IiAq0jQotpK8
3lLIuiXTRJQ+HDmF6zF4mqql3jw5FZyJLyiJHLa8ochSly2TsuLlqYQ3acH91ilBSqXu/h2Gn1K8
U53PDpO5sujN0wzUYdI4rvepIKz4dmbGdKq13Q96ltZGtqxA/vxImbLEmlNmCYaNRP99tQdi4gEK
/abj9ygg6FQpS+bPlgzFR07TEVd+AsKHSf9BG/VY5e/UcjEYDwE8r46W7Qq8LiomXx6LokvWRuKr
7jIvwPt3K/gtWPlfuWEHRtuBBrVixJEc/pPprUbKWmSkDS4GPlx/YCGlyq60H9NBBlRL5g/9s+63
WMnvxB2X2zHZvetjUojh6ZdK1ZSMxwedcNuFTFpM6rL4hI+oonIn2uzNlkctj3aC6Z1c1cOEXmrG
7pME6CEE1aE4JWptsrgxN86zNfePMPvyfwhs6Jms2dSTw5g1PSWBp4zK4DzA0lgVAC96A67aMRxk
ExOQQwXbxJd6LHsz/trujgIxBD9sB4WnGAhWLlq2ShrxeROsivJ22d+q27pSlBDWkbOV4rXFqha9
XfCQUB4hLfAxnakqjMnSvHVPLO9bw6xH/BRxeUr8XsJsMK9nftsVlf3x2Uu92iFKd7lzibPxu/Nf
aFae117hpTioqbOX4lJkEdvrHgf4onJd//reZ5LTTkypJiLNbSuK7/8gfUOEagKCCLaHFvGqeqBw
TJMPDx26VmtXvlPhk6wUwK9Niooj7kyYTIkUb0FPycH7m+ot55nrjRACGe52pUmaEnqkih8+I7TM
iUdUrDlFdFgRQ25j4oScETInG+FjtqK5dCJLiFWsEdMKXovO98rWUWBbs0fD6d2RA2fTDu5C5uzf
pRYlbMPWFzWzMH964dCaR4kHuA+kCELjBdzM0Q2LbLSoTsLjh7rIF0u7UpLkWdxjjrqDDAGMYe0/
MRYCb3ojQj+Y0D9YAdb54zPoH+TTXobzh7SVPi2/F3SAVzcEst2qtGbZQUsEiyORJycWRpG59xoO
HWeAoP5RUGdr3+Uwpn6xwgsE+Rm0lTKqi6lswSZk6OvH0EMeWcT5p1+9NoO7O/KbeON2zqtSQ+kX
pGu2Z8iTRCSdwBq38qn0Fm+VN3sqq7BAhPRs5a5SbgQidFQptsjeYD2x+sjxS0t2P03p1ImGBA0W
6MKBhrFoneDmXRKMeb3/rjIzoqKFck+QpgMKKPwB/lLZFAIKzV6xC1H3OXHBWh8Sqt87uottDXfH
F6iNZrsDtyTfc/uY9wLC6aiRWMnVrFw9d4/Ofbqz77Zl5wcdGEr8OAapsahClpaeG3Zg7qeTqCaV
NNyOe/1p6XQNxt80++Zaz/RoGKV12mUACUcu/gxTWJgtp+vLZWL3Y+BLsgiCRlSKyf+JTJPy1HSN
6VGy1nYQALwgtwQU53+bB19L+e6elJDO3nw67++KxBo9EJF+SVHcjQvolZlJrGb7LHX0QkTPPOE2
N36zrcej5r0iv6NQ9RSXEtXUkxj34c7yTw5ubtVlgWsQE7GYy9+xfhxzpEJMpBQhRORPjdgPgx5J
RZAz/5F+0wMK5ql4XfmiM23xcMeBTEumRU/NuMS5diCmZHzzKJDb4BcS3vl0qk0CmO/vtGW2H8cE
dYnLgqzYgsZscCT5rzLsDVVDftQRxHiDzRKzCuALsl5ZBYU538UXikI/ETIgcUnKPGb6bCnbb7sw
I4lQEbFr8PXdgNL5+4PX5/ULIL0yrsQjPfQCCFtgitkRqsDgOpVUELidxfKsxg+mL2DAXxXI12ks
S9vznkU7yV9vZ90ZBIxcJncafVVYsZdVQr4dlxSxT/xSPQpJ7eYkJ6lhGJlbjMicn1IlLv/mqFom
7nSv5fg750smpJ1fkOJHDqms4VPvwv8syOZzizjJ6PmVmSnv709JuJnGv8A3OPZYljr4h2XPOxvD
6cMKWVBGRCFE7iRBSkBPpRBJSn5fTVr8PKo61os9MigwrmcLVlbjOLLAgR7zT4pkXhUGkmNXmdS9
6qEsoEtYfV8Y1ZQflRLGIFYqXVAZ0qYnvH5mWud7uRKji7Z3Y8ShBOvsL4lZAqb+d2scOmvMo+Du
gqg+3F0fZnQOJYVqORIZKpqICTr1wCB0CoHrfYMxXJy6q4jZiCSsrhdn80CTxzoun+YZohB0FdAz
E/gUiczsvEyWtZ+M6gZlxp96oPfYxh9UQCzzt8gzTt1JO/XdrhOTC18jtSR4APITicA9evINUn82
mzkkYHJSX5qZLfpGcTHSRzdYplG2cdcan1jmB8U9nMcRxVWxC4N0TbvVH8iWxT2uXg8SBtKGJJzB
eWg9jG1Gm9LT5hyjDxAkf2TtPy/kBqx7FdJOxA3r5EEw35K2sotMXC64KWodk69DyKMew0jWdsjf
XVtZPMtSvGplUG9ETKj3T553GLfx46QiuZYOMhV3pAu4nN16ROYei3JpqGM0I8fU7eCgCOWt5Bah
eHxdx4k9HozlpJ2l11cZR1IxqWGqrERP4ZSTpQV0jTRADOwm3EhRmusXBXj2tJxEGKNIu9AjrMRp
co3Q+BUaQYVq6DugMy4QBGoaq14rZeq3XJbOffTx+HZFjVxvxgz+0COQjjP7Qos+KGXOr/gc4/5M
GrIJKyiIYawuW5TRby44JGnsusjXxbUIU5Zr0Im9k/YQ0E8Y16KqycqZuqOaeBH/RjWM2+qUdA5n
am3KOW0rJMN6zrKhYYKSYt07RQvIyPYNRXjExonzok7tOvJpEUmENYxFdDZXreiKcp/rsqKVSBk/
EHEdifh2NfKMzwfmzUYQCCTKaPBfzr0CNCw5cPAlIh/3FtaYRmiAxKehHH/n3qM2kBbONJOiONXh
mz5B/7zyl17u4Xrc7WwqcU/njft2o8/iBnWdJazMhBU/+ieiZBLrK4K5IwY64ha0vpq7+U+8MSy+
JT8GQwyf+vwgXE9cTr2WtbHxkIQDbGiovgz3w9TL3aeMTlKuFM2OhwLAeJVdrtXoJ6ErH9/Ag41o
2c1xYK39xe1h5S4YHBEeYGmlQdESDELYzZD5Z72FMPcYFUmhYU9r8GkCiLkGG2G+Lel9vYyl76eD
bNkI6f1B2ymLnbkqHtltQcyJJ1PwR7yx4eIU56+tff9aLRnMZ416UQmgowD052WpXhMwXlyjxBtu
dAKvxcA+tjRnW1d8GxgdpXcYIdBEPcsH+ZhV0AKUdofWIxIkS+5ibeJ8m0rAEEYzOq0hFIISbz0r
kwF59SUCEHPkTDMSkVTI3DQUqMmKA/uvjUNeFCgFJkkQPI18Pdc7YMV04TBfNpShec/XAtGUP8fn
HS4QmuJ34lcF3bfFUNjemxNmte4C1/6EPjUCMI2J4hzaI8jk1icJFnMttpVhn/CV0RBnGX6Fqv1g
vBTgt7Ls+QTt42ArbNdGVvFLST8q+rGQQY2zIDXRA4aQqngdTpd9jHn4dTRG1M1f6jUpf/CtYtHz
v4X1ufNEAxX6ufSOsr0hO+bSyDAii/nrV827XMIlvOOcrxXwM73RUktZpG8YbgX//mJ0ZEqM9RXR
FsdYD+6s+e2PDZYboSthJkMUVobTAObCR+RxmM9BeK4lQNDsptQU1Cyf6C6yJJym7G2sLVF5g/9S
63mpxGS40RcTXNQBvvXJ2+aQBw5MZ2nFkBvBgJRRidtCg+gMKFmMDIbF0ZH/F0RR0Ihk1zZ5NUCg
WAfTF4w8642sbRyOtinjRTHhi9YczGrFaevXmLgQrQJIOPLiA3KjMdUNlkOYJk/s/CfRQoMdaWCt
8kjXrP3EIs3cTpcV+o24PNxD0beu3t8tov/4s08IuNYrzVX8j96TutCAOnsDikZ9LmlqKhlTBPHB
xGqinaRu3pq1Wqc9zINN++smwGLXy8/yHf5YMSkVSz0ugw5BXA589RAVvVCXJHzjhAfd6STIAusT
+ZUh9LZ70PsQl/KwFzt1i502eCSLg27hOU/3FY79XIpBOzNA+c7YJnT03YDmoZPNG5tVruIVEgmS
OcL9d0DRpITFkF+AMXwXAHnWrM5oYEOGZ2fJg8LjI8Elt7Zf/XowVbk/sLJ6PT6Pkx/rwkqRRF4Y
mh1I7YFZ2wVlHSGqjtJVuJMCxwWpX+2LfcsV0x1lZgWB2+cymM9DblagKJm1QFkSCHxM2MMhIpQ8
3B1gCBU9laaBolHG69OlEyIPom9wxJ8R6xbPM/ePgNX6S1CXfvDqIwiw8qw0Lj07Qc533mETPRaX
k4SlZ5krM0NfU0a2mRmnkYoZksJK8hGZTj3zOwD46Tc68iBLEC9Njg7Mdk1IWo6GxCyicjOGlUya
BhCFdTtobkqVhZgPWzfog0wXQns77KGZhfTbdII/FOmDaTvhVb2rUhdnu6UIdBAcEE5+wihknzMj
Ytd/WUrziBlXPg8hbEnVO8By6+vwjx0SX7nz77qvd+dWP7CQWLMxIkI2OxUN6l4IRDWsv/nQuicS
tpkrlexNwfJT2buGnbHQ5WTf4tgHiPWznOOeWrOBHf+oktqTRa20rTw6CKwbbO4/VMOPN2JKAffr
wUhv4ohxRw3sPQtYzBcX2FopHIlXrq+nIV7fEl5OVNn8X1a+KagXmCBAydFQ7CG2YdTubAoo1w9O
ptqxzvAmx8RbVdHc8HtvhgX8DB4bsTGIuAXNHwpUNGNdShwRT6OJvahWd8BghyKm/8TKX+0PUt+l
IGvPy5wunzs3SUVE5cLvyUCVKpwLL/QIyMpKwYsI4ubjYwwSifNZcpEUPX1vCIwYikWVcII7H3fr
+HOfyQZC6vjBxOE3jWA0S8dpDobjrXuLnsV6zDQzcO7d6Z0IRl8na5uYffX/qGjDUGPwjR32xlpd
neOfxSVqlbk5nODmo5CQ6Ychz1WWb8q8uTCLdmpVoySrR2jXeAcb8iT60lE7oARA6hEeox/LnxEf
Azhb/YrSzB8gPsNQZsVAaTOhWwA0b2e1fibRtC1jGKHpewHlkeua1hO7Ipcrl0PmjuVTfAQDHJYB
6BxmAcVtCCw6ilYSzdjSKYvJVjfmzn7RJvIIZCt8tWldfwjM7rzEQ1sfd0I6/uNYRM+oKkSKEMhh
7JTJk3j3v6tNNkO7hf1eqIXwejtrInv3OcuUg5onBF2d/yuJqOS+3K0I3OCyAztHASz1mA839o8E
dyQ1t91pgF1TSW4XxY43sHy8gInCqlxOI9rz1ma2Tm0iPE/kewvsHc8Kam93TcjDlNSD5ub8alUe
7ockAIGgC4x6LcF3Pg2dgcuViIJevGTy2ZNK5OXQfSVOpL7+zhR7LqgviPcpq0yvW2AnhXRXGmTb
VBS7Pv18OzaIixunIxSMBZ7JmdSxDRI57Bb4yjVEmLF0gSqo+88Jy8kjd9fxWluXYnGFCz3zAx8D
+uQ68Py7mEbvaBgrE2g47PN4TYKFVRVLCSXSjOOT6xKXfZaKKWw/VvC9rokv5QX2Js9fjspRP240
qMQVJ1VBGWvqZa3dCdNviWTzSUZKsVpbPwmu3GlgLRFIJWS1bdBagbHMKuDsHJdc2pWmkbWDot8J
YQIL/hQJOi5oLq79Wl2IaMzozukeCZYu9e9o3dPWBDlCYVBZx1Ok+tSLkbh7V+OUwLrevzLIZWNt
p1XOlApx6KcYP8YHYTmWj/t0FjL52Z07KedCmz63EbbKURPVPhPD7ua37Bj+fC6gm8x07p9GYSYs
MIoqn6Xd4G3C+7q/1Mrz/0Fgh/xpa+hGZRPO8essm64BCD7LmpIoKINVEWMkcEeFNEIp4S5EpTZJ
Km3D5SVarmdGvvQo9cX17M5Xp7HM0TsPcJ6sxRdolgA/j5mCVUGM4/rPRxlZ0/AMJnkA133geDDr
LUuJKJRWRrwfbbD9JxqJyRx26rw0r3q4+GO0P0C9+YYbabRXQKM1MHFgAEABtfDswFA7N5RE1C4m
hvEtu1EQBPB1B808Z5b/mr/C72rZkiT+w+9BAD7SU5eYSwlDoAkf9EfPw0jBgXbhloHwd9Lc9kg+
R38mVs0agDV2OBr8VOyL+uKReCeM+laATqTfUB0U2SX+FRdcJFuzuMwgC3YaaQIeeMaAS3MpLkqj
JeEKG5fdGWZ6akwJnHf5dHfZgyqqOFwTCcPPYArq7KJGhCvxjYzEdA/ck/8+3GFmxtjdXXxcp1fs
vW/GlLJckRxIstGScqp+eZAxLVXRASt6s824MnjNPXFtsfiK+rcCRsLx8JSnsCofzOXLC3gvkJAQ
gvVllQoAwjEhIWO/6RMvQbe/o4SBH41gi3BnKH8t1XPmqXOYffabasZ7z4v+nz3jmg4O7K2rmQMd
pV4VhpNfn1Bd/CjcdWwq6hJouHdDYwdScfOKo0umYyURfOKLNt1IIirlVY4YlbSHM0gOhybPHBwS
/iVGOnvzrtKlQmtMWmekyIB+/O9TUfJDMExrPwldFuo2PyAnI6CF/TsfZELZ3QO88/WPxLfWyKJ7
cErLUvfLUOF7HedWCKh1E8sr9qcKFhbL1uYr5YfV2oat2SMM4GCuhqfdHXVg08NqaXy8uIRSxxgQ
n+Ebu935+ON5LEAfgbRDdm/9RFXV3Iq3pULuCMIwdV3sDxkv8u3fsdUIjJ4uw2bKLJirQjc2sjdS
uP3188QYZR0HbrpHLC+liacJKPtp5XQHRrnlkdwTMd6+kmx3/HajgB58kvzfwvmvK3fKHEZGaAjg
o+5g3TGo2lyoh7pi/yoQqDWMzAS4G2TXdWZzQiDbznCE0YY+MGpXknbDxy8O7fMtdEEyIS1o6zi6
dt8bz/UoiFYcutano+wslQB2ySVEtohNF/ETCzJ83m7vmQCGx2c4gKy12/4WacZdzUgQ9kVNiCm9
bPRZ5nk6+HmkhNfA7mPcaOPnoLdTjReY3epu7WKfYFxG/7czkqTT8Puy/jUE2g35JY4LBo4X+VYu
9AOPOyjNjwOoAWOzmM4CcWbvZMC/wEEfpMuGEpVkujJMHSYaU9CYmezs4W7fDZJ+cXMdzUD206Vf
3/yEpMhY1dNRlHlvm9tWJJzBeJZXda3oyO5v+BCU9VZaZDm7C2bvAC4t8vL/1d5NVKjasjBuk05g
vaXS7NMdoTkjZBY79RcW0q6zkEy4xO8kxZCtXMp4PQWrtcyFGpF9Yco7UvThbHhfDZ2fCPqX0unb
FmbK5GrhuJtPuYXUBtUttLz8h2vm1TwBjc2Q0/zsB2RG8gk805AZaWvekHTUA9uKRI68JFwGfJfR
b9DARJG9lMfKhc3AhgxoCic5pZRcv39wNEdC+PypfaoqX/ZkANG4MnZk6ifTS4bO2mXM1kY+Qvk2
VA++/QBVLdoh5EtSG4BqerXYres+PTMQoQLuthud94P20nxoE1MFRsx8vzA0VKu7xZJaks5a9ZW3
gc+QMJ0FWZBjG4bcZVYCtpKP5f9XHjDPSCcNQgl0HbCBunAJrMDHemv0fDXHOhOmPie+cZGDUKHd
5VX23OhN19r8RiOfS5fuhKso7InpPnGnjmdqbTUSzXi3sU3djxuLu1KHzlHKbmf62VHhFCrZt7xF
3UVQO1fkmLrgAtCeUIdjqNwp91WIohx+gZFLwGNKG4EhWqqMs8MWYzt3XuB0YUJ24+Bj2bZ0OeEQ
k4g8Y0DfLSC9e1/Lyowr5bHVyWJzc7Fyy3MGTRiHnXsTBzmxtiXzWi9clcE2TLOqM1VW7uHeTdWy
YFwBYXg2Nk2fKK2lKkJQTMOjLR3wm88q0vW0w7liirl+4sYnr5YRZv5+IcGscPzyBpXj8ACuxDqY
GcMPHXVMw0nIvCDvbUbiBWJqfDpNl7QfhbKkH72Olb3fHlY5JOOvi/FUs4s8WQ8Jo3XIYLLuv+OP
kimBLgWED2I0tyIVb6JQ6PJk9yZuCUSv/Gv2HUEPi4eqZwiKpWZGhAaBXZfi8/l3DCn9ATfkqz7A
H4J1POKKJUa9yPhKnQJmLnKlfENRERDD+RVF58dCiulnNyZ1RKdz1rUBFZ40ZkSQckt0oErsWFrn
Ssz6eCiGTkuyCZzkTJjKAlJLTKxvKzkF1FQrBEzSh/i41mV2Wnc6GXZDhphljGILtMbTjapC+mKY
r6F7+J4tMhgwWNYZ2VOhxIRp9Ugcpuai4nkdlN7xWx4F5NgOFIUUNg1W+8Nr4soxGvP7odPg1BIN
wx7qqBVFTB4LQxvbAwD8YCehTirlLohklX89dJXdJD1jjBoWl+fhKb7FYGamOuSwFGUS/QbBT9yR
1JXk3vGgUdllzuWL32Uo4Ixyc8pazkB8cLnhzgSfYD9L9hhrE3ZFWPxIIaKEMHa9RAgFZ3HIbi2J
8EIhnU0r2vyxgHyRLrjf8bjKlHEGfb/Rr2ZbtSih27hnwNCrNCQT2SpAEAqnw/hqHPL5hzC2IEP+
kJpx8BhlwJRNDiGWLGfY0In4M8kz0qzKb7SFpDVUwYGB35GI2DlzdTO161nyGn8nS4JsqsGADTQ6
AYo8ykhYgWWiM+xBWsxSXaqSIjh5xONPjNbm2ZCblMupHd//sB/Mf8DcqJxnnYjLJD1L908Zmcui
6OHfqw9BQ7lWIQ658OtzRYim/Sj86hBCzUS3R8nJugPRoq25YPQiK80nv2gVLriogce6YlAQABX9
+eG7dWrALQrkcBc3pJW9I38rXqxGmE7qW+THTQM/4C9U2Q+PwJq8Kr7g9ZXb1BCu6A38RwIp+HRs
OZDGujFDp0TAHq/Jd9hdYeZ4jX+e4Ux50aWtkZpWFCrMj90ZU8esoPh1wMrGGWgfpTtHP5OFGBef
rnnoMlLpKg9SVvDIbsaCXDNczKimw3iHj2VdIVtvsy4ktR2VxMKNHK0Cb3XJT2oSzl4eSkLu2WgK
n35qyu2IUOB17U+frwixwYoZ7GF94gtPRHiTro4Bth/wNs2h8McuFJ0H/9oqiE62QJiIMFuf2Imq
5iwnwDI02FeScrC6Nq6iRBglwEYbCI4aq1HROyjih/voaDylU5VCH6sJFNKiPeviMf6kFlBG3eNx
pgEIVaZ45tMrG1qAS28epWS0FKEBLzjia7eH51kTVRjllj1JcxczKpEoF+tP/eeEuuXpFKOFConw
29qPYko2okZMAxTebhjkeRZGscINjt5O4ITJ9MIr2xv5jUJ6oegz4s1xbM6ePAE+HjU/uwCNxX9d
NlfHMkiK5jW4h4h1hER2pcO+/OaKBvCSFZFLCrLeFUl38m50tdkCtfk7yqvmMTOLqNptJAKa8JGF
fbuFk+AbYNXBctat8z/WDCt9ET9hWJ/W1j2iQyO884Evspg7GqBcL77Jy6rm1lcwmEFcm8NST3T3
v0HAo5Of8Yk2DvPh86YZqqRHoVd9jt+5GqHa1XVOh2gi7C4p0maUb83PjdXavphfrIkphoSkOuLO
U1hHtByXixDd00YRmyFyiFuAXVstwX5+TYybQOEA01kdqJC03snJtNo0FiEjB8a4+Ps7iZMIH9gQ
hVfr/4cQS/cwMUBJhr53txkkypeWO+1/kjZbFvi20tO9FuQwJFlZQrZFnLYxzOA1NyGGyljOCTcT
6e4tcnbSpzMms4JYbbjhqlnvRg4+d/lGFLKBXOPWLDCsjXvHDtR8rfYn61qQPKvJcFqxqzb+MrzN
SbqnSqK3C6Rpb8QaHiGgt7zfyo0sn+K6w42cNGSozqZSh9/uyXtXP6dalz7bvjAXqoUm6YpDE9wz
kHWiJfnPGN9DADTXwZt3qVzsNrL78gpfVUzAkQHhws1rdJ66wvDeaWKRyhZRuLfUPTho7SpId44X
9flcjf1VAs3jm/EKBlLOrfbYQQN80S2w2SGOULQSLa1EBDRLV0LHYGOLGCndrPRZOVNIzkFbkIN4
tJmaMe/7yfc6Ga6kej0//51Z2gvJbe4L2r+xBprI9goM5dRVM4pcM2oyWwXTrHM2oERYuyb9tl81
brViv73Ib5Feo5hXslvHagI93PgyCT40D3J79TrDLX8cxmsfwD9V1vvsigSm5AoXm7Rmu9e+r1VQ
OF5uVsOa6plQHeqvtxZkiF0/96CqD4fTX0rjxq6iXNWBYJfQ63ivHGwqDADlglxddVfhZH0PWwtU
S7C82NRYf74VpqeeJqYpNSEzVMHy8NYiHXZfLiVSLthkozqRRUgZKAQ8WaeBEK+XmK5kDXKisTg7
5T3FDI3SXcKUJfvZriQzR/1Lc0oYScQwWZdKnMOKVeqbUco2zc9V1WCCRWE3r8vcvIVXgu5F4H/q
FyC5kN+YncBF1ZTJdhe7iUoBjuYTJkHgREWiH1qpd1MV0YiFVumJOnDLyOpbWP+VinnkxqDLjBXv
FGgTY0Y7bQSzo3bLskLwyjzp+ixHGG8xNCg9QGzu1UJ0nQC1tGlcs7qv+ktEC87cGglI79OQ4PW/
mNK770yM9NeCjCWLElYZ8LfeEbAknhcFjxxmmGibFBX21y12iXIAvKQ4vcDiuCzXv63P0Cw2nrfp
BasHhY5R0pyQLkoP5+J0dvNLFuo3FILCi/il7xrsZr7DLIcy/Y9OIZ28MnVT/kblZDy2W8gDAvAq
t3wzAPeso+rewf8plN57W6aVF+4tvQzFTgGH1c/iPW9B20KQ43VrozTE2WdfbSOWG4M+SbPM3b5v
9ZIgPXoKAm5fey6lC+aHHSK0PWr+C9w+zGBg/8oZBweZbwnRW7QllFDjdNMNn8xX3y3BumvjyJ1c
3M8z/DanJAnF8HjWvidxMDvQQUwKpEYUxC6TPvUnqfmSgDsMAW2PtnD/1hNLPEQrENAF0JlRS7md
lOHjNdp3dJiCIQTNFkm83acn0fCllEat5NzaDtuZcbqZ267lU0kO9ACTpBPUcqv6gv4VRCc7NyE5
Lh7ulXPnz8ZDkP5YTD5orKP82IihWmEQR/kKnx+3vIPIRveNF7mluRkoxXIWNB3e1qkc0uZunka/
eePOuPq4ravQeSiTw+r5lIUg4OgRUHA8uyyQ88Fb1fB2U2AyMLq+Nghd7/EOangXssUlQicjpyPB
IbAduIYoD4Pe80FUPkdA53hKKxxtKlFcdakYJ0nydUGy52eroCJRhca4acjBG+GfE6craL9O1Cvg
QNF8RRZxAKYsLoYAKA0pnoNQYkSMOmUPyIl0EgwWfIjDRla79I77W0IXTS3LdizaDgcb5CmQjoqH
dXf1X3emTB/zSeLfFQamCGYQG8GKvjUwKMxhxxxY6xzS7kNrCt/6GlQVi+XVvhWHX12tkeTeApOC
QRZkIvkRg8Kbpd5UGybwUoVh75xVh4SzRSF+gsIhRFbr61r71vB82RjYeAd0ZTJy0ywqinWFu7PT
PP3bOFE6cBJG1Q1AhVxXfCOfTTnE8hga3gYrzsWTSwKxe2WC5Hf/ht1NHPQT8hJ++o0U+gQnCRd2
QGwbWubFs6SBhljj5/uGC2Aw0RzMreFK/Yo4NKp8XfP5wYwZVSVLvvS1FyBgCdXfNYDyaRZkPb6z
NoPHxtZYTgHGEWeWt1sd9QvTENfwvwrvpYEaemVAi4QILshokhPRpeTdUOVS24TWQ5/y8tETzD/G
8yUecWyaa7WUMYlwPvGcr5+JsJfcQ97mYlkbHPXmr/5SiGbWnn1rra54ijlbj8/5URtPEuWXzmQ1
oyiqJVUkDv9hL0w+Yr8BZeOy2qNV+V+tCApipf6TsNVTrAXWrizdb4evsViK1uReEMgb9rG/ANVX
aM+HkbyrU1TG7cWk4Ok2GMb3qwgs3qMVGp0RGql2Wvcla+bQwrXl2w535jM8/niSN2lXvyvyLol6
AxOSfA6870O5pwBxtPwr7Bv4P14+2iTYqZem+AAIm9XOfCHTv+bTZIkpNQ6TaQwZK5pjvYmg9BYV
C/BfL2axpIvu/yJbEMVjFs1omd6500u6A7+pur+UMwMpoXFc6ttkg0syWgT4pOTtXL5vhbE0T9Et
enPHfiK32yhgt81p6QsQHm+TFNbuC6gme0dVYr0YsgEPe7ADIDgr65xJ7vUSxa+seuFdxqyBUVYs
HU7cPohXSc1bG0qTT2nK3/rM+pkxW/rFFJTj2Oc+QphQWfEfEmhfTeOUs9N8GgnOmvXzqYiCk4QV
Kt1fBtRoYaUaJ7TQD0PG/plAJgKsE+H2yNCxm8jvlWQpuBeQ31bBmRx/Y6INcqAdkaHWllYVezzP
ZusovlwOKl7j440ZLgQTC8lRqoH7i72kNJ1HP7SFHQNhN2QubAMIZoXrhTTFfB4+M6w6TNOCc+gV
YP3yH/mX+Z8ILXyTY4qnaLAblyKhedTUjBkVx4NnZj8pzC2k936qaVGRheFohB5qR0g7l+VDaOkM
47Qw2Wv/l/rJQf/SVuSRIo8RZuS+JwFBB1IOIuB3mjxisr4XEJA7ETO/aEP2meX41Zmvjm5hZu+V
L7WYfaLloBtxEplx/6Z9NMZDxGsDkS4NSYxLwr6YXl2mwx9VuKu/RxNMkCb5HfwPBHDGN1zIeoCm
9X0zN0QlnOoG2MOLH+tNF5DtOsYEfwD6jiW7vRdrqPS4UuajNt4K6lxSnJgE23cZM4DsX57pGbls
ccd8fsCHAuSVs7+Q+lb+1negX6qxRGqtduUcwS7NLKL5pJGb/XbBo2cmJXHRQxXjpBySQHqj4QcG
IXv5qnWjR2rgeiL2IutNCD3/2YubYaQt8184s+WRnlfXBQNCAlZnGkC6xmiyGkQ52o2ibWYvrO9F
jaCA4n6d9MbxGD5h24hZOam2L6F9KJPfZfL/lTdPpPaPGlQVsbrEVVMjvLybYscLrELWoodprz4J
61BZdsbUyHRe22tunDdGv7qRnLeqWHyKMhN7fSfeSSow/ypYpRwDzUfEjJbXe9pimt8GGjkKAEA3
LMa4rstPm94DlUVn9Sv/SyirZPhoYk2guH666aYtz92+zPwtP+SumOIJ80IxVkHPybFj0mHBUkKP
0GtN0M1kbfP2ogeuLBNp855HSH1DLqhPbdjsAfRVLGyVZpm/iZN9eybCAg3qyhNV7MtEH1C9TclF
tvkye9hK3LmjAPvaZ9qxYAY3z9uvaAJRnU7z1uPLcc37bVu6qVQCd0ALuGwU4djytmCjCXL2Esdo
+IF/khDsSVeiZhIV0SD21WofrBrM2zB7UZFTQwgNpGeCuMF98DsiGM/yUfDyzZmMnu7koq4nm4Kh
Eem/MTz2goAGdfFZ38dnAj2afJyYzcis2DZVOgcquj/Tz8AzTI8s0T9ipw75g6M29sjcRPZt+/lh
PoiPNXGFZtqz7Z313HE+yoem8u4WmZ3yFdCjOIRHHDbrJHpl2xFxU5kBcJPHZPAPEiTN1eoSYHO7
EQuhbzyAq/eNXLKtVYV2d69P7XhAD4XRw1Lp60n6FsOHiGMQpqLWRGY32yVm/As1ePMVU7jLEXLx
LMSq/4LKNYKwD1J+4SGsv/hGwsa6eSAhY9WOOvlXaaZBYId6PiHFKya9YfKiU7/J/rPDESent1HR
RwigxUpZ+Cx1ZrL44qGNtJilFUr/v990N3UvKciE2S76yJSw9qVI8QNI0HFxSiXH4D2omOJjSN5c
3Ypv/6ftzu0PUJE2+WgSwHV2ccz2Vuqk3MQT7yYDb5h2WlDBxN9nwehfpBToJVPD5Qpepg8KobUe
9hbQXmy8SLg8DbGjQyG9Fyog7JGreO6r58Qw9GXfrLu7Jecp68az83x4UI0RGkAo2/hLV+L6zRn0
HWDuG08iJTo7sg5kWM0/TVUcspQt0v8s+v3OwY6qHB9KaIqDXkOaeABWSI0ie6uBCNePCgsOp62P
Yq9hes7wdn5nYAz4Vq3QtXeAjpu5AC150JIX8k73F0UX6KPhEwfGnH7gZSJlDQ5fPQMGuqRX1y2p
vgwGHbJHWpIfUDJQ2bCilV5p3gYhea9uRh6RONMzujYIEoMgOp6PVOxxZ+X134CFjQMsN/01gouI
tOzH5IqndLnfexg/3T45pUqjuQwDdkeYTPPszjuJASUHK+Qj8dzFO4ZqJ/arln0HtkT6LwMMQcZD
l5MlSY1IDLo4JGpVDki8t3LqE2rjbe1AsNjAAljbhez6+VtVVsb2BK2BnIJnVTZmWZhLy96amZG4
Sb6liJccTPHoKkxITS/7NRU/h23oMZJnq6GX/foOcSQbpTN0BpIz43Ho9bTUlczPEsWc56x1NEyk
wCFnuCkngkV9m62NySJehq4s/jDORqsJ9cI8ukAhrxu18SdL9uoDpknBr5M2/1WXyhFrSrMf/VEF
dCinY4gDIuHq3elK2mA6pio//P3zcAzDdWp1oDvafjmd7H290JAbDDMpJl+HzwyMTgD9N1sjS0/o
nsEql3ucULU/A+mhU1wecwTic3I+3WP7Z1EQpvUnjQCXM9EQATvf7ElTIvhqtqIe0pzdyc+5o7Om
x0kDTOOaq1fHWdeplJjXDYFqv7Ls7glrBJva6i4yNhjUmzv1L2WMWi998ygT4xzR93RfF07OKgBp
F9vrXrzHlkv2kUixjKIT/qrwVJ9KF0v2T7Cp/tYUGseq/HOAj1SET2yr42DKw6Wf2xDKB1OXZqmr
9AqYrzdHyPtMPcOcbVTfNil/NZTJrsaWTS0eH5Fq/uViJ9/NoDN1EKnZCNM/MGFKzkR8yg/3CfOj
KHSVUmJUm1MIEx+YgqZkIR9p28H5nDHybFacEyvO8fHCD3YVFMeAMWC8VvScWO2iUGgxHOja7f05
0pC+AcOD39aZPjBLMkpdy1tZWApZGts8qgDTFrsSsO5qRtvxVBlBDSPuhxSrdNIz2SK6XR0DmCEl
yx39CCCwtctggCjH4hnn/yohzKHYvZcTQpn+y4yCA3CbaM3Gk/n+K0csxSDjTu4nRNXWC/GLEVdg
LhoqDcX+GAreH65eXKiUDiHoPcWD2WhU3yqBnwynKYbmqKGmr/7zSMkW958DnHANdGdrRPW7QvIE
V2I2u5R2/+aW6zE8xGsDN0B/EIktIpjpegJOTzWtV2JQI3FCdmo0iPv/pc8EeKHwDp5I5UJX42Pc
zOlbTstqalw0poS/Boao3PYywKiCnPbE0H0oaosCRvNWgf6mHQBDq1g0ECnB71ZzX78psNOS7Uf1
OPUbpQ6kLv5oOCU1aAHfUFYnhD3X4S8dK4lHPuO1cC7rlHM8gAYRccdbZBLdtTX6KEHxxt1+9GOp
ldlRg+Zn3/MSvODICGMJGLLgRmxRoIX5mFLuGuFZSa66rgE8Sn0Vm/QW6J8Rvwt6fAtVMyhZ1Ac+
jmqfmvaxoa3TcLk8N/agxy/rkeRnmMliuZta/8CZ7HZUtoz1sNHJmcaMW0gIFYAwL4hiHNUnfsZL
sjwP5Dt9xBNd+UkMnNjKwod4wMpz+AnPZ9FbphyUsp4xEWp9GX9k34EpjXoPyJmB08SNQBysZhXd
seM4phSUNz+zHUdl1AR105BrEhDgRT3CQ6l9QnqwwVAzSqWkTQtc83z+R9zcYjRZHsC4wn/qPN8/
wyB7XKKuXzbb8qJbTAO7kc6pLNqpn2QViVK/Mn80ldGN8IPzQFogYf3uQSQQVn73V5ewTSoJ9Sre
eQRql0IO/Q9MTF72zPU1NvhlEcHAe/Lx6k5YhoPP7c6DY2nIRy9vjH12PR1ilEcur3/A+8MP0zb2
pafZ9h7QPo+ua+D6JJDkMkm9iU3dBxZyTqmvGjzyd8BbpyhsmYuvUglLMDifytV74f18wJrJScGK
SwMvuuuAYfKCcpESoI3fMV0GphbnLDTGcQWXtU4DyCtm30MQKSSs0P40i24DJfLy4Hz5lW9O3Ykd
PEgX+WHri6H6TOHnbweeFNb5y/LwqVHtpgGT5H6ZqjUq4D7o6RIUgc2RyzUzuc6jWoOHlFpcGb2P
9oBK7xe44BN/Ph0FDbxlHzTO6IjwjCuSEAwgCVwUA6EL5Qc0y2lI26jRODck5RTfqiFAPrBa0p9c
65a+DYqk4xf20bOi4NoGwtg/F+AAYwNT+Rh1C3C7h0BPO18G+9AGURbv3sYa/T4xEnzzDipX6bOZ
ibzAWM8kB5N1HvEZ4RccMdMT2qs6OosaQ63Y24eLcJ387/sICZ8TiED4SmNqQa06UQfh/qN/CFlt
JSbfYnuFHFEYx28qw4AiZd3Xs46k+Qug/IOrYaji5k7/S75/BoxVLkgOpmjcMd+HKX8RNW/pcdVD
L15ALNBtFWEg/EfFZ7du8CyKzsDjIVVQ5RdHmRmFZ35y+xFFmU7Vj0B/EdmxYGhuSsZ2+D5zBOBC
EUCJsbzHBdLgPThi9wkqHtzwoqqvETMMrg80rDLf8FR63hVhI1PumQ+DPne0u6nCV8UUKI1vSY11
t5UOs/vBrZ5+gKe1eXbv/rr4+kRyWrb774Ey4w5xNB6yqXH2LK7bsdpHgmqozK8JAvZZoi1e31Ro
XOfEmpeotpUCAuzyZM7n1KiuEwgkL096WNs5/5fG0lv7gp91iVU+qideuGyEOD6az87jani18GoP
7gTMaSIGwFC8900iC0lwAJq25Z72hCatOA8tvInWsOVmTaYTN84MiUXYcpfMj9b7Tb85KA2kQdHk
fvnnt9tOAZn1tMK4s+SFrlthh2pvC5ARj5LRDzJIeVTsl5roJHZOlh17JKL+BD7qxASoo9jv41bf
zE/OWh1enzwI7Yi1q6Vqfir1lJCcOPVbMLv+hq2JQeZCj8nPwjL3oQVkdvnj8QjnZnwPWjY4umA4
/1BhQel3v1o8+BQI4jf1HYoTVa/cqTMfNb/b8/O0jzshoHuvxmVvcttAWfdXUO4vddQMB7NRQSQD
2smkls3/CvnFioQ+BxHlKEVFnaeCtxNtWc8WW/zftNfh4hJFplEyx1Iy5ccodO/eaOI+2ijTbxhR
osHNerdLI8XIK7nB+i2dKOBhC94+JY/qnaxjjzUj+1vB4mLHk0HEnPFSKbRW2bHA/6SUNPpbmzKl
YMtxvbCJdx75+UnwEJoahMjJ75TQcUUvJUODsNoNgMscB/TgHmo6Lg24cbgCK76+NjZhdEJrDpU5
c3E7Q9UxtwCPNpfnbyfDXhvXxS2IGPELK0wohINaY+A/K2VecHjh7axotNbLXdhoDrm595XINXP5
R97RMk3Apmb5++lS+d/GLuGsSKJPZquwk9vBJvwsc61TCNx9IYc+HsZY1gyn1CFoRTG8iMy6Gn9p
EgUvT9ocvd9LP9n/F/LHnblYbxuJNwqjk89HGMv/DFvanTLWAqzkrjJU2sSmZDeUOqe4pACzAAOB
LR9vsAizyIwrOgHAF0WgOsbQ65PL8G3njDriZck+LkmSmKV2H1U7TCT/Dbhv8trtMXod+x09lIQR
WcwugaLVwLNsphrdDpuELAfb//OiRRYT02cIAtYkFrBBUbQLpP1rYuQNR+kyg5BGWjt23PeQWXF6
rHSnFHeDxvKJyf0rLFJq8jdtilf/z0nXHvf90OJTbM7QnoB38ENiD93YBRqjdpbp9fWykICeSerf
4EAhcMIAkoRqPxWvIdRtIIbCnFBo10zexBkxpR/UixbM54Z0ycAIw/KwFQ9dtbbkEUgWg0mn9L2/
qujlhtKh+MZkt9POHgu/6LfINjahpweI78mSsn+gURQoOsG4NyOEYA9MBpMTb7AyrCxxuL3mggsT
w7MZPs8NJf4q8QXzOYFsDgLWqqkTeRJU5B7Wx4BjY66iKYQga9RR17YsDhveJiPwyx9bX6e30qq+
Fx3gS/41Dos9u4UoTAIdL3AoT2DM1dpTn5gZ1x57hlrgxtMBS6grb988YZgbdTVnX+J97YQqXayn
Nyu0iGB1+qKCKmlHwqN19RYneQyon+0C6+2HTD3l3VUj4/XP0mimhXqNpPagEQIc0x5y6sBMxgyN
hC8lN4JkRtX3c/Rj/X7oy3OfDfRjmLxJjXLa13uWnps55ixxNNazws3qIGRQGZuA/nm98S26wMQz
RubvsodTSavvIosAX5g+bUJ3ryehO5nc/t0ZhNrB2r+8SDzT7gQN3oX36dMnkmiff8Ik0UZqK+SF
XqZo9B4pjJxcmxTwMJtisS21GjH0fYsDk7CJmk6ttNTaoDvVDM7taRmXSW+Wq4ej9I4L1hclA31B
poBYtWLboy+hRPi408prFLUwMj7y++NCtat76JhXTFAMKTHv949PAn6HeRVTHA4pAQtpNXTt0Yiy
eXL4H9Wxoi8SrF5W6NCigmzYSWJD8Yl0n30ZE1uuXCuNoChiyabeq4jsw4sqAtCVJ3XFN1FF2xo0
3BdVKHZe2yC5dMBWp7EbRGfU+tUfJLWfZa/8PbX9kd62s20PhLHd3/+sR9/TbMcD6WFdgEfcVUjX
ocbT2IanS+gY9x9g9pdA5yBt6e4kvMGenZE4mgBE7bv63nBSvIGtZ+jC1vtWTPQGu66CvCoW7OCN
m0tMCgN4P9lVWWIqAg7ZsmsF5NMSWnoc+8cAe8UseDZikaX/AHubDqeq4BJDgr4jWv59hKqbtpSh
4km0/Hjat5vWLwSUROKn2srPo9aSe1LmDPV+ItnvENn+D+IhgDiQCeb9HWYEAC2m18DNs2EBr/+K
YKHQylUSMeS+IadnKUkcJGssYVz9/v7F1c9PVGFTCkCOA5aSVIECvZM2X2sboAp49HBjs+135h8e
6k2/CjDR0J20TQ4OmSjXNSORBQjpzNQYj8gSIX8EzVOeH/hIaoGgfKwr9BFlqV+3Ig4X6pQ6fXEc
pKcBMFv/esf1UOpWbS8zrgLz3i5odxMbQ0uPw0v1o5GmhQpypj4z4kzxpxxYy1u4ZYplnrfa4qBb
bxTkVZI4r2zOljZVx+g/bf6oB9BNRWKHhWI/SYTiNJ5N/Qincld63y0Oc4I5K8DMCN3vZkr+lPNy
VZPWolERPhF733NpVRcYzHlP+/RFiG3gPedaoI03sX+esnjCMsCVlUV4uM8HY3IpQQgCPkHd5lBV
rELuhHaPWqxpMdUaJLHPrl2qMh6jJlXoMdHej1rxtDGTKTsP14BPCo/mgyaxwjgSZssGa+B88Au8
5Lr8/uhGDv9foB136+yA4rRk7bbPPIp3XRWEntwknxuSEj1yZYzXPgpt8mv3SpEEC9C3ImpTzEwY
/dV14qyE69uW9h4dxaD1CsVtH6B1uEudycIpf1oWBuJWILwZRpzgpVBap0EdaZPoY+hwnS+7Wi0u
HpLTaVZV1uPu3SNHr0CKyWGsHrrQjkf6Q0bj0EyBX6xXvWxFpUQ/qVHM+YqJbf0y/V5+WeXIcTST
S6OrLRbMlxDKFgNcdx9VMOg3XqFzcS9rC/LOe0ohUWLlKMJzpe8cYSWUTRv7rj0ROlUyW/7wxabz
c8jSqRDqtWDGGM8PgaGuhUWrwIrsmKFSqDuM+XE0uAi8o1pCkAA1eTzcxTZMARnKXZfdGqW6W3Ew
76kekQNoPtFd1d+RQVzfJi8hxboWo5bhAhpWJPcewIIDLLS0rWxxy9cgvGx6sVsf/YmXu6XvQGAB
9httKwKuQ6ce67aGfrPxYYxdebakU+akFtEBQjy1bNE0BIKCS0Ehf7BowR7147oJ06YmWJiZkTi5
dK0YPdFhAG+6yJan/lkYMhj3jeEMiqro6BMTjKbm1I0AVLEsPquw20GkJWkhyNY3ybwX7iouMXoa
JOOJ7GV/pCblx6r+2Ddyv95Q1jbVgeedIznmz11G+RXpHRm5LTbUdMDJE6RHtxVVIn6WO20fXP9D
pU6K8Dk/DtXZsNUex7qpAdm4WKTJKcKEJaTOKzr/XaHcJVUuiMUwR7MAGGu1Ve3FqDgONRMP331Z
pHPc1lDIfmF8glVUy9qpXtpxhC4VlQEwu7T2POt2+T+UBZJgzhbN0hiv1WXGxeLkYGv7pnRVPj0d
4eJZ7DOMyIRt5JmlNfvjdGcPifJkBWJ5S4JYN6i8+PEv1FWCtdqnZMnaWHLUsHYn6cOUpxO0bG2F
SGBbXfahcYWV/TspsZPhg9QwtKYKaKnzsr4pmxRTop6aI39ycw81QASS5ktHknTxdXvzoOof8yEu
7A307GKiKGm44KaUCNwZhvuEAWjzRHqTU/Grz4nkRh6gAMs1pAD4fDpimZIMnBnzBSZwl7wGwAlW
voBt1d4fjjB09BI6gTR7djjQRyRgKA3nG3yr0JhLPtYLlDB8k4cuaDefvrT8EViwQmWp8WawvzAg
QMsKfOVbQtyJoFd4AuGZ1eVcv50Cwg4kx9bG8w8faq7Q5loVGieVVnPQW2L+VmruWwY6Q2xJdTa4
muBjxqSLGVYaHi8/Ee37LFhUu4t1XiLsnGkt+ntTl+DnfOsCxlVkkNjZPv+huNseUjjZbHt/DQ5F
DKRbV7g0zPM9hEe47KNt4+AbQlfCWOTzo4z3oLay5AFAT9PKam6LvDTXt7zspX9Mfh9a6Xc3dYfK
EN5BelYkPuKNyYQLY6WCzWZM7fXlkSlk3gh2ysAo1eJcwNSVaxpNnZflaxE+DU6nVBOpiCxl8NDc
zcxnnK/m7HxtbLLNkOUEczIpV68fFYDO/YTU4cMeJU28EXSjab5uEvIuW62DgNzIfSkg9bxnFs0H
ycGE6eEUzZbjPb6RRz4kTAPX1Yu4jEXYmuYacwtoh6jelykLgRD/2H5ZMT3mnQUMIaj48XNmPwi+
qnYdu2me9Wy+YKQVYG7fd3qm4CBcmnd/rW9J4NQyT+L+eZuqEskazGD6xCqBKTWf24xkJ29TDNOm
zrUzLsapz2RFCPIUc1yx7XxgKtlMo/sIYLLvewg60V0WOOG6v/7+YeSnkOi+k9ZZc2IuiDnEJ4zm
2d3wuICQXwae3nFTbiyIS3eCcdrzsH/KyaSDwD9ftWVWkVrnS/dBcwGXeLDAaSy1okpkxd42k/Zz
/KI4+McowJk6TkR6lCw6iLWl9xTWxNwXg/kCBwqbGTk1YEHvPPOZjMFyhJsad6hmSZnm5+m53rIi
6YYeLPKPk5ZnCS/aYvuJCcSPjbUNr06Cm02opk3cutcipEfj8U328KfyMjcRVLgX7d2t+l3BvRyo
MbOplwz7dIrz03SM476L9Lo3A5LatCxWTYutrV+FSyf95KQNwKQu5BXF0vbuq9Q/quhfhfo3eWei
W5z3qH/mY+bpADU0Hta9WT2zLgkJxZprC/OieeZAzxmUYwy2d/rJxj32XIEH8DHFnxOGfMyw+NV+
VOHrxZkSsCVg8FjhY+gVNjc5XoWe1AvCza+OoKxERslDRq+vfZYRnFiIjz+22ZJHOROMqDgi2kYr
jWuluR8o71Sr0NBLoAPdgaA+7ddYrHkWbisCRY/qNhtjeXaaUbX7dE5mbeLOJ8QeXVFemPVzCkqY
6lL1D1fU81JvzMH+ZxpV9A2MVSVZMnIHdqqwWXMuLrCiZzg/KkbIOWnzG6TjxDlzL1Oxaqic9efg
G+hMd8l2XeZEGiD3FWCVoQaDAq34XRi/l5ud7JRGP9vOjXqws4vPm2QyNBdDy+cD/HbNYwbeyxTn
coeLgC/rwlwUIR6dLLnWByg2ENLw9vb5PCW+FCbSN3vmqMYoF7RfCB03c+43VkBJNDX/H6NygPoN
Wu9+SVLtFethZNakyMVbj8VXvq5hmIhnrdR02mBv2LS0ljnmA19Lq38eAg51PZfn+c+hhZU8jaLf
8q3VfnVCVG2mlvrjUSJfhz6fZgn7JE2ncCyjlg8gSYYybtYgOW93fSo0Ig+Jdat7I1r9I58cVc+E
b5dSiOFfVPw1+j+AKHaygQ/1xpWcAexmrF9wG4yjwQcxel1LE+rbtEakyqIWcTSzoL/L40Tw5J47
yV2AjeWIKxIIq/1DfG9Gyq40eJ34ia5jFRDmyufdgIWJtjL95DON9NYaqjOFcx+SO4CKOdzYRmSN
IVEBqlkEtaMulI9RgcWYQfwBNiwIGku9tBn6bjAYduoVX/OhVJa3foR1Ef5mrXlm4wMEtv/gQvjh
AI7ccSuPf9FY2lXnzavj2HhBi1CSCVe0DhZhByoSznjknElrlRjWBoH9pvXl35awyT/uP7AqBtf4
EmL1od83tdyFH+qZkG0sv8aZ1NKrPyGQUzfvprHnBnmwHCEGODoit/tlHh2m6+agkbdB2Oj/SyUo
zo9LbnsiTHRznderCqu8g31qlhwQzdmoc/Y+F6kBlwX0XUyZrfnlX/ebNtcqwMz9Z6L9ZbiY1RD+
XHoCQY4q9At0lZinMRmVlPccCdXmbU5L73cbj6J9UmsrZ+D2Si+anNrXdnrkUBbPxJGD/Kr6urBz
gv8lSj+ALi+etHaCdARk2ZKAsTqd+Gnbadj5sOToClJCA+wdwy12omgbd2ldeOO4+gPqu9NTG622
j/EnnkhBgRJeeU7GRhglvEesfQf0iHIf+rM7bV58CoEVuTk9IyIamZT4drwKmzZXJCZTrIjiEEbT
9umxE0ncgxyoSRW+J+WE5OtRyTK1gqFsli3RyFvpz6mHAB2ZvcUVKbCjaxHC7Sq44WiSRdi+SUmT
WZdksh9qprW8hx/JkOhBDEj+hOMpVYD5iZuOT5XCUu7zYVgYnAl4TrEjjzHo001QV6DPIIQJd1Zj
km+Y9ljpWUqxW284+julnN3/pUpXfblqUL6Ky3dKZ2u2kXPRl2eAiSwe/ykYMNzPZlp44VAy/Daw
zHSTJmO0ozZN6d/37S+BoU+bOZA0wJcVwx5T6fkBHJPT9ltAwaK/Ld767gxI0WfcTD2OzND421qs
c054RngG1vIHpEQ7y7i7/p50z4oUf+KpZLLEVu5OJAVBLsi+o/KC5EaWMvfzvj4z+BDXjsPAEtdN
8tgrM2t3v0UVT0I5+FQTwMNYweCqSMIxg8uJxHOKtKjl/7LplXwx2z7F/JdoblJLnqU5eZHpSFEB
yX6XsKYpRwSvAhOVGoGibJX5OBw/CpujCmdr3SB6AmuzXq4xlTwNb5qkmh5Mmw7LaF1ZbuMc8Wm6
a7GtAKmPrWLzfEw/6rFXnx4R9VI+z7hQpcO2XpEyJjtACrBuWY6kYVeGR7sX+S9wOV4bVhPESKN5
299DtPNLOAI9FbzO+xmbcvihf7sR95kXg9aH7Flei3Ux8ImlZ7eJVvP5I5+n+LgFL6x5tHEMq1qB
6mgzZvvYsXnEsPMWLtzNem4GG2s9s5obqmUNsrz5TTBtaFYRlgmomyP8Qups5FXQmCnJkISuSDYR
dQhKTtLwS2j0phGafcz+0ZyS7afAaOSB0DRx9gSLmtHIif8/Ib5/lUYB4I47Ld2qQxX9SJng7j2f
fXwI2u3o7NFLI4ttUCU1Y7eDnD1LRhtkq0X2557Ln280y5yTvZN3V/h0QeJPVhKR6THQNTRRWUEV
q6twdUmgy8pS26Al2dKcqyWQFlepLRe32lE2G0M43/TZJo/+26rquYr0XeFmIl1dRBRGdh/p+yR2
hwJ03SAFdnG2N6yj0WwGz711/xazkddLOpCOrJj7mdgfj1WgGkRyJu45D2rOD629kbRw7x1c7xSS
DKzHOtAhLUGlrtmBeNyFCnv561NhbD5ENFlOSQFk5uaBlMB1j/ASmE145G8Je/HHwnt50k42aIMX
LOya5ALOlR9TLtVVK8bUC6F6Z1/rabYGSX+2xRUC0BBiQNRO/FQIjhOKOFK3k/USjp1LQrldHB1t
D3zvICxnJeOLjtnE6GHqyvlWIRuibmsF/PKaF9yj9CIwUPdWoNGXpIUPsZe2R9Hx0GleRCBdpdRT
6x+VhHTHnrr+qHp/TiDe8UDlYy/ZoeVltWNdsOSa9Os6x3oPCR+/17ukWnZEqA9Q+S9MvmQp7k0V
PtQRZutX8haUYiQWD+0ALRruma2I/bbzdzPYxPxyRhWDXDv1b1TWFT0xlJP9FVL2xvmmiuccvfsO
XuYi5h9hgLAqWnEXIGc0ydPIfXoh1CLGM6ozaziIYYLVrhrCfctwQs/eivDZ+m5uDeSPrXeYluyy
V8X878JCBK/BWEGmK+NLpZ1zUPYpch5vO9qZdJnB9ykEsCmxHtNcY8u/yg99pTYd0dPsYmk0ynbm
kXtNnYOAfMT7wrJVHhmE3w9ThKyfXhgRYOHehzxhWp/2Wc9dYin61f+a7TmQ+LDplUCPC0g+Whcn
SGPlr+/VEotRM+r+BWCg9AKfKQSuw1nWUjAI+VgTwSTv/5+U6hP2tQZqd+MUd5jDkkVAkkSLB2Y5
PZccRFfhxrHwW39+2ntGSBET52ShCWoEWNtXZnNVw9kU9J44qE8iL912z0lvMIgXXyWjYH+RoqbO
TL5pfuCEBCe7Tns5OEzZPeCGUVvcxKyiWnspkKajNlOSw3gGXzYBYwR4rN3T6PCc5CIjpQ+CzlHB
Eo4DqBn6FO3EM8WMCnPrse5Gdc/Yi46vDITBLKkuhcXDjq44Sh2LxW2OkqnDeDC9mL8UbZHVKI7Q
fMeQp7WDPDQYiInjVugCyHkPKYlkvja/wc7E+zvY6+Y6LImlo3xBnLDbu2Dev1RuhmfBJxnLDz/t
3KDkdvx8Uop2q8zcugQT4MEdjNXaM7zkTctZRKSzJuHSsD14tPoq2V4ua/PKGyHkdMsmaDyp2YLW
x+J0nsvaAvP2dCZ8aH11HyT/2zYmtR2yzEUJKn5mgpUkSH16fvzKTMoPuZ7jrQ93N++H/T9zr/XW
ekotJc/HvruHjhyqAo7DjcGi+3vqXBm0ttrJqrmFglfK1ie5usz/bKhZL07xd8pcDaZgqVogT9SS
KRCbb8u1s4/H6EEJrnZctSOQIWwfNYI80yypjWnDNjZ3rq6yLrv909i66ndEHv4/BCM4U4kdUph5
svSB+bILxIjI00TEUzZztUZEcZXW6PawlpVYxVTJO3IEvK+Bb4/z8hTtx6xHVOf6m5F0aH+AJJqq
Pp+Fg7f8Mhv5W86NgIVl5RRn54qbBgRbrjfzXuvHxyooQYDPLEbdBxOQkc0yahX3xIOLCo++NFjD
hnXZgkWEpccSD9ZA77aW8dUZApIkr5veQlbXuyzGDO5NWmQm8d65lTB+SyPX0inYLVDCfIe1S1JB
NcIV43D9gIrZIsVSlOE5byiYP3RlYmmsgdAVVnwpn6h3qQIe3SYLcNTEYc+G4zmDSPUQHviVXYdA
Je26NcAD+Vk0iqUN6E7vUfvyzhULH3hIA0Js7rx+IRYpN1nmKj4w/nh5RaTsluZeKyFaSpJstnZi
9KNgTue0OVJzSqhyfp4IwDZZuPbh8VU16pQicIyoY0NgM1O7VCI5ApAXc2ZzfyzCqhKdUtpCsqdz
s3odGVmaHx2JR50rBS+02cR2czD0Q+eH9gU2+qYE2eiAEgIPsfH+2N5wx/mwuGNPn3ic2VWd6MVe
t1LjqtH0MCom03ceXqh6NBVefsTHTimHlak2q409K07oTcP+YRho690fI6zxgycPt3jHNITBufqy
lsXFtVd6T9nCpoJcJGr3Kwluk4YADe1WBpZANvlOymfsOqFfayiW36cqO8i5H6ILMomf294LixVc
uYQiaACZWuVu5o8RcNSyczKfMjeDrq9Eka7ovIatP34w/uwkwsmfDBkr27lqzCSN2sadls90v+Vu
SDbn++W974Rqk9/xSV/NDcnvuvK7VeitBWBUOYGLHv/ORTN+k/1jmtJ2JWHn2CZsV28pGbtshXSl
Rkn54mVN0bSsXOIihy4pmA8rTqFqB9zXrgOMJI9SuxKTBLk4+BlcQm7RG2z/kgTYgtlQ3FsKznv4
w7g7lxFtsg4xLM0bqibzMZc+5JkizIOypy1/dU5ODAfPDBrSr5fU9yCwsBgdEEA3+jbrWHkLcqXI
N0m/b5hypPOrzmBn0p6jF32DijKVuMt7leMCNShSqtiL+SAk96JBWRH2PRo+3nSTf8nC3alhGdYy
h+pcTa6Dp8v3irV3dvmWaRZqQw6gNJ1PhyIA9GNa3A4OXk5ajoA1un0NbtDZYojhxRoH2zeQNsYu
WZRAolSkkkoo4OCG+WYbyOopNn4hLphvmPwRNkLpmeY9jhuDfcwyxozgyhKQ9K1lHIYa+a5l+4kp
lErldR2LnHZ1rybPHjEBHTBHBwRqUP7x+JVEtwYE3ObiPrijRRh5xnoke/xOZb49SZzCZo8YSnp5
dyi38ls6M9ZZZhJmQOkjbboknj6I/PiOOzMn8x90PypSuwKx1Aw4QfQMGcf8O5OL2tSQIZX6/mw8
CVu3k6vsUy4ZOcyRqVia8yI2Ifrz+cw2dIxKBnB+wCp6/RLX93j+dWe/YYEimJas8SExZ5qxEooT
vQU6rNK4FdpDqqJjBGHNSNqyGTRtTaO678FDt//zgt2yCGZJlqpdC6V3vKqMNNzpTd18I17wuO19
7kapDrte/nse6SihbK/5Lg6WTyH3jSspyda3ICGvE78uJqIet30wO6Cdg45hyFwr/AqkbaxNjnGE
jF+/2GkkQPzUbmHSmthGZK1YQendZzvHC/iMIrq3COwV/2PG55SNiCcqtst4FM10mjMyqtWkPvFK
ANXGbvH4C4N1MFCl6L2epK3w6MsbKloyyecuMLjn8DSOZy8Rf34YWnhfG92dd2iACziVrjawuPCi
Mve3oPSf+V7TBSwm9MB2xF8Xc0LFtWvi8X4WbgBOP/CxNGa7+0GIAN3c+T8z/IkMpdka5/OSaQJw
9H39FznoKRaw5nGX56wW4u292RYe1+TKq8eIGgizBCqf1bGQPcEf4QSc6We7op7Nrg6diIso25bI
4TwYIUKvzW1dsx7f6hr1tweLzX/A3Ekk60wF5les3cJIZ9XIV3LD+pdCUSyxIfwLN7KiXYqKDH67
RhrKHRh+rxk0cXbMCOBgSKN2oUyYVUpSEiH7btoNrlICRnAP0BPufdcDT3yG7hbfLg4eGceHeeDG
MspzW3bI3EePQZ5BcOMHjWDwbgPG8ah4SfjK1kVL3FbeEX9iJiymwM1q/um1FmcqGZ4ffDKs1dle
QR5xw2fbqXzVxSDG1f1TVbgvljdiQGhIABCtz9hFyh+Fvcmv00MrdimwsRQCuXeYvdoTpR/ZVoju
yu/icqZzQY3gH8UMRTuQT/ynyE/bCnBFAIBax+BeKnAS5KWJ/WS85OlBqyGsP3OB0ylmp51tkKcG
uqd5O2kDjEVV4hwRnH1/lhom0G4Dt3lMgU+gh6RUmV/ZoQLW01YFNCXR+OAO6q+BUWNpUotnBNxP
JmxgtTt2/W3nTM6GGlqXGATn6EQg9ohQT9+Ke1wocABiW2vI5nsLczmHPibB0nbGxUt4eqV0D6wM
+778D4EV/0MAq7uKEJeDLI+qaU5fgLyOzPrFw7MxIb1MoAbNHcATQ4ZIa1Wmx9hO76RNsi18tyh7
9ytZFHPzlee8T4nUYPYUw5ZaGcWxQ91CFYPxG6RSdOvIHgoP+Zo7/+6IPjtdsKIXPbwL5gF/1gXj
rBAy4n0z3cFYKAfbxLbq3zprDLGV0Se4EXyGS0P8os7wW7LdTWWSPnK5MK64VhcJAHkpqDC8FcK5
klSQyWAC0itPPHCgdBW+p28B80LiyhRpq0DtwVBJnn/1a3LWr5Brkk7H5NWavtVAfjjprEjOjIuw
yeiUODpCmjzAk/sKQ/JxF7wh4+0L/ULXh+4LamPFMMaOMDWFmsK6w7EtaF0RtkWilRqBkt7hezUi
ex7i1RLik5156V6g51lvpE+zHtf7o17v2Tmq1vM5Oo8MACXFBXNTnCkUjmrwFtUZIWWOLu9lrm9Q
f0qMw40nQ2afjYiJIt/O2S2F3oUTRp9imYuQ0bBJxeiTiCDdYjyoBKLmKJJ4H6ethcqI2qsDU40L
OTHCEYLXRowaJOwMDG6nwkuxSKg0zSewY2RAQCvc0IYMkitUMhypvqvHgeNApFe8vc51UFCE7khK
zi3wEUAPXq4TKsbH8pwHpcAJC0ukTVmynO3fjdky/6Fpa+O9WQuHGd1Agr854MayA8bYsMuosR4a
7ZSTdarwsUckkEmVwOEJy6jEe/gHW97be8Yw2NCv98asE9LHPtHOX5YaLZ6bPdWP2b/Hzca16fSw
lXYvRfaCFkUFcv0aA8pVwZ3mDYeyzJ2yLU1xwMiEo5Y+w88N25LigaRN2ifeyRoMKYJOaLlt74a6
ycj12HyhT9Yp1Z2Yp9IlJd2j3GaqtfrHGJxzjqMmkLKtY7GuorG6KDsOMz5XjTqnUeI3J7serFBM
dd/HfQ73jVNI2uP14s5TY7G8mjb2d7PSR522/pZwT6Hvg3a6eQ7kSumlLqarXAci00xLZsNKa6ZW
VSlGviFpK0DaP8OuGM3k7qOHNkvDg1ywtAdGqCAVyAiViAKojnDCc9fhnw+PdeK8+ueT5TqUMA9M
eroeGHcind5YZPDN+p8Us+wh63JyvHI32D5CLAiXTIAFRdcH3wqf+awyDKYNqDr8GpcD14wExx5T
NGnz0KZ+EqIq8J4/xuejDDkpaXI+aNR5SbPhcP6l0Ww/2hW92bh+6JPhKZmflsuJPoflO1QXBggR
WYbd+//V/X8bPEJTKKmrggjyImHGALUN7WPR9wH8d/zrhAXfWo5fgten2nMyq+mBLx7gsrkmle9z
Efz0AYnyUA0s/VZtN5Zr9YHqnPx9aD+YDiV9DVbbspJP1e0w+iM1fe2pe4zbYpud5Cnu4muUpIZa
oJrXlttwruyPNs50v37QBBCdV9nWXWU2BWfGxTQsT/U4BxgLjeHH++muKDdMHaUd5kRjFqYWdT59
Ak17HX2wrQH/gMUtUYG/ESSc94UTsQ5y6n1W2eM1QOQtiRtN0CCJ4lK3cNuwjMqdqaOrzv/KWGHJ
QOMBEs0liK37NbPXW+Tafc5xDwWtUed0GvKEM3G6cCBAJtdr7wLNuUYh/yP39pTvvN40t0Sm/rbx
FpQkDvA+HPephV3utK7QmDhaWwhNRjEesDM1ovdc6YqLHlH3KheSn+TTZvuHntaKHRWdfIdF7CTg
eeEldrAqX14UmNeolmSegAVoOeUWueONFdw1dU5tzQt2SpD+ovg2KGw0hzcV0ThX1qCdX69BlBW6
URmiMOz/ZE+DuY9mwD8Pe846v8qEMlG3twOnQ+e9VdkdoBAwfWU0ygehOe1wywMrSpK5eg23Vi1C
G/s5UHn3UfLZ5ZEg7n4A+FI0PD4Kt+wPxHx/rztyjUDsGzf7VoNcuZbNeEfxUM/5u8/8/2r7iBbu
EkI/VatvOSi1OFm1v0LHuZ60a7mosK4/rZiyhmwji/PXcHnIncEj/iv2DPokWClc+0yYzc1JR9EJ
ahrVLFNSwHasAQHr9D+Y3nizkJ/rfU+98DturSG0XT5UquOxnzFxevtJKZtBUYrxMKL+lKg5YGg8
rml3arUyD40Woo9bqFTThno5obLeXjHtIE/BVeL8U5GUgDqhdTErWCX8nMTLBMU5ZnzhOzA4DQE9
mbsVutRxbVeqEFvV8X1qXDSEYr6dwLntorxBmJ+eApZSQyDUVYmvQAHHrJrVqTQv5xh8zBMhwW0S
q0GdaMNuCJ0PAUFLQQXnM5XOz85+E0Az+Fho8+sT2yYOFmCHJaUVTGLq2XDj/f3w4US2nefnpFHM
ycSyjRmZ21VfKmFtup3Z5MfQ/4QRvv/WnvB0tg6+M/4WZqcgYnHjVc9yT3qjVlNtqAoYW4IFp9hU
PkAhVJoZcAqNv+FUkAv2U0RqTTk+S6QmJGaX+UhQBkpb6UhxS6mYrG6JgXI3kKjYj3rbR3Fexpbs
IvcE0Ho46SFTOVUKYyRIJulqmJV72HX04IDt334fKBI3CeQyOMyyfGcoZBD4keFQqWUHrokEdLCN
6Tr4xdFsoQSWcQi6yRaMyzbFYvoErPgac+52M8T7UvqurJrEtj04ml9J1Hfxp1HGGtMc3qzksGlZ
3D2MFSeVgbjlcdzf1Q4lNXXTPdJQR5h2hyNGEiNsoqccb/xESrfYswVf2Vf1641pLq3QH9IWmu5E
IqKrFkr1qG5YjwUH1dh0tEO/4sKNgjIKKU3bOrR2Qxw+SserdvbomdNnWocRrGnF/jvf84EGHKE7
z5Za8Se+k4RrP1ebwnzGT2vIoVx3QV2RAerQtCswsgO+a4Pt/ETudZqLmnfZxVuVtfWL/knz7Hix
b8RHxoyqpk1/f4aNyskua6gFbG22IILTO0d3l5Om7blFDW5uPG8B/hro5+PC71/ru1hzcI3cHjgh
WVFuv/8706B6aN1Tre3DJG7YweeZuGhs7wDmd8MUcbV3zdV1thZyy4z8y7KGLBxXAvbj25l77JMP
zut7T2ElfxwPJH+xvfuqVHc/WGx56tmgxic/mq1HotlejnFKc//qbhmNG89gJbXb/17cAm4Vryyw
SMjApNYv8oQvGotPIPFZ8js75bb+YPGl162TRbNox21x3aQXJfP2fEDFpCkfwYRwzd7tGFLKZeAo
XjMghegTRie5OxFxWbyVsYVYmflXiZod+oLrcqdlzWVdGZtPOI9ij51Q1rcb76EBFx0DxQ9BAZR9
KMymBn15CvIMMhRHHk6KcJ+xZ2WteEnI2q1vVrmYgDwizgfF9Q9fASTEEqWjz2i8BafPPuv4F437
Qa7U37tcj/GqmddAzuvcfEkejSNu17XHxzNxIjFnunWvuh2o4+qXzqF1HIRHMod5xqD+qQwBgOFM
v5rtfcbzI+5ydEL7S6AaSV4A3I+fD/dyUO0QJjdkJIzqTIr9omT6wcyoVqQshlVP99o9CM8jlC8u
u14GFRRR/2yU8N6LPA60zboiZxzPOLBQ+yuHUdI6GrXoi4WKZuiB7pyxvVSX98Loe0Mo52u1UW0+
0tPnbLPhTF/0XrV+fVK4TQ4N1rOD5sT5NReP3csLrZulJBwOd8/jT1c81mFIEwowXWt2BJnoU19v
kjmQFWThHQFG0inTcOrxhgEOinsmoR3KzjGcWdvfs2SqSr5eALDhehMYiA/K+4ZDzdUFOwe8ABK3
4VD3TWMzD4CR5iox4b8bcMs4CScR3xAbA281em/0TYo9+9Q8CwBWSnHMNuRlZmKT/cAY3q0xeV7a
IqsU5GkfCNq8xfbRawFwNYt1O1wJ4ORkYMu3cQq2znAEYXpIBvCLlgHPtGpW3jlUVUCLpj77u+Rh
vMF10ZURN8v6mDT0aQDQCriDkM+VZZqTW8qKEbMU5NMCjCR8oUSJ7BbXNp7HdO21r7H3f3pQaw+u
vJxC2cxH/fAVok0ISf/wdqjAU61be1MDFo35DGVLi0CA17W2AlAtGOQpz6YOrp8uAaghPFfzzGbk
unSpmzfhY5end+nfu+35LcD8XgbXAL4r1Alu/Y+YK3BvK3buQQNXaNoGKh8rURoHDH7QZaCLUx/z
Q0znN66ksgegXnEj0O9MFRT8wBFIPHEk4jjPj34jZdQUz+Glly9FFgx8gUhuoLwcIC43NXVJ3puC
EhB2bJ2sBn0i8yTpNY8kIgcmAPJTTHJHB8oijpEVd9lFdc1oCRI/DsQtdMgtDK0RlV3pct3X5IPH
pce8eLmOUyVm6MoNfq1qg+B4f2Iz0ghXQUl2p6WRnSjHzJRYSr1r9DpzNtjE4pzxBgKP6kG5EnLi
kbYYu/wGrbVKQYj2zoM0sw+7eUyHWDIinfaKhDBwsx7o4FEAR+rRsSBp3ALFEEo5UNoEIsQtAG2y
AiBst/CdT7sa3Q1BdI7OT/mch5R1K7rtdcDP9E+reX0DUxYu7RDLYwHiGAGb+wu8xHqAVIQ0Vx6G
tyCtk8BBKjdwTRGj04N174RQCL4a+OZrI3c8wo9mNWvr8uvC/YQ/xXoKr+nSAepxTQxXbjbINAJV
QiN1pvv2biYafTXBGnRM6ZsApf9tHn8WCY46JSEn9ASZb3w27GSgiNhjB94AwE1PJMJIwxRrtOhU
VDk1kEhJtXeFfeYIDFPe2p19QW7MCEizD814X9wyf9htj9h4W5mKk11qEBMhSaujEI0hNTvpfl/Y
CKoRxDtur7VO6HCs7oNjc3S3rgoemRAhuDd/4dtSFYbadsc/HXIhumxU3Y+xaEgsHoPvt7dLiLK2
PIkI2seAzJX4Z7kAZqe+G8yYQd9+f0/K1jogolHI089F/My4ls/hb89tWiHBD9hatrmTM57B5OaY
ZMVNDOLfeBGMVHDwxwJseZiQ2jN5h+GmzLCIb3i+4IuB89csFvt7rDlRC3cDEt6JcEflqdVxS06W
QNGzjx3w/AMxVNPbGSgYiCEDBgjrWPfjJr76OgzVXLwlq6LVRC94yydjGePXPiP3XS5Rn2dVm5rc
JX61LNjJS34vx4fMUMXM7+QkpjULNWkhsVI1qBpXBa7Rr0fnz3EnyLNAIM76EgyA5wfAXA4zUWM8
W7cW2ksL61bg+K5rsdJ6bz/5uT3VohQNzw9dmUaX22wIkgJTKHQdah/yFMJsJ+36RiyLIusrSMeR
t/VUmxztRJapKLuUh4a4w4ZmbthpbhRz/WsNK8BisuT3/bebE7F9mWpthB+NI2uwng0dY7SYmk08
eygB/oBiwRw+iBk7EHvJC0LdiDjIYessDgNGJ5163W2td48l8civItZXZEsH7sXwQxe6XnejGK6J
BjbaCpsNezIl8yyvo3CV8/W/EgysxzSdg6mtMYb1CGq/oCKTQ4U9dl+cVlgwrHXEUktbYC1y/2xj
hRN+fW68IIBocdXlOSOeYWC7Rm7LNVxjSpqQD6vePJczpUYB+FeYNhhrkhpsjWi1xfglqlyppX5Y
Y8DqvSl7VyLwfF/CnrwKyioCOm8oms/le3oisXGm5+/pSTfjuqRu3dKTTRlR62bFQwK9nbY5JtoT
413SiEM9XZwaYBZ7Z7b/Kbypgs8fzoVjikjuWDbvosmWrLpr8wgfIQ5JT/qx6rvcIG4Xz9joirTd
PSfBvWBsIM8X3PEMCXNPCowbpwfd5Svvg3X+EyG2LwS1kMNpBME986S2qXnozURBveWwIhMVIfXL
s+KjYcSc3hCx0F4xK7FJ0iQCLu8vKAy3/YqPxyBa18YBrGFPM/YANW26JBpHEjhupoof9oRSGqJf
O4B8jGEgYMCtM61rSuvfsYpjpyyRQ8UMjDtCTNQvablZbWfazFWu4Bdd6B79Mnv8cOKmmuUlEZFd
UuUTVWHs7vhfSn4dxlkdZA+SFVY50SW5EA0qhtpVF2lG7zGLhBytBfZL12XDUkoqECYPN3SZRZML
zjq6SxHafTmBS/m9/AySXci3EQhWwJD1fVmMF2yNId0357gf5fiTxwIkA/K4NIJTW5CDOhPJZIlM
JCvL15wMveHNthkkwtw7Th6LLabIx9yckltvpmZQAUc9jvioY7A0HKXNn7YbjbDiFpyAsF89I5UO
0cb3H+gy8EOoe6bdkGiMQbvUkarp6sCPFLTwYtsun19vIvi3RpeejcrfeUXarblPsviM43w9bb5I
kPSh4bYCZID0NGbtU3xKpujLn0AoRQC2J44d7YwsMiz5tBQanVa3r7vVmNJMGrV6hMQ/AVYe11F4
eMIjhiPpcbcOaeakLbIdSItuQYqaFiXGHYP3JC/FaXrQ7ANL4/1ZzyiAk9Ds/tfM6+IZvkOiMGc/
3fFJfwrh+fCgFHXreKlef963GQ79eh1q4vafeotLQ0QW4tE/oFq6K2CPl3twWrgLwND1r8hMmpmf
WDh6H9PeFtMeo2+ZStqr0lW2/RS2v3nGdaUXGB92d7Z8uT6mt4n3kHC4Tk5i/pR1zzo9sQvEkteY
LehoMJiouGFP5MDdyQ3CQdY2sJ9nwJfjXBSjaPz1suFQ2nT0/rKahuTja+lUuMObPgEHdYSt08SI
pHclhLvw3rogUqQGecY5VYM8kyJHOA+aZ6GKyfJQfgm0VNxOcn1M3BCgsmrzXdv7CrqSKtKNgch2
Wgy84VLQQZUrDkVpxjSsTvUECk4ls1L+Wmj/0JbwDtCsDNbdnZBI+yqLOyGP912h4TXxl+Nqc0sR
yra2mUODHkp5VuumdoWiYigpbv7ZSyL5xDnPDcCVJEHDfvbW1emQZQ/49BNDbtu1DyKGcBsntbX4
tKbJ2cWqKLu3Rx9QnKamVOamUpZQKJEM4DGnp6F4dg8MHa3NAx7HqNx3hQyXwSGbpMi+ZZWZ4NGw
Mk8rdU6kHV9LJTrNKON4tqRn6vg16bfIjEgsVsHDF3oFkMsNBsX/aA350T64VBEpjfiQmRiVG923
NlRjfOXECwFUPEGdAsCr/bIq5vXFvZ6zceM/SjeatBlY2BeZ370WFFz7Pn+FJZEuCerQ2abLSfBq
DiwPs5gCQPN2zKEGiHDSbGPEgmhMRSORA3WFstIWjHBBkjCpL0GkYbBpcnSlfPE6TEMJQUuARrYi
MUPl0GoOcP2ee8NuSsQuyuFNjxDqySSDjiQwV01vF0DR9REaYmJ2axKidwVvf9cfKMKK8hVn81RD
FMIVrw4jr6UMsQUK4C9jni6uueRttTFtkBONVwxRZgNBpxX5rGxistuDKauuFxI0Lhk6eKuhIoQc
QscSSX6A+HsDeMSDm/wLsS1aqk649eSVZqamPDYp/fB/gyPK1s9354r1hsNbOuRdMYz95TAihTKd
eRtewr6iezrbiehZ4gIgO7vUXPs5fdbnaGPahtNTvxfoeGfPzp3MH0rV2v9bYe7PPpwjdGYct5fC
ynXb2JN4y5BNeaGIdWJy3v2MSsFnkEfgMTjN1CRDygAYo01oks0zPYOF5qUcM81JSKOyZ5fZJa/K
qh+bm6tb0DyC+Tq0cRV0hBjHDJucSkbKDVrVQX/mgfGqjvIc+V4wyVlc2Sc2WxVBFJePw7C9xxPR
KIZJ1sUtYtLgHWH896EQY+U0LKZJbnZfJ735mZPFhG1Sl6X03FuMdWn/bJnsEk7B9yuF2gGO0bUw
+Lv40H7BEHF25W5+tgMPqMEHx8cADMddJ1j3IJxvOyLap0DQB0fg80CPtaZlyltf6qAczOn6xbrJ
zpFTqyVfuvJayF8VNhbODvpLcPzufz9sMSe6Q/E/5qxHzgbmGVMLeLPHoFOTNea3oTi5/jwz/McF
eFmd4Twc4+0zP1RpI1pTGcIyWs5kgqe+clhf4uuh5is5wA8QqhG/Jjxg8Pg3X4cwp8fQo+/OkJDL
g5U0tiSgnMWefE3iqfqapcD8AnJ1uvq/yC6476AeWoKPzyRoUnnKzu7mAE23gtMG5a82gOcXgwLO
UbHtRYUPb/FSSEu1kqedtuWSck1egsjHpyV2+vKj71bEWo+8zchD1WFckXQfNE/XxJrcS7HJvr4c
iWQunif5yq33qioL70qTPDQslhChVzvCnxUGHmoSg3AJ4jUZyezNqRi03IbwRR/QI8pa/dOSKwTC
CIuHjwvdyQoose2AMtPnqmH6PcrTgsKzCrv20ntyYdpvOV/tA7SzSH+/eUx9lkKofnni09uE6BZM
M3r8/3nqPUAfrAA6J0pYK2urxvSTAyXABwO09GiAmkilXrdyThOhc8+Cy2/7A4jK7eB5unTfWbdI
JJnZKvR9vrC6k2bRR9UEnR4LVVHMn9X1MWWP7p2hcUHKCd5rj6uOCWAk7plydybEZwHFigZvEHG+
1lIArqP/hEnRV1VvaaRTBfEhoh1RMx0z5RlW5RylNdkVm55IE47tkgIxrnZwhjUlSnkDOalGh8BZ
vWEZkwVPTgtA7Nn53FkBhGQQCJeBpGYarX9yxKflsoCOrgP5wHv3oSR2/zqccDWdrPHVYfEkG0iL
CfDsDZNO6LdzG2Lsclxrdd0hPfAGgj0gUvtaFX4tpvlBczJmhnHv7bkRKZJ8ZPKmVBJ5pXpNGvUu
b6ct7hyAVYP4T3krlx7PT5UMwpiSvdpa3KNm02RBV/RMKoY0H7YDveiYo5z83PHMvwzksX319mzH
AfjGfJQwpPHK50Gt6F/qgP8CjTFXwzE3V7BHebaXLUM8kIph7QNP6VpoAIhKG7ICfQpWXuPb3Lto
CrodjWDMU2BQdnQQ6aUdVKrdEFwhawiPEBI4hbdVUtmEER/FxbpA7nxR4T3AIh90Wj5cb5gyxTsU
fiW9vzuqKGNcAfQceyffxtGabthjZdLW3BbHaI3mPoGs37fNwkzVQyIsRlgzkrFFsdYMIemA92CV
cS6HyS9XZYC9jeMgXyGVA/2dSgN8GKDJ7KxLNtLR+BQYKdDGfDvrwaY+1bnx0fX85YAS8S8wZBWe
K6nVC4Dq+mtdi/HGqXPSx8a3whrMMcc8XXydHtKHOOFociChLS3P5QucqcRJv+K7kSXULaIPK7rM
jvh1V88+82L+edPfF650m2cyTfI3HUr2vIgD2ejTEdHIRAiuzWx6DFdg9+w89yDJ8LM7MTZkI8wU
78infr2VcJzryFtMBowI1zhUJiDs8tt1mkEPmVyAe/AYkMUPnddtgrWb6OkJiDggRUE2LnFvRq3M
WHTm7rDgDrVwwKlzUzCD/xTn5mPt1vn4nF9UbDNUP+S/jFQuwmhJuC1wCIVF2y1CZ2fCVRwT2ZR+
cnF4dQ1HK1kJwy7mY5qcTPvqolj519LIuYiKRwKABpmEkc8xyLoPqAzuiFj93YdaVb1NJ//7ZuJd
d1WhdD9gpxBS6AUksiKCwKCpQY5+rEwqf2TsecUqXcL9rOBurpIw2XbDV9i/5GBes2ls9aCFw36S
/9ei/YxVVA74b5tmXeoCJaUV0Ag74+zUyuXi3crerzt2a+UvryBYXqQTFMUk2AdRLS8PHhJ5Uc5A
tv7u9tyTrmyiWQy54CxqZw0JTUb10h/4uB0kDp1HzqLkv2yrgkx9qGWQ0SYPASYfX919R5t6VMzV
L7vx0d5Nt3iAhQx6+al/+j2WsMYlC9AzaV65gY69VS8leXv6EV6LK9XYmq2bxDD8IIO5GNgtsj+5
FJ+wrON4vdNFLpwLK+KxZ2Wa1CNtzhAetv2AjdmTYz/SNlEEoRL0IagSDSt7uBUf4adjZM1fY6UW
x80JFkf/oOLmX68XfB+P8zDT4VVq/a9jhHPaxl7WV/3jGLH/fY3+RJrif/abzOa2fwrQIgkApr4Z
N030LdXMNqm8PneuK7OvcHnAWcYzJMhDgnZkFwS7Nin3BW0ZQWI4UYfa0Km00HviXfeSUZj4gPcl
icqEitDVT9iTwM5hITIKCliLsKUz22L2//RfdcjS4D7mcoxmMMnDsnnOBJ7+9qANJQLm+n16M5P9
kjcMyGJkgIB0TQraZ4LltiKWTwhCXR+mEi+X1K+MTnJFZ4Tkt6CMzSzhoaF9gvdSy/fKf7JTLRdt
F4adWZrTttycHlCfuwrj34HNYospxXapYrVmvvsit/dQtoXjQTgdEB22vrF1xku/p64E0KcG3qM3
FvE6lxy7EmW6YrsovfIG/1T0AWxlNLXcp1o3o86UKl9z2aCq+bMu900afZjfCLC2eznotxi3XlvM
UqS4r+rsNA5CCL8g2fyl7N1RMAR/QWihY+keCp98fyL54qq2krTV+MTgbRjCuN645gGFyCb5+gEI
ZVBRb9bCN1ZmzlnRg/7vAyzj5so3tPskmNnzLPqhsOG02todIMCjPiZIfODHdNFHr/RFfCmVQWDm
6dooxPEmFfhmla7uJkiwL5EHO6GnwXcJrI2n7RvE4glq4qqCCQtiHGiyZ0wcae9rflzWNwuEnwu0
xvvc1z8fUD0eeiXfcfPXWZ9sRlh+foIjQJjgT+QPAUZ3B1YPouKUQd1YCiwbBcbj/1dZKaYP/NyM
coqj5eP59Ghl+56JgR4mx1dQG8+ZlfV1CQimGBx88qLXJhwzfrXYm7c0mTE3ip79GrT4PQecKfqU
I6CZvmMpCuRUsEzjPy7KdA/WWjcestXf3k7gCxJvkRy9LGXSwmAnGds5qpQ4cfkU5K5McKg7Wljr
yBjeN5wAjgzaDdVtITpGRiP5e6fOoRHxonULbd22I0zoEm99WQa+7YdP3Iu+wL29lBCi84AZLdk7
tIXhgL/bCkB209OrqPGwq5V/jTQDYErkQP6GT0oXADGZi++eBiOquZDzv7pHp6mtbHVN9uDs95pU
eNsyxLTfIfQvJRt3GA7f5KOn3/G40kBEqqP4EY8vvshYC1hOeXXtNmMc5wmL8yX0c53Jvt3xcCWp
FSr6gkG5dPGFs0jVyIXq8xVkAkQEjbJ7GrvYv3zWv8T8BpKhB7oGJWojGo6NliU8x28HQbmhgu2t
dqwYd8EV/k8Iqv9O5Kr5PQgLkhRcAqwE2BaC1Cw77LMt+cmnERttoavP2YZ5K97qF64lcNCaqr1/
L+NjNkJCZ79mrCLf17GBup7UAshD7ok3r1ph0Jf5/XmDi1vFDJ+aE0d0cDtcfCgGP9B8o8Y6ZXXe
GUwd4WZ+qnqvJDvEDIrsR2SeutzVTvcTu47C7HeQrDmHNzV/4V2yuR6o3kuxdy1so1ykhXM1LAyu
ph3vI9hG4CHab0pEpv9Nrw19Pb97TA5pc+1ojFUQSY8QPmflAjcbd0XTsLmDhkTrVBCU6R4L5k26
MypQOqZ8Fw4QSL34deBg/aSfihkBulzw46tclop5Oyz+N7Sga2J+jhPNUX7trrZ/6o3YmPws+uJD
MlWSBjwb9ToP6WkKxeIpHZPTTfJ+E45kZpYl6Zomh9pwexswJ5ZldOnc5W/tyFKnHq2nJ+n6orZ0
N+ZAx/cTW3HfqOSWl2fAiVa+jUmHHsAWDFnglA5hxPpeXsOqGFWxIAT+osv5z4Xv3tmLsnsKB+Dw
88IQBBd3syV9lJfg4Kv1EME9BZ6RuEJqNQWDW+k22TpA1UFy/VplNben6MOkqrwtW9yrHUD0tQK2
ywPB44NYME3iFRlJJGen8UjRPbBec81kb75JkSr4cKBVajG3UBivr5KFE3308WN3pye45mBM81eB
MESAO3iqNALM9QHFhQcjDfqiE/jDa6HMJJamdHUMSjhjmwK8fljHOkrFrexvnTDY18QoJBb7ldGR
FliSYvGokmbsseJGZ553pQYODKSzxduZSFofkBc8D0jfgej29WDkwt4XfyGU/5QQ1gmsKWrUKBYv
+WqxsWWKPbCDTp81q1b94UQ+px3MQJcUxyKuq3s68B8+3xfrxdK9QqJaomuwz14BsJe6kplWGJj2
8Aj/laAeUwfSK9SmVEZb7YGHq5zZsUqUH22tjLYlkXeFgJcvQ5uvtxbYWGvYwxlicf83SWp6x4lv
pMVBN57c35eHOHSQnZeuOnbTXGg5X5MbnZimHJ5/qfC0QSFWQwTeJzuycrVQBcxZq/RJOoZ4y+Ij
msS6Oq1Wmb/j+kpqvgDmkbsFxOut0Q4mKZ7U6c0FS1SO8OiRv2DI2vwu3+zD/5nKqY8+eTg8bppN
4KTw0JVOtlGMeNmAddcbc2At4/nUWffmQfClEepZrue6ccRHRUl96IRF6da5bcBMCjJgTBZjB9Xi
GDMP5d8pm2kb7pO9R7puswNJt3KFD3Nq+20gGyundjLNuQ3A0QwSlT/ED82lKHrrOkMmRZjLYJo4
po2dj0YKI9J9KX2r4Ht4r4aiWcyedZ2z7jfOFnOE2vR6NkYXl13kOh1upRKjTXi1KivEBSPlQ3BY
W9KK8E+924k2pfodV8O6xaP+fheRPf6bXDS+ChftzjggZ9eiBtIaHoDfSw0rXXZrUwQk87NO/h+T
Ai2J5egC/1a6UqCMz07Hvz+UpjSZSQYZhrCMSurvFhKpkqF4YEUl1q0ZTv5615Jl0Df7whlaLZY6
UPrvGAE4D18KvyLxQLC+ZqBaz++oK9/P1xYjlWlhEooBStLKnIE3/oVa1X+HsGrNq+XvrQcMckxN
VOny6h6F3w97E+kgvQzIL14tsapzl1CJdod+9CbdeavXNjCGo7g2vHqJuzcEUWXM7t8s95wCWymq
JK3fyTsjcZGOrilM0Sgf3pMmGEqDn8JTeuN/nKCLFgbfE+Y46ilpytEtHY3KdATBSnztfJDwtAUv
0o5MoL6z3srX1BuTj2VRftr/lClg1HD7W4ybppvoa+7/DB9uJhTWNX7Y0QCO3k1ANTty3Lu/3wjE
k0Gad2jEZKkY9ZknF4xJb0uQTYC8ye4i07utQOkuexHa+WyfdvpyEMWv0mcdNSIIfH9kveNAhiMS
W69dwyFqIXJUBwou37/UyDopGHLFB64ZDLfDvGvR+35HqwoWSrXVQeHMzPwtDJ7+ZGsmQ9pf7OzB
kBWDkvmmSv3clygKhehxYbmD7ytCIxhVzhKFyrKNsOfe17ES7weJmm+ljM4XvkiCPpEswhcXaq7+
9Sms8Koe7Hso5A18U4JOOFNDgrrK/rxj1FoJDl2Ld6ANHh009YvscbGqkaKrbATj2K42RescrfvG
w2jKwY150NFabbzkQSQfGIzCvhvMwQslwDGzg475Cw7C1nzR23yOBCX+HeERJW+yy4DokmGD5OUG
JRA+HYedvSrWd1PEiHHg5KpNGQUeaRERmQh+0mj2uFLa8lbpkr+/UN7IKifn/PufcmJO5bRdETq4
PxGJKiZhOlYuWAkoT6Y8G6I+5lSUh3ijeLoprkELa3QgsdCcoG5Trib1S48F+Irb4QhkJLcmVHlR
/VNZ69OhxVl1y1uuuxGkpwqRIGJZnmEf72aW/58HY/fTS2sRAn+PmusSIJu/+kj2fpCTBE9DSzyq
IKG2Vm9HERt/Li8QMuNM6XZyWBYD3PusIx2ixFRjWtqJNUdRrUbslGxi1NvZHETlVHygUoktIBbc
mtaLTFaBHBPHTuK4JR/Jn9pmAYTwXq/TlVMpSlkQX+rD4QE9v6MsdnB//yx4BkcAukzxHihI/liL
1eceeUDkLWToRT413Wv6vbcgytsCpGhzQ+B3WR9luUDVvjSWO0vx13U1eaF4cIUgPfCLLDvviet8
ARpa7WGxeHE04UWyD/8ERTcfyQVI012bmH2tRH/l4NmY0dprm2pzm9IzP2Hqy5eIa/O7ds0auGeV
71hwUNEJtzGr7uh1IJV5XhEk8prW3wYgQzY4jO1F9Oe4yr/t7nAVBRCVFAENYhTM1rz2woGBQwbE
ntR5a8ofaE1rMaCvlTOLdPTijVEyzsRMDCyIU359s4LyGvo3/ef/GVV4cNKY9zXbRVvSSr5UhgPj
gmmPiIuFn/klaDV01+CM7MkGOP6nfS2k74oX53AQViIAaYEd72t9v3hLMDwjIj7wr6IwfKk1ggAH
xV2XLrmyUerKXED2sSmI1jMDYwvzazI1DvVEQM2ItH5xKwaueGT6OLCAXUI3URpnUf99kZ2k2nl8
Z5XWQuFoiK8gu/KzkTLgo1fd/ocnuWXvvOr/TgaGX5kt10Y93zihfR98g6RptZXGjN/sh7iX6S3i
xwhr7ot6++RfdSV5qrGiuOdPkGdck1nTfrLumEuwOafVmK+2fEaS37Pf1YLvBJ+NDf9K3QG6IPJ8
A4oC0xEvrvpRzS6TEi/W1N+fx4t3soq0+i1uAngsaFhOQxRtjQOYJ+hdYJAC5BGEB2LwStWHb/IU
n5fQHfz+sSGiTzjTnS6aqW9nijxHJ3mF8OPsxop/uw7Q29gNsr8VcSljyGd9BKKzJP/NqJV6nOwz
N2X6L/dKCH5S2cg4hjoDAqcttyknXThTON4epHQQHvA5kTKPOpR9rwrDr2NnOsF13aZLiUIyqMJz
QWD7lXLOiPwdAwlKDwwpv3JSRiClXZrYV7qweqXwxnsgdCcMvOUpSVqNdXhxb9n8ecM8c0FucaQt
b5eiDTISHJyj9c/0UPmmaCEA3o6nK6wR/SIjbLbypdw11Yr2TYZWg0btOBAMpR4gO+Iu8+Lx/zu7
Tao3ROfyc6YlkIWPsPRxQP19dg1+TlDD+KTuZMduIIneFW9khT3CJE1Oq6urNL3wQXSVmH61V6nO
s7zxNTJJQsZAX0y0ZQdoNF0dLM9IYbK06NoUt4SCq2cBz7iDG1UvpOO7NZMQueniMY33d1CJOhP2
Aq0vwC2fT6d3UDVSsV7eHrM3zJo6tAFTN+UX9uuJvwyxcd9Ue60ItrHDWQGx6XUpCl8Kv9KTSw95
IMGOSIJXwlMCfIwjRJBuofLq+F7zeddji5QD/sT18+mI49OZpVgTloi6X6jkr3b5ivKJouT1W1B2
1URXRMn7ve7DtylwqkwfICcx0+zsDAY1FyDGeD5zE0XzZGxdlDKJg+ZYjC50l93ascK8so5CL/Zo
Lr1NrPBnCz/lF60ry5NHuIykb/4YjXLR4wVYvRwO9ioEZHRh4HBVMSrhFEiK/vmFxbq23wdPIaSk
+Lv5yXhcTUQBoC5gCfxZMeleCrHOlBo0c17/IELcaEeLLY9NKf/kUOsRBzq3oAv1e1gTVuogUZwp
R8/FDrTMXbns1CfY4c31Hvms1INkrRx5QvoHqlT6aTpDt2WpTLJwGtom/8/fmF5i+ncTBozsHGwW
9/3/Q1kaGwReE0/NnJxvlGVbAx7120G3RlrMIrA30P+36gKPeGBAT1434jek/W2E1SHEKiJyWuBR
glPNc28qITIY5slwpBOl/LerFSzPsSN5DTLD5jXSyQgflbHsbnwwEKeTkAyflD7jVEIyoYf4BfnM
vX8Dm+V617HtJahh5MQKG1etZQCujAvCLKTITkN3uSOBIE+HbPyNs06cr99oniI6tMTcQaZqVaFy
f0WYWhWgimke+lDo71S04CNlzveQngQCvvpOm/7Usm9yfNIDsRauGhqDH6kvJH+Q4Ic5Vg7iNGRa
uCFaHgVgpU6FizBQGallGa4we8kVU+FhAaFHV/l7UAUwratOrZV78D5rCPuR8y6lyGvKHZpaf43x
jEVKbcN1xb7LAZDIO8gk2rRyEP+602vpIz/HrSHg/G9Abnljs8OXikbKuQ8neif0rxyXcwLrNtPf
IvnN+lELHBvsaw/3jYtT5PohXeMtz9xHIl7uTL0jqjYpAc2Y05jR9mpHa3A5FTz242WlfqXliLf4
LqiuWtExPSNr1m7SLw44/EsqYgA9zuwhSsToPwANx5EM5zyUQMFtqvrJqUwBbf8L2fSzw6Q+T7W9
q94+sWI08dgHElf/oGbJpJC60tU5v0A0ybXRuZlkocftBa63lSf+KSKO0Y9RKCRbgKt335myBTlP
ntPD0GUX1bpUdg6H3PLzTM4M55WUthK7HAH79SskorPuBB4xX37nA+exXhyk9WWJWbD2s4IE3y1z
O8SsNqT0wF9/HlKAtnkjWs3G/e9QQvwetHgG9KmxbSJgU8rQVFMVIGH0QmXkCTNvXujEMNAGM/V5
ITiI2PkWRwv6r0rHIeNeRn4Cij134Z6oTfE9AO+LCG3EOtcxHUicddOM221Bh+7meeMkyT5yDJ6B
z7JhEyFaySHZENboS9DBbRBL8ks27fnpWdhg/IJWH1rgmQDCz0bLPwRIsAO/B82VrDsndE9mM+th
VswXoTwcA1Osx5ew9PvXsKzFzPcFsASD73wJvtW90oUHXurBDu0Iens9iwUIIiefd7CuwYCbqBH2
fzp0ODe02g/qp2TQeWEaisixus6JHAUeKGeDzo9h4oDM49f+efn/Q1LsGe7qXqzxXavg2GXXXcmp
9KiC3wghaK6wOcjK9sgjmXr/Hq1Leb6NUubsABqMjpthcl9NIpTUVIM5p4DTFNoaT5smj23hb0Qa
atcEG4FL6EAoM6tZuRO1C5BkcFcn4ZUCLuRRu7K3W3UNTydSyrFVEVVDrbJrahjbll8slM3w4U3b
0Vw1j1orXRz8agOCV/yPbLMH159JG7/MdAa7XxZARwBMp9fQmdR+EG3ELyg9nS8XgYRLskVsujot
KySqogVeF1mL0PFxmhlkPtQF7zzb2nRiUAsijE6uQrN7g4KkuLqCVOCOHZPYHL0OcKwnBru/eiWA
K4sANqYWcreq9AhhYSb/MpN2Z/gSV0XS6etdX3MOD9X+i2PJX3fg/sgTdvCwUlOUhZ/WfKUadcgl
JjdsnO9kk250S3kd2vaeoX3f0FTA/q5cADiXSWHZmB4hRcAvX83DwHBIL+xR7eK2tTnvc8fUoCgk
vdaSPfxZbPycLDYun5x75IlnrklW3A61PzKbE6Ej4ZUs8Q84jb6yUA/8bpeWRIFhRtmI5dW9shih
310tS9zKswererF0hydotKkY170wcvFc8uwMoo7hrdPTv8yJLwpqGf8LVsgMTBd+Wdfa10/cDEnm
JKI2J54oWjuMNhrGpDJaEoMupQOTCvqVoxkCSWey2RBm47da56krKvIl2obmYCfSDTvBTUU3kg0Y
Sj52Tk+CVK3nnAn79Cx6iSNEHaO4CtgWFYayDov235FpEm0smL803WhO1VGEIGHDeoW/YLPATmuN
K4WhGhZyAvvqO9vTB+66oL1hbUmAZhKtzLjp5E1nx6ScGwDBs+EpCByxFZD0s7b5dfKFuVDAFndJ
GHLO+B0nrIZv9IWuUdQ8036a+J6XWwukR1+55ApY0R0pzD5zrAq296vGAZTZBni1ysjlbI7OGn43
QF3o6MBtu3i/NWkTN5CWPa78kYPnYtCG4BsyO9kAImnqeslSR1bLWcC7MWQ8UIemlzrFvMrFCEX5
+ZX7JVhtbJ/Tezo7rwii9egSoLcLAWxghosmM667gVMkQ2OSNBUr/3Zfy2Iel0yByKowyJOsVEEc
gsspuJw9B1hfiNjJmWVB9krJsttc60Gl9TtMl1XjALTCv1lCx7g4gQ3RSaqZ6pNkIMOoogCKWsd6
/kPMYgjZwxflUpUrDDPijgRGYIh1J1jrfT9ctayZn1cEkSPVpSeM9288cXsBsPiIYE72rPyxil3N
6Q8pWR3jWmKilGgEQ8YAHsf2rMNDs69s9jJHUFYOQBI9D2FyIaH/DpTMm5w7EcSAgiNZ84vhnz2T
KjYrfNPutnc34EXKeKnIpPCVAwlnMjKxR9UK2pL5/MqkqQYNUJFpGdpi0lXt1/1M8+3xpPlAvYyt
vy5rUmcHjPsV8ZsvzyoMcdOQoQKRGAHRcJX/5i05iRmt13fpoFN+jMcJz/6g38zo0XI5e0y9P7YN
6eOW0K6Ypc49+QGE1IF2izimaIC+EQQJKLYrZ4uZCjy82MJ9gSd8xaXUSeRlCSqELwIlaa7HHDyV
C1cNCtcaVTpyklmA6AtK7CUEJlFxP+eKCiKZxXDnMVt7kHe9hDsVhmqNThbPy6GtwJVUAKukdT39
9SGlopNp8+tcfTeZAkSDHqaPoKF4DBK1LsVI32Nq89qNS2WaG+HD/V8bROXuONZKBxCg0o0HQYVt
nUeqvSs4arbXZp+/oRZUhq4yypttR6PUipPiKjh1NPXgs8eJc16DEG8BHE1TklzEv9w9u8oI+LzK
2gUZIXSyAItQzGN8K7OMzNyNCj0GcfqiouRXs/jhQsbZCAZHbwiseAE4/19+BF254odL8i1oslKU
fN54pT2V+pSSM14pwedAtclCUtLGxm5TK7m7M13QDDeUhxBhtCIcU4aMSUJfeOp4JlorG8kYyP6B
11DorlsXbFz+XEhHYi1EgUD9IILmLpat5QPJoZJ8p078AX7GnN4ITg0dupvpES3jUSYo152k8QCD
FKFJ8kflv1otvpaMdhHDVDr6ECxldLTz38AkAcUs+tPTnUAUc/oSV1T9LczPPGUj91mYleZ7fXqK
Yh8Pv24tio6ou4X1pdB2KWqgl5mdfm1+A5ZxgdI5LaGSkRD3bcp2ow+NlQIXYVNgbJ7EazjPIp+J
iHIqx6xNA5+Gi5bRtXT5cxWiFPL0tEasRQPrWqWFR/eQsFDlBiGt5t3qFff6iwtMETZpJSlr6cvv
fN0AIsKzlUuSuKx6cKAjWWM5OPTaRleuKJ3EcWbY4CldmM/tLKvlUvSJeFdCN0DEmli5xQ6z/8ZA
TPiLdY+bi+2pGSwBU2T22gW2R+Wpq46YPnGwGVcgJeMaapGB0EikZL7Ei2L8ZHsHXc124ylZKnTQ
6b8vNhCNXi3UeAYJdSMENgNsP9qfDDbfbIk92T+BB8f64Ukv6IGkeog4w0pZkNPipVww3NX1WNnh
QamL1bL/dSQL/YG7ndu4gWxiw5taWcb+UrLgt//KFoON2QALFzR9xj9zy+T7+B7x1Hsy6o+WCoAp
PZEN96VALlzYsmMTYjGnZzPH4ZWl88w9eokMG9lg6uAjlTAaaZcwdfHeppSiWMbEWGmTAkSGzh2w
fZYXsHZ5syv50G7hOZglSY3dUiZ002QTx92VlvXcZLUCNrgnOd4vhcI74ic/GJn3hweuLgTEPiFv
+ULtfLWzSHKVmWBODJH9ty0mWQT1Tw4RwNp+nyKpM7WlGAU3mOqc6tPmOEgZJrqagb2xwWC1egKj
olf7wX9g4KkoYAzQGybL2PSz1uJ5g9oX+PkAHFvbiMZ4aIxZXX+6KbKIYilHhjzT6Be3jx1zmip+
zHl1r80TddaPiZVY/t7b7g7mP0k5s29IQ5V3uMcUsFMqiS0qgnxdMExxjx3AgENQbMl39ZO2XkZy
0xwlALEbhx7N+8ZoPwH3raZ+xWgQwS51GU7d8eADhGRxzYBMP7e4XuLe1oAxsNlTE777+a2bmX1x
EBzcvljc8llyC5GX/19U2OQ6/o5PqzKbCe7jQ7311LEXhiuVaMx+71YgbmWxh/8CPe4iPUwRsMH/
nbpPY2r4huQk3USueEz34ppfbhbvSg42jLZXgzSqJfGTOGG8XsqOYZ5B6UoFdBBWW8uAE08x9Qdw
YLXz/VMOg8RZjFHIi8IbtAicwvYS9Nm9a0e0fTMDn2QRJslGYt0Q4OgV0zeg6/8rEt/cbTpqc2z7
Gn4iqgidjveidftv7Uz2P1AhHl/HlzNojTkMPbRLJLXKKdhwxqPCjz1WW/cgrizFl/1yZQzD63cZ
KIxvi4Wif5pHWw6UwW2j4V0sPScTHQggclmFs4RKLPThbFrMkkGjhef828MiZcuLax/Gy09h4gTK
Sn34IXpf13bexrU6TNkdiY60oqhrEPCUopTIf5QfjgNUuS4+x6Kn+WsdCajW7nqTIklRnPZPZXlK
t7WuOlpmjtOqqmgVeXluvRV6Pmo5SSLmxhwfFM2vAN/FbCXP0xGr02BE35qZmpJVBHVstJbGCz1m
GvU/jkMUVNeyoTzz92itQ28zgBRsuII8cEpKwn5eqi+3tN7d7K4TA9hV2FEBVc1uE5f9SNomjTrA
D2t8b40+nu9Ze/wh9GZ2ZedUaZKBfaL+0F6tWXPPi+PBhqlb4P6mkjqrhcaKBwgAnKffnowiXUrw
vY2Ons/Za01aUv5BedxCECPiIGX9WlXKBuAlaZlRWbogwiIiOz3kLByH8sfGR2XUbk2yxf7NnrlU
05Bdo0i4gWkndoMtkmp7iF/M4rdryZRNeGu6m9QmSdPWk2DYGJjVz9jRxhDRauYcB/5IDpfvD9Mo
c/zzxViiy5vJt0dJy1UP6pS2//jQhut6iBBiP3qhmVCIMI93fPXjXyaNY5YVNbu2boFybSgG062d
Ipu+X/XhezrYz45twejQpMKcrLRM/p88XhQ+fwao6a0yf4AMxAoR5vuH9Qfyt03t9boyvqILT8uH
3uKyn0I60sz47zKMnhkjF9e8ibyyy2iAINJYE6Z9d9AVl410SAnolbKsShYI49MNK9+noqI3ZLDa
Eb+YUMM4nftWw/2itoK6bv2Ntxf1P/GKcx11K4OgMVm02I+OE6Lsgu/mqgSpZN7i+amiCHBYmOme
0Y7tQEpPSk3iK/+qpn5TgWievHhWN6nxa2fiUmGLjILl3gnL74KcgfOq2Ufzcyosv8IiML1Vi6eG
O+C8Y98D+AMLDDhqGEDFc9pFzrq0uIv3Ki1/Bcc6697yUoUz5M/YDQSebSc1Jvi35ASXfCJOXAxz
K/QPYz9J1kdXWuAn3axIE+B7LbZGHc+ZRQqDUvqRJamaDjxOmvbREtZXUt+9ILNNUUPtwuJLPWUO
bWQfqqjpzkVGXQ519T4ssL8jjgMeeyOm/xC42PaaGnzO8//7KaVebCI9gz+F0lPDNu5Bnslmq98Y
uMpphSpf0zBsgSkaVl6aHfJqX+2UrP617tc1P/2qU7cpiT9fm1nfHamPGqDosY16oH1TcN7nX6qb
3T38bUK3kD/No0aY6cJCpmJU+WE2/KWfxP4xLO23g0dvu9CPT/SkVC8Sd3ClPpLc1KeZ8R9O5j1r
708lxpKaLI2ilPKlf7rxqKwqrrwjysnsvaXXwNFbyn34dIP6J2ggm8nA56cM9XnQOsnvk+nFZpiC
ufLCmmuE0vZWV6JteNbUdkeSfVxVxF0p42kdZWVmK/ZLJWFGJmroRAb8RdGtoPtfTWcNYYtHvhxx
wCJ62tuMb3PJ66AoJsxUSuN7dwkF0UUdFd8LMTDNotMnbnMrX5tskJF3OarDITy+jAKBl4Cla5Hm
22NC9AvNr7PHXhJV97dHCDH5dC1ZM89wYR0DbvLeuXDaANfwXV96qoQ30lXMxgGQI9ySuQjwcMRt
v0CdnfJs0I419gbmnlE000GGUIPF/sngRJXWIIffx2y898VeECeLBgKP+dXla2kUXVzrtSubdJAt
HYVbUpyNYt31+LiJujXxGg8mrAWNSTAsCOGL/62M1OVSueL8QdHWAFMsX7h2MJBPIpdP2DkNtGWW
lSTX5rkSvEzEpvsWFuFAeISvKsGIL84Jd6ZQ5hxaj3eltJtFKC+EEwJbpqtBbgILH0pFOf5xRCnd
WI2omWHLP8W9Sg0CCu0useFMVPYoK8u7hUjomMVaAFT32r43zu1mPz9d9bZO8oeDqyaubBZscQ/z
sug23npiCr6WN0OMyHN/cWPLUXamalSl2eT0uHLD4mFolAfLeNHny2RBaKU7D4bQvWit4ZcFWLlB
LdOJM0AWvn+ePmuiojVFcP1Zg1YF2u2LzMIwKq5vbR/KBmGR3WNfEcjlcTWG7QVKNNWlKqFIexfd
ShHxuhjLJUYgQM2ZIqlSLJGEzNAH4fmMaeq5X+ZS/eKG2sxUFpGXqrPOyR1Hs57BYUo55jQIp87A
DpfwMXgnhh7RoOof1yLo57qyUBbbEblxOciW1WG4kVHBZE9wQmbxmYrcbDo1G5WYGmN/9EGoeJ4A
DfrNYeMhTFk4GrpDQh6VC+30dtZMtN8neZk6aod9Bvww/jHPaJ1xX9F9u16uSCvddCC6ycvVEoE3
lF+G1SapLE4kW18i33j+4F4AwJ2syZK1wtM4V88x1w1nqrpplrI2DOSxmK1FOtPC6W+A/7LO3I1j
TQJUyx3F0XdWGMsBi5JRssJfEYkEqw+ksMIWpw3yYb48JiEajhEJPjUXaRdhnvwWX1KYbOy5Vedo
0ediY84mlS61kqKS3iHjWmCcccSglHKm3qxQnhCUZ9TcUA+UVTPJx6G6tmHRjmUytDj4pcn6qbll
kdOPLAVl3YOFqUazjeUjlH2BgiAs3k0Xo9DfH6gicjIKrLX0hqTsB6GulcWln4C5J7+NMsjcmzXR
EC9hiIPBLGxc6k+SNDQAvruuKlIwvPGVh2cJinSYcEoqkDcP7d4fhrizU9p5N56AN0qC/BSPTMvt
Kv04+aGdFrpAX5Zz7ulcZB3S9Qojy0GqejxMVcfO8pthc0AdhHJtXfNstOaVwKPZjIjifMJX/syw
wIAHp8ivC7LoYgCIy7FGtikM+XcBG9o/sxLINMqiudWoCwp9C0tWNjCrvYoKZ0WqZ06S7LlDTLt8
3za9uMvi8gT2FwTa4WTK/1jmIBugpTZ68T05AGHsj/JDqbjE19bK1anCRMAAtJJ0f72z4okbziMo
6ybVqD98oReC2PP7vYaz3uVpmkV27aBAzqGiYe7JRy3ncKQjSVrS8PiYPMu7gzI9zN6/sRrfCj2j
y48Y+c3bS/eqJf03j/fsfY9z0e/4CBP++GAsK59IaS1AY7fTv7kT1gObvRnO3J+/jD7a6S6pdiuf
HIpN5/pu11X1UM0UdVR+n5qz44U6ATbwSqYge6uRpyFkiXNUPu5+LXb0Fz6t9KXg+oep0KajQi/H
pkoep1quFz1aL3fqYXjH/sHxOtySbP9tlOGSb3c4S0TFtdz7bZXAXlTUV3znL+sySmhIdzy+F7iQ
6rtZCswmBDU5FVCLHyP2w60je2w8AYT2zNe3KI+ccapPuuAGOVCzN0KcEyxYu2Of1rhLfkMLP0nA
/kWPadiQ8NauVSe+8UsWG75LAEz4h/CrDTlFInmFFukuqooDTVnaWaBz4gbsYHVoLSeSO33zSn1j
ayuSMku+TzW7tdKGWzR3eF7eNgBwn68ujOOQ/Ie3RwJ+8EfMIp7SY3hiQsAmWkq2b45nPtZAewqq
7NX+E/ZTufe5Tsh33y9WuwFGnlW7NGzezKgtRkn5xLcjLYfY7Hcu4wDmw5XWAcgOEXHblDDpc8gs
YRQ4Yc4rHTnt4kuz+5AnUB9CtfK5lBopW4ygVsrSDH6eotFE13Vv6M9MowbofAtKd4VGn8OliZJf
pND5Vvd0nBzwcACQQJbpC0v1EYdqprn83zluMnSgBsgc56/bC5QyyvHTDn1ji38T7XJlIW1Gcb00
4Nlrn++T0aGc6uWDK4abZaUNP7nAldXtRzsGNQFTk+MaU/ywMfsyS+1NRPlTvdpc+FbP+hTiITMO
cMdTO6Y1P8oZBJxlxwDdcWtMDv+Mv1VDbc9VRv611FPVr1KgsEcjw7rYuc1SiIV8oO54hkWQSl9U
rrFiFtIpZi9QPRNJKBpKaOYet/g/4Nf0ZdXp/igTmGDvW5oZZ3eEILyoMY52otzEmHzaCJPwx7ko
J55whgcNSt203CX4pgPKLtK3RvMbRczv05eS0hcft+evr2OWmtIj1/5ZuOQQHipT1AS63d51wIYJ
Doo1GXQzrsJld2KdAtHjqI5fRuYNlAXS98u3mO17poY+LPelP+HzsrJBj0FA3KT6wBaKrOK5LKdZ
NgIh+Bp5uTXHWL6re9na1pI5MpgE8VpqyD+lFQKXNqf7GgHRUXdE8BxIetmW3wF5KAV/tpf7Z+EE
2IWHl45bJoUtOLmAbxYjjSfYe1MdMR8K/RP1+HieiV8+rmhhlem0leQtyDEOU6L3TUz5Lj/+zzH+
I1ma/Td8RJ/YNh8Nobal/yIWAWpggIhBh9jiDDQtOTRlKfiiizmlTRrGlO3sdVjBs1xAZJTW/pa5
+IEyyRxUjeqbxG7ZkXnP0AdRO5VIVTj3iIPS6n/IvPBthEoyovStqPCetsiUrcuUbZgTdi3h4NOw
NDuJGKBD8HVKIetdd3pmiDeeoBZasTGASw8f7m26VHndpcEWRN2FvPlWgF0vWBKNMkfUxodYU0Kh
Xvkav3V1u+qDWQPf8N06MpSM5GpwBgJPlhrfoHf6hcYHgtQP3BqZ2yTWPC88aCI6eDvQf0dlu/EG
dD6daFLCVrgq1PeDlbW4h4moYBgBfmf/+ZnGx0w2z/wPn2u/WpcaA6ygYzOggL6hpiRasE5RiPmT
VnKh3JMImwWinDvU70OCrze04w7ozL8GPockVxmEssKSDSmSaE1Zb1YoUVdxKiNYQC5JJHZIV3nN
s/vtcFtOfWbDrobSua3PwqxQtHbSbwLRhsZgmOuRraqpzPfK/UPerrnAr2ytB6NpGI6E4PLipbYz
FS4necEGgwYjgpZkVrfHYX0k7QwNsv1p8p0Xp/Jffi2tr0zEQC4jAg2CE/cY5bbvY6R6Ct1JdlIY
qL3+bQMSd1CyOu46u3gWiZaldRWhVhFqo3ZEoDXaimI6tkacHoPaBdFV6JsNDQeZ/XpqwHYqtgyY
iDVqWQC7ntrGtDZdywPpuAVlJVYalGF3w0r2m/Khyu0zC0fd7gb2RBt33JirWULQv3ZkGdCHxnY3
4sSlrGXcRM6eKMTDg4Bm67EA7fvQW1msRua1+UO+C9mSF9NK70FBSuNZoFhFuyxEOWu+nC++cSSA
SMboMO7Jhi4wzdVnGTM3oKrGyRENuMruGNKbPQIKMGd0OrgPNXowP8miJlySeFB683y09oE6+lLJ
94e3xI0BK81ytXiRlP28to65XMR9/P43UnQn4T8VtHboco2/tKwjedVvdduKWsmLNkfH4boZYiR/
P7jGfOYExZ1G/sHDAfon+XN9/rN4aA/SbpSAQC/cfDsC2YuHoc37uh1tLMqflOMIpE2yrGcT97FX
LbbQyz/a5Bty2pFIW+qxkPWpoe2tc3c1Taqmp34f+no/VzkG4b78uFD9LZpqlMTqeY2T97RiHbA3
fKah7SL1aM44tB9sdF3JWtz5KpBUX67sn2zzrhNfYWd2+fV/GiZP+rJZTNwOm79xz6/whWjhL100
UuUooFhgp+vP/vDTC4tuJDH0xDwqJLq6v11ds/jEt8A/DCfNT5N5iykN/KHfmbv3h2na6LuViw5y
ccl34P8HXWUn87FfVec9am+JrBekPwooa9wtFX5wO8GNXWgdnwWzzJtXBOB9Wat/ENy6rZCSEchY
z9nuSqblHQR5DvB8qnJRDnmrVCCT1pPkNufShitOps+s0Gp1i9txYBo/yWbKtS9hjcb/q7NRuIX/
lIAfY2zvrHFWwUYnIYw6oWC7AVrcf3iDDUyLItZf5WTpVJyfrW6Dd1Ev/t6w9iURxTCv+jcyS742
iiGR0uRPITKw02CKg3FyYYOnezzQQYH/hR/FgMjOSFiokEI8HNo2Z4uumfQB6EK0SlwC1IVdxdJY
aksY/bFmDsbswXJKtfrtrHmhHYansqSamlQo/ia9NvjO3zdzTQ3Kvkk9p/jIAVBsHix6jmbsk0zu
4/wC8nd3Vn7STedmra3djVACatoL8EiLX3B65aoEKv8gM3/JSs/rYZI/0VoS45ckA/ALZ+36y5lt
pceJ5/seEnT2hAsBbTSW83J2Q0y9hxCd2BwmJhTHVXBZcTr7m8L+y9Br4x1Q4ysr8SffqAiRuoCl
CUUUavgveaHGglaAi7G7dE4jbYieD1XWsq0P66NGVy/nasrGGGQtUJXJrcyh1fMpfbEfjK5U7qiI
my/m+46KcuCH181tqILuoSkdZfQte5gXPxdK7dDkMKcWMhl8M1kN2PZXX527icZuU0P9It+emIIa
4B9PtmalH+y4KfSi7rCseMOFKnyhyt4R63Hwl/aekcYR7MWu2ohrV3AiFjW96yZK1xJqW0koA16E
6JAF6ZNmrSJaYySgR9G18L+KJNfo0fO1p7dqa556CsDrWVgKEDXIoT2ldRbiBq7oPftZtCUWIYmw
A+AcUwah4oJkKU5NmDpJsoeoXQaxSV9NXuafdPxHRCrMW2XJ0ZFxbOlTLh/9TgsIsYJaymdgT9jp
zB8fSAqgBhhd08vShzAh8mp3EcoDX+yPUm0wlWZqVyDwncHjKW0RuaK1SHKk46Yp3o+zrDOw6xAh
OCm8v51JXLFBvH0EXf+6eN1y0nGq3UI/42DyVaQF9kZVJLAoinbDowVo4sXCfh5HHDvph/WoPrDj
DwI5o3zJDR6Yw8L8UvPOabuzbpQW6fYY22xPia2rJGDDEFcYjk38Z95R7Fn8h7WYYyugJeNTlR7x
XErksc7xEcbzCpMydviq7axhPDoH5/LjhS1mVzxGIwUpKUlg6GbpuebaoLVtV8Vm9FCewD/9purU
Dab5z/9Uvuu+8M2/kGBeRLid8bBrtTOSHq7UayhSts/6pmkY8Bp9cRtLKDkdc/jTxqHQGAPwhf9d
fBOKhOdKemnvnMSbSqECcsi16Uwa4dyZZcLmlELfKOZ5lvQXZbW2InlXVp9Js4jHcaalh8KYPKxv
0Hnh9UOFttvvoHCyxf6DmrpV6uOnTSHWcsjyZoI/C683klpJSMiWyX5zmWxecuBRakqNVHYPfiS1
t19y/p54wMD/RwOkJU+kzmy4UG32OBN2hQ7yeve9K0LTNvFZlSj3b1H0WVgONbjB6DVQQD8QGEgM
ycZn73JoFsFeekAcqhZup9HsYSfxmFVcgkc8rWJZvaD2wCYk8C8LCrmR0GuZbguh8BwxKpo1/bCL
NuTtmmCrhHTP6voYtV+Osps4YLODdSLz1ihUikdSma0tJTswSaYLVKMpCwntgH+0pmWKxlv9177b
jnVRqE8CZt/qpnzXVTIe2hRS/+g7j3A1QCqYHda6dtD8p/fhTVf/JnR2899l72VAAEm1m3C4ys53
noIM422wLkJWWsB6mR0jRiVleP3T25rtOYIiDU7p7zXHd6IN57+pYWJpy0VSYJHx7CSODgphEnhn
zJilG3WQl50+kh40K45yIVRhsaK00W75ZF2l74E6xicWZl8Mu0X63922VTA0M1E/EABycE0Vh9wZ
VePxMhLQL/tYy4fE78Nn82DSnz4yRXNKO4IAxhb7nooBxaRVs7dRV+xiGtGhqeCBY0GbDf6IOkHQ
8Le9atpcl7w1HQ3Pfi6OVHDK7ppo2ELy9+y4YU89QiCqsEy/J78iaqvQ9OVAFETptZc0f/jPjwv2
5Q3iMlPH6F5sM9xSllXGqXd7gv1ZBfO/20TYDGTopECWa7Jvlsm2vBIEy8d77XdxSct0eJn87FRa
Kfeky4PVO2mponu92O5nqC2kslED7t0mDEBpzth00Qet6y4Yzle0krdaRBjV296AmBf/XSifUBYl
bEAgIvcUBG974ic2RoGlHfHmBRXmLw18geyoyperhYG8YkJOXl3XYHIUc22xiA0/WQRF9fvyASim
59Goddt3vJXukMK/WLd0vSLMyk73PYyJPOMnhizK0Y9jiiXaUz0V3knRrfL/pEx8jo0wi2uKJjo9
xoj1v12ztFme10S5hW+zRQUpmZK/ZbMqnXM+rnZPSiPIJz3gOD5loftFawvowWbD2/W0r0J3/3Ot
f0uS+1GGiKCkEznfMKtO+5NZgqrP5f0CWI68xEnRKXyYuOYj7VoC4pdN9ea1tKfwY/OE9VZWQJNx
cZ37WF9rmufXgfQis9eg7yabC5NOx6VCsx152XqngZt+TV7WVXMlyR+3liNCOJvBBKx53Fgto7Z2
08KewPkFYkBlQE1jdyS4bEhfjUpsWAqbvN0k0Pm3erkphpU4C0K+R/CGtQYOp/LhIDz90O4Ol1j+
Macw4Yfxu86v5+hawRNWnUvIzTyI8KgtMXUPuAz5Q1E4oXVS89uiHg+5xNC1B0qbssmBQZAUhb1j
oCxBuheED4PxvDntziLPGMvdWRUj4welt27k+Lxlz3CeOmVlYw8n3R217jPS4pRBM/WET7jjCR3E
bG6xt/+F7wa9EwhsCnplD+9YLGpSo4pggoiKhblddRp/gN7uGI9QyYSUQUhjBWYkUmavq7rvJNKe
YFOdWA2RKLYBYA7y7HgcooUc9+pvB1D4S6vVfRwkg4kzCGGY6/moKTjh3OWNusX3GzBgr25or5dV
HSWQzhBL446gyK1ETF3L7ufgX1V0aj7riO0yryyTB4NtpV0ZKnUlXeA37+ArGx+bmgWvpQRHDt/A
vYfBY2plWjhP31tvOD268yrn5HzHDDM6hdtBlGD9V+WPCGUhooowQZYgX7LDeRjlvDM8ZyKExl4t
9hCptgaqgMEnXh3O5ZcH4l1Whz3EMuU0vrwgDRwYmt8mcVZr90NSE431EHhQoaAxWtNJZWlWFipk
RweW+CvNA5Gz+UcponBZw6RihZPtbLvar4tthdfC2P5teLfJ/0ziyiBXNXCwkZ7hkvyPPAPvkZUE
5+kQS3kkAUjUG0/FkrLiztGTbBkRIA6lC/BEhDyZFWkWXskKS3/+WxQk8DumiQO+MtP3+YBswAGl
s7/nYPNjnCKHqzlQoThyR1H1x/W66sLI7ZfgITVlc8HGci+2RaJ8dCu0m2orSldsFFjtzzv4hTIC
HNPF1V95I+FpNa136wIs79kIiibR2CCDkBpzUm4/131ipXdPakIO6ry6jrFFjBffmwXptyZRXR+J
uReGwGPpwv4RgPn5y7PD6lW2/tIGFCBIN3ShqbytmQ/fhFYsB3vJ6jUigkw/oJ7tpP6fkDQvzdKN
rByDLqqbOVeMr+3zEfAXs954cllE9b1NjxvdN+6AV4Y9m1/1SzoFNDExZ8MC2RnoBWRP/jYMmJMv
xJVyQEsVruVgKOYwD/WZXnJO33mLKOhRxh2FU06/c+rEi+ZtCzNFzmfdqUOC6hs+B+ItPAsw4f4D
1okNhbjPxE9O9n2d5Tyl9l1H11Jw8Mhc7d7/0Ox49ChLRT1VN3K07FBw1GGaCkGhl3qpwTIsIEco
e9VydELtofX3EZe+SsWt36oC+TUobIc/X9IYL2nl0vJxu+nWxzbzFjnV+PptitKBFc/nheIXVT1b
MzgHMec+zDbhbtMYDBpGzKflXGXu9Z5EMln3B1rc4dIpZK0mte8V7pZx+2E42eSi94qe+eSbukTB
3iNdqilXOR9IRwj15dRPiZZ8LL8gyHZx0pLQUI8XImuQicXuAPTeVK/vtXEVZUckPOBBFmIChIhr
ObaNho2bIrDoDGhM4Iwfn9ZGOC+Eg1R63z2U7AC6n8Cu/GhMvkg+dpjbEpK/nqNOFlx9o4ZglL8N
JR5h1SBU3k6/Ur37div1vADKl61vxzzcAgeTofHskWaQSSgiu8++8so2l08H5empNbPHjaOhlt6L
4LuRE6+rs/+/+EYQ9Yk2xQxTVqBcO4suDAOHp+OlIDW3iEEvC+u9D5vnSB/PWGDnO28U9ly4o595
AFva/k3pXVgm5H8PJ/z8vzGFKeasxbp10zQaFO7ImaPD2AGkEENgyx6du5+PQBqziZHqt1Apjnsu
My5253qNODIqoqdne/wk4GJVBX/geQy7vl8WmRpvh9liIuwEdTEyo1YjYr4v5x0y3PKj/Djaif+f
k58DNZtUASJKc0/3GIq+//GNecS+mkJUX+0QMpD4e+287eA/tcMS/qD27iRMYrJ/gR02gdl+IiZW
D6kkSx16dHnI57N4cI+9/zvx5ZoX/l5ckv+SNd0j80yX2FVkLYnVQ3Yxo21c+aVveCupNLTsrv9r
OvexTN4VRSxbR7r/7ubm4Hvmy5ocLU2RRhEg2/p3miFcMTlQ463ve4qTdlaBkzV8yytxQvPtVqk5
nynCpRu2hWhsyn2BRGXbxYII89RAPlzAXcvffVJqlBjdGIQVRVagkMTJvOGP7AuX3IghMwGs0UK7
cyIv0tmr+jwmTzcy4eHu0hHWAFFrlPlDTzKOmKuXC8b3A0e1wMasgD/UQ6C5PsuI2XjNI02vhPWR
pq7fOd6OP90P5KZjRGKgrZeL0+PPnOW10kYuaI6V5IC2784TypSC9hT73sxaMAN7raRAhy+zGWnX
aif0pkcqhnSGgHrrS6Iqn+rRFCBh4AaVwxs6VvTg+2n/sw86M5rXnWkLkCd04Ux4THFU7TdJ8eWm
bi23KQweh0I2cqzM131vUN/mQZYuM3DKe2OrmSCh2VLJFFDj+B0XtGPBUkOQRTf00pOB4siG11aI
tJAhSdxScrpH4VuqGHBnzImU8XNbRrlNLXpCGv0fYHZyWzlOa+fKo3TVyftg46ETZVl60SUBGVoa
4qI/bCzArQOk1Fm2ILSRQt7qNyAuJRzcozHHXE7A0Xe+3+0+0lv9B+bCp5Mxulk6QDLQjyyqFF+J
JSpQtormcM/pKabAS1NZNsNF95ezGoGZSlvgmMVuNbo9kHE2WifWEiIewbsvbi84O9r0ZK6KQ5X6
L1RRas2uEqfOw9/+xV+8yUOrSmcqWpivpnTB/T7V0iSrZZtQZtyMnjIGisljIyPp0kyCzWKvKfoi
QXphXWY6PCSs86yifh0k4Sopb+c1yCixlTI8ysLlpXrWeXisxriQ9hoXP176rLWbpXjR07sssw4X
jnWdhXImPhbWOuFzUal+mWERpdcTtEuZtdNLxJzpH1p0q6clzD+7BoHkJ2mhHrjMQ4bLe39V+Gd8
f+SoMHYk5SsMFtwLKlKXwQ91mMn0MdrfW054UiQK0qcWb0jHTAKM7CXdl3AUzu3+cfvN0UsbUBco
BUdv6moPkrBiPaj1HBryMCJ1BDlvzC2rCCYf1UCgTWejZ+tAWMKKyl8ST+rmHDwPYU6wnYiQw9Ow
yAhwftCLkeuBN7spcA5dvJypiJlE7h7FTUJmM9MMf8GsgpQnN9KCyKk3QGr9zK79DPhZuFMA+8t4
ON5NETqsmcYjzu89V2KgOZTtWI5MLIWUMu8tTtc5VGkcFXIa2oG8XuM4EitKC7vN0UQ3qf31yneZ
SvJW9TeyvaXQXCbXkjJWnratXuCCzVIIeMxFYO5EfPpM9iNLm36ndcJ+6G1PU6ZjlyrByGQ1mSi6
CWMS17U5W2Et5aHoe2SBEP9LoHpVf3e6KXQVsvpdLt+tFs6af5eomRXp+/38q64M2MkALAOP9T6T
4hy+SkEMLFsTvs2ZpcwMT8X4rF9IFH6yHCf9plLW8BnPXrMbGDmpMaiIEVMZcwqDD1B0nMzClNxA
fwM2gdCV+tbd9laLAICKzjf/RXoU87m8IAczWuHKqJMRsYM8QeZnQ+BlqjdtGV0xoaNhemTy0P+V
NQgkmoII+egQwDZ8Cmtix8JL8e/aCmEyLzToNLPk/SWMGDboys8Am8TGbtraQbG9/QVv4mFdsnbY
Dr6DKB6VDtrx4cxVgTuPy60cMxoPgkeLPxjRk7oHPq3wH9dEdo+zwYlGBAI/Wpr2Fl5XBgH4yQB6
panwwL2DyhIrMkVYD8S9dQHEO1Q433tpikbrZRl4aEQvAqbzQwjYpoVcd0Yos8Y/TBm53ozVM01e
l6qVTeoJ8eJUvMzeDXxGyvk0qVCo7lhLZkRUQq7OOhQGEwrBEyrSEuyiB9bUKNQbxGN5Dmf0cehX
LKG9dwfhXIVnJqclVd+bHqnHtYwqrCWrkJ2T+l5UAaSC/j8vIVIgVg/zgP5YnffHIzgLljfi1zWn
X1zKTFgdkk7kOhxMTI6ipYY+ex80a5wXbV07KVBl8PrDn6e4iWHZ2JsfGzF3PXC0RBNscGKypKtW
tN4rBqgAeiPLIkfQ+0B+5AiEjk+aZUCJ2qiLAiVne6viKs38c+oAR0lPpI4tVOtG0kzglYVGRXdB
TJYPig4VDRF7ipNU4kFcROYM4mcaJu/F4/O1PtX9SwfP7f8Dr/mEs9IM/Lh2S1lD1AWiAE9Mxz1e
Yhl/ptJzZGzgBw/v0hZvJmG3kDx4MWv8KGvQn1mYTVKGEx1h3ACJ+V0rBZD/bTLyGeHCP2XX0am3
oD6x69Ty3grl1XtMaEN2PhODNvQwD+rxyRH+GIFRauaa3E9j+PhuS+C2rWVn2DTQF+AD62AO5eVJ
GxkUrkBPkvKfynVWi+Ric71RFYDJ4PxbI1Z5g6N4FsWJOvwh12Xb7wjdUT0R4eyTmyejXI7U6/Cx
Z0ULnFHkez10PM8MyAMD3g9wz48JzsiuTwgtYVea5sxkRE3AvWxet8yMclVaOBezVZp+6qsLw2dS
Oqug/Z3D5Y2FL8G2ieV4rJrrGHBSASKDrTqcgu2BtQDcNv830ajUbcvEtUr60SYTFNnppDrDG6f6
8TbOR7XJZGWHAa6/mnRUJTdThAwz8TdbWht9w6WqzrAq+3/El5/B0UFH89O+1BGf3GYCy61beUad
VSfW4MIchWTUVgw5qlwJW3KKLB+CrWGiIIv/4Pq6jCP9DzXJo/SIvB/LvrhaooAi9UdW9uQmFYsp
CaHFMYqybbmak8OWQ5LHEPZCFwM/dBS9kfTi8TMK8gznvFOufAmz2zEa4deDDxCr6lwyfS+VbdOa
iYkr+oUpaxY4AbNKBaa1YYiSU0t1CWzZVhkuvCzFl/g5bseY+fcAxKrlibXx4GYugfnWi9t2wNgj
8bYyU+bhN/5xTfoINOQH5zvdBXZJ7h8rWp0N+lccD0RecI6fWUnrPBka4/sRS1d5k0SMN79ISNSy
CEgE5zlFiOOTv//5onuGXLoitNQvPDWH6/WRsNTLnPsG9PCTzCDCjAJ9BdtY6VXPtJtZu1jtj1c4
FQluxA7f1ZTKabPeyrDKNxeSv8/i8xi4QLe00z2O84UNOXEpQAQcI9x5BCpzlQMWz2LUekjF+KWP
ftW8r7ZusHOgBxVy1lVc4YqkMnQBnwyZgMaNItURmUY42z2be0Yk8Ku8ZUnUkijQVa0n8ydG2daW
e2SEMPdnI+0Msx7Xj73JYEHsk+SMw88+INBEu9D1ngdupYa2Tl2GaUHBtPNtFUw+zddFz/325IW1
zhFk0DAXjlZpj3QeFnZ03R1BwZ9ULXSHme9uZu2Iq0h8jXuBCPJgkiVpaKKYDHiCECrtrEwZqT8s
yHEYRrTKIImfMcwOpRpMlVs6BT88PUDaUrZr97523VYcFFbhHIzzf2OWG1uzm3GNhCj4vyPj2uZn
VphvWpH+YKLGPpEs06UMLZ4oFuLudj5AnCSliKh16d/TS77RdWixoibio5kZE3GCBk/shqKhoE0n
+PZ35WiQ8qJ5IuUSnOMHvWFkuDZLzFHkDUj8rdvgM2g1uMtn2QJsLTLZHH7MDztm8UTKUjPVMK0D
FiTjZg8HG+lPRIv9GGAxExYb+Vq1ifO1E4igdLoicT3BXjCgTI+rUz6DRNaTb5ElALDwslEGfeaa
hnxQnIyOLJFWc3O4L1dSfcpTTktVpOR1UiMLTCH5yjFGuWJv1EUBOXRGEuRClZYUQS9J/TQITni5
PBrnTXtyI44YkYH9og8xX6jB2VK6+5SPkr6XA9KrP1/gj8KwGLvdtnOMIR34AhvTbf0q9lbXYuYv
cJ1GSwjK1NkF5f7loBir80M/wUXcjP2fAaaTYKn3LVnwuZUkx7ho7rdepGx1WFr8+Kv8xy4riYAq
bdiQSDpfZVJFrYCAIFTxCrSLQipzKMi3T+prmkXMiBe0yBp+8IbeWji1aytuBbQb5HYmS5fF6hr7
rZV2HktZZ4KGQ0RcWPhIJeEXseVuMixK1jYYCwWWAKtX/jepCyCJf5Q5Jf4KZHW/LGaGvdnXbRqE
9JU4IjPdAUgofjvGxmgvFLFWDCOC1hqao5CUxG5rlqC4Nd76Ol+vvIjGxfdlsspFS22DPvq6K64h
WOpXUN5XYyNZU2mx3a3wq3lyEqHrMo8MLShP053jBT2tGAR/SAYfedGTiBY7tEy/hIMgzf1IXvpi
s7aZKE6SEbYUyJal75pbO1UyfjNMvhcqRRW3XFsOMbaMivbxypmHE1HESRlrnUtokxI9EDTOKDNi
c+Sw3KVDg6Wj4qj435PeRUFPq3N2nJKE66DwO80HTD9N5j/vf+aT3beyYaWVbwPsrXPoTf9l8UYE
MUMYimX60v3+1oA7ybyPoXWVKNjaPGgt7OVxe+2kMd/c+x+3hmKPwpld53a2Cp9aphllDivt1tlC
pcBXmGPJendNPP1L2jOSmHloMifAulW8Y2KQSgiqy9KyubFkE+mBLDhOsU7uMfevJZxJu35oDfJk
FbrTfJQfZETOv/CBcHwTLRdoHud0T4dXHjkAuC2+9ij/+d17UwiSKyN1FoyEt7vEGwHnmzbeT7y3
cnxmrCOp2BkospuxAt6DpPbi0E5ulNvP0h/36lxxpEqYmbC/ZIVaMCbSGBrCQhqJr5A6BAsLVVkN
To7evhSzR9CmEJcNsrdjQUw/k70w8ef4GzKvr2QKKcXQz7wUGHqZP/gBotr1CTog2O4u7F4DUqjA
JgSQeEULMuTvWS1O6U119fzKVKtH+Cp4C3z8+PTipmcSKMLTpdEwyi5ZK+oUB80hJSB6pX2zQrev
PX7TXgiijwanNLm8jnlom5Z2OuJJb7rT2LuUBWccI6hdcITrCbHZ4vUepKFqPZ4fGxb9OTqDfWrR
vYCOz54/SscKy5NyO0X7jlWnt5YsCkRgryhNJId0b+QJIp/yYqbtjsFS+GcP+XftUm8Nu/UFhFes
AdOUDZodK3vrQgDtKinDAYW50NTLlNMq4yRXPJjpWGMaEvF1a5TGx1okptV1IFQkSK/0Ii3ji7jY
JI18ZP7RB7hrvUclOfoD1Zz5ffCRWju1tkS0RscCVdDHOOu6av3g3BKQEQKCh6Sau57VCRF8eu2y
864U85YybOA81+dOPZsRtl/I4MFwvLIt+kfJRmJ3+79Qhffq0RcjZXsXyF2dM26IJ0AQcKjo5tTe
L4FtEGUut/sTnAaCuEqfhAlT6tN6OjBSrARUqfkU9HuKcvZXLZKAmLIoNJSfaLUnPadYShteaAji
/9Xd6MgylqmRCRQOQn2avIufpwzJDz67YB0Gn95n+rOPguzK9ltyWkDHeD/rNCi9Zk4/6oRQFnHp
NQWgd2fYSGbc1rsHVMSKxKbKfBoDfRhvUrJmElE0xRioBLy0aM3IwfaECl0HPj21AUL4iT7g5n3q
ccgysxe4zYQbP/Q09T/9+DBFBvb89ldh0P6syHD+HaVbpdqeSzKwx8U8q90ajnlqP4eJFEy0hxU7
dB9zNP/gq6wm1nr/hKzFCuVZJ2LmWRkre+J0zmEvs0D41MFbAGZTRZmR9S1WzBs+pWEdhe8UkpP4
TbuMWxu6OaG1FPkBIAphOnrBLaINAS2tTrKb10x8ddYz7uuY+IFfolXt7o7EWJza4eLoABdfT3zI
BepSPyCMBvAjTF80lC90ER+sXe/6KCNmm1egw2S7/dRz4uslEND32ABaRNRw6P4PWi0yx4962W3A
QoffL6wVKadF3cUtL+NZj4+X3yosQ24ac7W3ItlUKMiTC7a8cJkui3598W7xqCcCw05rrounmqnl
xS7ZrHNv8DfWay6Ydde2KMzlF2nh/aSmQyrgTBP9/xi7L5hFrYEaHInR9YZI3LRRK/ZzrblMk0Sl
VUlapHj8LZGmvTLGMAt0XRMhtBJhxKnrwqAL9EEp4jf2zHUM3avNhqufIfiikmtbn3IhDVHqUYo+
xIAVXup7A9ueckDeOlUL2V82syJl369O0CxevSCtm7JYIfVD7874VMACZRxRojIQ9xXPr8/8Q132
PbAMDNLoqGM0Gb9ERN9KclW0C9Uocn4PPrZL7unsVbK+KevF6pJgdbeqameL73iYWowCg0MOEANQ
NCAmRnBJhWfr5vKNYjwtpj+SuHoSlpOoR+SrRVB2DEPzNBqNQvwlpZOe1rTUgqFuIXYTYMhQILji
XFKf6BO8UWy3bKvujb2oIsOMwD+1WCoC4HwLElABGRdE3w7k+34zPowJXO/BM6SN3HE1hkqDf/zc
LCGXWqgG01/S7FyjNY7kmVDLDBBJtvdfOh2CSXanfPidj7IFRu5WI+rCEGplx5B5KM6aVSUu6y2G
MdpJApnIMpTWhiZYxEsM3yc9MCVqAusjCiBoO0sGVCCN2eEu7opPPZwuVV0fWk8qxMdCQCSjngZW
1L7+VALJCzuvlqd+Zm/HKQFD/TLYhLJ+9PcYc64zLC+Da8LogwEM+X2eJyrqcW5V4uqWyB/sm9dG
rhBsfF9QC+PFYar7+lNC+z2h4FjeDp/wTlNN99rOo57voygLuWVrBELWKxviuE5njFWA4MPGpyXj
Nn7s+Bqa0t2oj7cw+vyZVBeMPTR4qcQmYKr4tfjD1zht22+106drj/fjibgsSSBoqkMyw+b0LanY
dzHR22v4smaEVEznHlBLP6r/DjOuHMpqMtSTtAtN23ZqetYxbOPLDJXd/ea3kqDiYlgJnGTMHi7M
HE8uwZQDT1/fgb6EWInqqpuRkJgyfIUgqgbqidq/ZyK4H0+MMZhxqwsI5BZmW4/SDHRLLpEj7ExV
r7lhwkj/bH7g+WLuCSHERjUGeyWsItkmYnNw9s4YdvDVWv1MXQFD6ElEMVgX2gVOFpO66FFHp/X+
yI7dFg3FleDFqokHvq8VQfhZmvAH2lu0wT+CL+JUxGGdxq+XNcbcDDLhtT8z+C1eIFGk7KGouJC9
1+N9dFClq7SFx12a0wpqI6EmP4GNP5fO6ATDib+4mL1nh++KWtDog70tMzhleRLRFTcXvXa6BYy1
BGRUDiX2A89iB9SEYD4Sa0wI+n+UCYHl7eymwRcaDbQfSZ3WoBh/YkzfSFag0tB6bnsLvJBL5ewX
Y7/Yb0nINE6p+rm1EYCI9UEkaYu8FZWfRPBlMfpxPbOUyeehnEpSQkII6B1J6ef3pL/0xUt9YYMj
OYk1t0hQiCmC4jLMDlaWJviC0k0tgK6dr8RX2s/zlNlyJ2G5HshDlULlOUSsOWMmKUhBDAtNiPxg
oAZ0AaKer3EJ6+lPkZJTujzqcR+r9LKytUJTPpg6h7yI/tLGxGns9rvK5Gch6TLrChNEF2GvFdaA
QmA6GFk4k3W81vID/qRk6otT50lmAqeiw+ArByDNqaOYEwjBOZQ6zgScPG152U7fQpIv7NjKp3Iq
Ta39u2OSJCNfKjoEun6oZ2gHaY3rkhU03hCaNCbrldc7BPNY3R09DOpZ2lMF82e0VKqVBdAOF63Q
0BB8KPakOxNtn0+mmLosrmrXv41gU4AI8Z+cxi7RGKrfJPDkbtP7j+pexHNKLGpVwPIUYbRSiA5W
qoneWQgrkcmJTtwhYuHc2trSIkLozJFyaJhIX6roHVb0i1+l5BI2wToUpMewE1ut/FsaIG2SkKBf
Lg9GJyduiC83XYm9c6Xmo0+Lb5lR/imAB0EQncfSxLOp9/ZsyY9G4JLGWS0DHGbzGwEu8GOX8GJ8
XMfh18LmSzpLNJ2mSrr4awiS8AvhBT7L2xMgZIo18EHdoR+VvhTbLl4t350t0J9vnzixm4Gv2980
QT1DDdu3/9QDmy5dvOktOvGgW2IZA7Ctqo3VrpJl7/fxV5C3T18PukNyUO1a3kqbVZpB/LCnyg2w
ut+AHCPhhXV9qu4GN7psR/l8MkKTp5rG3wnEcJ3BM+lKKjiiYLc/aoLUxE3qsMtDI2TOqy2K8YHl
lu24y6QjuPokh8n0KRkReHFn9sPefsRk7WBvaiK+pI4M3B7gJNpK5MvLq1TOqfwWGbNnp0ydOwBg
fMedxFUS/nkh1WnpFB5k+ME2RNb7rHHdWksqSi/bXi/icVlzVnJHjhD2hNEiV9M0ChzgKfO87FjK
ydyigDmV1t8b8fnxG+yifr6ZR4gXBAPpNUOg/YI0gsiv4UZFh7B1Bhnk+mwZZNMLpa1qRNjxHKDO
hm/IGHzJR+rrUxS4T91ujWvd/R6S6H5M4skV3bTDggBcxX0DoUBK5Ss0qcklzH7crxTWwOITHPDp
pdRQvxVcKbJNoEj2KX6LKKunz58zdrRXdelSiptCVhRM+n2pbTqBMrDmMWyjnO5Lokm8x+3yy9xq
c8TrfgOYLkNCC5kcEsQmtvreN5cs55l8CcC9DytDdHk/x4hxQ00NC3I3R03O63cF+5YBrsvDaGSj
iSjKyhE3Pa/jKylbbDuvLTuvfmw72Ebh9sc/VNXRH6Cz4qapC61l0mq/hfuJpwxp9oIBI7JWVgV8
H+y+iEUkHcmUWUzdLZcr6g3BXGXnwNGeS9w8CR6oQ/Bc2VgadWLmy3GT9D3VF31uCy1MfgRsNmOM
rXEPlmjD23vOaF5StvzqB/29OQ+SN+UanWw4CwiRxYY8XQZb/Sa3pl0OdPqkIawULLihjXBYg5ui
X2z3cKevQnOys48tSqJyOO0E+GqtljfkLBLKcCdcEEfy9hodpv3QDIcu1QA9mxezEnrCoMq3ja4w
f+XV7OGmC3Hc2xWlejYkcqfAm2KuAFcaiaEVmP5Fa68xkqixWcCE29W4y67cViPZ1ncJc6GNWbjg
+notyiUrRaJZqCh5hSnSZrd3pzgp51Vl65+4oOLMMsoIsD/UNfDE5p/SIZMzcK1Va2Xn+zWhoQrE
B/BRTiGFpNtS1uAig2GTeKdcDA8mo0a0h2o7fhGmj2UZ4mxOiLH4YU+5/V80R5UY19yLkstdSvX1
QfN0st36+mCKL+6+NXiYHvKtymwPTGdAsToKADRAuCel5tKGHxeNgG6zhFWbyDvmxbPuuOswfuOz
Iop4fOg60RR96bWLYecU3+rvTDZsBvhKrWvdxHZUP+IRlS97JPt789UsIM4DTepgySFruHwE5xRs
LsG4wXcpJ88JXv7n3JkjdFsZB6BJx1RoM9JBtcIE0SBZ/fKswtXQZRVWTI4520udOdL6OGl+m0jj
wDVMj3FKjUHTaitG91QGgLvAhOcwaQ8K5azpIusPnlO78Qgr9LQVhLcbcTSElgqQqekWlewLpcJ4
1QP4ZiGQJwtTCqWu0ZHWyUCkrxsm6deiRMTjaxO/tRU97napKKwrZMk6+H+hOV0Y7IwBjI87S4Zg
p35wxib4sIITZ/pfjJMpDI120jG1OaeaI/SaYqQY2Y1bl/SQXhtxdyKKun96p4jz+JnjmIBbyqYn
8N/X70/MxQ62o4+1ek4jE1zXgW9plkutxCns+ZC40gRgG4jWoQ9YWAdGavs05A0UjXwDpZxla5D5
6jqnlsISJiadgejS+XrwceT1JHCALxodt5g63rKMqMIGLrtjYhD30S+pMUIh8s1TrhV9RJ+ZLs07
ki4F4kxgeyFRXSvpBnTGxsYuT0oRjLHlangsL1t/U8UMv78tpoCySudh7WmJpT5a1YDwjE1EdsOO
0CWbeWFL0eqEFhhifc67gMsLdVe2GIvoedd8V6kx/mbfiH6S3jUZW6oZZbEPKHiIwcX146wCo2wp
lxb+m7EeeCfkEQqPmqUr9ZXgxZ/XsM1+y/bawXNqWuiNQdL3OrUeDgPpoR2/WMHOe2O8qNT2PdGa
Zyvj46OivEsh5WVfevs6vg5GCOumFuwDRF5IFMavNg45e1s93bZtviH2CWnrT4EE7JGnRd6mcn9w
f/NZ3+A2WKIUtGdQXE0HKFu1vFAvOdKgz3J8by4xSlx0at16ZncW43L3cmJZZO7/L+CgkZmHdw5C
nq8NHltr8078OSz/NDW3Z43VDf99Q6HQesNG47GI1l1BXH0oVkbPOp2WitVht5iLN5uXv6Vbf7KJ
tyyEOgOJO5uDkHtM7aFuWlNfOB9Kw8+juaQQ3ELsKPqbAx2x0ak8obOtfxHVwxf/w9pn+C0jzp4G
8Z15U3GAFL/0Zia0MqYuTIXRdDqiXh4lIC+foSKmk5qHvLBpixvS8GgkkHP7A7pdYxVwPPq/Y1WM
sQxPCST53zt4C7vzAfdKfirP2hxNekHVD9R6lA+bS5FDI6tC+aBapdY6QUaUMwbdzEMLADuY7MRe
y6QoBbX63+BiemHqpehHxGFJ/aYyMOqRVzTA7bRIJWd3qRjfDgY/ua8yGzXRYdQ/uiFnfV4ATEJh
2I4OhnPzmhOnOiaFlPiRB0iU1piFcO+13A1v3FYlkxGrUTGKPs7DE3n94v+hUSgS0FvtyOQLIgrB
eO4h+n3ecg4lDlFRIz2fcFeumdveWQASqjT8ZEYDXxax3u90Wfu2NFQOeH+QFuW8xPW7LJ1FBN6Q
kqG1kLHuqghAqmFiBmU6QKY5tyxIHlU0WchaNvuiPu4/aj2np8+etFpdqM0qc/6FWzCjvYFMEps7
A0SghuJ6VZRClZYe31DGtrsXM6RkFCt86AvF8RNK0RJVACpNxnKrriQsKfXIK5wYtCmfAkl3lbMM
6LGb3tJjfbcj8kfPpT32bS5iljGGH0aV4V7yg7OToPkVw+STAYz1ZdBUH5Ahz8sAw14mQonPyVsS
efrG3HCxIDvMkYKpwQMwaAl/9hpH2eFqOv3RlXCoiXfhYDFeWcL02z4M8TLQWZTMRzaACVx14hCj
1OHvKTmOWSI2mwBZedXKqWd3AcJbeQ2hqylhmgrlR/8taiB3IxVvTCZWoxUTLXwtQ2uUgQDzNnOl
4hzcjrE17DBSd2rv1c+cLbHwyw7IgbZn3C+F+bsiwxjnb1BwHAmz/zbhh2mXigB/uB6M2Ano96Qz
/W731W7alOgjdIUc7D8V22DlbAZchYebsGXTWV7+EKJjpalCx96MS1jcODB/vMV7A6PQMUlZBcr7
Oxp3/YKDinJBGIQHjNVvszuF0VWd0qVJajgnrgRnfKUSh2kzjEFz/6dfgDZhpc67g8xXJt56e3OP
5O6LaOJX/mkd7pnoMwoRNtBJvYjqsczSfKn2S9FBcez57Wsh+cjP/o7+uJGgs+l3EUTNjO2ptvfr
m1iZE7oKhXHqhUJW/JKvgdDwuuSdcDeG2j8CR/qcsvDvXtuS4CSgtuMoSPXpt3NZQgwU0ef6G4mH
gi+cNkGVxYRMjK6zDI2rGbd78czreI6icoJ6uxhAKytLKCrRrz8BF8ZrhOAWaBUUOXNWJ1lZ/K0d
rHmrCG+0oYdQjoJC2ig69fRBpGA8Ib5o+xEMwd85dsqi5Wnvcj+YqfnFVeBszf72G9qC06OCalFQ
cnSzi+SJLAyfjot8rmduKqahlsgqo+XiuXWD3cHzU5ZQvqTX9Vjjm7rgKJKO2jWoxgluFYRfIWxa
GvxvE7apfAErWiTTzfXGoqsh3JKSh5Wt4vRzfJp6Wo69dQMIv63Un5+wl2e/eMryylpYCa5phhHN
pekKWbCgzXZPB8cvjkED6FhPDO8AjAjs4aoakd+XN8zDbE7oHjcwKa5hC9Sbsk5Iq8+H9hCKySMQ
+LJAxaNqKggX+DGAdVL42jvf4M53Pj4mZKJ1oUOOfHL6BE8haBh2CDMR0aAQ08VOf/Sglb0DYFHq
WJWEnIFDH09FAamJCoZ45OhtwbnSbX7AanWOJ4IcsbNtCQxA3nUfI4Ln5rmpT32m0842hALj+dCd
y4e8gXetUCP5gPf8UxfZsRmrQh40Od7ZKVq91V26/DzNEXqixJrQzRhaQay5l4F3+2V9KAJFK1T/
bB0USX3hohOukJ7c2/yuUHdKT12tasNB9GYGIGaQIruhIRx0XdjPwKMuAmu8gAMBM5tuXarHdN/g
0jHogr/P3k5A8VlsnffBUXSyTTE/H/y7yNYhH3c2iZRXn8QcVHB5We/a2u9N5E3dcXS6gbfvZq24
zSGQmPEZ9hK2+RECv3Qd5HhQJ5X2hlUSaiRGREXZrK7pbCOE5VRNonxRz0dJe1LOnznlyeH4INRC
zYMCe86I9clfUax4hcDcmj+8DYAr+Xfpd6ax2zURBV3lPAOznfKLBdqTeyFc3ujb940Xo0wmYcAg
YGBHW5u7CsmoWO4iaG54IDxA1IlouT72nm4PD16gBiJszY1Exs9qzqgcHg0UVwmPtiHpswhfdkmH
eI2OOD7yiiOTSbtKnLp3qmSv98Y88P2Pn6HEqRYeNByk6vhtL/HQOGzmLKGtAlu53BNxFAQgpFD+
eR6BBzEaAaSXgocK3oP0nQKylUnPjBWMcnwyo8GhQWoOMnb3dKxjpjjswJ3yXmkZwJP/Xq7oOjk5
GmeqEQEYeUzjJ7NRPGvYJ2GquTlKgWEOPxBE7ilIqliS1K7sMW9qqY4YB6roFWn/TODtsHPJyCaL
htlCJLwAgyIu35HzypAx1FOhlcPAq2L13mRAh+I7Z8N+D6WtYexmyyMF/8Cjf7+u6wOvVkv8HOwY
kKDLlMv4I9k9TUWXBima0SW03SyVzAG5ie/0oa8XWv8zTVvz0T/0ncs4SjRacHsbYUpAINTrlsVh
iKktuMhgTI6iPUv5Ih5fAsdJf8Tj9cNVC+Ag8YgH1CE9q2tWTcvmbsSGbFP/obuD2uufYkK7Byvo
QsrI+fROcqio6bSEFDg+GPmMdXcjhDmJ/1Vlv65/FtOlZe6OnX5UHmHz85AVZyAY5wlwzHq7mJ9x
sNOdzLzwypg0lqabRbjFx6/UWG6BOUekqgUplmvDw+KLY33hJ0b/Cr+d4OCH0mnwRyVgPzMh1JBX
QCMAFmqqyiHfPHVYtrGVTkropPIL7muUwE8nw3wtaQI28+YYBwV0L25X+6egzfFaKKjLfieHfJ1p
X9zAktm5pShjvUSvQTTzxapUW5xA+FGiIyRjXd8Yl6UP7uM6Bby6FQIniFaG6SDPLx/mllaMdCsp
zIfYiZv6+17NKx9ICNoInEZUu34i8EshLvgkmOipSHv+MjeHCMIYrwwahY9EwKRaJRie3+N5sT4l
3uxOM5luILPHfVRFH7YR3MsfBPHUZ+HUJyd3E5mcexgJrSGvE0MlxpRDnxcqzaMethXBAzpQf8z2
BmLW7WYGhhExwy1geuONoN90hYaoIFWDDNesOlwHq9A+xUbtQ2XDavLSN5Tm3RnGWbDvC0+0iPjJ
WL8E6dEW3Y5ICGmN9hb+l1e8qudL+VdhzYvAZ4t1BJUsbFa+k6T4S0NGGTJVTyYm0lKLnEPx0/Hm
tJCxYdLl1jMh2wZtDO9vwlPmm64cWMW/1jYxs9cXSN+2FaWWQHOlnJWIU8TbHMtd3sqiYsl1jkP7
9iMu+e8U6y2I3WLWqgiBh3TdyyRkzvkh/nOhqa817+D/fqjFdpW/dfuZCnTAs8G0LX74lYWYZUmB
cXWNphU6XhWOC2F0hK+YRP6XZ8elwfnpl09w7wiUhkk/gSaSeK8zgSxIlDe85rFzDNd2UeYVXRjx
2528bCvm10qw0CHSFBpqiYYq397aMMoG4mvEJXDygeizg/iLJF8RqSRj7K/U8ZbWoCFXD6+r6DKA
/EZtWqrKlaC5CKADBL+pN9sqtkj5CILzDxN6xbSXiqzq1SOAYeK8kV1/cDl5Yu4SGHf3L9lU3+Qp
cX+LO5sEig5fkzrndH3TXeK02EeBF/ZXpOe7Ktvltzudr+itB1sOayi2QRHeqNdFxhSTFIM00UXn
C99+qsXyOqluVuPWFZxWzZw+L2JovcIAYOnyJDpJOZ4kAU2rJLP7ForEXyJ89XH8a8ZpegYHSiih
Dv8BnNZgmPZPsLQwEIB2Y3pYxt0xD8Mbflsh0yzT1RYfEEXWnbZARL2/oUSKHzySrlP0LhD/hwrc
d105yXuSPpoHLvjgnmTMFLhogIobsV5W6L1RmHenYPBzjtCA1Pca8Ydq9n7E8e6pl6Pxi6sSXaW1
ZkNYKwJk2DJruUh8qr915lsiMjVdJx+2cXQpwNsJXKfxM2Og8l153lSXFLJ3Msokb2Vwcf3VXiA7
gPohjWoydY0TeyvvKwOTQhC9cDtm6I3kWqak5oU74J25C5s4NFWfnAspZAFcB8iIWjqFtQW4e7A/
3n0GgEbHa3oKVNE9SXrD0XgWl+HrMWWKJhP9BVbS8ATGRrVXWzZJaM82YtWRjTWBZhRy6UT32R3h
biFgFkUCvqzKnWLBQJ54J60oVYKL+2iyxr2v7d9d4O2dYByF2c8rAD7plBptWencTFrB8KCN0Umw
OR8Qwx2207lF4hCAHneYyPqsXOYi4XR1B7H6zImT8azFp0FYm8R72DJQ5VWLlk/StbzloUUiZegu
gTPBXdEin2He4yUxxCsgDNabTMQ4HDN7nEVxq+fUO5ddbgVMT2/ZXHknR9ec2CkpB58PxurPRIL+
mtKR5J4AJQvClQf705WiFddV+F2hgGzRA9ZZiXJGk1/fX+r2g2zSnB2wXp59lfCHdA9OoRDUthYm
wyD6Srab1pAEmgqO9X06D5g/DdBP5f/n85AYowDehaIJWymzAfsDzt3qpl7shXmXxGFUmvsMq7Mn
PM4XsU5N/yvX1DlQdqHzjVP1Bd6KAAINFP8ONppwhaxmTFeDxoddlC8+t/ydYPUB4g8T693zT05q
x5EPk2Xav7ZVQb11DCws3tmkSDWav+oL/8svnDLDTR3Ozmt3Tj742VeF3MKeWyRqs262n8PtuVKv
KNIo/vfAok5OhY4liqTEb3JkS6BiCFHYPcYhXlg56w+vuvN3uQTLRLxqxLt0nHRMMFz9TAu8oHLQ
OgP5PYLWbdB0ZbjRNz5JJ2Wta3N65IzNE9dpBTj7NtmAkVHrkOQZmnkrBAfux9UYPU3utFiZPWb0
PmdDEqzJeeGGOlfG7Sepqsd3h6a9ZybIM1/bzdyPZHg8dhzEWlomxcfKiNuqwV6X8Nm5Hwb4PPi1
XkrZX1hTyW8D3/lTdfbRW2xDdfuU5zEcTGMFDA6ox/FLLvn81VU+A01VXiAP6VklAySzj7iX5/Q5
Wj5+T4k8YVSE7CeLjwp3Q8xO7B+Lc79F46d2tCUUzKWyiAVQRINfVQezMPID+1Wg3/umktXc21h6
ogcc12pGk8s6elOVGQZCYAKEIe2T3tHwTmyQqrJMVI1kAm9sxffU7nzWPiO3mEVjTb1FcpsfzqJ7
m5lteYLNMZ5uVBBUJBfsRVZvRNZiANQTLbqNTxf+Xy/izyYyiB/uN4dA5W5I1m1sHprXaibrNQRc
YzpMxxCIOzTZubE1eWxx8AnP+VIyfowxPdJ5HlWnHcthROSefL+ruU3lYX3G1DITXMvDtaJalzcA
dEtc/xjYJLIBiwskXNy80dgH7wQPPM2PCEoadPz0S6V6kWd9ZVT7itHcuBIFVlUWr0X0V53i/2+F
BlZjOzs9vxkqR4gSs+MmL1bDqzqhL8cFGR1QZUdHbDpe3ZDwTieu48Bz8qYHSJQT5huhpJc2FNbI
3/UhPtBchCwHfqCBiCYRxyRBU+S5JDvpCj/wWkBk5k7KoH1fAgdq0ZHNcijIZCG4S4tXNWEBCAGw
luo9mdmEVLuIQxMFzYUTM5qLXVBM6dP05IE+EmDJqCKbOE931KR63cFZbiN45GmSS0kmlkPqgzwA
B2tVc9hkfJTsHHIWbilw7x+eJHjdsmAeT9GBVrLvWRhkBsvDSR7z9hq4PHyAxe8YXWomiPh29oo0
Ehyr7EntX1+aalmwCETEjIsc1sUlnNuR2ipQv/RFSpXKv902tmj/DB4ssbwwKarIJsDTcp+jJp9g
FppaqeY0VKE078SNYQ5P/W+8g23FZBwiLoxlcvqmvrEqnPMFIQw476uFNvpTBxXLwD6YB/74OryV
u4ZJod2tnnbk5p7cnqBPycjg1/L9ZLaIKp0AfO8n5sMsV8uRKjwjwLARLEWytBKcIGizDli+E4sL
rs03uYRDvyyxQHKJVgHmHQm3zUItOdS5p1unZTKFLRbY9bxWQNxeGuQ/vN0wBedYiDIpdRJAdqXj
KeGi3eu2WajZsqraR3nF5vzHDvdfzckHvBDefNZ39jevUNugR6qUm9H3xXOePMNFdoIviGnd+l3Z
H0tX1eW68PmzTkrVPq3TzpY5hw3A1R1IHArlggsAGGzNIC+Rzy/7gf21vaXdm8PNJKQPm7bG2vlZ
y89Q7wOPm5EVHBBepmpHYToEy+uHvKvuP3DyRn72j040wVoH5vtweu1U+UvOGgIrBsHaHDPUHCMe
6wMywDKikvhB95sQPQAOsahgab/n1hlD9QJ7tImgTYKqhKgAa3U2Bw6D7FFO03oDq9+ty4/xO6gg
0J79UWTCunyDM8/7FdJZd3C3iOOi5kJm7qTkDao0zJB8j3z7BkjjjRETDVDcScqs9mzUCQOe2h2g
oDrprP61sX8lU0qMGB/bcVaUsCSR18pmHhu3jNRUOom4i14Z36dFQ4I5jK0ZWHJkRqHpR2/aihjF
eMI0NnWYS/Yx491/w0azJEwrf5RoYxXBI6fy4x8jTlnac2Vds6OiKlESqF0xx21E2TtkHzYQaTvL
qiePPEdTjUK8CMT9I0wbOycijSx+LzCvbgb15ynO4+kLu9tXdzD+kEFJ5yKYfYHLQAZYD9hHkqMx
1iRo6vRFsRVr7bhXQZKArDVqCKv4DBuI/f3vJ6LoFya1aDN8U/NRgWe97K4GuxQacvjuEkGu0jG0
mKq2U3RBrRDrzacgiu0KoC0tDfdiwnWCzwnc3tbQFJi84remUwPq0MHUsgukb3zHK+4/K4sxetLf
dYTxurJOAgbRp4CbofRser86amPdQe82EWuz9GtzyoOku4dw0hyXYGq4In4BPQLPtXepnGEUiHjR
lSBTxQtVZi7WB2kEW+wWwWO+ocfR7Y23HCHwKEGrSIzGtSbSIhGJ1F86IfDTux18exM20cfJtUKd
QcsXCzrHnzxbn2KZGZkek5m8pcJaSb9Wt6klFJ/qxSnwB8pi+yXu/59SJYDXlBC6s49yAAcSIi6M
+jBnCdYc0el/wYlzxBb0sv1SxLhmQmg70yN3f6xnmQsPRIVQVk+AisN243qHto1Vo3m6ek/Blgi1
3tTLK5t6zc+kldAkdel/au7ZPrcVoVHx9pPO0X+Ywk+ueDKJngK7HOIpV4p4+KEFI8mQg3QoE73s
w1re9VBWtBfDCN7WH1GUl9X1N2n/BhRH1DMuMjl1O9ZPxs6MyOkXXyWwC8G31VzviF6lhIwJstlQ
YzT3/h16gxDqlKGVHM8D0M8tnkP/t1JYHKhBroinTkkr8UReohR82t68RjgaKtLHwXMzzNIfEs1D
JPp5R8IrGUg7PO7y8jjkIXzyf8AtPs7qLLR8sX7PMs9RFBwSSXpRQqHCEN3KbmDuloRlG+qsn9jc
pZEv9ojo5aA47ZjssO/Ce0sYFCfzl1YMizmWkullNMGARm6pSiNsEoNt29EiXigCgqbfJErWgaVq
E0VVO7QZLPV2QyX58hbOtEkL3cbXeODhWR3ZME4wHmrO4aetgnzXJlvaP0lWc1e+lQRlkpsdg0v3
XkRtw52itaDVI4yZA+mltQDmBxWgDMSKWimRm36H8cLOJtMbOZn8Zpf4C9DrqwlP2mdYxnd8q1XR
P7yTW5cp9H3DryRt9biHYsuIV5YWvvtydnaF8kxiSNjMOXkey7nyKRdLjlg9fELRFEj3o2ZlNPp2
wjl9Dadf0qtY19dDgsrnO9z/6SHtBq4FMOv9M1EYCEXHcqSlAkT6z/sD2Ks67VcCfWXNi5GD1Jyq
gGeyzWzz2f+mZjdaCGUucUTup1gkCWbavbYuSx/gtJ/2MMaoQankVjBsxRF+X3PWy+OHHYlQO4zL
uNLHwy3vK+h5ZtCVAnww+YyjZWOASuacP5LpaCMY9nLTFJsO/sp54+MIq1D5Fo55IYeB0IxaPh1Q
vBW7o/HqhKmkeV224u9TOyjiulEOniIGZ9fcrMN+/iVzmGydt/tnVVgqWVcORMkczGvHdW1yI1D/
MznfScMzxNKCefNbK9MWe/M9NDtCntWGNpRoxcHBTHn2MKtismwgqQI/MadeitrzSNFEC3IMTYPK
UnBrCGDOfoCxUWlJGCs/4gy9uFzV2aCi2RnQs5nKxxUWuvNBBrTI0jSW3K9xoRimz9FZja51AjaM
HNKto00naIbxQabHqLdTAl2vAvwLJ9pG8GrqhseanrzPNtpASOyLQS5m3yDsZ39z2exT45Vmo3XE
oZN7BN+oNoSrcpv0tNIVB0V6ipJ4zHsknggPPyLVkoysiNaJqfUtzyaeFdsorivsvpI+wO4PSL/K
SLgbt89A51DH9ZobVhlp86QCKbKpX6ABz4HPhZUjr33yxES283PCoZydio+it3Wx2hTDrJvIudLp
rYPeGkMdESmf5Oa8pqWXelESSOC0tmZTKTv9hNiFb3ro7kqjLhuJ2iba4D3OKzENAyYMsFhDWX+Y
U0wlQCOepGCtkN/F3XqQtW10pm8t7mX72BrNvYFJPrKxtIsNTO3esBaNGVP4ThadlcPzPsKyqGt8
cfE6WhvfnEPBQyUT+0+K4hW2prCs3J5+2w0JsnnzQbqp0JdGA3AhEmJMM1s8TtHkVmLsrbBC+Izv
z9+bFs+v72I1yTc0XNXnA0OmB+0BAy9lvNDepYdbI32mPhLr326vDpJMgdWfY6dx6WnGzk9WfB3J
OMXG5c9dU+09XTwOHw8vMdazainIN18xVlOGjQL38lLndfd2AxezWHmfcgnmorTsXwel4N0tYXzR
kZFn2hTleyH5Ynr35WP3YMc8grE5UZb83di8kyB0SxVh02mxjx9HJ5zroNli/D1DL4LM+GOgtfTr
Mh7io958SDh29EniCyXbwLuXkv/zTUwrZEaGbzQO9xRToMC95THvQWzYtuhVNwz8iJ2MtXRmau0A
hu83q7ZIP0AGn6v+cgRiG3UytTjdclkDLcUi/W2Wix3CtXObyktyBdOmecS1nvzj6ZsOXxMjvj6C
RCrCLDaWMFmJMMJQjKYIpIO7A7V5kkoDxpmh5pnOXtOi6sQAeunJh7FckdThrrzHKgwl955gA8In
Cr8eBZHdkVC9Er7zo4FUZvISHTCY/CBtn/GkCLaNg4U1QuVkdN2EMQK4vztwHQpfNizduqlwpGXS
oCtr6Qcufol9ClWeggNMZBG7dcWo2uYTYgOW+A+YpUhAk/rs+UwVZUrLTxHlLWFLzKcJ53nk5a4u
Uy2sklRoUxqtctt7UiSxDrid6Q21N0/k59I5WH5ghJd768Qsiv5Vok9ux4o6fuw6umzWTOTrVlmt
UJ6p5WmwWy68TL+WwGnjGPPKPsSpZkoh2mQKf2+WI/mReIBrmqlgViwstNpir1QgJbY5qVpv312G
Q9vua1sVDPXDUgOk1KwY6ets5Nlp4n4kLRIOIuMnzIQWkTPdv2+6pkBWB+d+AQiKIfcZpooEg3CC
FQNBUdEyxqQQn14P+rzf9Bc4H3k4I2nIzyQHdrdZLPAfhtkfdxmhBSF2CoBwOhrq+dgGtNjgtFEx
P0Tqk8X0/4Ak9XRkeKUW3Ho0TBI2RcjpG31UW3ppWtVp9OE0zp07NrS6/T/fi/ncIaOZrdSFfXT9
JhAJEL/RPEX1FzXpxTyLzdn6vx7Ry8GjPeaEB+CjqOVH0oRJfqQdggfdpf6KywFdmT7H7Eb6MA/v
sTLIZaCnhD7hTlerbSIMFouaXCxDs7vIANUWeJ67315ne7YTsQY9xM4JquLtoCk6LrXxgkQz2er9
qb5OyX9wY4lROWr4FyS0pB3Hka6mtl1mwc5LvPHWWV2OeEg12axiGMYTbPDevKkvSDUxypLE+lIP
WtvyyEwXb815PtOfuswiXLP+wU/V01Pqd+Sj6ZjwWndidZExzY7Wow1qSnMzm8NaD8NFEP/7TYC0
vfwJo8O1qiJ2HIcIYVoFFMej0Ip9sINGHo0HDrtNCAJcNQkEHS+2eYIJnpCDWU0iex3Ca7bGzhnY
YLVegGmmw2MT8tkJwErqzvjg2yd/KloQcycIWPY0PzmtqsmHhTB2snY0zie596hIkZtSkL1rlZsI
5+uSw8Ah9N7+0J3EbEhvrjszOuji1wVroXbVZKf0QC988UHEnPxoHVAAE960Cn1PpG6JLbUdiTMl
eJzQIww4vb02psmQzuRCZTXiSNOoArLo7bcO5qu6IyTfulknHk/kf7k59KHoZId8+QyKiuqwzLq1
WKy7oHvFwkeNBsPSk9NjHxz8h8Xn2rH63drI0/ZhiH7jCGjfyFtU8oBtkLXFTo9UQte2fNL9iKKB
bET2fOuDWjEWnLPtDk7sPoGrPZB/2i54Ovf+fWhQn0U0o0ilSe5gdoRycvEsbgxY5iZPS+5t/pOQ
LSO2GzzvZer2NA3a2m1cauP7cE8Y+LutRNOP7jVHdXlOT7976EA/Fkvlbja/dXOjmnq/aVof/ECs
PQ0sKmop60QvuqK/Zs06IUyiPAQRjZgVJ+vytf743lxXYWgrmWjzEdbUuFrMs+IXCAVKGSPLUrmZ
zUd+NjPCq1EOOc87/BUsXiPc/ruLnkgmks4VaIzuZp4VLCkkeuUhHfBOVYRVOoDuTYGuzGGs5YKK
jnA8QBDZElpHQdp2ZEFgrfI4ubMe3PqB/o+qw1P/vtdJdwHr2JI5UrvfTspxy03HyINzjG/zrlz7
0q5h6KTzXuyFi28lxN9J3UrhGwVECJ6c6CKU/8eiKv4lGfYkFVzxhkahPF51nmlvTgWbdmB/sMdL
DB+tlIzITCcI/0nuJcVEkkVsLj+VyABWeK6JEQb4gOJKaQAGipRygSCyIsbdzKAf785d1RJgATKI
yviucsdUngRaD+aIOJXCXNEgMb/55wtronQXUtbHrrhzVg1ELQfKEfPaRUJDo2pSpk4DPIBFJavO
3uOnSTaGSHHREevsqY6/N5ZFro+3wqPFtduvet23DJ7xqxgGPshxRw+EkTkT1L8oo0LfTjDyz48l
2ilfc26NSGhmNOCVu+bTej6X9lC9TeYDGFxeX4w0qcGBU45XS/HJg5i14UAPwjnGbAFvsgDEWDWt
yvk4/FeyNlpUmRu578OKCTQnNCdP/vYpBWWyuAdQw5lE8C++27nmHMNQ25ECNSufWfA0rnYHcYz7
q0oplF9swDtZzxMJ2Wh4hcH2h47N6e4Kg+7iuov81bPXpmOZFZlAOf6DrYRfPPwID0QdYRZRPDvn
cpFJeL0O3Fn2TyQ7uX6qqLxSg6qrqEvXdxB8zXRBUvGnvX2O05u23gpxBdqOL+EI3QJZJxiIAj9o
d3R+XdFFZj1+pQwtvlcEQEqlv8emoMgQU0qoIYrr9MBAhqZMClrgpJpQrwOiOrDj3JgxnABt47Zu
VC+kkl/brH6IB+F73kTLsGSp9V/N4doOvg8PK53LnOr7EwoHgqBV5xNptuIBNCApVvw1mfw2Ov+n
cyZG3DzKOzopsdoOBs6RZFnN8HCCNfEgSf+eAdhahFNCTCYchXbW1rPAjjmWU+BiAbP1yllnAoFi
+00wIcdYVaUiwqn+XmMGSpw0fssKg14iLSn3w+eJXqFLpeley4FQWv6Z16MmgGHCeEc8dKlnmrKF
R4ZrHR8ogO40iWP+cSdbpm4SZRxpLTugwE13xXZTxdoO3F6g6F0WKk5za7Sg6rptcJHn1vZVHolI
CEWky1UcW5g9jpiTkZlWLPKcN4Q6dl/xzGTTuXvHEuwBfMtyclg043W+fa40321JOsPOA0mzHRRB
hQeyP3zFVh8+EFXCicPfirE2qTWHVUDKc3I6N2jB7xcxiEcdAfPZsLKYJPbKBtYq1sX40txW5ou6
wIl7S/uG6noikvHqq4yvViNPP+5OshfWQheQiZFqpZtIseHhxgmaHOQtpj+cuiUj9yep5P01vp/l
4+ZXKfZSI6fJ6smQNSwGD/rr4O5bB8ASKS1/wnbVnKFfdAXQwu9S8o03/zCxrZnu01ZAI039loq7
beqyUpTLi6PBDm3L2z6aXMKYC4fUF+8jWo1c/Kcb0kvAhEKuj4uP/T+embZCLyFWFU9fwMjegJaW
RXp9O25AT8FnnrCeH0AjiExmjZM/2yFKJOWGs+/bXNZ8Rrr8Kse/CN9udDcVFgWEXAxBA3M8pwP8
+eCbjqpjv+hLqSvUYT6ncTDilFUUifSBODdgk0UKk3WkinUkejY7eAnc1gybjHx1ORvI2yfRdoUE
RYYcSXacfgOMofPHpKVismb3M8ONvvVLtCVXMLEwEuwae8IUCYDWOWOaRVNornIVtQ+JHLDvfKmg
Ebjwsh84I7P4fR82+Xh8fWzegmnuIRGzKTZVZ/FBIo9/MBS/NB78BTcM6mYixJrhvUj257zHL7hk
GOhsMICCVOOSIuC+aVmJzS7gqxu7MGVdumToarj3e78r/Q++N+6Wre/gcJvg5n2GH/WbjTd1i9II
JhJ7MJWml7f5HGc2Z5j/xgpfkdt3JQJmg6yViySqW5n9VEZlnQjZRbyAzAaCiEHDpfelaHgUezvN
QGPe44JSPItINCXahderl02kkeq5KVyDQoA8W4HP/2QinI037sCCbUvXAuG+iWLYDIyuXMjtMJXU
R7ldvp8hJBxGWbnSc6R42D8jRwHyL1tecJs+++L01mQaIV+KiWgkWutvk2UUsVieyX8mzcE935bb
CKXcXGOb7rksN8Tm77oS6xpa3GYjFua1Fb2dhh3Y1hxNUhU7Ujq+UQAiBwlqcTgT5fbwadnjBean
BOVvgw3BpbxUMvxXcxaqaLzI5+e59oabBcMeOalFXyOP9XG4mLgKYgN3ALRWYml7YaRSMYhtICTD
wxplrNrq+CKCyS8qO8xHbRl7iIJdZlIEG8YWVyjBsiYjABUYU8aOsr/CmzgaHbdefSyid/jPKqk0
2eMy9STTLEGog/gDj971F59IiAwF71GY2DF4mD7Jwv4GKo+P5wdrG+CrZO9YN+ruO7O/8HM71C33
XeXJltEk++j5Ba3BLF5Fx68tyVSnLBie4RiCbPePu7f4Ul7A9xnykXu9Kg+sqAlzkjphjbCOBh/b
5/0j7xTuacNUDdeb6ZQPM3oDda+AFsl6WhfnUgSXV0vGUhTRk7NJkRangk9bkndNH6UXQNH3rFnT
pNcHg7TP6QAlIx1NQXXwIaDwNfs1HzLadZSybWjvU/Wc/rAjKA4ZWlFp5CB8oZhYFFskhbj4Q9op
ZGk5IJfcCA512FF9gGKF3prQRRYsB604bXF9AdCWtA/oheBxu87A9nIfW/YEjZ2iIY4R6aZyqs5T
xuZ0S960L4BU4FVB6QFnEFrIrblZLzVJQOlYqEuYAKi37M/czuLMMDGElR6f+DdsTQdDkZFmVJdL
ocxJDkZK7XW0q/hCPYUvMjn+HU1+QL+sXqjixB84bRGF9nZWNYsiiKK03Egee22lCH6LOWdueiuE
BRM1qC7QQU9Wh/DtiQSgEZJSw43vtbWE5NkjtVY+l7bKjb2RoIvkCG34zusj3/6MAZr9t9tSjfxK
P7UrOGuPk3UJ16PZvwUYxPKsDKuwiUZXm1bL9Zq6nAY3i7XrmZdVH61IKlZVOG77LCo7tpBum3Km
+NMgNkcm7VqPn6z58gBRrlkf9trE99r2UekmnggD6T6CuE/8gHudwbJtN+5exCtdfAR4douWadDr
lpunEoDelgukCUmrw8kvKU6Lu1Oi/mqwOIiQsVK5d2F5zMZZ6Ca3/qKxL0ax+v7UiMxv/9O5wV4G
yUc25vmhMWnEX8r63fAqHilavceQwwSG7jMkTazVVUUWFm512gPX4ssXCkN+XQGZV6zPvDLrqyAk
U+d4blxI27mKK3LNpRTDZ6iXVnhMzA7TU6baB7xBQvtGONGZEJrv7PMj3LmnDVhFI3FPdOD2pIMU
b8WVmBTenaqwh5LbnJgOUfABP2fwyuoy04fIw3YT5jT3isGAyRMH7wkGzIT+chOdsXXR6vRIEdEI
9N6oBg3icdRz2LUG0gyNs8aH/hniu7O8tAG6dS+CHZSYYq1WBxWJxJIb7PHurhO8qCphD9TLikp5
3qnBUMr9mW1CGhgwmUViChqphhlY5vqEnaUgKmQjIaWGaDz6oI4rpWozIhAzEDg3OO2Q4jhwKFaC
Ww3eVoBPTSWkYnv8bmhdY5XFE/rHNo4P/jau1WSRh1CYjlSwCv83BkIarJ57niRTG0Lhcd/p8+/f
Q+RG91uSmEGrW+I+ey8FLQkydS3XciPOY+10DNvfqC1t1w9Tkuh6TsmPF5hSgyM8xDiANCsBQxLh
J7iKcq7dxF2OeR6hyysy99x2WJF31xiSBJ7qJS84xsT/RXo1pKw+VL2kHI4FM8sDA7u9hlpiC3pr
2PSc3JGpj0sMrAyqh50oKUhHRRAtozks0U8o7Jhez2vX7L4D09JR8ygg0EhtxCCpnUNibZwby8Ej
AcEMzGq8agH4OMvGWVpmZlJPEedm50RHzawUtFJpu8nU41GZ+XiojWhuoljg+Bs19sfN12zG30sO
ezlDVS294Q18Mznwfns6bUyCinI2HSmGMJr4eUI6BO1SUoxXa0dzDmBQMXz4trlh94muAjxaghYg
ZeaeLC9CS4NmuHApY2HcY975stCfIgY4lRGRAj953cXTe3l9gjM7kqCDzuH81HcKKBq3owTIaIO9
z+EX2SxXuF+6SBes2Vn4ILo50f5e8EuBaaESsgzKIMHyP9X8xTVzN7tBD6tfhTyEF+kVP4Hi7u/4
7MbKVnJ/9uc18YlqPrj1yIyk7p67QSMHY4U4/T4wKfyORBwFRmz6ElFWKD9GDjOj8NGwVWqGh3Sn
C8tvLSsGALNItMEb8q32uNN4x+nk6+Kwpn06EDw/VDky3PTTWg4FWXjLYgqPrFBQQpzxJyNih/EW
jKbatE0ofPmdCkTGSUgZFvkl2XsaKjpjX+4aoEldiyAtKFa/5L6AAfJ1+pp/h83oVqEDzTZLMyoo
9QKfna1tSev4+9VP9AYuEozM/2gtmntD2Y73SEJmHWuSxkM7ii6hSTOSwMArvvOmi4xIAOnxza0r
CSiSnCoJOS/iI2D3wDgS52Rlks+ufptFr8MIua/BtQ2U29Spg1aSTpohgjGu0x06p3W8zwc0Pony
yudKOborOg1Vuqg66SznN4nC8R+uaBV8e4aDmOysACaZBeRFQcKQz4vt+bgWtFipnzQ6GXbp2tJB
y+1H8MMt5518ggiCjn25espNVNAqiL3ATpWaSdHoQajgKW9f/tlV2rwDGcoDDzusFw/LdcaJ1cF9
prLZTlNTAQSW3fIxoOKWk5+oF4g9lV06q3FNvZpBJgjutgKe5XkegXzsmrTU14tBZBebbuslXNfJ
oaA6sGMQ9ZB0WY+Vl1Mpw3TO5JYZxB78qvHMq4992w9m0kKnkKNnCdqxtvGVSpqQcZgY/jxQGAn/
A9fQRPPAwN5zWFsxeY26r6xDBj1RLS4tb3DWJN2PXU1Gp9SHlpA27PbV1Tn6/coay6VCiwd0uJgc
/M5l1qksnMjluIlzxp7nsHTzzcuCDTdDpvx5g+Sa1pY6s2aH33bcluTCHtKa+DfplPPePPS1fuM0
FlAavdagD1zvNyW66cUIcripzcA5BZvzoB7e5Wgl9v2fmvVscsJeYOSdcJzfTEdxV5G/Y5WbIjkb
Br+2eEo9QnXz+bSnSKw5SVN1eG79qvQeziH6trjqZlxSGYZYKsKP/h5z5bKQEDziPGMXRbEURD4O
WB1IvWvaSfyx2Wt8DoMRwdjTPATRffqZ9ZekIdznyFv+F3zSVMWcVfmL57mH1q2MK1yihJeftKVE
X6KeYLnnT8mX45HjcHR9LF3h7QGNA0m9Naufl8OfV0osr4lVu2xXf/oNs+SJWEFqB3GWVBP3cNVn
h9Dz+qXwri0cfQ3pwPtS6gXPsZ+sAl2wEMHPZkhb9xwFE8Y9ifZnnrxO36s/TENtT0yo7qyl8YXq
bdjZTPB6DwoaP51wqIf3BdO6TnZlUPx2Y3459eRjhPMQEF8EMp6u/DVWCGk4tNSq2JDw2jqR5oTE
GExjAr30MBLNBs1fSFywcQdCxA4U/XFVS0vyWPNzxA2e6kFX1OAlvBe0V6n+NgVR+NL5OGKckjPK
5VSBoEql5fGf+giXvglpLSiuphE/uegAAnCEl7llYqzKIzWJjXV7BiBLcRhFQS+tGluHAIQDMA88
cZrH8XM+1WcUZmbtTs9Gp4BbylOG4eIK+tSIIMB3sXlnDnk70eDnLKr45U8B+cmR2oH/6wVYqati
1vX0nL6okQnyEzhpKvPOrmpvf+LyMocSC96OY/B2udpw7FWbMxRVCuHQ0l4WHwT4FnrWVCrAJFso
n6rs1iMYcjwtcPfO41Fj7CWe26/9KdAKk/Noh+cWiBlsz/CyrBykH8fPwmrX5FBvSGWpFe9L5HTL
TOfasLPK6okEK456Wegql4a9ZupDO42gEjqWt5Cwb+GJxYzyme+alAv2nWp2ZmATUeDBTbtAnj7k
R/HR1nYV2VcjpPYxebgltb430v9KasBeugemG+Q72imquVH+2pN1UCx9vaVuhxpF0Yh4g1myrKcX
WuHmambnwu4aCBldowwkk4Oet8/katACEW9dgwo8rp4ylSPvnTubIXD784pNrDAWrO0lDrZXZ++K
NAx7doiUksXgB9jTrlNwgyXCOSTg7y+zKCXJ4JVliybxbrK8B3KCyWiTrxfyu/criUsPsk/Dg1MW
PuZn/wgV4vzmD1pusP+PTuYD/VUqMkalKIiO3/EMG6YZHidCZJprPItLzvHRagqLlnLrhNGpIzNk
14X6C0w6wSkXV6hi+UQL18KCWtGTouDwJ0mLgTWklyRrRa9jcwPdsPwBLEztPe72OgnpJ3a2I//y
vo7f8BnJ1NOzePL6GcBEwR/+2uKyVKOL1VXNLP2MInotA/AnBBhUdZrYJLTgjRxs6CpqVxTV1cUO
Ns+XJk5aFPbtAzRGwQDlmn2sxIegBNLPBPKPbPjqVY+xM53CAh/9+OGIpWH0S322aUQ+DR7vHZLI
CTW+siFavKP9C5KQoT6I9IeMFFGdohzv3E2e584Sc77sGXrZYvV/MYHrzReNe+rhRJa557SkIcU5
G9T4nzI7L1REPE2G8C50jxMTCZ7Lt+pYzDMbk2zQBQacJjkm7VkhLbzVLUBJ9rDVthbm4eeG6k/z
iSfwc0txHACaPfFz+36jNrYdkrcbyBG1NApk9vbt4bm1wa7bzvBQTqDLc9xt46ECajA9WJJQnVGE
dOtA0yWn1cqgiLSsGTI8IQNANnKOF67TEJNlh1udXCj+SFC74tmOgbjiaQzc4925acTYL76obHk4
rlfSLS1nlJXqqWyrEoDEIeQyVhohBgKM+85CDzyjSbADNCtsn/4KL186bjDnNDUNz3fOLju9+nFk
l6yZyvV+dA39lvLltYp5uZDCK/6H4DMHmr2EfJMnIWO9ZHg7ryxRCDxFeHW0exyslUQBb6IVr0q/
ZCDKWjsBZLm3YjtSM3u5iu3d+FZm2L0pft/7yebIFgEbdzlU5+cwVa+fofhB3BMcrVpKHZk35UBJ
8kz366a1fWn9w5hIxpGv8LTEZNizISFH12NACv63fk5yHG/EAoGMC0sqNsJMUiTQ9eNwu5wGpuxi
yekHcGYYmMwrB5mvofy32/5hI12wCN6BEvnm6LC+buc4JjKcnYXiKLzW/OO+QVFVQCEbiDEz+Dgv
m7N9qCc1UoNc9zPvLSNpsPWulGiyg/qd+JA5OnfLmKTzoAm469zv16Mzez1MjLpXpPEV4vOtQefh
YN1mIdC2krQ1pZbMPhwz1PZ2L424p+jYFYcPyhkyZeAdw6XxEVyMOCCxa3+xv4P0eBJUnX9hMEh3
6q5KbCuCLYoz0vwXWo+nDVs0YhlP9T15zYCliejbkQQAB7YO6Sxa5f0v+70SqNbO5R/5vweQw5pR
HeNSPZWz2eRsFX951K5SNZ1M0O9ggDZOj4wl4rXxG7r4h9WY2YjJixTMm7rffy4m6uvqnG4z7RW2
Js4fuFBMigOSUo6OxDfeAtHDS84PwMJL40I6DaFDG4O8JuaFcJjOlrXTvdS/Xt37ncjMN6cKMrnB
4H836ouUtR9euE7v6aX4erJDiQQfCD241inDDm8WSki1wmphLFs6G88jBLsH8SEHorGFfTiREx19
8FSG/1KpJg4Tqc99A808RtyrqLFh9686qh7herqcCG7/xXqXsu3kZMJzPXQeoOzmYihX3Uv9pTQs
8ZezKyiFTeaIDBlRGoV8ZNMnq8dVfp2cXzHUftzS/uROUHwwSzAJ0afCrTEG5XOX/B4XAftzCmJD
5/PeLRzZvoAVXAX4LWIpqY4e967EIz9ROtOFsd5XR07PuwqxFmIigGco6PZ63U3bc1QFDVyoLhST
cmZyVgHIJPUZERmoNg4UtFnnigiQMSiUya+kmtnXsQWXYAQHrNJ7Bpk7Iz0+4+pQ6c6Eo/HnGmdB
LCBrGGKRDQVeOT5lSVtiQop1c4IlJexMABPL+zkKE+71mJCqQEcrVWi950Ae35heFAib8sKqFZ7O
ArxBzfIA7jFccmlW+tc59BI5GKPCyCAL3wDS5cYFvW2NBBwkbiEKzFSDYE2zH17maL6lf6B5pnAn
qnCeFRLoVf1DZbDtuo7UJTdClDgswt5bGVKespozhKR0nYs4DjHRQZmXbvcfLFc4XoeOjNaL7344
yQQWC2C+aJhL8Ak+OpA08RvAomO7ZM/gTK4UC7fRXCqo20wq8nZZmB16JCnZuf4e3CG8VrFKBFXr
oZ2soLSCC5x2eVxErLW3YfIwLoeFvNBDZXItU8qBfeomx5ZDJcblCfLfqtjH0wbKtLg0KmhmF2to
BTDNZB2p18JgFP407uhXgk0JhAgXUI0gqsDBbz0WU1+kJxS4LCqo+w3FA9zhIThRJgciLGyg+Lb4
gv3q7r+tBWoY8inNK3OU1Q2wedtcICVgCJEV4P8J7Q9n+z1iAgKMWAjsg50TOEqILjB18tP+XdCO
6TVSdqlB0gjgsnn4It+f8hYYovZRdCzGyhxLtFeGrGZf204fdYQ7r4zbhc0CMS+ppSFrGvYATlsR
l8pU2XlMceHpY8rNVc98ww1YX9foiNp3ZrP+CulsUUtXtVEZNq6hhJXITwY2POQcjEfVQOCycnIx
IBeB03k62v+7YCerQsZTnBf3SU6BFAlAUrEM/bGINVE3TFcVDLjcyBuYZtm7RgMC0HakE7nP+MCr
nh9lJn+KHgIbSO113CMj5otytgj7AK5zKg/sr3+1zrj4GkmfdUjo0V+O+yNrd/TruSYm5vHRRcyN
RSs01TUk5BKCVcYcnrhCMg/kG+YFb165sPaXElFkWLXalhiDszyS4CklPrAIRk+ZCxoRORvX9iT8
S/AsKn/VMvIHDR2xwHRfKboKFhCl4mWrxQHwPdoBStb0wFLwzgodYPp+pnFbI0xfGLf+Umr1an/c
mzpk60VLjHtdapsWIL2o01GLEsiDz9Z9hMLQW/M4ezCsI2pferGRSL8ZOoIMZVAslfxAtbKX9s3N
NTvC8E0iKBh9HWFvGoo1himgwk6mq29mLgXIQQp0H2y+QdC66JjdI9dRtRz2jRHGbVSq9iks+PpV
7P9bGpvgRvQiXV3r8QY4RKgwBc4pGPMSPEQYlkMt4hxLMiwhuoxAPRpoSYVH16EkNvLU0oA7Z7Bv
xk8gnObs1qCnG+6qczYttfycZfH2QoCMixQgpm9LrO55rqstpNd8+B4erOQd9QYtyGQdgwqJGLTR
hbYAjWjVca3oq96QxGdv95dfWKpoXrbWCA/GrKUbvmBvQXFlC3NMIhb0bX9dEnOIVgLDL8DACaHu
zmJq7m9gXytupBYer+xJpV55MXekyJo3OMrF+FIX3PBcAQWSaV+LFTuTg2OSWynL7hci18KlE4ge
z7cByHkmlMFI0+ULacAjq9LAlYiII8ohKd2yye0g4QhnVIv8HzF/jWht6IBAaIL1Hwtp5dkuX3nV
CSa080H5sLdqIk4VqTCplcMTrnYV45e97jiyyWDJHzA3IWVp8LwFAsX9h6O1DRSwtHxCtDPT3btx
cYAxEB5k8dhy1e1ofMDam0jmqVxJQorFatlgUChWYvkMp6EajI2H7z/ymQFFi+WpLTX2vgEgmQMW
OB4OQRaSA3gc02r0KfpIpimtot11FpUe4VjXhgei/+pgOXRs3/wVe8GUnWYRBoSI+Eclci++Ahox
lY9I5KStPyZ88E+H92z8QEZrInje7DhJKZ+JHr3V6eTMoz1Q5GqB/gxxY5Bi/hhbfF0QL7R4Pp4p
aigmyduiRy0es9AE5iVoco1zfq5RHzXqxF8rgSZIdGizxpbpvmkkbh0Cv3FsDEP4+I08DcLeAOf8
7Qak2e0ttr5Gmwq8zBxKYDgYcxcH0KD7hUuMruJkzZswOKCoyo3AJ6TSNejna5SpVaGkqphk8rMS
GDLIH78dcoxynIkmF4TbkA9XIF5x5DKQsu9/ZztOVuP8mTHsG+c4BJVJvwOU1DixYzGs+PLa3ocg
r4g6VHj5XpDLZj3Mbw9YPm02Th07+JKgShppSgRD12M+9ne7zpnHG9uaLTxBmkFM3OWOY7SU2IHT
UR51F20h41aOpXpIo0E/48YCvo2RV0bdSKpTrE495+EYNSriVSB8Twf6dXsA86O58RFSmTq4IvkS
tXEzJSCaqyK671S4VjdZA6L/GFVm36RTxX4C7i3FTyefNSPF/bEGVl6rJAKQhkm8ae79FNlnshwC
LqU3etmeTHPSV/pLQsQ1Gs96U4gFdNlSem/mozK1oWHb25FkXfbXGHzrrlVRG57wAfbVNFhNrB5y
YTu59mPc7s5niI9ArwYI9wFhgC++Pqk9/KJYAR33lAgYc38YMWP+QSSFjjDwO0z6W83oGO2TAQo/
Ut8IVU7pgB9a6hh5rSvyRiL9JBzMzO9IKzHZwLhD5diHct2q2DJ+Dezo3tEcOCUpMokbsfgSLRXt
oVESTkedoU3QTHz6j4KKxvnr9Y/3a6XA6qHXaMTMYtwnMugzpkMvLqb/B098OvKs5bcLu+Oz/PqN
eVFz39SufR825Po4690UmzHjymVmofyUQpDdQODy4YMmoclucCDxSN46GGF9iTkAUA7ZGU5TJlg9
Xw6uYDmrIROs+yAp9KvMo5Tn2tyCdvDn+43ydmWWxEKEX9O4jASgjxMlehZktPlHYe4W0aeylCDm
asNxDrDKBGZX81ADwyZmFhcY6P7N41+I/SZugV0RtWmLpgUAxmTw9H0CEyY8SKff0WyG48Wnqo1/
5+Ip0jsZSJjN2Q22IsryM37Bj0dAFDm3182A14kxn/W63KmT6PW8RHwcSuV5DidFgwdhfXyqvVd6
JPukd0PAJojJ4PPqNHoZwAS76b0/OgUuquPvCk6/QfS0MtxilpaZMYoADYnb7CBLm//4BeCjvdf4
8RkQd0bDBvSXeGXjXzoX3ckpkFjR+YXtrvYlL0oqeT3Xdx0Mh1TOQgCjAf87wol9GU4EFpYYDAzg
ZBVajkvt665qP47G+kVM3cDVe9o+DotS7G1aae31q/SWhV8dbY+RcNGQyEv8E18n8VvLGRHIs4qo
4Vyf7Nopu4x6SrPwCiB8dvL0IwlY1+Z+3bDVVEdTQI+PP53wfvr1mg3g64I9g0bAFe4T9tgRNv37
uN8k8vlmPjLFrmtUmf5Bad1TnAmup1t+/LfSH81SPnkTgqMzQcSv5LaMrLtpS6OmI5/ksiF3A9UE
Gj1Uu58zcyRQyUnbedgh3DQ0CeWHEWZYGlsK6fFEtHxN/d62jJHmV9sZSTXNvlCxHWt0J8q455n8
PzIhAMtTQr3qGm0Z/MMJI1XVls8cd9PBneKDD7vr21UZfTxJjDLvxJ/DmW96XLOMS64iC70i5iRT
eFaFyfdwsTc6c8q1ECqKRTN5JlboJWPh/x6H/NKxAQcJe/uAbPXHdirnAUIQe+aO/LXiFD5ciarT
PT+T5wvAuKzprSifnugbI8zxf65wZO5THSSxr1kI5YGz/snGDqFDtbUO8bPlxVq2j0XgzekFSpu+
WulDj+EujtmuOQQ/7MocyvIZTt7qR6TegGpP9wz3yemT1+OizwjI0MkZ0o8zVn3Qfe8qM9knAQpg
73mTm8L0nTJvKQrRPL0hg+Xj2RRw72Dg1kHzr1BkaaKd1GqPm71wiBems3DFPenCyAocyysGxhgY
dwKTeD4Xt2PdVRKO+GUQHv0ssVu423Q3gNypY82rLk/MsVHPWKZaEiuSlK9mWlP9Rk6BR6tLMBCY
MP9IsVUrONOBhPN8cMTOVG84xKcArxMca9/MBaVDjKTWLviuCIJJYj87+OTOlji/41u19jFaVxdm
Nmbro5JQhAilKpdCnuTg6OAQ2z60vTcHgvwgRRmDDgre8MrCt7vEzl1IYLyW5IB5RJPWa+G42dKI
TApIk2BCQWGl/5A+Zspc5dH23CvvAvF21q/iG4geQpnrM/Eo2CxtKz8oGzIsn29TQji8Xh5fj3Ul
b6VkTRXUcU87yLFyDZzh0/72Brx+sBcGOqadOmzHjN88MLF7HP57rnz7JjCpYQoKBO66BVSlBvuO
znOLPt3i8yYUJMmnxehJXhjDKZGKzmWoDnZXMSJdwCNLkPvs6doQFj1Qre60NVq2and8OcEKB7fd
i8s/RsBZkwLhE82KMuSYAAhRf5dw3VzASqQjBqGo46Kuyhzm0epjtTE8M9ZBTdR7ik1e8lUX5f/A
wMfaOFRhKWFHbV31VHuCDkkhfCzPu8HSdcf5PkeCokyE93qZtH9yfFbQ0YvCFxm4urV2V779odjV
09yD9Kt05Va6Goi65Htfo5xlIaC/3UfrFDGCwrsc4P2/dNIq2V/TBQpZAa6yQpgGShmBrlsSB7wp
FrBQJatJq8N4f4Dbc/T3iUam31jUtPDmDhnlRwFey0nrJoQZ4S9nI5GoysD1ovuEEKUKFq/mWjK4
L/ttuSz/qXjqimM7lmUuj5YFQVBvd2ZUfTf5eIw6tIw1MA/SYuaeTj3ZiaUvBV7MAP6v50NJVeI0
0+oKekUu1J0LkkleLUmWWPxgIR9AbO7gNJeE0CuLlDtERHXDzczKZO4oBjh303TQxxrer6Xm92Cc
jCPC5SErWxzO0lGGqi+YkRHvXrm/jEqC3yacVSJ/g1gZw/Yn7NaqIv/mwcDcIain0+3CMyqW4EKM
AjPojeQc9+kpJcwy9ncz6hny52H5JzFHwE/gbz53UfjDmhbLeufdGIlHnViDEVFivgO0O94KDv/d
yTpxLV8T0IeaviJ1VA5Uybz8oO1MymDE4xjGEdIjNh9+IDX+TjpMHaUDaGwfXw/2W8kJY1nfZ1Oi
DZhpEgtWAxeddQ2zAJ6EXNymMHFE5299k/6YkgqGLQD130Aozn6xEiZAi8x0KM5rsSk+W2T46zrt
jkmxxhRZM4S2XRs8EDqRxHo5IXUzsTXy7aV/fL5k1uwGQwcBzs406zi7nT3/c41ItRM7flDg08yG
hgyC9f7w5V3M9XfIjJAkCaIRW0HEerwRG+BNLKGIIleWK0OAYBO+kuV+qvV5pVytULkTBVIaZf/X
BML/bU1Jc1PpsiztvNHeNhohQrtJ40Gpa5BqhuqdBw9F1YHnp7BkriTdn7q5907AbczSTJYssKsn
OlQERNuROlICheSY9ZrtJCseeCeeaZAyhAHTllC7nmxCK9ep+rounPodzw4yXYKd9SLc/tb7AW/v
3+K7cEkypzBAk23pTEn6cUiDMZgVEN4CrwW+zlhO2kT0QjQBNW3SetImIY0wXovQnkonCu03dUE0
6SUCrCK/rXaRLv8nrnrVw5XUzQQqpRUiViKQ5tRP7Gu9+33WXbHGaoeORL0fx0MXA85bHV3nWU2D
Hv+Hb8C9cML8gURGvMNSEnw5AQuxvK24i1YW8NVAVzF/2R5d/y9VxwWnwrurp4YrH4+7rWEbHCgQ
ytElNWhY+vtXD4aW2tVsT4xcOtsOACTw7os8o8HUdHzsFnX6DQbIaNSpcCoDavFHg2sskDRA+/Im
exXXox6QhWutMv+Lkt0Wec+uGbHdxC5yeao0txgbM7y3/jqrIsiDEk19L5yqSYt3xyPQoPy5ty0l
NIJzmqnpMIPyhGEfRUL1kwQolkn2D+PPnoHANBu7y57HPwDiK1/wjhFwMtpfeQx4wQA9ueFFRRHi
G2kAlUr6skVwVi27WHsMTJCTJpx0Lcw0OunO8DhKkYimlSAZ+EZlUJ60kQ6BkcX2zbi6s4J3IsHI
EZxPL1YoszPEOzUHNrhLfOkVLD0F4cN9D8i9/aty7ixICIfU+Qutu5M9ER3EC10Q2cgAOtvQlR/p
cf6WgoU9x5cx2Xdr4pNyavSZ6Cu8/mL6xaMbPT6Wub4PzgIPAaphiv3F2KvCGvEQsRr4Q9v6E0b2
S90bOpbgg0E8JjyKfFTsT2x+XyBTUkICSuwbeDL5i7oGaZaEwng2czU7co3DeiDS05hQEiWAzajl
riCAIZ27ivLZDD2O7D8XgBd0H4/WJNjVStLbbav+4eRi4SA5T10fDUZEVH1gGziUQxXYdCtey0xR
1hGMSkIG/7hAGWYSYLzF6ZX4vaGOPRZFM5yw1OYy49w9E2T7KGBzPZo22SADZsRZ9NA0aYNLUWzm
OVyyXRKX5JB7aNhm4XYGpQAd6QjPeLbMj92sxu8mrQXwMP2SZkMBXzOAkcOhSlniZVtF/Re1L3HT
Jh5l0GXzhZx6dQxL7bSTOnp1lYas6fzQQ5Me+qS179rJy8Pd/erO3w3BDeLTxbdgTNOf3DL3wC/3
8FZnbzJ0DjxMGBRJC7uKNmk0un44WSwi2kB17WSoLRibvihv7RQahKA2o5p/StVL8yYXicLDaau5
Xd5jdMe7di8axeHMk4YD7npBpkIvivvrjK3/9AFWBvbqFvZJ6eBcTL+J9gmOXRaJEzNo0Qrpx2b/
SjDQdhf4t5BRotYkg2HTWn2T3bh1PBDSCmIvBPJlzViLDsv7FVQyUYG/z8fZfgmt43MH2lquet5l
LRG1c+CRIJgNDdcMCAv6yRBcqu5w8ZVUtDdBFuttHAwVsuSi0IH/DJKSDPa6skM73CxWrl2E+bcp
xZfURgs4vtVxODDV0Drb7Hl4WTzJteNVP0+qL6uxfitcnZ31mGXQ12BRRyGrw/ZUco2lnzeAnLCq
qyJKHgiTSEL1gLRMhVf5vFanL+cJGJWlfJGE18ltL92cD2YvRtq0J25zOr30WxMyVXWwup+5sfD5
xuf5Qg/BOhJxSAvgBmsywYm94pH0yn/DVtWiFk6FkqTcmxqLPwWh7wN70eNh/vlxlZ0cyF9RiKRs
y5uqQGr7JLeQvSc/g/BqdBIR6bWZ6IXGs66QOjT1RL8EunHKiKk0pYlJt4ii7nczf9MuPNdA+128
t6HZ9Pg1YEndzFVTFkGFthhEcT85+mumlJ9/uQ8XaIxx3m3z0HfSNog/N9fAScHK/r64nciIuavF
6qxgcVnBkFsYe5cP/BvijOnQdokD5v+2WZ/GayzjjuCjkTrpDuaC0ovpT1wfOqOdncFNmT2Qsn/z
aPo+C8hBO/vQR95/49398b952RnewRLjXIReh+QdQpk/jtqRItIUo7am69j/MgcGqMmyrLZKzLLZ
Wb0oEKMVU4Bztbz6kckM9IG8cIhGdcx/DJWmRlu2oo1Nqd9u1IijDCaq0MS9Atk6oS7D3JABBiog
R9lNkC45sgis0DNajLJw4+HoAbacnfY3n6eppQ6ygUuL6fXo4HxAzSVO/MLg4/5RIN8urzdUsDoU
t/w/fiGvowO8T9TiFsGdAutVqELCgEmX/MRPRMYaKrmMGYb4awFLWm+JtEahwl0Rk7lk1fu9G+nw
HYg+dr177Guieis0+kL795RTIdeEF6zpxV7ZQnMAm5FcyU8gpfmKSIqVUNe2hhWB1BcQXCTFSW8r
xsk27loaZuJCAZ8yeynkVa9CIZEyasHK9wSk5tbY+2fSH+PG0Gr9jjjzh3tW0e9mcoSWsANlVPVZ
i1KiJ+A3M6+FaJ2AgvbiOfJuMo52jtaPERW1o96MAfFfrvFesaRs6HaeVR0a5WM/MIddcwbR5lrg
l4ReA5VomJtqENLoiR0cK7X2uJ/BWTJ/YkEwDrCn1dXEqq2v0gV5wNn6yS3y7rpJx3y1/uW/path
LaRk3vmtq6kIP7xgC7GkGHRKQxoi+H9rF5KP6r98h40CHFyz1pg7xnvz4FvxvWLHisRFWXCNHekr
e2CHm4UyRhtjDBr03917oLNaAAlQvUdHl2gN1XbSMnIfY7OidpS5KNz21xKhxhGSsXQZpfa4oTBd
tWWgQ8vQvBF4k8qpx+bySjxf/DkIPSa04kPy6Q8vxI1U3YD5PJaIF86RjCqPcrd2J5uGZ5JY934p
DsxdNBCchTzIfggd5tXE9I1gyP3GvLqDYYs+rHwHnNnTHOXfy6yVEyo8aYY+nNB3Y9DA0L0ph5fU
vFfgAnCILFIl1rpQRgUE+KzEZX7goeSL+5bFDsQ5nuoeNEP1vmE0LZg5R2jvOJabpLBsXMSQrgDG
wnnhC2f4nb0YI0o8xQeW/W1d4KSo5+tQDBbd7FeLad+1Cix3FJd055HrJCBLZgDPlpSZM+kMfjLQ
3+e/k4ITJg7gWQ4DxHhfHuYn5e+ugHbRmTegcW0tnbd4RF5tH0NV4BC9i8Scm0VfcjpD9IhtRdnM
bLUeOjXl0ZJM0Di1reme++r8iIvktWW7ppeCnAmcjpAcLlZ9huwMHs6syyuOO0W9f9ouekCOPPtw
VEPGLijxBLO2vrgGnA5MSGp+LAeA6B3KtgIyVxUSLXvW3KmWUi1Ye48R1rDRxF/k7AZnAcysKuQB
JUT2PfzBHdGBWJ1XvTSjtFxy937TX8wqiLlvsDvxxMUzKfolWF8plyf23KzCE53JKcqwP4WXV98Y
Ul7oXboStNr1cFIXC4mDJfez79INYTToy0XRQK5Va+w1nNGtnHpdM/pdMfqQr7vrq1KEXEp8fkIm
0owsK68uRl4jFuXyHUYZAeDLJLn02HRiX2KLkFbi/pBqtH0ZZt9nOLCoAMQDZKxfLY2Uj+MNnmct
lNa5krqhtX9Mmf97sv/i3Si+gjWOR9GF6cTnvJgEhSLjjqXSALZbGAjTIcq5vQ7tzHjAnxbY7/6Q
EaZRejTwKezq9Dkmse/Wzizx+z+NhKX8HtmIcGnl4pF47a/yBET9XmuDTXJy5VdOTZdaRa1qrKTN
nC8dRZthK1aCDyTm9wQNcD/svtClRtrwYum6FAdSDTJ9/RoDY6tozKsw+mD+bhZctkmbHF7jhUHb
2CPzWHLlUpyM3cEBGYkJVLSi33dozeRe3Q7qV3IbqcdpLgw2qyniA6NTB7BAd1Uro1lwI0ayiUaM
xvKghEa9K8+Kc0uuCf+/yjgxjdhmpp9oRkuHV2OhgCfH6WqsoGG+n1oJdehsVTLJzbyHpPJj8Tco
eZNlnmMfshTL/GTSPD+YUFClmv5iOIPfn54YdRURzzcl4vLwNZIgT9Epr7Zct+b+7gUMadaLGbmM
UwGfTjKAPecDM2nm2C5wuwS0lY0qkKO9CdbbYQtHWKurn3UleC8h8T9WVEhUTfUifvriDULyZGIN
bSST3VRSMqmFa9GghhjN/laGvZaMvCDxwrWZb6odXMpcFKdccW3yDsBnnU5e4r2EDj6O6kv8DiJi
ZXGP6uCibqP04kBuNLDbo0frqt61/o63dJXoNKv+SGikgg8KgwfvLUZvhu+x6si2ycvzH/hMGDJi
0yr84d+a5DOPqy4TRsXzlGtqii5tf42twPraKIKZxyUHSjDZKssEUKOxEzLtYLva1cHPGxnUIL7o
/DvAjCHCR05+wKZYde/01ul4faZxS841Mw0DwWW/sA+j8LaZmTLJxD0yP4+t2z6YEKQeLmStsv2S
9KZr6zuRxFIH3ZHujiQPh3LkDm5rd4zuWv5RWGsiX4ipsVt7JKE743eo7IJ9/BtRYHbyDdj4Atza
g9qCDkkWTfRZyhO/s/6lyIsFv5yVpbPvrkdfn0F8SzpgZUkv18D3jTk6IoV+mYlbKBYDhLj4+DS+
z4+9OT6wzoyQ9UNIWMEJ6/yDyEpIawCblNQN5dN/g0ksqaZSApdg7L5DTuxTvoCU68J53aRGfESM
Gc+kx5pTJMabFrhZov78Vv0VTkLLJcZCOvXQzvSFqVJ0kmBlZi2qe/+bkDnlGnqLtBEfUPuTyBDX
GSNu+s63ub2cyeBAhfp1+WowbjK4nm4k62UDKQR8AnPKhZ8HbfTaIJI7pyGmp9X+RThWvYuylJBB
gFVGEjn1mHNj+v84Kel3faXYtlR9JyX32eZmXaU2e0BlMDVnnKpBUBH8oODKxo+1HQ59kE8a/9zN
FcHM5pJcu+nRjqhlrjmK3AGlzJC/QSHru+3xrXbrCUkVyphdH1eCawYxpiMxiXfyX0No+oeQRmiy
7P30zEyRrz+wQfy3XliL8IQO3iebV975A9MHiQiRBO8uPzvFf/a7IIy8bKuDNA/e/ImVHPD8kfYu
srrIADF9IrlODBrFx3jLbF1zuabhzTvo4NO0fu574jmchsAgpQH8dpew8gZBt0vhE/fp0h6Odwlb
r1XS4kDFlKTNFHn8d7hkuBZjsEomz0xAfQ00SuEAQHe8KjDpWRlaKDghNTnIusNOhVc1VEqLeRb8
p8w3lMbEiIyd1nxp+DSFkGb+B5Txa5W/bYtQ/qUTliNeQl8uvBcvp/+FtnfdN45aXd4JvR2tnRJ+
oeiLDH1sUi14EyblcfAmsiu/uL2qjUshay45UA4SklMQaWpGfFf/ic9W8Fqn2x+IuMAogk9IanQB
KHZzNgBHXvt1gtSaMuUYwIq6bIEqlON7lJ/zd2qpYM9ttE6g+Xnw2C5WKVecJXwjWcQgzNk2HRXr
+2tAvF79PfnD6M2sDM8jc81e+HdusqJ59eh4IRlhTW3Y17tc6BsZbrmNkApUDrNOxyzBV+6+pa80
kKNIgbjHusRZhcqOynvznmw0Uel4eQXBV4TAhyiLisW0RKM/1a+UULtDebo/7urFFPJJNyHiMKs5
8QHBqPZH6J45eJk51ucpbIi2QsVkOEQkPp2wgVfJibBbX2qcH3RzaBccOYp37oHafNKXu0IO5uU8
TA9JPBOl+l4GgqWa6blRLsh/H1ULSwRNU6E4l2hjXmtSxdeVzGWqbfabsUHoih9acHxCpuLrFXNj
YqJebB6w1L9GvQZFR44Mv+ZE57WuIm+PdEjU2JMey10L2OWAJNiGZlvZydvajSPOBLgf64SEaeSo
/v8oqqEDryga5j+x57RBg6xicrxHqRAG/kGkTmkddathh8zuvT/8akwN6+4vmG/kUNFd1IUBKQb1
NVf2dpiHsM7w6Oc0zrXEDtP581Lvu56aJGlacNabMNgVQI5mq3mjHCS1VABFOGDXmZ00GSf36LK3
Gw8CN3rRKqH46PWCSAzwSDk+ZIQLNNikWf1P5CW+bGcAaaryZL1MSqazCZqM4Md6z1o+UGdj12Du
YZDLBiJrg248KJrhbac1fJ28NbUx+cAXKL7tZRASYFvw09S/6pBG6owQ34Pc3lWKzA5zfv2zXdMz
ZxRkM9JwivfYx8VDpsUAq7FXP/YrtYthJ5Va/NYqRZNEchgsZFqnZrT1OoEKFyyNlHkw5gvvggv6
1bAHbYX1BWo8p3I4JExNi2vv7+b6FiKUkq6iR5q0RhELi6QWRgBg8CiZM2TgvFZ5Sn9CmB9jDWYg
pxtyjB7y6MnCyiXZ4lCHmIb4d+sXot+JASSDw4/Gevs9Vn1qDB2TdbO5/UMknPt7S2Ny1OJrRyjT
BzBFzIyMQ/tYEWZjF+f71xYHkOGpTJS+1UD3jNL/NDl81OhukStnrGeh8DIcxNXEiTqOFUSN36i4
j4zxkjpSTSI/KH/HposjQnIITMwhFvNR2HHDz8UhV2RyjVQ4tZkfoACUKstXODXgXFVFl5xGgETR
DiudXjI1roT7X5aud3bCVAKo1ey/BY9v2Xj2GdwzgMIG+dS6+5hoXVSzPiXTAJblf0KKMG7BFpIc
jS//pHyy9fW4FtbCiopTFsl6IQVzliJQ1djp0sCocPPasus/A0QXhWZUYWkqXlZ+VJVFTmIndIOY
2zwEAm45XBxXr0aHFGviN6C+RlPs9GLcE7Ig79HhfigQFEZRR86lL6e1KkTzJtdbXxw5VfnHaRzZ
xjDxm6P6qXkKg60/suGNhp/+TvFud+fWf6KOvyEfS1TTKgQ35Y5C9gkpmaasSdqzCr52FpKJVxe8
0IY+mJ2AjUx4K8n7KzvMFmlL81Hdy+b7eEkJVyx09gTzdjHrc3xVTANAgu39N8JkgAOdfzRIZI0z
wWy6b2dAi78/8BxHNHs/YpEh6rOzxMs1dmeWRsis8HcI1yyrKKd29R6gm4ek3MqWNk77kmJjuWeA
2TOd4EziDANxrGPQOiviJhzUAb4m5g26BbjsRLVNltTuARBAiNdZt0TnyRvmYeeRCNNm5bFeAlBb
rBXj7lAxaIZY1/iPWGdISUORdGLGRwVwiC6ztVm/L7adDheEub2Mbs1n8cyAcI9fZ0qFSgBTNNhg
dl8/tHm2VVGHDho8hCrWUCWXSte3MdYi6Ya/48PRlXiMfj9DWT9CjIq5alwbBM0Vvt8ddDz2odqJ
MLDMHiOunyDI20KwqTypH23XVYsyv7maMhc63vhD6S2otaofFiZ3fwiJUyxyGwAF1sJ7NlrSgVNf
T4oxrjT8e2hLABrK01mQk3tTH6Vvh1/a6JnptIfy6NQwh2j1rDbCT8vZzRZCUBQfY/AhxkO0oXzc
Mv6Lx+RSAB/yWvBi6e/JDtjPtos9eKGoFJiy7odbB4U5KRIIxed/nyDpvshv7OT/T9lk4BWRIAQU
5nk6kGpP13bcpN0nUvcCcQsUDtkWLhJamKFc2+h3ydgwDE5AJt328FyGMNkYlGoNsOc75SyhAuDG
46j/5N6Liw4JDshEBVPdnx4b9GB2MGxOm9Y2XVweZ8i1KWcuoKDs6E59tQU5FW6CfoilrhOagpCs
UCUtpLQJm90cCe41z+hs3mdIfCU6DN47yEJDnlO6LdzrtmjJyadorjo746CZyq+jsU3y8UObIIBg
RqXm58xWQocUCdargXgqoKujNHkvx1xP2rANy6UPtcvvpl5y7eznBN5H4/Mx3GSygc2XxY9/btkI
m7FpP1BitujkqM3L6xnWDaSTF3AEhQLDt5Fe6UHKOFAgbE+kkwxWO+ZYsbgS/CrYpAdXZY23Yx2J
+QAfvwxiWvQE+gQB71/SMnHqUieDcC1oFMgOH0bvdfPk/B5+AwNszoI4tzp/ivMAW1IuDcDo4Z5W
k3kxX9OCrDyDg2kJ5hsIWwRwEZqz6ldAfs/PIBa2/LwPah5+K0gWFk+t3/tmIEfHBzmg6QaB1VvQ
AJf1t1+2r09FMbZ5sjjqJD0IqNUH9JX/4aLWUiTPir4uO2cUrmnXLJoTDMncO/U7wcaAqQhxAzXw
wsysYHLNwyQPYPTkSfgpTMshpAm6z+gmPs8tyj85fF3Zggh51mD48K+jDQtQ12iPcdjq8Gh0Sj6Y
oRcVx39V82utiMV+Rp3Txph4bQKOxSX2FUqdi0DCikI+SZbTDYAoQqoUjIPBqoHCUC925kEN6jrC
as6bEuARgCIQItYTKnax4lgsXNnbtpe5Q/V6kAjYhRJyDwXFgeZIP4pcdujaieLvXSH0KHrmUyh+
qkdoPf1ufSd7pORzzkcOJX5u0JY1vxbC9tQgpx72XLcXCwN9woMx/PQwO0zbMwti6fRT8kIL9cqH
j29ztXMUNEId4vYiF2oujm7LRMmUuF5pv2r+odFmxQ6828zTFvUJzu1fQrnmpvn2ZSAZzMq2O0Gg
Fr/Losx+ePVw9XfzwiciVbnLbnJfuaBYdfz3EfnXhETv918oRps7/9Yv1nS2GHqq1VfC6+B0uTzC
TWLfeKQTdRUuy4oKR36GhnoMWA+nVCardBnnPumcRtyRyb+9U9LyR7UVvaO02EGZyLhPiwLgd92n
/rgmiIKygaDBClw0viqAzBiuoZfWMgdcmB3LUcUhVmZ9SnxS1Yql1YvMZiBK38kV08ZOKDADG+N4
4JDWMAUWZQWrz2KTDZe68iaeXCE/g+neuqRHVwUR+CnjU1SfEej5oJ5o/z5girYHdsyCwWyfx3Vd
A5r0uhAa4O3V/a/JJ5IEfLkHh2uu0soA6ZKMon3hgmyaRGZY1UIndZ8rM8sVQBH/cwkvYs2RR6+6
sza/WWFpGbR2fED/L1C+wKtzVP3QTG3vlALkYH38GvOJlWiews/9YQg1T62JhMxwYGS9mu5BKvw+
s8xxGmHFcKPROWUrOAuyur+0P+mnKD4f8HgTfXCbSMlIW9qRGHtD+OtDuChoaNk/iQt5WxguiN9f
3OHJieeYtchTx4TIU4uzrZn1CAH0df9pLawDvVnShGXF5uC3OPJ1feIc9LNRlpV5O2ATvTW8QdHZ
vxIz9Gjh0+b2eyZjp6IuJx6EFrenqfsF9WLcKJGnReamck+FShbdvYa7T0ysIhGI8NeWe11H+M8O
R01TygQhk+iR0zfcziOCiOiooS3KJjhLzj+LjF1Nco19lcfzauAENDDUz4mYid2gNPYsFbxgHtty
9uPpCatGMFAjKKA2olrfcynQ9HeMmY/P4MwoFgqlar3N5He3iVPQxyoovdxAMaSwfDY754XTm/35
1m0vB7pxBKJhv89VVGB6qFEC5tceErQ3e4wB1BaofBCn1IG0TqU2XBYrQYeExAXmg9SeypjRVm3B
pVzOTRxWYm2AZt1immL1VmK7xocuegqV3+ecknqgvFc4Ix40RCYRYBXaL7BcyBuxmSNtYNwQAP04
2O7L3BpY3nbMae5GbdAZ2Sob32dD9JTiEkbzFHqU7uwTAF3sDbZGLtboKvpF364seCcP0rBxowuJ
2SxT7nfmp+Jj7SnbMCMc3Hqrd/FF7MOlPGH/EOzpKAfyGob9s8kDD9f4+PwASUY8J482MJDgMGf7
sl0WEa4VwQjES6qX2JltVsxIjg6Tq1q4xNqDiBrdbp6dZUNssQTUtQG1qayGKdFz0LBueaJ2FZZX
MIunNSSMsx2Xjdk3mB1EWIc5iQIlgSkE6WU3M7T1nQ/o8k+vJa152FQ4idQCG6yc4gdLb20ERO0k
wtOa9b4A59kaHXBTau3pJ2OxjkiW7/wX/RE8YGj2Bj8iXJeB1CTknj9uRVGSQtSCIDhkBtvekCKB
8YH/9pLRBccaaazBreRJidardka4fHzHW0ZcwPCNeHbqQA7M2LwIoNwyxDf0/HrtKyyVFPk2yRjN
wOj+YWCjPGUY5/cbih0WTmAeWPhFK4mqJXVfJlN00+y28aNaDjtcVrl0SSpq2EkeqbXRwEbWBUSQ
OzfLiVBlPOjRx9E3KTtdSgHoF43nu5JjVkWK8U/1DCPlJ+YvpAiVEEjCC29m5i/h8rPEGwkR70Rd
hP7F75UnbD0KctqBBkXH3MnJp34YdJSBBo/6kq6rIgeRSUnvzFkbmGAHWtC0yQQwV+un7CNX6Wv+
Nt0ZCnY8j5QLIc4WF2cGG81OW5aK2xq/DylL7SIH1lL8eLq2i6LfC/v+HAZVcPPo/akRNz4hCQdn
B+Gubt8V793S7U5MWyKm5P9vnJRWufzJ8LYE+LE0yqlklb5H3sHrxK7CFLEBLf1x4jCN4NNJfsTC
BRCbY1ae2uSpd3wAbq6qbQ4vx5R8XxXCwc04CHySEkgBtnSRqf3YWsHjM1nrb2tKXIgksl5SatB7
x1LurHpGPmYVhfsW/4yHfW8F7Lx/xo3XI1L/lXLHMF+MIXeEgaHhAd3zU6U/YE/UYY202fqlPBNM
uLw6asYBxlmJf1RuKC+oL/z55q1ifncbwomMsAPuOSjMEQWELHZWRkBl91o0nmRqfqGt0q/sf4l7
BMUDN8mH57JvK3xu0ddH3BewYwoOakcW4BaO9k1V45iK5n7Js/kcLb3rP3mWpwTnfLvID/y+nA3+
OnIqykiTdG94XIab/HhikBOLRZrOdDKxUXBqMKlsy5Hdx+BjEq1ivSicluVPYAlwsMWdR7OX0iMg
UrC74PG2S8W3klIMQ/eBiiuOfdXHgIunivkPU3C7/IaKY0gqov4k5D5n93HBZRl1qWXmi1LWrYoH
49uG4mI1wBvkcwe5531Zonq9M5uWhq7IBqGm5RnYaTeJREAzOaZH15vGVrs7khYJSABSje5gnAKl
Lt+v1RlE32LW0hKkDIOJbwLwOYDCl0y3s1p6yOMm8f7u081lAWbiiVsdcaFRnBskA/ACElRuwuSq
SkmDHn7AjkMw/CqQjSAEEM5YdjNKnTT9bBlGN2oJdlndWoIp9VU42Gpez/6rZVc000lIRbamjMNZ
VVzZKpiX0TV3TPXCVcq9ugQeoAr6thZzOo+vaTaApwd+5fmrVW7O3QvjDEONkalvHNoQ+bcbnBC6
z6J9WdTOu7IC8aCCyluD59NsVU7i3Pq3eEgcMHaOYejiMsmg+CZQ35lZHnIVifQzJvqte386SvyM
7Qi1+ig7TW+Jj39H8bhTPfQcSSRBL2JMNaFnzgytgevmjYRp60N6hLojPIdqguqA2M8PHdbsEqYS
rvPcfqG73jGrdnXTl96dy6EB69Abuv/okVfaY9wIXTdbRUVyS1sK8bV8HghfvkAW0yDkbP2gtr85
K9Nde4n2UTu01K4Vle4711A0OTRo2CnAb9JMmqMG7tTPf/eH+xR8sDg9AFBMroolR295FQgRlW7Y
MO8AslGMI4S4xPgUsGOpFMrZL428XtP4Nw70KrxnuGwFJjIJwPqRSYJC6lq2/rp50/C5F0cb6WHQ
XFrjJ83Pd23j4GRiZsporiyWen6jwCYDle8MhoGqmJnBrwEXQfeUTTn8/PrTdI5G7KQT4ZxhRv3c
RJ4QkEu9itxi5Fnjs6zOoFF1jr4eGaZPDogar9DWGDoAknl2YowsWODJtt5H2ymQEuHqkL2/pRFv
TvoRuErA2lfxSV8qRpEljFhOypUCIAqXYsbK2oNgwVonRaI8G5yzvsz4g1L4cSzf3Wk75ST15SQU
ySs1ocAQvv6wT4EQ6WR/oiOlkI49Kes2dmlevVGm6pru1yVsdhLdiN8B0cr4tay0F9S4n89Rd2xd
NMdR6LAWuV6tLMNYoh57Z5Uc04fIYNXPi5aHoNcujx6PUGjyeloUpIcHH+PKt7IkEWqICy8a5z8t
N/sZVOdIydHWURjrTsEBGsG9CZPeIl8yQypkM4nj1XmstNWDwHxpbtyEHHaTHHV1CwKhElv/upqf
rut1Ytsiif23KNU+xieG9aJOZlk86D/1IUdMPbmiWM3GxqWkU/cuKVdPvPRG3YDl5Yxcg1EHLN83
ucC2/xiXkxnlgwBWaZCZrcKcG4ky46BMSvomRoIm85Mcwzm9QiRYMUjz3Go+RoVOBbeFdiIG2U7F
T9KgyrJt4O92I8BeNNkmMfIS65dsztGhq3CIQAQStYh9ckydR9bFrilC+iJOoBD8r8MHauKtltux
ESXTpIieBzYG5N7frcECMBU+nTsOl2pIzEW2v1E3IoasFQDcAWgqqOlkxznDQ75eNkkDKO8UIGS4
LI1i6If8mlf57LzTxbtS++g5x0jTpuvRJQysqtEl1rP+LTOMdGDC5SLu2miHfjpA0Y+hXJ8uX6cU
PGg1ANvRcrXZmo6loW5GMGawAHm8rmq48t0GHfGO5gn27KCRBoiANOtI5HA0b8LgW9ObI7d3QycK
EvwvKKeI9OsQYgpSa3V4dy8lhDUdHSQwiz7C+IOMsSMskccwoI9LXWPzbbzLvSVI5t4t6eY2sKiI
bE33By22Pve4PfRRz7XK5tpvwa7iJQboUdkDxEeW83q9jrETLkV6mjf8AK1iPuvtRlxzbmSM6Zao
kShd5bi2QVJG37GlfmVoWyQXm3zmzOTB+DfE9uLrnoSmFwUyXy40oZyxe01UfItPB0Fj08I9Fm4i
Fp/qWHYx9H5lbLbyg4IeM3F2FjGAeT1y+vKuoUdlfbA8skPxKxGUB3Sc8h7YVE0yXMNOzEHHkJFm
0xRbcDRJMdjdt5DPF1em63RUDv/hQHQKSeeG1EGaBGn2vrhAWvRirL0Y0UuDKbTs64srzSZO/oHF
b5N3cf3ECNTY5EemBqNLw4PQZfVgsb+XMH0kTGS7H2BOdTVZGuNpng/Bye5ZFLnBrxigO6ElU2Np
3bBep621KCFif+mARJ5d6B38O0HKDQ6ihPG4ojsVUIPfwWUOAdlYuTfp+vNx3PV1YqMcr8QVo9B5
G5XGU6VfCUFg+0l/r2AKRnYV9lOC/snoV1A+WhYY4xxjdWKGMzUZHKfkbIjrD5DrP168EAVwPzKG
4BYZ8tZeWCGiwdMJ1R1CjYPTRNEmbiy3vQ1HZScMeslO31Aa2LKLg9PBNkWqMic9QGlEdQB8230I
Mdyt/LiuUEMVTme3EYaTcC1Mu5dqSMcW10Kdsstm/EYag8hRs3vEA0Sq/+v1/0xKxW1woysplPCe
4ghf0W6W1SlUvRAvO7AMhYajdzZq0zf4uxk3YEnQPDr4hP+x83muz6XFrfPI1dkNOFDUCLjrlkgz
S4URM3FYY9gf6/qho3xABqTaHpJT9b5V9ENwIxZZKHiYEWvLX7TiKxdU52zuh4nFioDhhnuFT8yk
f467Arjm6StoycDX6sEtywO3nToDjxj41FJ4Csbwu0gw5tPi1nmlzKNRYLwuahPkEwe7NTNOs0EJ
+2g/e8/Ap2Tb7JvSGWt1zNHCVVV2ZCK1CAOkhmRJYsN6rDiX1yuH3ZkRky/KwhcgCtTPsAfvNvj1
F3J64j/5oEOEzQZM4mE3z3QuJ2R7lVn0JKQ32qAzPuRDt7eb+yEw/xjUQbv7KdcNJy+Q03jESsE8
7bowA7syGfdjgbKo+IV02pxeEsX6gBuCPkw3jkQpVahYbackn10wQChaG6S5IaDDepSU0yoVl76y
d4fUhmAtUuc8aCyhzVxkBPxK7ZW/g1/PfWDV50hN8YfzkwTH8OHeXqMVrqeg0y35dGAvncCnp6nE
lKEaUCxcOJiKh8Iq9MENo0/z1LUDOL49AcwWMHY1NE7A6rO6td8Viiqn6EeWg5H07uZOyrZypIp/
215RgvhARTc7a8MklcDUw2EtbSeNodtdlSeXtF1pDQ0U9G8+zwgijrt7V2y3s4s2wUlpBNsZpdk5
n+QsmcjZQoWooG810VjMkSqxkEgli7z7cTv2a9wL4vi1IqS8Y64waVlKRUygS+NHV83VJ+X3PCDM
NlD9Bx1Wtl6uhWyEdGB3gOu2Zy8rpnYhKKoEB5JV9SUuEpyoPCe1hEJOdj/YBJnZPvByqquiEgIj
B8c6fz97l5OwanPIOjajzhemcIa6nsNWyt1vaYujS6biKYyWP5PPiRNui7bUWwHHTr5euNkpKRRe
ADkqsJtJRwAz31SBwZcY6W2sN1ixc7ETxdyrIRWpSY+Kvq+K9AOPeqfFgyHYiqAgp0pzIRaMN3kZ
iaCcIxs7sQHW1JKpKVJfa1Kp6H5IZG9cA5ew/mChkkZsmR5Z0uO3uLxHLGX86pYwIJD1f1sBV+Vc
a6i7/FFInzCAG0GgrQnhQL+X4SEzsqeMrqVEoAXggH5YxQfC49jmeU8KueFPtlfig7KH+DFZNAsz
uEOBnv7b3tfTOcqrSEg03KAQuwuM2gXSaa2vf7PloB0xILQ/zpGBbJKnaYASHkY8HIWfBxp2Ysgz
3yUkyEd1NmaiPi6zC4KzxyDKxv9AgQW4CYDO6zxSWbeMOau2UgJVP9Dc7uC33Vy+Rj+m08z466aC
yK02CY3z4/Ui2Ml6A37qc9zSCAM1EdQDtHDdG0f1ofB1rSXSgmGoJNalSWrbSNcRUpFRt7Iw3f7W
CXU/wFQ5ckxWnXhr9MpGI7lgfarRCGP/ZT9zUS5+xAx2490LXD+TqMcWQdJ6Asst7ZjfkLnWG7BC
pDCq6uBlZJS+6HuqFqP8/CEvA9EXxjhBDqWWCRd7tddj62UoJ7DCoWc+zDonalXpLh2HHIGWEOYt
VFZDsbSlTpwXvGlVBLxEyCKS9MeU9JmBokTXQK/fQshm/0z2jkYFYLAymTnls2sF0oa5IRLVx7TB
bZzALIEYBKABeqWPrGXFe2k40XvcfD9Jkd84L53Z4wl9HKu9jj+R6gjKYPHYY9U4jIEol5pRtQyf
e2Z9kTvTgTR5XxO0Mhd6Um/vWjbrzhaAD4IPwk9UVyjgIozhnQRmQLVXE524fkD3d3r6jVfic/4q
6btjq5hRXV73ggn/H50pM2Le1mkZj0ych97BcBHiGIzt89XoFVxR3p9n9jRqAi1bucR9AsJYttcL
TrnpP9XGDAdGOSFzHw1LxoYheos3LUvGKFFKekX9AoCPC81ttJzu/sTfWA/82JrcHcP9nDQ0LApX
jgWiXoro99jtzvPapzve5ImL4ftp/4dAgjG4kgIL07f4VNGEuo9Huk94V3JFwab8JcJfHwHTTpwv
+MX+VNTqRAWZPdOOHHxy680KALxs9Jqu8RMnTFPMzw74MBSufQXlV7zRrr6gZIaFGihpapoEAzhD
7G1/KGg2BSso8A9/uVCpNba77MzKeUBdRUp83UAHnXiQ/Rc3B5iCf5jyYhMcaBXYmOSXiuYY2hSb
u27xSyoAP53mJdiJUREq4V0cBjU+itxK6QCfU42/So/yk6k/7To5Cjhl3Ss0Sd6v2e/SBwJ84RjH
Rt1jgfwpVPG1CAaUHPB4sikBfkdTveQbxH0dZ/Ra35nsCmqEQD1OYQ0oBzXVD7CuQIB+C/aHUOcY
QumR+yZOAb73XkVmwdMSdOevYyFTbqlkK3gDgF0bChPZSVkEwFA+nPoVoAo1kyIlVnMFBcvDi8WK
y+sVUcT7gHxUZYnwfzkBS4ELjT9nkm9gs5AP29pY6vMJDJlLl4Xj+IO37bJYMXMmkmO+aZRAvZWR
S+ZXesTd3ITHV+DTIHGxByQTdwk+mKi8yFjvYO2hUAg9rEk8PwWTsBMfITKNyY3z2uXn/7gWdViM
/9tqtQSCQnL775rzZZcdhy7mlOTAPLMt7kt1gUOynhMK9WYKpmfYpNzk3Wh0XF4HP/fUq6R21QXo
GXZXXkf92FlHPJNYQkYiQy+/O1UZf9eA4974JwMklLeZjMi3H65PJCv2OOalZg9p08nuwr+rjgOd
6wY3GmPqJ9QLU2sxs/PERdyVHUML60IikigUF8KniGaZP9trO2VDAskekoPM9Oy7yXGpCkVTYono
406bt06++5nPO4kbH2JZRu8sFkMEpkcYgRCPpp61DvR1UZ0NQ1tcxWQrsFGbiuNH5199L2ESuXmm
HIFXfhMk/RYw5Zi1uoKP0UivaXMQhnPy7XsIUyF06NNgWDncVWOnuGG6MVHpRBQhBoBGjNeDHBHr
YWFLZJypaLyvyvXGB2Msl9jpRnDty9Y117IXMNAFdwNbSe9+OhN4g5ZWk4itO5FogQbQzGm8ZEng
WQMVYewKaLlE4SJLpiXb/cAurdusxT/3NppEjPA4rWc6KHREH71fz+0Vt+j+MfDhviz6a+6+rjYc
6YsbPwZhUxLsZP2WZwJmigFKrOOI5+WMzO7cuLzb9ntocwTmGaCfgLzwZdDy6TZZSSjfTpcQPLNd
wyLyWciB0O70ocG149ylGPbdFeP3u2mdqKFGhgkeuRL1JsDUTg7edmmUrElxKmYde4edAW3F0oBf
ppCVe3EtsK+fLCV+JPhnmYfSa67+oqvmWokwqzXsRyriQrIpNcc7zl0oubnf03THHU2vlrtmSj7f
s+pC3/yd4o43GedsJi3dGFNPq3uZ7tjwb6HM+sCp7eCJ1p2btftx5xIgIpNPN7YwCcFUA+eqAlDe
HIRmYbn5ts8lk8xSK6KE9NrZ1IjULuKTP4k++yYVknGa4y2iyN9YLI+loVkRz45yr5VMof7H9E+z
fh+ttbCHESpFK8Iqe4/DMfIKfdVdE/G9hKwaLuczxgyMKSWyAwx5EZirSDWoqtsQScrWBlJPQViE
AVDAKx3YaiVgqM2vhgzk5rnIA3UyR79yaBgtSMxUMkt4vwTZRMoFppEnrnN+Ug8YYfhfE0IGwlK2
KWfs9QqSMx81k6CtMGC2DuW6jpsHW33huBpbHTF7VEEX7TOuqKGyE2+qye7+ZX0jXzC/wbersogp
HJC4m5iXABga+VYa3zK5i2gr+ku5WHCInzuEvggro4wkdDqwTwbQ0CctAlmQxvOMT79tIpIKq3/o
As3ZPQRmtiYxKQJYkTLVO345nds5xoxBUujAqIPAfAQDT+IKdEa5Xc19HplCSOmXxybyB2L0IX/B
1ID5v1J310UcLuYtM3Nzaszt3BkRucdtJEmNnaBN1PwaI672t6EJK/QdRCjVL82s49iCSQaIiJXL
keHQBi+6dauSooVl9cPAwN5QRY2+04PGJnzaL0FsyAeQsYtjXDatCuejuGThQHPZwIceBSIENBCQ
BqP7KcD/Zb0z8M9W/FmN4EgpluWt8X/v5M1U62+sC1Yq864Ebu5RrsY93MPju2JTiKllqycOqwUj
nhPskJTBIUrpmFyL5sNGKCNQwCNeib8wv/qEkffqTFtFtGJ6r1UvOjS+3LeCsuxN5DIYlZDaAbsU
rvi7eVnAPbDBjh5p9Gifa0dtDCF/LTOF7liHjb5adzy/zFvE16ezdZsjWq83ba8BCYtNQUoXWyeH
usOCDxWxr+aT6ZTS5wEDyztzTgkWwBNMhulqE2bo4nIeyyxjeKXfoFcXszFq/PhyH2/0QQVJ+ha8
22xwyWZNbw++c/8ZaMeCs9LvVOGJU43yyGM1aJN4kse5sKPYh65H05f7mAx+aKRCCyUPmV+tc6EC
moY4yQhlhSfmdn0Fdw3nTAcZdTeYwkxz3VGkfiO+2No5O7HQMOlM33FQ24pLfI+Y4Cd7QSBljbmZ
TalcfHYhEg4Wpu+CZscsmHZ7g9cMo0XkavIShv3irSSkJQU4lwL0HEcxqT5EBdYW0ygwtC98QNmV
BPdpHqPWfwg95cF1pOYV7JF5y2qv04lF4H/JMS/K1Oy7VLdEdvBskaM8pyFsvWPFMrSkUXzFVJOB
xr5ZYNFvSzQ+QYUo/d6X4/KjD2he6+43wq6A2BeMkDx/5LtPOA/fY2zgGTFOrZ1zNqXugYJuWoPJ
PSz2Dvf1HPXkizutKfwzd5Z7SBidTuj8odCwB2cbpMkTwMPlUcLCCYZGOnwrWM5vOgESbI+xeO5Z
VRJ44KGasS8UnAkxJyjpd/8DjzpCJDmclAmE9Ancb7DGWabnnVazr1fgthyyRpFtJ6sYI+zx9DbA
GO9UHUzwyO1jtrbB4um83ycgnKStky8BUa6D/Gm5chVEVEPT1yROstWYm3HnE+f6p/gN8lNbKsbT
VdqaNx/UgCySCKoTFC2rfmKWlIMa1iv8mYjHJ22oNEmlBS7DKNr6NQZ7iNWMD0r8rYYPtWFW3XUT
TIdhvaUgfzY7fajVmK6iXMmZyZuzgAUL8RFCMn2BS03LQA4vomjPMixSN7uYOs4k9Os9ZQNrnaoz
qFkhaVUTBbGmzeak/1PZXJMPi+2kAPd/+P8BN2rPiyIlJJbIAiMGgkhKdHOOfslvtyXmBd74ivq3
hjXzN+GiDMsl95M8Cd8S7lGOk2VNiKkUQx2owpHTF10/2UsZ51RPQUIguprZ0K1ZOud6LeHW7foq
YgCnc2MOHTQtFYTNlnE0rEpzMwkkEt+PfrUf+GVaFdsffoV99ohM9ITa8EGT17lSMC6eEOc6wRcu
Itt7QdpSOshMBUH9b/eq3XfflRTJ0Tu6VqAQiRBQWMbGPAD8KQ0a6Uear/wiYGuK4ntScqew95GO
JaugpR7g+Cs2V5h5/Y1xqMjneyo4GkH5FHQc4QjyWt7hEXw205K534XP/Z2IxsGoujGk6KpRQp/+
lh6kt6xIQKqUjjhvzA7ZLCSrVK19n3XDUUYNwz+SaXj5FVFQ84JFTbAAv4of89gfl8PHh8DbdBHf
12RNR2MLHy9VC0WTnKwp2+9oGF8w1o3aKNBlcxOXSKAEjA4r35j3GQYW9zASexX4nreMkVbGjBnx
MKsZ/r8xLdfEKRjDQJ0vJiltRKYtaY/cL2w2dhcW9QKX2cWhhD+q+IZtxWzqyNMpxZ23NuRqv6ZU
Fs3f74HbENBvPk8wc0LJ7fOm9+WEoPUq1A+ZGtOFRjWlDhZ0H63q0m4MrEm/FCBfY/WnBBuYsXkm
yS3bGfXtEdJjo+/whQw04LktZ2V79ZY5SHHUOBYAqMbNlW7Ynl6SUoqlKqRzI/QLz/3krAfjpt+F
tpY5O7zXYRgrH5gPRidtBB6dnza+1wJzgaceiFZo/nZDAtpaVCOrRIU8I1PT2HD28KM10WhXzawW
DuGADDdG+7dvGePJKuRh2Fh//TbZhIKDsdVkiDLkLmnwhYdVQ02cXOnKiojuZRIzIagMuO+5FZco
iIELY8CALNqY3wKxKKt2XIp6IlzgMsJ5MQbP9OV+o3cRQ7yNwWB7yNxEBJq36hn+vUmDyFPIpOo6
SrQWwWAJI1orIP6LsUJc8ryfqRBMSRFnhcdGELlEqHyGulizmh4HL/lmhMr05d1nhD/itf4RyOot
btY8Ap8rqUcFQTaDGnqzFzsVeFvDd5loym1k274fSh1GoNiw+dKqxIiUhZlo5iIFMctu9kTl0Kdl
EW/GnB1Qc3t9KIrTeodTokQtqL47uiNSoe/8tL12LdH18AXOZEftx7DQOvrIDS4sFFnN2ZG4NdM/
eSdsGufZSPp2AWWfdA9hl+vqSOkQGKm7RbDHkv6A4TitMwSDgjop3ksibiwt0mCYhdrnRjEeK8Qs
IHqdGTb4lE3Ss0bSDSn4eNNRNId4UTvhiS6wU/jToj667I33aimHBU3K5hEPPtwfmhJ+yBbWBx2u
jcPqOXN0HTYjJeqBDeKWVlyGCiMhW++1QD57HxC7KH8PwiFVhtgNKn8wRcy3keT69mI4/oI/vBQP
0f1zrtze/BVitLRj/OU9mnj+G/15pwQVllr/JF5h91OhtN+C6KLaYhPjQpxrGhRl7dUc/lz4+xsM
uCpIjelL96alWPnLvd72dyps70EpvqfsWk8WPkQoaH9aQnCy9IULb17qLstqBuN5gmGCmGDnPhQv
oCrfqphBBoCfn406pnWBn/JgzXx6OP55RUUZJLOyEkPJdqioz6iNNAF8xa1wPHhflPb1HAo0mwyH
PdJt1JnCdL8Tu+Xz7LP7RSGqzKsycqJ09dCV5cwWYU7YNyzh/wDD3g9UpDzjNbQ83+Bc1DxC5YUo
7gmIdSWjS+AL+ngGa0lpbcRYuv9OwCkRezsUxFsYW4lCbQ5vHvBvQ8PykhBkr20sbTH3FO8PXAxk
M5ql4r31KHMAK0ecFD9e/m0yKfjtUZAWsmenvyIBOHSXDW2K0rEVQnE+SCGUyy0fPJmfNXp7fUA3
e1f9D2rws1ggdtlNbkkmdBpOYRfgAIWq2nY5hl9eC6WVF4EHj3k3p2O8/3SalRPYQZtglkQVq0um
AMf6y5eGlLFzTVXosJlrSjXQYsvlaOEpLXs+LY980Pt4cuwsZhhRo+OPfcPOL9+72lOAWZpQif1d
27W6+VmdSXBneeFvF7dE6mN0/x3fgDblGcA8jC/Z6nJOeJCntjhgunh3NLEdngF0e3qDjcF3Eu0I
vVBsbCf2QF/bAzvd3yduT8C3Hj24WOcgGc2hzFplUEDHbHP3R2qMDt5f/INsuYxr1bTRp4sOeMO6
a9uLqJTEHYzMDRIJsOgcoGJM63786HWZ/+/8v+kJEi5Y7wYfU0fn+GP9NuAFn46Q7IjRTs1ffyuM
M+ggddgcctO46mQKWsYLaaPOT72+st8kG0EKhA+O+hpAuZ32xh+HNa0nHxat/Fjg3fUg/iN/UHuh
roI0gdjldHZVNyxWUBJaazQnHkMh0PfQFNbG4aR6ZMA+LuYau0kJXD3MCaaMmOVat0azJ1KJbBH8
JhU+8kzSg+p8BrcCQGgOsk7EQELIILVcs+fh0vzH15iEzGqoERkMasqzyJNC4JTjpCh/71hbG6ZV
Pgv6WjIapn1weeGNBYSNpYv3qYux6EkBBKmCYn73kxAUr3U06OzrsQX44KJwvM049d6ecAEzm/xH
spLHvLb0Kje/hX9GOoNFjtv/CzVcYKwrYkK/hEw5JDebiju/gaxH2+qI51r3ZGWurQaxa8YnOESR
MpL93VSZaDSNI5Oe41PPTkel01d4QoaBTykuwfb/YtF46Jr65EiByQf3Q6nLd9QHfYmVwk8uh01K
HMy7ArB2L+JWOlO32OpzYc5lU/fsaq80UNr0ud0pavH7PlsTON0//qBdKe04xQqM4ON1P03ZlPoF
buvmbAGxhUTTTqeSNg4ljcSFRBW0jY6kVCaMBqY9mQXIsHJ9Fq6wO0jhj86XyMW7zc5Ahn7mJQB/
WUW3cUdlZduJJiCfU4TQscVV1FnpNJDRzbhzFZCKi0fF9VE2NLMhql3vVm0BrpGCwEX0f8/srM5F
ZwZfp/syMa8hKOPayIbwb/Mhf4SHtnLEs3rbdumqfxJdnH00baDTQVavpjKqZaA0uXybxzeXGgcD
tmIfPwSGazBaMl55o3Q0a8gD1U+wZQhB1eQaNn68mzJcVNsc1xG/oZp6XMVcUMkxjvCRxc4fRGK1
ye8Lmdc7lgJk4GafmgCaC+iSQTb6kAsv/BuN/fr8UtHTZP2xrfiLkfsxu58P50WWcWEj1wzt4il1
ZrHDXY2bAzoqOEcuBcHlxWfU/1qiuL/TWMM79uUSMwfROAuBnJZVJ526B1i84mE11v+VATatt3N1
iUnF9HCoz2LJQe6vtxajHzpl335yFKFUzUHK04Tq1kqXFX00dAZ/lSKrboD33RK5AQDp6uax7vbe
qnkezWOwMPxETqucNFeCV4NVYsvsX3Qxc4ZDCDYMLMsk/++Og5ODc4CxIyDTcw1Q1lwROIhonCky
ycVFRLYsiudnVNsTbbXIpTQzElDbIagf/MXToXcEWOVPQ3hhhiD5UNKaX8Qsrfj6I26U1iT3hUAH
NeVAikYqMVL4t+QzfPgLmuIGYbk8fIspb0P9I9bV9Em0R795YeDzY/c4DNuXN0RxpGQp+Qo3VyRM
xKahZB4PUcjbtZHiJxwNP0b7m9ipkAbHFXmsI6PeaLdQHx6Vu/0EoDYxfqxhv/hxBX6gsbNBW7IJ
l9MGCovUV7cxthMRFiaZSflfL1vHkySmbYhRBWO+OstOGI+pQmwhGChcL3Yu/2iRx2+m/6F+ZKJv
FCb8yP2isn3opDCJZffQSL/ldu7+V+eFrOUyGZrzIEaokRldYtxwccQW1nrIaR7V2Nl543HX4m7Q
zvqWfQco11WcaBY6c6Gzy+NU1x0x5NWrjTzOPPsQ73510UyqXpJ07a+po2XG6prD/Z2iVfNs6BL4
o8b9TnfnASO1LNqK4nZhPjIgDTrsxqerQ3e3nMCpK4z0DTHvO2f6ta1FgesYUFt8jKQzzTCUkZzK
ll4labSTpMNXwZdy/7cSlVFNtBFChuwsiyhb5ZVPM4wH6FwMchET7Udl5Q2OrW4fH6lkGw1mWJRB
uF5wqlTNxA41TTmzpsnSpWXHqt7Gv8Z3zPWHxVjfM6T34whl0ck4HlQ8kUeuRWfh1tLCGC4gxr/U
W+Qoan4Mp2TcMMjRrXIHL3XrzBUJPgejXwIblHmbdEoH1SCOxxxw7OVfJvbb7FiUnW91uJHtsHjr
nvPqe3fdnBvzRN+fXuF3SUsjFf0luQg8fhitGxPdJE96Cd1r7Wlf8+0o0y3AMlK8eFd29EMubJrn
dN7G2bxHhUtpvnhcFAXitW1RfJXVMc4MJPWQ+u8KeRsrtL/tXmwPBpc2qKbPgPGWqRwadkoNQk3w
kyrzBLG8jKTSX3H2GY7Hbv03EoohCAYDKCnQaz7kSQa3ts5ZFNfjCIdhJE1i9TJ7GZwzCZXd9R7C
vXyx206fplTb1REJ8FDwy43lUecMsxK6FnyHTEzVdZ/8YGrefeS+wSjkO1fNgUZErl01/A0YwBVD
eEjfqBGUlldu18iGw2yx4jZhKTAe8I/L+oXVG/aywJ4p7kWqdsjMH1nwzmkqu4gGfcWDKfaV+JaS
Py+wt+tzOb3qP2epsKeB+kkfCMKDI7VXF3uCiGxQxMUiE6jdKBGdGr+psE1JjPuMfFYG3/pVIsao
ZDEdV/PSNHu+YLHwrSOx/sBbiHQaA5aCm7ClU6EGQE4lJCzKYOIgTV+tYa+XYF1iaWCO9SPLYxNz
x7R39ipSE61BZbnFRmCPDE5rMyF+1E3KqBSYkDd6qUiqOTtLdJRdPKmkoVPLaQg6EgiiNnil40Zb
9YXA5qa604sOn6Pxb8tofilE3FbA3BtD6tsgxM15DbeZ2w25FZozp+E/XD86umOahWgFZgW2i2NH
PkFrNe+5utI88vq0pyGCijZZLtL7sH+sJS35xH2fO9urPY5nQBIxlxXPYPKbAMzZAohVuEpvMhm6
T1ntsQIbqqMRfdBLKb0Gdlr5m5LyxrkarXvUpmW8k8dV/FR9aawL64/ZC+h9ZKNBcklXoYzhpZmZ
amC/nnx1S5cldwrC69aGVgP3E/qAohUMvL6aiJg7ecquNF7nVP7jv9TbifFxT2PDxDQCjCKOdE35
kNelS3sJ/PcpSI/F2GDsSta+oByVVpVkQDXzAIJBRMdRI4RE1gnkiW6ryZ93NRIaykVCY97wJAKQ
Ozs150yrLVKKl3azxZJkYnnG1tebFaz8apldSsGjTvbFl2eadFl7R9DdM7tkggiGzBkLmm18xZC5
QjMTu7zxrC9qocL45aIttasA0kDwBXmcLMG1EvugrEx1rNP1hKlgrZM87D2Drukt7upSg2W7SPcF
RTXc+5wnTXHtH2rhiKt1/Mlkd//IFSGUxAtwMhOOQYeA/vivczp6tBAdqecyRabRDvnmFI3xN3Oo
0vh2LjE0s95UVLB/6QI4KDcyU/WX5i8oxxKrawaGBd3YY4Fnrsm61klXKe7RNXDvmK8ZOoGWSNNj
J7JXLPN2Ruf6SH1sj0pF4B/CPJFsaJYuuI1VHnD0lspJaiRLpAy7u/hKf1AXMirZG2MSPrD8h7EE
Dlx13VaBytgnLfnUVQEuypJcsUZqyTNFjL7ldc/674Nenfr3FUoDoYQJLLuctfGMtAU+NlNKdeeX
VoPG/vodOtDoHH2b21yo1tX8G7bLZYbV88eGtjMi7g2/0l4Ss89lS96An6lw3QbQ+staRFWjcRkB
HVHhxPsUr1v12s02efyhb6GMOdaXoi/JDQHS/7zz+cCi1y+97aWIArKu3qSWqVgAkH2irFQpaMIb
qSjicupIOTWe+O0xUbw3EOMuWZxZxa24p+d6tWuYAunBiRNEoWiVvXpcx872IJ4K+ZZslFG4SBhd
eeCXXuwUd3VruQkQXXdkleaRn05jNxRsG6tqzl3Hop+7BCq6nYV+Yyi9quSi3MmduZXjP3077DoL
5q9rjC0iTmB1EOoXagivUPn+10SHEi7ef7+d6hV03aqF1G392wkNioLw1yET8ezRgicZwGxVa/f/
CyYmebbPgF/0vtgePHx7tWT5k2ufxk72HdDqi6hIPR5cKenAiw+FHuWpoN2t3hr//XVec2i6T9jF
ltpIaTJsvL7cn1Ht0/r+Wlc60QlQ7k5H/kZw6caTK2a+ZAjmS4lcjdRElHojPJuo29mYKmwV+42t
GLdd5GVAJ/t3Ozx7Fs43r2vlMUjZS+1snZJGqwWJTGP5MGr8rdrg0tP/7IxQsUjUUx269mBjDLdW
3eSdepLFIZFW4/k6bYo44tIJ4Us6hD6d7GdQgJnerDhZbxYxkOSG7V82za9TFudKiN6ai3PirApi
YQHenqWf+dAqNvQTNb8Wtu3hMjdIFHu2jZ1Fyqk91tYb0DERp++L3H+DhtScNMR9jPdj6up7g2n4
8pXm9sOPark7LUAck2WU98OBRzkSdt+oa3NI5Eb3oecms8Ir3wUjHT2OwhvufASRv79e5nMdu3QX
5IGCXz1YTJNWGFAyuuT1qhTTZ1M5walfP65WVbyB71UQzt5UqVbHxlozUC/JBRkGNk3oNvnQNuDH
ZwHACqsxJLvP6w0iU5c7MjLWzhjR/PGz36OAbeG/C1iqdO/RcqiR7tmWFD1P9P8DFsgtJX1T/ynj
+rLo7Ww12YTDgRuJJe/O3JB4r/iAUqw5ZaE71eKc8v2qt86Gk6br765S6Z7jixrcMkZk7YyLYlo+
azVegqgoa1htvluo6/uobXW0fal0USWqmRbqNPlQ4X+h/XoN1HJnZasKHiGLvpdKM0zj4G4zf9U/
zAOhC7j4aEadzonFsG5HbeievHXhMSGL2cBAIXP34Y0qYcJc3cJSwGO+nQZu99U57/NlBqhRXsel
ykz/uuZeTH4RYgZpF65wSJg/3PTzQTBxCIoZu2YAfyBeISpolG5TMVznrdUFnKGTspqtIlTwkQ60
n+F5LnZH/hUsxOB3T4Ld7YELhFebz16ksNWIfYQeI0bLfJyrsuleXhbXSJ98NOZYzxvoxpATyvxf
MMm1up4Y48KdLr5Z00yEyZx9uGio37JvJ9de8atDBfSV2LgsKZs+tdstI/GJUTPvg5rXNEtQGYan
e5BKhXvi/spSJNqlxKnuroUlKU/FEvcaF955469m4wCRSF85jEXP7h5le4lnz6TSDNfXEvn1zbQl
zc4WmF1jA5jHVGuqn73Ka2s8OwPjwhiB+nhWYtEnzgaVo0VPoeOttLRtU8kEmb49AK4m+PrEKJwi
nEiaqe1IiuQ/SUQ4tHcdvLRsxmih/1zUBsJ7mkNYSpqrdWC2v+6H9b2Kyyvt59AvnEkszEzTyBzp
Hbwd2Z5mre4TVZGgk0F0pCNbhHIFFABbx7z+qStocYsJ6K1ktA+Av3QrGewRX/gOSmcKRWy5gqcI
KHopfghEUgHspuob8AdHBe8tvHeHukChIqLdIzgsGnUZY9a7OX98qAk3GVkQyxhKqK4AE91LGjLs
ie75BT3hr81/7duV3Lz8aXSdxJaWEAw7uOb1vzYzTPZpXSkG8a9Gq5kMqqLYDffouoMhDE8Tsnuh
zlx3yxEV1H9vhPjRJIrgzF7q5eFA4VLtOGP3uT7X4+IB0ebiDDQB4jO1PISxlF6pbfkiwVqgUR/d
B1S7OtVD2gMKt0aE56nXKgoTrToepBxE6cUykDMeBRQfHFj7DqJkRHX+wpz67Tl2h9JflvxZH6yu
M1mPOHqQtjLKakJJt+7obZN8ATzAz3yPy/GfdFmsSxF74AfNQa0t9VT5LZ9cC/8UL81wUn9R/noo
7qcl0BmMlp7K2Y47Xo2DtKsWpElR2Cxj5wXrQUDjfo9Dny681RZpchyN/NP2M/AVUEVfJA6RJSIn
kcec6zttrgyOyohgOsMxXHUocfZE/HYH6ecYbpjMXEFvQr5t1tx1Cac8kp0Q5BDBzfQcp5zD3GA/
nSJYxiuWm4yJe3bQZ6PEUO3orlZ3nfdQ6iN+EO0SjLUBXs6qL53c26bB7DeXnDeHVieJ013ThTl5
0B064SKe+ENoyYU9BtcaR/hcvHGZnit2I8t3LaNZ3kuqWXXZKOIKbX1yfxoIZ2sFdfWZFII86mvC
hs8ZNVZWpqG3Y3waoaru3r9QOTP+TgEWfCiRXb5/FN0J7DUbNrsPP6Zi/KWLrJIcpBfiVhK9jHJl
kM98C4Urvje/+D3DUPLod1l//iXiVHIxsxQZfqXabZp27U0LSKW2EImHiQzjFU84bfDnaMqEUvCw
Szo/9LdiFKSqLjCgZG+Qe6GXGo/uPH9zEPCuI5muHEM667egl/Qy+/fEyfdx+FfDhUyPz9AHQjxa
jva6Z8BOP0E44DEtIT3wf1SjT7iMX+Ryz81c7e+Ugbbpq1hfabWRwBZh1LbZND0a+bJlmzhmIkEP
mGtoQ0XNVtFPOhfvOWBsdAw3uBbYcM/IXeGLfvYgtgkPvcxfqrXctToZKsDTcWkCPG8vQp1mYr3I
eDVp28tB3w6LRJsrkYVw+HVTUdu06yZ1/cSP2LN+wXw9EVYUW1bjwCqUVeqDdifCva/ruK4jS3NG
w45DY35Oy/N3W3+5+06gP2DRavkTZTBKULOWGhFLsSFfF+TTxGa9ESfzUc0o9q4wFwjZ+tieEHdO
1WmTpToipFWBujkVNr4zFzkYmem3NyNmuSgu1Hc1CEl9RREYTLfZ/+UWxQ7F7HA1q2uHH39EWJ5k
so7LrMDTOncaCk/XIokpaDGDM241GTq4bSfH0IQhkimU0i3sdUCESDFROWUpRt01mhef8Whmq+ug
O7VQEqJktOs7HynsVAeSe/2OrCgmJ2DMP8qVL4ub89Bp1hLl4T+1I7mx6I1hfgp/rALo9atbUpwN
2gX1pqQHXxJYix6e+yy4XqETwqhm1LvNCsQZF/A3WuyCIqENcHEhRocq0NfBGZ76/wNCC8DSgu7C
VqZaZXL7JND/tMg1dbf8Ae7xaQs8CUk95nPAGNXv1vHghLMkEuQu2tpp35qLYL0C7Bvx+BvYej9F
ScODg4JvvvpQUTeLtWT6KwcLk1qwCqnNlxvzuGEIAaGGCewaMdLDj5q3uBT9rZ1DCq/yFT9+Oryb
6A1+UVvzPwMs9LqLeu2uUaqH062D3U0/J5/OC3z3OxDF4JtGhc+Ul3zgnmJM+lklOuF9qLOWAzLv
pzB9KZ0WlitMxzh4hTwL7LXKb00ZBhEVaqVkXeVb8+hH8tP7JWf7/bHDWzCtRjg9v1GnLfx7OFoc
wsNJFYfd5J2TYFb5/hNSzDaLTzcs8LSxY5VeVpBINmXvt0cJHiLZ71EZ80BHHDjO6vj45SDeDiAB
w6e3m25Yg+VDfcpFR39zuRY1sx87SeEAc+2sDS4nHV7uUb5kySE9YfiqNXfialRvItZ0sbf3FUOu
I9biHdOFlbuxj0fCtF8PeOm8fu1Io/2LwKWDtlyI8NaQPNHuMUtUonwEsyQomdGQzmXvHLTg48m1
c07l88NkdX/goUoYFmLxdjov/5N+5uK9dpMBMF9ZQbjJYYVLGPSj5HuNxiIxz40TXSBNjUEWLCj9
MJkqTKPcvyZueKxute/S2kNGG2fntg485JPjQ/CJH+uZxzXGGXDTf9c0Xwp+diQJfQgnyv6dSa0Q
QAoKC+l4ii6a14PZW5cMAUXq3Y3PQLWDLT7wousGYkWp1JkMz6U3ro2HSkPmkZ8FDMyFG3ecZAjN
QW9nMjFmjhLDCLPxCU5UcXd0JWASGKiXbfuetL5uYbfDfw79FrlxEtmjmy33yN3kIaVO7mvvbC80
JWNuRaPF3Q/Tar5EZwtEv5MEEEdbhuV5JPjumKdoJdO1TPPGhkZF4N+g3h2zKKyIB4aBBXfvX+EC
l57cnRhw/yLbMiXfnxtug+5tRdkhQGnhVQ44zL3PpFlLlSGQhCrzhpsuaHZbFhlbZaaHKTWTM3SC
wXoZQfrDesbbjeHAhIEavG4EqMxSrjKDLYfCtcvQjEFnjPQaNwB320MOsAU4Fo+IRrZMWwha2TiA
Y5KfkQmzteD68dpXHtBcFVENbNi1Alo+9nr8oAh/jzuhvcD9GSjEZJaOkD/bYYMi9FzWj7rhY8P6
HsixOuAdE9EMLUIEpxX+dQXV7tO55Za9iE4exePjAFc4u4gbZT577x/ROlPx3SABoMd4tNXSD7Nk
w98WWXdwsQd42ASCmVKwefl3xDqPL50FwTR0YUJDHi6nZNsFfUA8zEufGA4fujd5leYNuhpebGte
z7Sq/7y4CKlp2PUOtdyDLVcgKYeQrCL73fom3B8TmoMIokhDQEV+cv/wJ/i7uGvOMC3LHihIwk5i
TDfNqks4FXJggjPXVemnv/dOBAkMNjyp5wnxu6iYKMSe4wy9BT3WlXaPav/7ZX4UbcB4aNCtwAWm
AZkMyWqR/1jGcNz4+JjF6B5daL6TklOdN0c+YV6YRApX6NPfyljUf/7aDoUwIopU1n5NlEanljs2
R65e/HbyZlvDgUzDVQzAJKYs0Cgv17XwC+doSTBUCClvhjSO84r7nrTRSJEVqB0F3OGzZz5VNhu3
GLq5lDnOjJL6eCdK5GmI2FIATo0AEKFp3bFR1a5LfB5KUUK6hHxCvuR6ewWKMO1DyVstLVdzJOqm
wbzj7a4NgPYNv/b9p9ap1ECWbTJD/7X/LnDsTD5X6BWE8lmVYyj2TYL0NM/bmYRue8CMRJtI+1ZK
BfeSGqO5DlXMiPOU3QJ+Mi5C8JOyHzs9heBcpT5STw4HHiZgMbgoiktBLxiCzeZSuBy0emOjEjmR
mQfam7BkZIiabNQL/8CZurf3oolsy1rhaalUdikK0rTriCXpv0p64J7gC58CBSL0xnsFqtQ+2dQg
9lc3RpXuCX+Qt99MpzMoNX/RGJqpO26rbkTOr5FRVq9epSnp5h5TVH/ZdTHBbyej2F924njMm3/v
wAlcpQHToqkemB9qh26TO82KkIIYVWPZfw7zOANNJ3gSFJY8CSNEYlG0MAAjtpZJsqTOPBdIIHJK
JTFN1Ww5YwfdVkwVjn4aYeIpPISgoUm0SXmNhRCGwvC/olARI2APnmCutK82hXOZxkymhuniUXsp
gRxChDxV+ivCPfvsqm08/sLt3XKK2kCZyTODt8RiA73edn9cPwQ2sentYoBEFVThvITFui+HfsIQ
dUqAOBb5sWuXi9kmfAFeCuASorZ0yK0zVjObApmMxyyLPq6WldGnlV4/puBsItnNwS7a7D+Um5oz
u0bmNHVV353gz9kbXMEldPxIYcGfHn+G3dKzudv5sYRBzaPc5eQDNFnLtQ4Mc4OfjVt2ZOa2inu4
AUyJfnbq/UcClSbTd+6end8Yr0Bw/37DfAG1T3+wG/dKNFSZWJ8jgZbi58IfxybkOCVU/BStQetn
BgHC4TjkRyCQpb30lEC4GhL1QLc4QSo3ELr98cSQqmsHVpsr/E5mmxEAl41O0u2Hs0i0RcqmI9WB
/SiFV7EyrcRJJKGCEwnJ5jD3h1CGkcpYcs07AXbkgiAwmp7G6OG06ETipLOLxeUD8XCJMDZ5f8rf
YQ2v7SQBpU6OGYncj8KKpOSrD/CnrlpF2iq/3MILyQbHpLgTJ2icY0fc8AbGvMbVm9FlEThX9/vy
f02YfrVg1aM43ObCswwJJvfB11wzUfGlC3Qccm2pqzQyLGblCuKGmbWX8ahQWCsS1k8n99f/1zD+
ImgXjBECE2wdPilbj6lAVlh6EWna2NbOeQf6zT3sBOZ4c0/NPBQlAlmhJTM+KlQdWXRdW5Dx5C7c
w0wyiEzmsM5xS9QP90w+ssA0N1H3viqn6oKZAeuwnOzL3Sm6FqE20sQgLd8FjUB8/TM65oIsFGIY
2IFlQ2vLxtJkA8X6YOFyC+tIQKSzINsMoSY9W5+SUudx41/U2TCI4EZgeFZ52bqvH8fiMpAWUT2h
dtCNVAtsPxQTR32NxWNvBON1ZNSbpTADupQzj2NVf3XFx9GMctzryIE/5gjFNhumOG1VtvfpIG/x
1VZhGuOZK8Cgy09lUUURevpheszEMvPQrKn16GR9eTEAUa2OGouxaaH9wXdTlI0ZWjR5SIU43M7j
mgtDl6mm5eaRZT1bCQmAi3PJFp0Kd57A3p1r1GxHgHP4mqpzfEKJB7KbSEeSeJRmpLbVYwNjeL9Y
cNaZp+lzJkdo//Ub5Wf3qMaJdUUBAh8fUUr0OLNjxqyuW/ggk/Nqp0jZw8fxXthLHwO8x3EvjQjL
l29yz1M40+CT06wspe76nMOqTWIVwdIbLaKy49i755QIbPIQNv8KYddjFPkDpIBrR0s+ABX9h9zb
4owUx4Hh5ZBll5bdwm3GZCPjWIdPLfsFW2sHfW3Kdavdon1WEk4MmDOX1bTnUxNg5mLYGuwSj87M
Lg2UlKM4SYpLRLHCFHRhEZyW8UcdQdoWmR0H8xvO8SuxJO/HrQXsEDV/8tgoIox5cl3Qwu4/BuqP
zbHDVzK6LF0E2Qu+OP4WaKiFv6jNQw2zrYoMXTLcTTlIGf/Q5eBzxsN6JJCt49GMj7IMX5fBHMAX
XyB+HBbmm3ZBPAqQ9TsmNHhwRK7V36JWWf6HRijwbN3KNRiG29NOXogd427BUw0AfNsbydrN/Ik0
5eaMm0V2dS+v4E6wk7UsUZ/d1MKtmRN1omj3GjgFod44NJsGA9f8M/bjxnAFCnLcwrm2pcrPZkNv
Ik1GEOayKbC3bZoQwX5ruNb/fxieAQBWYS4SHSHNgqmbR4jzrhi95kRcq8G2Ab7Xv/vQKogWCzPP
GUyBffbHkrBA26ifMaoArRIaMjbM97lFiSVJMYotklRDwIsuspFom/VdA9mOYO4LjN7VJfQBHFty
N2WcSSf5YvfFqusmshC/jOE2+u88MUuJ64IRju+SVeoXZBWjm9jUVD0k+orc+Ip/8/Wipdja+W9n
JUH8VUJYa3r9AJnFVM5jc3VoZjhHV6+hheml3LGXrN2HlVzkP5W8bhXb2WYX2b54V7/tFia0lYt4
Idqr/r/5hGX4OfaBHhrYXFxLARZgZNWEDz9P3wYPKGj6q8Fjevbd+87B7qHSe/QOc0PD18UJubo4
IoA02L8Rvbxtwr9GNqlM/uS9aL+YVz951ywMCsI4ujvp5YAQ5Fb9/jBvzrcJXnCm80cmlH+JH2gQ
s4KoyQgdNHy7yEdyFUpIrmZ0OVBW2fC8jiq+Ldddr6Sx4CzFYRW1vrqpQXnoicGfiYQTgmHx0zcB
FcR79S34+C+1VyW5VwIzE8Wnx1QO4mANVYCcy9i5y6oPCzzJpjSw//heNxyx9w+QXCqDXeaxRq81
D5APaddS3UJSd2a2JNwPkNrC+ZlGEXQvz4OlvOgCr4sp97vr4RAPJ0Y3Jo5tvPFWo5LnwnKdqU6A
AqnlbVFE62O3OpDvwTQWB2AhXxWOPrfSItjcBC+DMQeGIkhOruoOYPDHEg0KZ7fZUcQ/Uzq41czV
k+IHjYth6n8FmHtz7DCc5/F/rQIcRVBplcfJwB+T7tphZQRDzGrRKQITwVbEH+bstZHQid4wR6Ue
IDEYYsqPFtcc/Qkn6LSh5b2nCCQGnQHfL+ZGZZX4PVq8kDFB0RAMih1ow2aSsIfIN/CLlKROPUzU
pBIgSzeWbGF8jJH5Y3GhLd+b3j9FhPFyozYIuk/vsMBBP+o0pXSLDZ6os9teud6S1EBeaneW4Bd9
KLn9g409EOboKqPusIAHwja6RiR7AJC2eF/ML0BwrTNsv/1wmGa6hgPMg5rw/0bHMMKTvfj+i/PI
gib/w7x3TSdX2awy/lXiJPz07B5x2QA+nl/oza89NhRXNNsGBcX70oatmbTlop0lyOzI+033UcFZ
TYMkkcQPLITGVpcfYJ+ZlO5uwBLzt7cOf9d/LP0jgesQGf3kbSEr0Jy7IfVV9IYpVTaYIsoNPsSv
tIsxP4Qqn4M1SphlVTZo/+qF+rfbYlXW0DXjSd6c3smcNS7Q7LfRcrEFevzowTdzFnYAg/b0E1D7
4MiuX1seeeD8QP57ALtqh4epUyBp0aYUh+tGyaxXis3Dt83sD6pfl4EwID7PE8mN9TieFu9uZ/Z2
17rSU6pnD2NeB88lQYvVmrJrU+tIrU8z5PHLrm4cu4yzlvuh4VNrXFdqMinNugZL5v0Y9jqxyJbU
s+yhaPT+KkmBJOHN1BJ5LE4XpJ9hhXDuUzasLDWc/SS70zWwRUbo63J+WV0LpB9O0zfQ22P4nNEz
AlU2P9XXfqnZTbqfITr1dUYMKJuNFKjUJP5SxE4NCnwJJ6DLe6COlQhb888M+7VsbnLkkbGFuo6/
wW9JM7RalxxigGr0Y12iAjlkut7jokpRuzH60IQcQpnYHN0EzYt+3LsVhtbJIdrt0LwCXs0dFU03
TSz3qdyCPJ1qVGXLEewR3MgBUjw3GZtQp21soDscyV98T0fFKm/ocbs/uOAMZ2yS8r4fChqIPFWY
d0pvE/Fvv1dC6JrDFKY5f/qexyVrFyxJ27wl/9BrsEau9+YTd5QMUZaFoaJeLCaPfXKw9TbuFmfU
5kQrN2mKA64Rg5k7psepsLIkgqWXANZq38/Zz/pk+6grQnaQxSWUTo1No+Q+0l2ppOOBj7pljgub
wlM8Tp9gsx8ShD3OdzGRtP1aTycaFSRArINnHjHrT4yi5nxF85n+F3I23Pcn0KSVkbak4xFl2exs
j0x0Qze4K6ieqAbQXbWX+0urSktgMq26D5ySRE/pEY7XF/iEyGJozt+SmUnB8yCGBp2GmvyFDrk1
2GdHMPj50VDpx4Z2Qv46//4+E2x7TBaAXwH+gA0nfzZJtNFHYE04qbs1rPW3Ex5Ic8Uy0mj4Dl8S
vEdfE2CGt0s+wwlT7eyxzfG8YFhB3/EQxURfwPgcn6fK/F57gUePeTqE9O8xscQFwbhjVzbY2htO
wlx7QdjZSr27QloW0w36MIRlR9LILMtRYUk12p6UBGgOHCdCCAcJb7pVs/EXMvhzeZEVx+Vjpwp2
byhRHrBavtwxIKBoexGTm7CbdlLgPIqm/hrF+Z1G63KKhCI27APGcXDOZzHQgfJztHs8WHeoQTEo
KfDg89iLVFjCpVaBYxTvokkGPMulRK9MpvOHyIga7hrQ5G6p19EHtdXnMLA9fB/qpooHX7cpe4pC
/H7V5tH7x3jMR6dCmL2sqYLiKlbANUxgblDyLPTJbacwPF8hVhWwMKlMpiGFsCl48e69ejPwEou+
lAVbMIILIilZUev/Fd43hEJqCxoW/gdmvehrN5iKlTy6hprEM8QXdxe4MatPQf5F6LdfhsR651nD
XOEtplqh2tpNJ7Mx5gVGoWGzJgDXG/MT4UsQMimB5GGXifVM0Aydzrc5w8hY8fnS96JBuV6AymRB
TwZpofrBa9ziavugrg6ZN622b+1+iypK7v3IfP+njPvjTlP/8/R5sXRlm8N36bBDYpwZ1DCnxwlc
QwPZV4sOLlbs8hvtUorIf9x4jIFwpXE3u1jWn2P4jr/cDp6ba8sJsRs7Hps+gDtQbI7jiZeTGbXV
WtxEyp0f0a5QhPQ4Y+z1aFmR3hgFkn8rsRWgMHWaQG46uJkjfDfPrvdtvCRKz9GUsIgZYSSF9htL
3o0+VUSNCMN6NPjVB/DSlENbUPeLKyjCLfa3fAOK2Yvxmu/vh1th4zgarlRA7vRnkhOePEKQyMbW
0KUWilFOj5iSIYHwJZcbsh2PZ8IvxIdtMorZwYxuRrcdxU4uF+a3BMn/c2wZPVb5rM+St0jvfdD9
IL9mpvKpQjGNRSEWBJCCbnHwSPJT8F29ibgGIa9K5oH3zjpvCI8XmXtM6/xOfWN6II7eOVlLnRW4
XAMm2RZGWZtsSFPkp+n39dQYolv59IxXLR8kMAc3eVV8+RtX3sVFtA/8QX/5dQtFbrzGMVY27dT+
SQN47eqv7PCF3NxVrWtPpsMiUcidKq9TSZEmlWQf0pTBpcvrQ9Y4xCAdrhDGNrTMxmMcK/AejblP
eSRRvbBmlGg8X9UPv0yoQoNtC5Z2iej5COk0A3EBtLXMTug6JnSUBiLZaH3VkC/rvSh6sySWAhbY
XQV/zoRPD3JOPl0rwJOPA5LpQJJ6y0kIeDZcx/ocpNh3TrvLNRnE5EAuJWojNhLausvPeomLbG3i
lEaWp5bb70iGMoh5E7Srx1KV5pYzcclEJQ0JkdixWCsqYsugBGaM+52dhjr3r5mH39bFkrJU7vL9
E96iz+5cqgN7qhGw2mLpeqR/FlssKzVhvNh8vtWKmaIFSbdOtWlqtViBsmNk2K6VMKcC2AxcVjYE
YIRLnZIPNM+nq7hZZ0XfKpBRGwapANYsp7v58nthhzv1SaPdvc8omGw/7iXvqnUkqEZ9Vzq9ZasG
umHb9ctC1UvxPfb3UBPbohgpVjXeXpQhi2TuieAuyQq7spSURRUEBZsfmJgi+snq7/ZhKsDIGqWe
+NtRVxy8MpSlLiZHiAL+BnLIMl7m43notZc4ajl/PIl79c6caIidvWHMSyNSanslz+Zo968oLG27
n5BTB5t7XmIS3IGZnKEBHZ9ywjm0yIlexaDX8+1BMigRaS7dXmLNTOn+GMLdlL58d68Ed9UAw9KQ
2kbqZr1g8UfNJd4jX8Y0bDQYwEvJYFPjFhRsBIa0F2/7kIJace6TQbUm2ibjU1OErb7pzkbpaLCJ
7xHH/W/mgYzopC8wZS1lqmaOiO1ACfGI2IH9rd+CvJOBgQhOx2wv7jUH1zey573elpRVJb92no8l
P0LxcinyoB9KAq29lc6e0+VAxcftvGuZCgyl0w+5vcldRrBC6sHS7gZAWJXWNXR86D4WLtT8aXPb
sf+vCVGzfYie5qB8/zN7+Lzf77TnWV30GxO0fMXsUHYvG8C/3Dqh3ItBNwBWHkGbHj+zsC7FsShi
TrtC6OSMP3e+WulTnNKIzfE3Kow7KT6ZuvNfosraf34ndfc0RFaqKUGmxL3jtvqzlFSCeFRmeF46
xin34UL4g0/18xqBZ5AAQOYjbjQm23hbnJAd2YhIBQPSQccxDLQBIzcIjbv5SYtNopf2JU9KUpXu
cJiFqqEvJWLDtzpFmF5HI1yNHAfrgxnpyiwRL4z0JgoZTaFIGL44XfHJ6d+mfT2iqbWufpOFOcfs
U+cScSh0WV+ZsxuNmc3b17beIDSo3wnU2n+OCmjkGvlGbTFgSBMsnGJarIqYvwRfPF2pyR6bcb3x
611+GU216s3f2KeUlSyEt6NHTHKd48fqC5+aCl/Aj/6vZa+gMai7mPLjDFCWGFVXVPCZO67TNy/1
+SPSHrZ4YzRXRmx/pY28s4LehZFliHDA27OLDrvie49ALfoSimJN9V6+yWS8rumP1qA9UAn2gFbp
4ujKsvVGUEfoNTh/CzyEWXUy4xH0eIdszf2aTYDgYZ6/IuOxGg4pJY3Z68sampCXE+56p5TrP/7A
y8ptI78NKjlJaoW0usrv5VoUC5w1p6HoNeNfPQtiYM640RdDR8QsH/97Bb1UTPP6jcUGI1cJv2hv
CIh2TNe7I7nxzzFlqCoRN7uU2WuJfxg/YPbzGU+kmIlJXkl2w/A5+pbjik5BC1nwIOzVgXQvM6Ct
8dIdYHS/qZcDLcYBY+J61ofwOazS3m4UcB3T+OmsRqdLZIvuxhlumeda1FPqqq9C1egj6z9vRFqV
Vw1yrISy/hZMGPygm3ePNVZrLpm9kdJu63SCoolK7e0p97jGpp8gadU+l4pf9aEXOgxf6P1KGglx
EEV069ArqzK65grvrUfNTQahGLAl5JhjoIEcP3ktaoS1ve41brYa2XR8AR7tOi1n4sRoyIMcGev1
go9Ol4iHWoxkv48pxEHPYplqSeDqAXZCoSpGHu8aHr1Jd1hmV2U/Gy2WeZyvFHcNSnDlgePzwuM1
Ue35WV4GMHEMszebd+q7V+w7nmZq4Hj+X2oMXxd4EDDgqkTrH/dcwxnhDSFZy1ACk24yx7UcU2KO
XG7g4sOpoQV0KEJV65PCjLNnQb+Fl0AENd2g+e+1M994PlOHzrU3w5Za0Xnion2+A5DSaJMn3QQ0
g2F473n4eBOLVlaCcv4IsLwnhGVnHMIvGjgrcY1n7s1iLtHFusvXg5XQ7+Ll5LcKhcRk7fLRFV0V
Olwylrz9PsFTlJbmQEyTCw54HSlq1v243TYU+Bv7qxeORjNVVfL1959SuzcbEIR3RL/0StMVT3Sp
Vmzv+pBqwqCdiGO2AdF67URBFGAmnITDo6y4tWOYGbZM4HNlsrizebpNwwoFtothkbrBPsDv0ynk
QTnYsFP/2C9Sl3gX4WG4qZv9EsoaQjuJWhOCQ7zsu53ICkn2khpMegjC3T5KpB8e+bHSEdksKajj
1/noTOPmFbPxkGu/XeO+LtyxOSQUQGGMpp3MVCaeQ649g9EwQy3OqIFrrUydwSYSKgFb+TGIKuZA
j4QviAT854uRvY7a+y7G8KQR6G+LuLm0WfRZtzGJD+2R9HiWb8Dd0ujO5CwCROwcbZi0Lv4Kmo++
tP0F8oRDSVtCR3tOhDUN1Besi9oX1W92nosV3NlicbNB5IiVrpNpKNMRyt1AYBKReg4eGjLU8t0g
paGpunCWtuzuQc1tK/0mNWGxrCSd31PSufu5PpWKleAVXTaYtXxvUrjkCTURDORcE8NqcEVgTVj0
wrHhe1+JQkbQX7HZS0oQYeCqUr/oSGQjSlGgiz6WBUZbsJLD9+zcRQ8YoNNFylK2DSzledgD6duA
td/VUyBjj2Ds/YUwCKTRxxK//PBg7fTMc/JNj98OfDWLrgDCq5vaFl0zmoWomMgSCxBqZLqQI9ER
SZSJysviuSqj4uKUS0R6CMQqv8e6MPdrGMtAoQ0+Cm9Vqa67izNPgPol7NoJUwGtDSkChNsQv6YI
VLfJgtr94x4oaesY+R9o/HMSHpEuIoIAwTlkCR/iCX71RMUHni8SW6uVnHGDvdti46heowfdneTg
1mYU/hgIwIX3is3sJ8pLFBAmy6S/VAU9QurVBdxOhOwseT8pZ8Su0KlUC43AbNJCtf2FpYBYJRxv
t/UWnV36A7wYB9WxvIZRvhHe5LxNT2caSVBMSMEMWW/GJoOOqsDYbXmW17Z1/I/B4+z2qi3VUmdx
VJl/COtVHp3z0h1xLob8maNhPXKLJsrAlaniHv6g9/SnAj131nDFpJj1ppfYqmrxqkxnT/rZrXPU
rYjTfL4E6wCy7DlB2E+Zvt7qgj/Ic+zmXVsIoRxN4AC7KXomTr1zi4tSvANWhNyB1yFBifSQRCsq
9HvhZAlZ4Ky3rgd6BPfb6dr+uiSO+ZPlANywj+ezCQkcVGk6wujUMmtwT0WyJQsYI0a3jNh/RcEj
NDO0UVv/9JKOfS7tD/gFHs8s/s8KlJjSBqgpTivRxdMhF/DRoPtpmDerNOPJ3fz3GxcBcAcaVG5f
+ys3l9wtVuLqvHBMu2/zIwQTFyjSduzDFIBQK9QoufKugf5jHCmum0wmx+v/XmFn3vKe5yQsUi42
upEQdW87cZlZ8nTJ4nDORWV6A07G1r23mIz4fjtW4aNmBK+bVM+3x5P1NvplylCLfFtYdkIKCbUl
83gPTkdILPDePj88XnfAjpDw8RcMysVrTVjfx9UWuJmlwug/BzsfOpCxtBrQrQNZBf+7twEcCU+1
gDKVQG4eYmPWUrms3lG+wpk9Cw0gzmNHUHkUo7zHzhcKkYGwCz5tbHQoi63QubNxbexxm+grzpVk
QBZ8BGCPq4EZKvQ1bIsrP4QShCMx52wuZ7InrShzlYNL11o34t0CpblFJL7oAvtiuvzPoV5vehBB
h4DROUwbfX/oQiO6TTsJoVYVJP8CN7w4v4D95Et+bIZXndemoglnJK2bR5DVTLh1ViSFO1K9hnG6
0RnE6o9uBmZ8zBj7c2iO7kxN+f5PnJ32fEpaRmc1M96OWhPYxi7DD6o8b9xkVL+pNyUiLwZ4/39j
/RQwzey9asxIT7vwi77u98AEDPiTu6KZs9WP+EtJCjuaYdsZSZY9jllC/LTc3oWpKpsN9O2j31LQ
iV1K7riOmrCoBsLKAhTo9OcffRvUx/IBMOPUuf7Mn+2C1Ms7F+bHwwsfv0vO0YbAngjjr1Vpx6RG
hGcLVMXw1a+troFDHz23dMr8ajxQvviM8ABZe9wBg1cZ7XhtUGaefqZ3Q/Fb/YfSbpwaUK0ToBOQ
69vVuQ5gLH3s3oJ5hviOe3N+Rdscm+mBY3rf0gtpUnaTF4sxea71BFyA0F3BIuOGK8MZGeB+vwrU
+77CXVFjwYsBl+1uVTT7h7Q9uWWx8XHt8qOjNix4jPeGEOOnn6XAhohboFaR3rT2L4TSvjL9CJfn
y7UxVm9HWmV4pJBlpvV9MsOKYhz/f0LusIWRubDsGYh1uFXzP8QkJjQESz6wVu+sC0d1wSRoAgMW
h4afCg89Gyqa7X+nON2a6B+q0EkxDPqMNqIYgzSbDs40hP8ApBGx3u6wQ8P46CcdhgGqPU3WWm6s
6/D3ULIzR/G1ayV7XbDA/YsgbybQdHnu7RDfxxtKZxvGa17YE/1zhaJ5iQ1QKnmP4FpYLIVdZZjB
KaCBnZ1Vza1UfuBqhC8yw9J2Qzm4m4xrTRPk/Jbkt2/1mbnX+bqLXzmRbqabvUYKLxgyl1OFakTa
WSFx2Sx3S4QPtJLtFTltv46TKJ8HFlHRicxLpIFQXwybwhGrxQ3JSmpOUQvehHLbzoCTvX8KhRoK
0+2WbPmsEZ27I1wB4Ps7xsTbK4z/MCWlcFCOKw4iDeoYxM8naGbOUya0CctVnihnlmJITYN35eqZ
TmyR0HhKKD7gEHUeUsOQ81M+hUFex9wX0U8QeyxBUlHIUekNgNQT1MGXsq6ZFuNgh+7URlhJNLvy
X8gCr0fWHmvMGLeRYetlGd+9mD15x0mpK3OnoJMmETSK8wilOgYNdL0vio7GyP06M52q+FRfJ1pb
Wa11IG9f6oQwNVbeh2Mc+iMXbM+ivM4JGnUi7tq27UJTXSZ3RHJ8OyKuILJubUCCsZOcIInXyiMb
VgJkgQoR3KA27INdiJSOWCdEVc9q6uhqop7Rx3ttmjo5TbUeNx0g3lgxWCWVgMY3qgG2nWmBvquq
BhZHRRUUOMEDVKfRWP1CvEQbE2/6AzJ0yGXCMUVCZUNZty2wh/Nw4Jfa+RuRfofYrPBwGLCoWbQd
0cbjdsoMpo8wW3BBWGWLGQcN8q8GxlzBfOX6mO9sM89ZVeAm9UrOEUkvJkH6ZT25V3iafjn16FnU
AoOcYvOOAc6uOn1Q66tp6RsN3XbAfHZlq/pUQ9YIIsKbTf+rP1qxOcvGHonsnMtEMj/WcFEyBskg
PWHOVKiKj/ZoqlhVemLJekuzMrIh2yvJI2/YWHNvJRAwtZT8JQrGKs2+GkDpR3G3xUIZd3VbsJnN
04ekkHZOEyyUM7EveHHytHVpxANb7NAU/cxNuXp00hccmSFiSJXiraqO4dm4ENqu1AaH4CEd/EGP
Aobc381i83Vu/EY7yUAZrEnmTLrNz7q8/+0ppEA0w/g6fTNnQGmHVJeWlbtoYh3v2HUMIREkCEu9
yblcVKWy8OnOEeGnpS9QNjfKwqSEjP0QqpEuAuaDIuuxeCYOEUrGy54a1FQnSCdokfiERadXBqz9
6XFA15P/RkjPudlARLciV7DwB1fOdPLNqMatGkX/tPX66N/wk2SVsyc3MIwo/dyu8xswun+KeIWO
KGekyCpJrvflPKs/IKf2Y/gka6YTbQB9hfMEQXV0mOxNI5o2HVEjtm0tLuplq5s/c2fCrz04Ai2z
+iUCtvmUJMRQNeBxzQ4d01ayltslC7gAvHSgoQG6XEYQ1UrBxarRkl8DDIFgicpbv93XSQwXK+lE
bWuCDnbhzBXIYoncHlOHAfw50sMiJB3olPUi545BBeTXLfMtyu2GI9rPSCuIlsS4/nw+jMX4kGgw
/3sASNVcfWMn+9axkRAEf6douNucFO/1jXtGQXNRDC8o48WXVDOwz8wy3RlnN9c4Obleuj2VVRHs
lyvlH4HDOwWOVjpXa0ixbbdkvb/WwHWEwic4pcaaWOQba5hq5KjZIY56qsuNmFhhSYweXt7ufeeL
O1j++KgFcV1T0gyLYkpzkGdWipYKrkdwbwxUiElN8T0/p3GCwp1O3/xvasuEXxtyCsoU+UfpK3lD
Z/Lw7qFYFdaZUnj5Rbt3+5cUa9mcV6l6PWMRoj2oP7e7ngC9skiqoy0+acV4smGHY9mI8c68rXTd
y8mIYseC6ZZGlA5eFxhfSr4/WZwr6I5bFWm5Kmrb5tECEZWM0jY3er82KKJynW/vhI1J7A3QQHUp
GoAQlgslHXuA8YFk64I3Pf80tVLDD2kUfvfQBNoD3ch1qyZc+R8iMqG9ySPbe3wUzqeDO3ebkCTn
jA8GuOle/fEXGSuZyc9nx0w7p3rvvgfbPXTg9aE7rvy2U49tUJIGSARHatjMyBk5nzK+rD8KZFLK
tiIkUmLZ0goRLxcLYntP5Xjstol6shiIxdzAXFvSvJb0peKe/3bg3bwNtLk9Iu5SlZ1ndMyBPPgj
T/dk7ytM4KU+kEJx99nOjVAbVMAFbO4gg+r/sc4jHCWrzKPL4B2Ie7HiD/dJcqBpKmsgFo7vn4Mg
s99vZKV20/pLjeolBdJbqvEoOjsElCNaW/p6SUbBPoHDswH92OuKg8ICC9lmQWtIbpHR7o1avJbi
7rNwBMvrlK++2o18o/pVQQjC9CZ0+mslPtru9X2rMoqfhaHpDN7lq1YDDOM+a1jfBgeUQ3tPB2tJ
B7YkpF4nrnKNKCOw4HYvYNE6Dqvf4H76ejqv6hxRLHcP3IwgbdKcFjPVFq648oIl0CVm3vLYKIeZ
tR1Q9dKZSVzmOAXki2UYbURHQEyMXFvYh5GWLbroSGrxYlHTkT08moasGzVV3cISGCpCOM8OPPqK
SouzGZHoXvMK55RK2xs959wPwPqVJndBUQFUj/C22V7qBElN68+fVQkD0bnsu7jKyIYF/OcdnV7e
YVpjw7g56GvcBjfMTTJh2sQgz5TXlwWSyj4F3rGF4UEIN0R9mKZunA+Z36MAuDkPwqiLE2hHD2+c
8/YNu2BzSBskjMxofUDUVgPR9lXeo7I8cgWIbIwsEJJ9ySeMLeA43GLxINn/njXsHBCjMBay+qUk
3dmlLTNNNcyIx3R4/D2GjEazzIBW9QXmfhlo6qYP7ZLCTAGbqLWwaLRKmjtt1LdzMacfiKGTKmz0
JN4dDP0rMYyaxMkabHl9FY6Z8QeITdrDLdjz/KviZ3VyeEw5sK1Arzif9zsYDSR+g37EbiuwChkM
obLQDVVEN+BaVaj3uNubWHf1M4qfXW3V0wBDCM7k585f4ycdfZlnsuTSZeEa2ZZBEaELCY0An2Xa
eiTralQfz4XXGXS6KFYfjP7Tz2ayCV50qEGQaT6u5w4N6s5ER1zWjV81auMXgtof3yl/K91MLCzt
e73lrwCjZN2X9nBgrv+J0yax5ojd4Yb4be//02A//hRVL64pfqb/Jpel48P69EzuBSdLQAgXxQVY
aXRyiwo0OgZfUXS3xm5IGAMHGTwkPUBiCPTGhA1B1oQFmQvHKEguov4pveB6LcDQKi4gUqNbtt4A
6HL42RD4ZnK74Gam+pjjt1SRqdN1PHkipZ9ssOuqAsJlIYm8teKiT7AcckHx1x4/kvCR59X7CmSF
pA2abFcEUN2MPQ0wtEY08wLw2XzD5ljVFBYh3GdZzdYSTIZaOOuyTkgYZjzPsDYwqj4c3NTW2bvg
vTNgrfK29U5UWBThOuOqGNv/mNEwPSnWxAC9BVsG8DkJY+JO/UYowW6DAXj7euLkeoGmY4joWoNQ
sKsHDgpideIjXofkRRy2kVlmL2BtTeunw/giyBl7vQ9MwUnWU0qP3HutP8fBHmM1P2309Kqsv1vZ
sOKlRKAWsKcCqLaAojJTqbyNJU1f2qX5/f19cziPi4rgtzdUA6uqUoKReRKNLzYleIepgLs//6Al
nDUIUG083x9hP1etypTYK2WKRTvfLKyaC9+8Xc58FDTajKZUzuGSpitDQj4I0NArmKeATYMdstu8
xuMjb5SYpdJ/tcnY4K3s47ZunLT5OGoVqFIx+y5MDDS/dSGsTWKRfWi7S8LLG5XJ5/O30aBhfYUr
KMjrydzhMweb/rIEkvkDPeNHa7oirPkaBNB9EntdRfBEK9Nb6l2CWoadVTmHKjfxeFmb7q5MqQ+a
ibttTNfp+oWKyeF2hfjHR0Q3UuB/dAPMAKLXdxTR4WJJStd+T60AY0Bra41V2bIhLkYgwGK2kj/q
v26vhQSiORElfJey77hRF8l6iXFYuekOp8Hn+avDPs+Psax2idnagp/20A8hVfSuHKdYY3+N1VgV
JeQDA5pUrw90Vx763/N+FHv8jNF3GmuN3SjWTsuKV+n6ijQoxcRkkywy9c9VACK3so24rCQ3y/rU
A1qizTA/Mx0l3q/W0AL0uUoNLjJ3vSc9ZVZgG4HYSXzsPrFdMt0CQRrh90JWReFmhqyxOcriYzUw
rXdemcPjDxpLZtvxTR+Fh3b5E2m1ofn2pumGDEc/QcP0HhI1EsS1PzYlTJTzWoGHQTKX6U+AmThT
Q2QgUCj4BuKCtVnieSeokV3fhjIAMOfb31qIz9oNnOSlleSDwgcO01SJP/NfPiH7b7rYh151yUGE
wMpfUcF2/fSDuNtBjUhZhlAEKgMtxn3x6wlB0+jIsRqi2yETZTlKq8vmjzhiPA+rR/lqg+I7HQG2
7PRYP2bUWRzTzmUjjIXiPkeMc7LJtCFVZJARrBPvwm33qdm2c4k4qPOImhHu8GOLhrbblSKtXnqR
RETKjHTysLCr7pvXOR4HIp/izJbZmivGEeUbF/4VbLVkESRPFzmhGiY9ucn68mTg9itRm91NwUyH
1HuIJB16hjuUtD3wbJ28mi9aCIlBfVCdXUnfRwBY3I1OKsN/01bsURNTY/J+gLN7iMm8AVIIqzJK
J4pnMB/OEgNqLqlnyKIUXFFhbAAVfic+IMZ8Qtiz6nXqxQ8jaGDCqbR1eUq+D9GJiZ4u5YmWrG2s
AGt7AljQuUxpx2RcWbr9NZitBWoPiz2xFjubBWp6oNt2sRRYKQCWnuxZsZTuJRgcrwZPjr8m88cG
bCBxhvDAEiHfZbSWS6ULMwECbfMMRDfc0I/K4of900rGfD5ZCXE5MidvxcQU1vzMrf17G+p/FNPS
a1NNgRNgTjQuVd3pNgr94jWWSoZGWgV63XDi1uJosROlx8EWH2PKwaH9Tx3ClEnfZkHMqWkqNGbW
DggSEmIgpmBx7tFJks3k/DsDHmET3greLpF/wHruKfLQK3T3tbKuAlRNmt7LKgZE5MP4QInrUzgx
6Vra5CnsUrtPn8LdHTfaWDSwo3l5Z3Lrk3nL5bFN/6RJ+rGOiUhCDvHttLmHPxTtkNtSc9SorgVL
Znj2BSA4fmGK7t9xbQ5bc3VIGKqUArUYINe8rrqlJlhtAMPLkvvyOKGgCmeHOAT8FlhtifZcyulB
tuZpfvc0bEBGX4bDv7PnZNsHiU9ovbv11FVrXg8gyfOTi45MP0A2vN/PUKElzK4LzWbNwjZTniHx
J4wdxNXiMbzxLMJY/cJ2/kICTzSxQNbI4nCjdQrAxLabol2xnxwehgobkwPf6/uBSHzrCayeee/H
ivznpabF1rbjL0/c0sgbtoJsItPZIqqtllafDXtNv6k1lKYMorn+NQdf62FBwGC18TSen9VBVOyz
pUlPNiQqVEhJx3FYrsTv35ISkcWWyHFoAseXCOR0bsOZD6gVtMpT/r2N+kutuiFJZlXgIMfsUQl8
slk7Q6G/Lup/y08JL8ELw7RPiFIFN7a6IiGMwiERDSIbdpyhnx/CLXDcCbtdIAU3Jg3hFyeNqvo9
3xq7PazoTtewKNS7yjkvROHauyqszv6G02xzX5BOL/sG8Th3B1yC/vvOjn72VrUL2e6oWqhtV++v
PEyNSx/YDf88hjxLaC0xUJgAHvFeAd4oVeCAMdK31CIt1ydx5NQEoxJKprVJCUe4KNwErjj317jC
8533/JrpH6fPxHc8rfJNym5U27AKVVgKfcgDm0PgWJKNCz7oKuDDmn1/2yfc2h4OkfoTZj5//Gp3
FyAA2isir2g6U/gB4P7AjsWeXAZCLdrwXLii2mhKxV94mYfPt6fDRtifzGCG9Fq+PtcKWMLxkkDb
KS/W/7GZq2l5ryAIi4CFPqqong+SzcSyqt7Xb4poZP6nfw8QiHXmrzme+YqhpLw741HLUmuNs4qJ
tyHqkHaTP1ty9GPSNEuQGsi7DZPfD4f1EGcmn3H/KvB9yw5uB3wrWV9yKawi0GDLxXTGEJvx7Xv9
Rd8S5t1OCcpdpPpyYRqjgvpwUZTTpqMmH+axnt4xWycScPMgl6pXVtBWKkIW6p8JRZm6MSJATAXA
HMmUZsu/tZaidTW8ilaM8JXF7kJ28X1jLPAFRgfnZKcscovNgf5OuIlEXEJguAkfFIhRhDQguCJr
wkT7Rk+PzMbL5Fd7WA+eo6fDXEGhMJXaOcAPCnI49hYeQCTARHAJmDU+iM1OvPKsAUaL0sKE+lJj
sAFms1w4cQG+BsMaYwxc3L2uiwBwlYhCUmPmjLGiqqMDF40OxDeHf2bgr3kuNEdVLyxJNUnrD76P
7zS/JM757oTusn35Oi1y37yh0+OsGqfF9cVUwjT7iozramsQzYBKO2ZpwX02Jw2aF+NRdXWWNPbY
LirZadamD50OMQB9jxOT3IxwzV+hJMCo2LLU3RyXoKyNGd/psM2wKBSugwfweCcEk99aFGTubhkN
EMLfHxVUsz0W/iIlYWi+0ywanbC0dxvssRrlr/w+/JPIr5XbCFLUOdCD7NQONuVPtI8msznX+9oM
hxlbK68GEinNTA4ZeFfkGg0jnaEqsoPFcPnhh4HBvPDxMDv2oImPpjFGeX/XO524OE/sP/zqJrMs
s+NzMcf8WUSEEmt9nPZ8v5cxXhCmr3vNJoF3+3AKV14LiiLhzgkhlD3SFMhz+hwzHV1x6AUktiwh
v1o0WT2SEF2BLSfAe44OSmRY3czmPzSnSyiNQ+HqDyIIvY7g9ONawWxzEGMBSQP6j/DYKmEmow/g
OJetUZgk1uM1ZJ1I39mf77FDnb8Io8dZwWJduJoliYRzKR2zSLyuro832Uwnmqx3C8Pr4QG2r/V0
ktYI6A+b1GryDMt8c+pMlRj7bO9nK+yXIj1Vnrmsco2+KDMlG1Eon7kppZ3sSiMan/MMBYQ8X1gC
r7k90dJwp53Kd1mBMOVjpbkFg2RujoZduQsanMThJNKIfCvPoGlTqzuVE5C1Y9sdEWhpGKAzVXW7
1TPNEWLNgruy+hIm5vn0tIDfAzlZf6OoUDcQM1xm+m8Uz+X4GTfkidT7jSUwZ4gFhOF93+fE4/vh
396S78WFHQLO1kA1+5g0ft5ZD75lI42ko+kgDY1wHu3LLrSOMeK/zKkIevRFFDZak63OcyySUyyU
+J9I3coz5Nj4A3xL4QgjK95mkfacpUEjth3+LPg3wgTzb2Zk6RiHCUh6OZi4FjFD3kf59plFkdOU
EDpIsQEZAjfK6OYZWLfto07wSlevjQz1SBSiwfu9vhneOgFlbWivvV5kk4ABOA0N+s3YE2PYcYjg
r2sp2QJYG9CzYGcQhgrAa/sYatZXwotY9fIuCpja6rx0w+LKM2QuFzoj9/OkT2TrRTImdA4CIaZb
fMmvRdd4HpIVnKeovosVIJ4E7AbzFe533CfxmF2cHcDsU/X9L6AE/NZox1G+5ONrNA9d9P77UvJS
BuwE0Sxpos2vDgzAaAr9aOmuc2uu8gZoIXKOHpvmhLjymF3GkA3vi1I/0YaxX4erDYDNAc2j3ELl
6bWFkAhW6RB71Kf41F2nAb4K3kvC1h0rj8gRreM8Qk0+aBC1TR1fpLkjqpRF7LQkth+u1AF0osYm
3wRGdolQBiF/1M8wMzUFpYPkjfpwBdtx5biaIyqtz50LDd1YfU9yBs00MJbHOKXYn+H7kY3hCxh2
9meSRMG1LTzq613yFaGqjlnQIK3zaCIMiD5WF6IQ9VvVC6E8RujvV/YcE5Yq8SgR3t5bvczP9ATl
JP5nEvQxDkxi0H8050LVD6j1GJjkL/ktDsTzK4qey3nJzn9vM4JkWOKRaW8zh4s6P0HI623IxjXR
s7QPdjsLqq8LTRDAMvH2BAh3wR1vbw+3WpD8Hkxj/7ow4YHYDTuxvUu0UN0jJzUdSBLHlwVuE+dR
r0zgqJdOJSMF++Zj6QgiLZiotYrSzgpp/HL4Vzy0KKXvwCOGh6LVFXdtkBPqlDiQ1vJOfd6rtFoT
9EZiSSzHdizhtB8LhHOpXbVYTASrJ6yC+SQWcDMqEklMVchh/bdBVZohTpwtiAM9AWOvvsOGJYhR
GFAlyWzo24J1C9I/NgTNtT3dPINwMIuZKma2fS44LajFKeDjn9pgkhREsX48mTEzP1TBQ/OpRUOs
t/NTtiWwFSNthp8FcKET66s1XsaZt7qoRc83dHT2LYGEURgas4jTp8KQrqEMalT81gSHQWJL9WMn
8O/UJHe8Ut7fqSdzd+R7yqYx+k5NHpLilQgH3X1kGhsU40wkaR2rTacrbQQMECZhWGjKcfrxZHzB
YIY5bfOW7skixm6Z6zFGwJ5yABVTr+O0q64iZ5N/s3srf7793fC6rmC5Ab4H3w83XovU7l8UYEcU
6yxN7yOEhKkcyEfOYDbwvk6sWndxQaUyS9RXgRNpXczy6H+MH+rkPAR3ykVHn5lI7WeXP2ijnSHT
91GH6gmqrNVKbPWNw861Qr2TENB8+Gs26XyzPt40oaPEYUIxIuOLb7kqBrHAARarjHWC5/ZzJnWq
XAfteq8ZG63H54N+NgIyfJQDyBdqcbDvl29MsxoxPiTaoI7ANnA/CslF89802tiFiLmQOJfLIoQS
TF8rF8rQELmHfRvIBw/3rjs+9nEZfqEAI+yrO0rZ7+lu9D8cPo4Kdlg2MEjqQ+2PaTTyHDgdKAjR
YcXoOFbjkJ78Rzsmh754jo3QSf7/ksYRvc2VbK3a+OY2Pk2X7EdfFkHqRwMRP+hS6hcR4YMGuQ0G
p3NNdDax6H2vbaQyHNWPr9t4cX9Xd2zTZpnS6+B1VkP/W95tF66Yz86Sc3rdNssPa1yrCObz2Hje
lq8Hx657MBhmFA+QyWqy/DNMVth+/MJd9DJmA47IFz3+oI299E2M3bCK8DysoOFL8p1xFLKyB+0u
ljBb0Pc+wAvUrTmrQB41GGMVBsLzh9TgfrIa/QmbVuByqypJz0UgVQuHFpkJcI6qcC4Tqudox97J
aNSJYTT6/ct6qAs3OBPTlDGAuFkZc7NSXBa4PPbHAGWwn5ZWq518tYB2aHGvSzfwCfmBJ8BU7mRZ
8shasggVgBn0QNxR7htebQjlgqUubsQFhYa5cuuCTm1HuzluTTiLnbTfY7cLlUXXaZYphzvwFXOI
7YMvizdFQH+J0r/O4vYPwajjPIuEdcQ89MI6ngyXYPPupWmXPbE168prurYnHPSzNsJS5zApR2Ln
QxAWExGpuLP5eqHYHKXkXmPNNAwQy7kpqsKSOKa8VhWqUs7ztMohpHfa5wyQx7R1IvpMZouTqbi3
FvsqCwEwqRg0AyHN5tUYR49mCcfDgW56Db2olK5hj99VsctkYbYdvGy20iJvCAdaIIw0UmG/MSS2
b7pioRLscgYo/1Gnt648Yb7u1hwphrPCAjdBXpWmHsKdMvnZ55uCq4l62Io/MMPyDPhTYdLmGkhl
cnStoMIoANItqsuLJxdhmrTTa/Xlf0LStDBzcgmZBqr0C83B21Yt40ZW0P9S9VNZPY3M2TNZaIGK
Drm/yAYn+sP9VPIpj6Aia2IN7pFCsGHI/2/Vf8NvQNp52n8+E5Wg61648cqx/qRizwtVDcFpZIn9
JbjfvWXhVaXtSQmQaGNDJQFFhr2NLFAcrVN519K9LCrtXOK/0rHNM8UGl2oDYyKIZo+/eynw4NqI
AvVlGvKoYhSkehB0LArMx4rzELKDLKBxvtiOj+95TQeUPOspWKIBQYsnysgLiaLbzU/kud8rC1Uj
cIjAvUNVzDv5mHy7zGGkstcyHh7aQWLsafhqWfG9uIuBfxfC+CJAGCX3WXu2lORCJrRMefm2Aisx
B35A9CVGcKGFL29sqaElB4VzAtjm9U2l22SFMCbf1+jHy3Be0J6yi9lrnbV/tD/Arm+KTn6WV/Or
ZvKr56rbQGticp5XSV6uZwM0lFfuxD4q/nV25va1a329sy0gKO5/eBZhdoGqBJCPC/LT3jFHdN0C
nPYQjTQ4EqvpejqfsNyst//QEhAtntyzLzlg6Ac+grGYTFMztN/B/qh37YWsUMB4CFNFi5tOHJXD
DOY+yj6IhlUSlsVGnqDSL7y6F1ZsKnXqdKn3LBRBLviy/4HVsl10jcrXwOO6V2skcmChgS3IUDXN
yZERTKOeVhlqJDcplfhxCEvjV1hP2NYCBH+g48DyCymOna2odnOvttHrfaCc7ycoeWujqV5Vxk7q
8pqo/QNGIxMSK+P7HwrQCCPPGB1h5YUC7cpNeQTo6+WKCiFKe1jhAF6Q4Xs/f+RrcHHHpC/yRtnM
ehBJ2LQNQfOS4QTwde0LFMmqVpoxrc7kxpBZUXnZqIanNDyuorl+nYDKIZ3LJd/+TR3rvS0KI0Q0
cRHKassz9nuV3OhgFDp1laP6SfCpDe3l49l9/Uaab6j8DBc+IVlW6qytjnPeyszY9iFBBjKy/jMO
PTsvLzWsMaqQ2xASxNZ1QGEhW4JW3YLNL1+hDa2rW8SAY2nahQhvi7DVQQ4LAhr5hAVZhUVTxLjA
WEkuysDOUthssiH4CJyiAIxmrf/6EjPTaxubQBH0F0PC7CjQUBkWb2TUm7azBMnvQxsMii5d5sb1
2t+xx4tBavMKvVnQ+iPFgiA5iv9vp7J1NXfjb7rjKI0qwmV/9aWWWC/rlMa7tY3HiWhSSrMp/rU1
Jz33Ydj4gvFXp5Ztwdu5PwF98Oht7VNzZPfSbFvNTKBu8dURzSukxrs+gEX8q1O3FjYTuVZMcYVT
aJqwr6DckPjRSQ54J8DSaDeQCXcI9EYx/j/o2F2KwWiGX8xQCDSK7aT+otMmOaJxWOveFCPz09UY
xB03QnE1gYA1JLcZZ3Tbzm6VQTkvGGDoBdQiVEEHNSwNJyjrWXDLvYye0jA4MeCd4BXb/Bcyzcc5
G8mwbreaDuJIHyVQUY68cWbB/7ZyoGINmX5s6bFyfHgwUUwDuCLreFapBqMpN9Cqm5c3zZB6RWtQ
S3JhbQs8xSBNicZh+eAIQdQOCi5j6cO0q4K/HJrP70KhDO8BRvbgmmtl7IdM5aDoFEmTxUp99sRs
/LjGuXkegb0H4Zq5m9GvHyuFoANA5+XQddbqp0s+l3QgqIN9p3NxevqIMP97FRBP0KHti1roM9/x
o48nzlqbJwUKTAylo1uXPYNgLFyRsvL2Dsc1DDkD+7ycYjYixI5Nm11opLb8N1/CLo0awzfqQ/WK
TS54/F3PS7FTbAYN0Sl7ksx0NdeoVM03DXDgx26Kvpq8bNhiRQYj6eRTE7tZ4/3gb2HY36JRl+//
MpIIq1W9zhRNm1dKZQ7O8qgI6bsv8cVU8T9VxgyrqXqHK+XhcUh31IfRDXSUAenUKbNBynNYJuyq
8rVYrL9f0UE1kQ6di/ajF1tuJ9u6n8yG8FABOgA5smW9ZxnI5BNn2X+wLQm1z5G+BdADpoFzTH8/
9WYrfOhvOOlhP2y5KxA5Q9pLKMpfLDJxMUXx+Z5FLjxNocPQDuMs5sk8ojlBaucd0XKCY62/hwjP
Y2QNMPTfG4DBIHH40VrVhXblMPs8+aLUqlvVVvq0WwSKEVOwy1KVt7Vs/GSNxcDFREur8NVF0+Ga
m+OkDtUPVjuOMgjv0Ra/zhzkhGvbRpwqXZ0dPOG5dW9IXpG1g1ypnYjIpf9nIrRDF5FrKvEH7gEY
p7jz6X3Fim632LCVhyIAAzHm5u6JcdcrPfuVhPrAHEu8sk62gSKi5oPGj6IBBdVvggrvb9Xkp+uE
9v/ttg+Yg8AMAeH8NUFagu0hvFLWwB2t3479YHKa/ix+UY7KTjMZY0e2bbn3NRjx4vsv/nLQFRWj
yQ8muYAwLbxoOQViW/pKqWdZzkBp+UN/K/WbQTXfGT0s6lxth3JDzOBsNTu0Qo+gn4YvjVAqUuqt
hpwThXW9EbqerjU9G/mHPlPIoKE9vGJOtcF/cTt3o0heqdwjNvFJb3K87tio2P4RaCcHjsdf/Rxy
f/m6PCf1+MCLjBYE5+4jX9ReBtRN2Y5jOL2GNCN85IZwybvIm9C/jyTO0whss+HL09LiYsmViYqJ
JgnfyEy/2Eu2LEl8Y8BOuCL/7Nf5QZAy8vJxaYVWgId4741l5i1s6GN/EpEcBcbRdA7BYcF/KO4n
ETnDh9ldFHn36agFvf65NcfyBJiKH4hNP1L3cg3cLp/QRdIXlWbeF4i6jZjZhcRXISB6EZBKJCKj
CZq7Y7RNQI0vnB8d5dVdGbcngtnyuBMfnA3E/pxTWhArPqIFLuyZPhmQyPOL11UQR7nfolgRZKcn
0/FbFITeA3Cs3xidEgYVlr2OffBsPHWctFSsGrfiuB7jcILBCrPA4jA/nnbRpFwuMjYIu1WX68T0
1vwlRgEEFp3DucKLx8/N0mjQT9KbdCDyLFkhG9mTOL0TwK0r5uzBqg4zDhzYAlgg19GhAW47enI7
tInAn06sAhG1NvMw4mWCue/YJmos1FRmlRtzjAfK0mA8V8i1t5EGQ+gkSUalcGKJ81R27auuIcW3
MEZaNpgv4Q7i/JcTHA9PwSKatmT9dkz1FWjLZ/foblIN2GZT21h2E18HAAMlUDFelE6eNAiar+lH
tfAvJFiGcXv9FkFzrUez+XLvzeTT9vV+dDbkGCtzrELq10hSFpTks4UztxT2VRR7+kRBK6C54HvY
EQtTa2QB+xYVOsdC4ER4Zn65pyNdtBk5CgRNjMZFvrP8ehuAcTFyNFWmOlu12DaC75KfyyWOn6A2
2HGXDrUMhgTSAquW9s6sXxOfaAHy/zTdRM9CgWhvAthuEi3PGapAC6KAnvaSA9O6TdMb9ba3Et0g
l6hnElyCqP629f82dhTOa+BKiGa+XpVGKRPM1HGrVR4YAgSko02rMjIlobv2zoTUgesCeC0TJlQP
GUXAubMB2+DzoZ90ILPIubR89NGNTKiGSqCHCkO8Zpt9Vx7GUpNIr096r+3ES7nIVF1fbfdAAN9r
ixyKzNWjN560hfFuCpLWdCo3UosCXEzcQNOgd5zcdyudzdJ62e8VWzUWwAx4rjpkklS3Nm8BTn+C
/x11KPDZhX/+v9TO9zocdycA9BqyOIB7YN6a+kBRz0ZRtwqAajbGtlnWCon5jV0QOkdC97F72Fek
Zk5SQOPucY5jW3wYjmsg4bL6BFT9sn8GqsXi0+Sq1RYjEnHWbHm3u4fkRnuOUH7RM4Ybd1plmVoF
TtJrKNk5RTGs4r3uohJhoWt0u+pcXi/MdMmQTFf+4tpQ/64KVqrQho6ngXkWcXiF32ZLXfG2GxHS
XMwvTGEN+Dc71JmkWP9y4XdyiT3E7pMIqXzj4foPId9Ba+0RYtj02y1Dh14JfzGTUCLj1cIl9mWp
Vo4glNZaZrk0+2eOYrMwpr6RXcwi6Ik1vXsiKd2h1hYh0iBlfULuwiPVjas5sQCCM7CtVZkwK2y0
b4kW9Tz8G4etC2jctZoGDSRg0k35TVmIqCkUt9Ik/M5ngxHrHeJe2EwUBjSW3/h7TsgKhKx11EvE
djOynarzzw9uxSWqd42Op/2PVg8Nph8IH1+iKaagEXKvVtS45orlGFHV2y5HDt30ZHnUMxGeY9NP
v3fVfsyzgFXGUm03RGBvTAAnH/ceaKllJjNT1z/H2dh+NMEjhAmQpEJwOPu/YpRHadBZvyUNaRXm
8Uc4Xf1LoNg76LwDJ7MtQ+sRdFTT+RaOOUSbTei2jmno3RcCSXBhgSp4A2Q+Z9o7YeZYa1C27CX5
VscHy4ETFfF+/ucSPNR5Y/wVjrAsfkcyJQ7A6xVhDJOlveDABZ128flGC0GonZLkoj0/8WQ4VvTt
M9aoIGk0MqJbyO9vtlUAmLKD0gzg1mwNEXCtmUs746kG8uKP43iNjSkFbfUQNLb2REhqrE4+hLbh
tK1UZAlgzVXqSBscMSZDZpoQrPnpjUPIPgS2vmve1EiuQnw6tepssO2ICfbZsHMtAfaiPPaBoVCR
Io03ZLRVW61hUoXE5qG4KN3yBfEk/3yhO0T6/myQM4uqx0YGLIcmk+3WHOWVGpveGk0QQTE3aFiV
w40j9dFnUS0LBp+rXY5xh2iMMwwavoQUD57ljFeMefCAiR4k5pf3Yeq5ZOnoyxoWUuk4Xf5JH7be
OVV/80vnZziShZEVreh4d3xtoCpwb23WanMQ3F7YotYun+rG7eVtqWV+nfJ0tgeY9+8V0xi+rSNE
MMmrOnPST2CCnM4Rc7QvHDgqD3xQVaq27yTdryi/Hc50+9jjeovQKrqMOhvNgNy2dPjAP9mWRvyH
1ueIUv8s3YGcrunxMASwVjdi+GHsAwKokdHUObjeO8yBFXSsNVre7ERhvgR+ymhB6d+SA0nXfinF
L8lBUQrozZNTXKrpxqc3UmGjbgOwiJs1k2SPtJjZngp8oV0nrUPJzvx2MWp2iT0yUzpI09mGWqfk
1KhKZls0ASHAAq68Vc1714P9e4WVHSz40FwG3lTEYjSG2hr98cDheo5ZQXCs0hTOhoNyNX9U1O8L
0HFfbNNg2dUU3AGwxvf3N3HlsGfyRGBbXBQXJelSHoEj2NGNRQZNYJ9bGLftp531hGAOyYzrXEZy
9jHvvtGBZtGh5zcFmyaxD7PShDqS7rxb+Y1H0QdkZAmIUVdQhs6PpiZlGz2qusnr/6jc56vEJ7e+
F03q6awOWqKEhtxyIt5X7fOoq36okjBwZS75RJsipUglFnQ/jJdbHLq76RL4K6UJah29boNYQEyZ
LSDv1ykHkr18shN39ly3SbxTCbHELIIMVD/BpxZY+Ff/QH6Y+hkattW8OPhrf8moEOHNcow+XMJJ
6P6UrahCMQpYMF0epO8BqOdbzyksGwPZBVDUTrFvusxxuut0xPV71q8udCWJAy+E6EuFjZ42YSNz
MTjAYye7a2LvvkW0W7nq+9BDpBELPJ6Pki1HhWyCcRsUFeKmejDkw8ReNFmrCjyf9SIKb+pwegem
OcZvtkz7MnGqtRvnu8+M/QzQkEQfdWyj46s2YR9B3U3gIq/PsE7DwR9fmRgW37n5mwX18GgL6bUj
bHOSP8q0J62d1damzVeFaY5FIG/iW4vsWy+wB8ma/YFagkJoR/YzGFgBNPOfVIvtRpgsxys2eiEe
1KU4XoIYmiHWUutlkCOyDNTo0Xya9DzOXkb6fC7+OnaORfXFUvx3IgpL98cLAlvV5jcE9MJkXw/G
EF3OsOhx20pWNJJS75/cOFZmguNGV4lXCqpoUtGLFXMuf5iWs9i0v8fz5GLG4u6aZcUtyRTN6vve
uSYRba45zns4yN9PVT86iAjxksPafbGx4QjjOKB9Cv19otsmimOrUEF9yNniVbDejuOmJSEPUZ4E
y5ZEhvcyfloH02E+krfiN0yKV9nah//KdiorlGWWmPN5Mzq+ekX3N/vL5DLR+5nOZ7v8V3Yv3OSQ
OesvPpFbVa027HjqESGo7dTFJu9zjM3t9rLgmjWKwtaf8AXBF6a1cYx4qjnyKWXFCD4plfercuW+
phN22J3WJEfMtvwnRh490aDJ+6DVB54odKBTd/VI9NFQXusuEvVbl+3HpI+3rKCFN4A1ZOWRLMhU
UGiuMR1uds08lyB6DMSgRnZBmVTfVmBVoP+xGx99wiSBxuA7e4oOqll3XivweX4laj4cbMYNpg8N
TbH6ktMdb4DLA6xEahjiqx7MPDzfrIplpvhtDOoGKWbzN0G/fPkI6EiBQto8x7Thc+fwgp7QYW7b
aaPUYJP96oSOOPJoULEO7TThwZo9WWhK7EgVd2CsVqS9n3D1a+9eWpXOuxaTjkwQAbQ8nbg/PwAq
1d2QqWCC/5YdCf2fmvwsmeB3k5d9iQu/tqrxJ3vBnGOKL2VrLonBwQjV1AuqAQDVVpGAxlJ2yu2r
gYgeUbh9d086CX6drw2kGpVuYcqw/FW5xrrIhiy9v51rtRiCvBTMukNycF4x0UrTWbbhs12BQARJ
v+4LM8PJ39WCs+MoJfEoFWTePfS+EPF5+tgthqMcs49hwhaRe+iBUqoSBQDPIiCCGDymnMsDsaYM
zEbt5s+V8AYr53adSAmz7BRXVftYWBUcD2nlD6iuXmHZtsqMiG3wcOrgGYJPyebW1iaB//oWVYWx
IcSm6guounK60ajQUGECYXw/IdtMkEaDlX5shh+VnQ57FHvVvM+UyTsd9cBt/D0qaGNBs2K/jOjB
UFBUPLFtMEJzWnVuOUVAXwBGtFrjRArVIwrT6UsLsbSN9k6ZuzDnlSbJ0h4UsJ4/tFDyu/0uX5VM
JaCHYxpstvqnPjZsD+rXKPr0UYi57XxS/guiEKKp0Anviei8iraBNhPpQjyQ2Jl49jsRgK4PgWtv
dhOwR8JwFcRyihjAPul81VGEVpl7X+g8VKRWBOTg+gBQUJc5DieWlM1pOBubHfDLRNRwdgsqWMTh
vT8wyc+IzY7GV+bjqb+uDNNBWDM3O3Msyu7vfTe+55L8G+9js2DrKmEN+njQVPVsmzPNX4g29ZoX
8rgbcCY8Y4XTRTDZdqjN5w/pz8TqIEsSxoo0AqcIvLVESLRmtS9a3PvUkoFgnvvVV5BrpplDL9Bw
zlG2pRI+WA1gYjkO6Tox3KLXToWB/8xbl8Lto/0t4E8KSfrwQl1sXHbcfdpTzS4Sxg5qBawzU6N8
cRFdFHTazwmzNmxWnM4qoBKuOZXUy3YY6lE/5FIS2SMsyqaJXDzj8M9py2Cuy6e/CF2Rid4wi9IU
hTiHg9bRSq2r9XURKhZLTgEd8WpeThuqbN5l47d6vIxTtTUxKcB1pit34dM3FxHohowadfPa3u3f
VmD/TsxdEZKPTRtPnole5ZY8aTfU06t+o4uE3iM8DZOOYkl79WQsmE6j06//Va0ZZK8+A6UyL9Ch
qqCVRc4dhxenCbyQ2qKaKci1po4Aip82SetZKIMrrKV4AcmkMfTcw80w5ftApBHVUr7EHh/Lz7zK
HLlBWmhrydX11dS8a2rEP6z/IJBXfeG4xyx6RmyVd86nk2yTDU01x37TdAnW5Vp4sldzZCP4jqu6
usF6NVNu/0XKxLdhc4YsqVq1p9yyA/3/EwjQv/XzJMex2BPPpqyeRpgkuoN0AZYmjH7YbC9jAcOn
FIu0t1cM6GqjEkCg4agG+8xTtvD2uWI++BiAE/GMQk0f0Jb7jPqjFJ2fcb+mBSzZeg3leKQ7yDl1
9twFgs8Hqe9SUMBWOJ2bRK2BbusNCJLt02cM2ABv9tuen8II88AXlr4Erqp+M7ZlrueDlR3tdNeb
Vw/7M9KKhbNjlwjl1t0XwCcWkQOQaoLEmfnxqdt4quXGql1xGSo2OHZco4wwvtUYvMBkv2agWRMl
QQMU4sNwVdqPxF8UcX62wXJ7SH7aUhQ5/ytGq4YUQ/aX6iCgDMaqVtdBbNaQGru8HlpYUqXUWfvU
cvJppy6qiyhOGjz9aBG8vWJZ25g/ZJcAy9b6Ow4TOiOb1W/5MMZIWdpvJ3p2ERmcArp4CaPNiXKi
LMBlZVjNRjjJli/yHN0UHj3mytCerlcEzzBS1+Pfex0Dy0ow+mLbhbYDvh9KglsxtIYa2upvCznk
hH+syf4QwOGxRiXjc9p7ekVPGl+Y4cy0P8O7/hbkjHCd7wMJ+r6oZCrxd65P4ODztCScwhqBGzG1
Pxg6QagohlAqG4KjBnV/HxidMXr0dNYONYqqcjue8hNirzm/nJdtMST6jrqXJQCUWMfVXpfCMgER
DuHzObe+YHa1YXJG/4G5SpHGttofvhGQG8ekHIj1Mg1E6RTr8Ada8lvUENjaVrglaTeDdyR6fe47
waQaJnU2sj4jStH/F/f26qR8qoCcQ22k7KeQus8QkdF3LztW0PApFFaQwyzPPjwyqUwR5r5mD53b
ouIWiHIsAs7DPx1lLU3YLiiek1W2uURmQDgS+4eHfszFW8GgFTP/fh5LoUYnPgdYgTx9lIdlDE/9
b8/2WoPeF90MF0uhMFNhPeZz2eMZI7/5iazQcc2Q4qFloirSgnM+NqboExL85rwlR15U5AloXTLW
fYp+S7qAR83btw28SVMwiBoYHyFKzeI6t37BmEnuv56dZJvNgDlrzhooDZ8lIqqvyj3DKgD3XabS
ODRkxkHs0YIm4ELClJug12zLZ0OzDH9kn86sQa2+u/q4pgpTy2Fn/0OU7SWcB9mAUAhy00IP35P5
u44Aux2B2+Nb/fZD9z8qfdXBuY1djKQS9jvx0I6GOdn1UcJtFl6O3GAYC/ubsOVscBPaNIPwanQt
qxU1+3Bl3rcQrMxlnXXVtCL4hcqUOyATK4BEzLyaumCdQ54iPYIbxoD51TufHXYijIo9Sh8WPxbH
pZhekyMO1XPFr3Eu1lDfxRunjQNZhHD1X+nnPiAbuvYtAtR1S9Fp+nhOKDihU9GplLdGSg1gY8NI
p9KzvqPNe/KiBdvRdDa60PUiZhXCZJgd+g6Rcfz0FvCAku4dy+Id1t/xyRnoxX3ikINQCHCreTSL
oJtl+JkyUQ+052bnBb1+UtSpOy3hC/5ChUMU7T3GtO5L8Aq3v44tlHJCjidugJseKf8Ea3KOI+cj
GLm/admqFC/fg3p96rH3TSi/tBmaD+voa+raCc62VUNPwcTeGzFiIBlM6WjKYE0Bui88tFqR7WEO
TkiGiwTnXHWHftrrwsjwmMcQ2s1dpBZeTlMmPDs9XG1QvsCoeB8DrQ0aR30I+4KRfngrkptBzQac
V0ACX3IIMuEvCCkC8nXZQIm/OPO2L88snBJ+DlS4+QbO1c4hmqbZryY9lyBO3kauLNtEjJ18TsD+
HLnaHEVIFz5aA/FqPj1+45+jI66OEb0/auRJouk4ZG6jvD6smAOWHZ9FNy++rI9wW1uI2v1anWHd
5+0wdmXgUovcriVNNHR4jjBamzVyrDeFZIc/nwpMDhW6uy4TizL6CN/QRIfZz2tF0UwyuM1RjcW+
azkVOx8igjnLBs+xFy8/fdgK6czEveiEty6hNLKvIxdh+VQ28CKzGf9dYbBQnEdq5Hhnr56EI9SD
EoaxoeBYdcVKGFnqIVDyInLy9MwBNQcYnGcB6tPNui4a1akBmqKHg8xXk9cS+Wkl4nxyexmQW2lf
U5pQ2iGOEGBSmHUncUE1kxzcidiO5xkz2RXkLpnytqrwZE97a9p6bjhVJ7XhbKXq7nCKaWyEADKE
HWhn7uwxLaQjTpr/StN256Vao6eIR+T0Wb4IkS9c5xsM+7St5XYt6jQRzeCA1ik/ofNdbyOHc4wf
d939qkT+jBhHz6LEKjYyePPa8TLtO7u4QE+4aVwmJMTBe0NKEE1ln005a4qfSdekzRBYDGpwaePx
q/XfdjN79dyao2H9Je0WExqPgfBtTDohATGj/S3SX+mHcdPQoqEffaolsUsrXsNwX5NqGuIlmy+i
lfVzDMaSUHc/5aLMznDeRQn5QrDoMVVkO9AcKOTWR2JZl6GjuHhwfXudp+TpAzc3R82MyuqKS49i
i0S2DmXk86HQ7GPxvGlIj8tz/iBa8L3N19lG9mkXUQfT+110+DNiH/mOEsKtWyMdom//bqTAycL3
dqm/C1lbxWYC83vG428VztumQo/sbMHsQ21F6UmJn+JibOxU2vY1eT2AePBuXCRjN56Rewv1Mzsm
RFGRUn5spLsv76gnJji5Ep403+aVq3jZDLeVuRMzY53tnDmdVQ6+FV/ppAULugV9CpTHkLwK5RNO
9eMv6umwds4mIECpAcOPR0vytOnZ0X9hI7FwP9inQldE2np8AJW79k55nZ4CGFVeZBqH2qmgWQwh
TGjs2QQAcnBfdpkWvzm4tTfellh/uXMMKErSJhKlngsxnSZJ+hFhOr0qXQ7dl4slk9bOIdpjd1CH
22XYPwEQnKOTFt+901YsabA0d4xUjgZgjXMVwLcnjKfXg8i6OKWpij28fTHrLpvYJzARnUPdozkI
J7JSkSFktajdyUEDV/VPolLsX6gBObvAAX+YRpzMhSZjJjPuEEDZ1dHE9iYCF365Dy4ros3uWh/+
uE/a/cvPps49G/wwJFzS1DJDDfuX4FOgOn0tzVYMyrQN19KvTGAe3DN9+cQVWabVZeWKcRbYowbe
KjEgyyIl7yZiWq6milZa7fls8Swe45xMNWU+F0HwVswmZErMaBvTNCODGSVMHrwl8KINeKiBh6iC
RtoHxWmGG3v4ukfnbu5K/FB84l/ZZfUGErK1UPWb3fyOXziipCqkuSeOd1o2N5zwTrwWMiFL7F9t
sH1932L+BIH1eXw6HelO2O7sv80VXguV2/UMsZbo4mRhAPMIudVWTMR3fMlJbLXl7Pv4j9cJTo5d
JXU9IZgNQtEcUQWdJ/SiminQQeznoBnTrRU8S1sPZgm0IDmg+SWh192mfFN/E1KRfEl8E3U+KqhE
L5LB4ptwjDRvVcqFEalKsW3ulbMImoA89B/2oyCI4eYhm35oTTy/oN+d0eWtsrO/jLikZhq8AO6F
guFYzEJt8pduKbbyBa00xnR2Rj/CacX9ExLe6Gf/9C79VJuvh+QEFqOPXtnAjQz6HUOygEVUPDbq
7uzHSVJ0CWWlRp/EpY4NTg8bAlIaicQJDzh2uyJbUJmSzC/NaviEWWvmq1WdeEFzbWLeUD3DB3n7
b5bwE3mlshbBRhlYMedzeAjwmgDpMrwlPD5gMic4hYiLuwU9UO1i+kzgBByLRmC3PQ3ICvxBG7ww
O4WzLVD5UpokUY4nRmCn7Mbl6rmFoPjAzl8qHalcrp+9CdsYpPACrSV5Pgma70FPieWwsYJdJGSE
Yj1ekc8oC/GdeljZ6F0i6pFsg8bzkZ+8i0us8No/5uKi1Vd85BHp3rYKBEh8mBh+OIOwifod45Rs
scSwmEHXR8twYmTEPEIuOvH0AyGTWFZEzJdfE5zoJpqIVYMjzGL5A6wca9yvZiHLxYg7MKSZIjKh
cjmIMSJtiCi5zwAPo4+gJxnpQCwmhzOF4NLeJTCcSug5/QS7K9LHrJIxfvBmw8dOZoVM8efwBk4X
HDqXeATwz6Ea+gXIstOn2AYRA/bFLC/aZkzuqWK1z+/uMMtyuMbIxdQXD9bORATZckQW3TJNp9of
W2eM0ZWX0QQpBU8ycCuZ/IhFMK9bittHqJs/BQlKAKBNNqOmTehUQqAljJvOGjt47FPeHFWzyeCZ
hSRb4JG83BxopypyXm5/rvHrFnjdGF/w+Y6kklsTeG35nXojlAo8tB/s3eihWEjPTZlFN3p3pYx+
ebDeQUlufAb5br9jMtNjGdSRmcCFE5u6Y/cLssuxv4sEW5ftbGzuYEyZGQOZg8WuEqEKjOjeN8d7
zd0VKmHQFZPqDX25xqVnMJJirr6IrE2EIJWS1EljG+EGJ711CVsjo96OgJ2Q8s2K6YSCdH++q2zQ
kO06455DvNW41UNUvIcyYz/QGgqYckNGAxqVSSEJcZg24zTMe7I242PAnRYVvbh+QkbjzH6l9BXk
pkcQxc7MOZk4nZ4M3+OEVLZ0TIA6QWGLL7ziFfPMWKjTj+PohujJX3OhcqKb6JdJJD44B8MHikP2
Gj/+QMUBSmTsblAIZ/yAu8Gyma8hh7t5qyG6el8z89NlRE+cO4TyrHbI2Tg5BuRS/IBfv7BUvRYe
oW0Z79BkpNv10ClwCTOvtPLi4iCDxDasOX3TK15TVPmjsNVv9aoFL1c8VmZ4FlAvBC/QVDEeigU+
Jii9TUbPg6fhrbkuvedWRLAGb1R/uQahEukRgrqQiOfhCUJYakYWIdnrDNlikhvwl7RxlEXq1rpt
bnMhVNMLk9PRS8M90GxsJBkaHl647NvYRJvtjT7eHYLvhBY21ASAAWj6+x+PCpYZKVo6w0AeMMUJ
xIpxnDcjQSv1Zz+XTepspHQxIS0bHvdZdQRj5Dsn/vmBFhxy+3KS7FdMOkqpVPB+lvHWe0DfaXMv
HcjhY34MhA091xnOPWq352NTN3PmUXu9knsOyP/UXykMszJ0C914UiLDJMP09gPjBUeTzN347Z23
xp/YIGY3NiMUb7S/4LrfnFqaqUYfsnkj7VopvALhSBVzyWWy/n2W0+ymPOW58oX+FXbclfZEJX2E
CJW8R469Traqg5X29dQcJPjkHG0dip9YhFKcdvTCqPdeO+2ui1/xwSm40DpLYwfIY0rn4jWh50SN
JC+alt/l6gA8qeEZIqB4NZ64552bXzAEN2iUygf3WHcFNtQ9e/i+v+uodB8SfuRPSNeygQ/gf648
1nBibVYtYH7K96s7n+Bh8bKukM2WT2uARr16lKX04aql4krxBrc4iGbWXui53W92yqyX+OI7HlgE
cxIQ/dScD/lMCtm/VIuoywBPO120Ip9ZioE3NTQ6Z3kCDh0rxdfP80YFf+mnFQdol9cScUEWM0Ie
x7pxpdRSa5hOV2w9weZRn3UTaiaxQN6d8Y5kEuFRhJvv5wFWGzE/okp4LEtaCoYHEuEHUNR9+cYX
zdSFadg47dNrba3IrFLQ8Gq9rXD++QlK68H3zfnifdbe9MXzaIc5GigSk2UdoCLw/k/uF4Bst2GD
tLruaNMl+oSZrLeSng+5gNXpbd5ofRnnTRZk5pmrkMkaQpm1AITlfDiiThG1eJITFAghjmoDCNMv
XtNW+ey0D2A7yCwUw2aWnqXPZkzpBwr48YUg3QKLawfzn3w5/5MWOvLcuHdmuhODsRGtsYWtBjYx
2mHeWCjM/SEreivdgnWjSbx6tfRs6CP+xWDv7rR2RILQBpkQ4NhPf/QBVxURPL0sVWvHckDCO9CC
v7dBgSAjgGf027YuZIptblDUE7JYiGZWh19XiydWrJ+vBzZuq1ehnITpn/chXxhSilEAHiCV00Q3
Iqy975v6P022fG0p+mN5HqFH6q4DuvtRAlhl/ybIE0oH2fM9itTkQy4efaH4zYGTNciiJTcTGaHG
XpOVUB6MWmedD8TvgB8U6qI9lA4rbFw0wKujV+3v8b4Z64yzg8pCqIogThkd6fSfBN1NvWbW+oR0
rW0y/g4/xV3nW23pzHL9mPl+EgFDBj9+TRDuIz/53NjyClIR6sqE8Mem41PtG6wRCT2VkjZ+o+KM
etpjiQmjU7UeWxhPu9OIqgfdoRrzCmqBCOSJ3YkolT3Bw1p38aVyechoUxYYEOr2NcwDZngwxhJQ
kYHoUSmKbv+920ncrNuIbSLO/PPpFbC06zSMUmAmz9/6zzXZLnM0Hz/m7zFDKGH0HqVjhrw4dsgZ
/vMHN8eIXEG3EIy7nfzRt+9UXB6k6ySYSmn2IGbWk8J2GyWOQnoamrR1Qr9EjKqhYtLeePxipMSO
oCnGVw37v40cNC8JsIW0GoCKAJjg28Adsby0JgEcVOZXyQFOehoViZ+xJk73MmkgDg8jxE3pW02P
RQCnA1N/vH9oDxFE9psO2LzWvflXAx/yJ6mKQuZ2rHzCO/y3aWnc3f65OdbtAPXCYtgr7rt7/IZF
043oiPkUj3gFBHSteZ7W3FViP20uAG7KhEdBAEnGOmRDWaACd7HqgijOqdqufUCHwNr/t9BsHx8u
1j9ZAJRQXiEpeh0OlsBBFRnsZR0I+r4gPm1PTnWw6XL3yCuLpq7D0qWkDBrCX7DJwxEdrqZDiOLg
8JZDkx6uxW268E33di5x/M0Cthyq2VJ2cXx5lALzhoO12ytLywv0OlghjXSnAsLk/47DRDh/6AhR
puRSGlSlHWDVMg/tUJakKnbv3vXdKN8r6sROpAlm0yQAHsvIFpzDVr8pKjHMphIYwvWOHt48kAMX
LwEu+Z18Lpo8FRZouekAKgmnCGUbsPGiGCwXdseNlbORh4ZQH9ioRZZXRfdEHfIlBLQUc9lvgxRw
O4Op2W4hTrb5/IlXrEyf94ld0FE/ey9A2Z/D+JVIbXOrSfhIEyAe6CnJYGJ4Ah2LXfW9JV8cOVsO
08ERFhrCPp6BeX21iXfRI4NgPe4tftYsX5BZtR7VsQL9V01VX9rayqrHnLlciNOalfC1cfsXFftl
YrIk2NJEMD60jMg91KoEfS2ZFRfyG0IKeCUpTmQmscAozgkxMZfKGWZT58zTRpUrUYmHHeYdCPGs
329aAd/Kn1VQzWIy1/Bh1uIvISoqPE1YdXjxMLyBBNhG9DnyDt/GI3w+AabtgCQprIy/PNp2yjRV
CJdYxK3faUTPStZ6be4zQ64nFVZH+3OSBtcE3fFMFpjgUdvwKGHhHGg2A04xpejnHPnzxFjtUNmX
T2++YnZ/NDlPKI0ak1L+RZF3/hkX7yU0jSeeYVF9xraxYMyQYpO58gKbQ0vtzvG9Pb7dCTFaiQKr
plcFmn03C6xGITlNJbIOO9uT7fIBNGVKzVaHpBLsl5yN3u2vfRuIIXh8IW63GdbJOALu06K8pmly
QpF+KTExtP6ABkoJ6pCwdHiXImBtcN49tj8vV0rKsPRmP+oMh0BJPf1awUxw9aKz7NorSaslRNTy
g4BVDTaR/tobzmKnRFfHH4sqsLwiPiayeAxz45jl5Rh5KYU2mgqD1vQUBRAJ4EwYwJ4GOK/xT3Lc
9WS54ZY4iERsm6+z51nyasJX0fuv+wn7/UYGpeIik3SbTOcch9HvY82gWczbbY4IZUedBg82aMpX
VpmneobOvgq1qjVBbpKVN62WvNs2ug7WxuI+ETUcN7xF4a91636bP/9+kFPseOAJQr6clawO8qyr
EK0jDjguHOjokXscVgs3kdBGlQim88z7scvPoeZWWLXEtBa7bjgmXnsArjlPLtGfBBxnbouOw/73
nnRVIQjPt2xHrWdD5XLWtuPXwZES+6jqE5cjsrlAdEnfyswbInJ61i1Ed3vVuQLGgul8y3boxY1L
5OirWKZRIzpmB62qe/BDElygVQdFcI4VC1Bh39FU2EX2NXGYB/f2zAoGH7oUZaFhU4S4eBzxmvAa
I5/DcsYfi3xHQsie88uoy9ner9NmghSkqB6iYU1shLw/vITo3MS1ZNHSIwK/FF/k6rl2yndZCDfR
diO4enPhFEf5J0+ulqymFZpn/DvxL434wzV9zhCpl3dHXlfJFuofUPsSF0XEZE3XM2r4Xb1ztfUo
2gp67jgL4w3Lqj1pfo87TsrqboLFpF23hwPZK6NC6NglepN2t2tGq83CHy7d/OUreOOWWM002kJY
OiXQDOQBGw+qImKtDUmqZxLHOK+MRTxdb8C/lJcxpe6ldIEcfSr4xxKQWVFf2xMgqhyC0axrum9D
q3kB+IF+2WmzFPvtPQH2VNJhRJuxP1wZzyVKmQ/DjPE07hVxMXmmT/n4paM0IBICTQS8I1vQxIl+
viboslQH2xSlh8NarXRPL44nc3yyFBcs94T91gUGVjTTtxLSlPGR482nQG6xbtTexywFCbFRRwFw
163wZDffo9soqd2wSs7Uwoe1AI7O4piPpxINWhV964yRHDoqUYypLt9buoV7N/QyniB/gbNaLNk4
uee6XPtJGLkfMak3OhoZtRLvTJTcM/kbG9Us+UQi0DgMnB6S58ysMayyFxc7aeuWQbc2nupzNcgH
ieo1PakEGR7Vs2bdIzELpBE6MDg2XgU75M3Bclu/tVaELhhoRV8JbQO5dakX/TVHCKbeok5S4REY
R3VOOTPd/khdsSA+9moGbqZ8gxkZUoYPWVTPmFcxHTcJ/B3w5LRazWriDGs5SPmlVNNxzS5ukl5l
kOiZPbeTScDA6OeFxwlH6C0IFo2B7dG6i/UucA8MsPpcpNy1YV/kYUvWNuT/lq7u6ldYD0buK9oH
wPtoeJUl0kOlPV07+aldNdPEgKx6c3f3MzF/brtSOnrZSo4kxa7P+Ss1AY5irN66vB3z02avR4rc
WGsWNlaHQSpc4OInYgYg4H9WhvwzUkTTNc5TFDx9I6cbPDJa/0g2T+2E8AKkFi7ky3hPLIb0l036
gxy9OCcuQOqgCPfih5Skmt42q+qAhvAWKfM4s+q9Y+/wypZaFiDPczwBKVeN0zP1b9kipt+6UttU
lrSgJmIwJqsMCafLCpMz2IKPR8AF9tN0BzMm8Dv8JVEscPLhXcSWE+bKUpJOmkMPqHru1ZSZth7R
IeNuHDZaTkP6M3/HWLxxsCHX7dVeDm2kvQapho9KCGb8FLmfWtrQmzVcuYDovXiiUJA+pUMx10rQ
Sd2xr3ThtSPq5gk8yVSq10cg17wZDU+KTsPNwTdmpkP9xgysdbooyfQsFoFpYxF94YHIGQcoFeMX
2fDIRNK2yvUhWYqaOotg4pGNc9Wb5pHgG7aYZjx8fBiTBmKU8ERzZqqlyWzhTfhgbR3L5rXgg6UC
1oFy0vjLCYy7zQt/ho/oGKqaEdngp77jmySsSEePyAEXfe9TH1I4OtXCLdbbs65cqV4V7az5Ib86
lsr+lmsOrfyA00BusB/FZITHeqk1wxwBTKkniMKvd1mRkVo0MaWW3wHGl2YMrvmANFoaFKA4hH6n
tWnacONXIu3P0TpHWz2h50iCji4arXYu8tXo4Yh9FoHDacccr1HLqfLKswPHCCDksR7uc/GxQoiC
5bJI4PES65GbfTRZ4jkIIt1pEDa2paqzfxItSY8p3iDxliXQDTzfOxEK8JLqYz8dq1k5tCqMNCZg
tTKKneue5oJ/Kz49w8RsM8YuMPfydDr0ryGKMKkfiFDVdY+ugHejDegA/bOeAQ5ZeyZa8YQIZxP7
3aRsVnYySbXA+0BiXQrbl2bPpFHOHrVDeWhiGEzo8WoIgRe6eWEIUK+1eDvmFJKOks6tnGI/rKUM
vmx7EsMODWoOGZhdgNOmcnOo2ulSxvTwth+5BwIJ//Zn5v0MvJF6USic1LYJbmvG8jECCEGkzg9X
9BArXA4YuiE/bdsP2w0Au3u8Gr6d5t76ncsUGsfSuMSmwCIJeYDKlcTpiovwdc95Iolf9HTdsgP+
jBr/xhBycaF8H2Kiiw9kjmKmRPlnkvbaQjbD/H80/q98Snyc/GZldoukxj6lJXa8tA64kExYu1Dd
rfOwa/ZodvZOalp75BXQloRjm0M/2j7QNEaHm18cbzQJYpP3Y/OGx59Q8Heu8u9WmCBd1gPCaM+g
F2mlqwfeih4tYITWIHQRYFTCPb+0RL0O1cZ+GYfj+C2mq4MXRBzr7uaz7uiNtEcfhAbrMIgiXcmz
AWqinZIxqfJviGoi0MCN8OEmgj/6NMDANEhLe6pbpgiT3IuJY+yqaykRNGoaVHRjVBfL0uYmctTV
wRSsrC+wQtL4h0hRSj64WHDZRRXJX4lzV1sl2gxL31NhDggDLtV+yk3ZHcEQm3xxbpTs34m04jlC
FGD8xSUYs3Dk7RJ+s1yueTn/toPdqeqWaPWpoO3MJz3hfujET/AnF52DYDBHo83OaNhAwmErRzm6
PogbjpNQsOqPLlm2/mbhZsj7JniDzVDJbsggPgYStd4lNnyRZYZ2eniNP/byA0Nzdz81ve17W/n7
O+v6mjoLn9iML4IBXc3PQLyw/3XU0///nclO5QkIkk2d+XDjgk7FGdqvMAPiF8PNdS9tNqhVVWWo
UDUg2En/OBK0vfBZEbS68kGHCafc9mrzgBr8Nw6LlfvB3bYmKKjXGzHCV3ZhjxkrB3PyMEW/icVB
DivEOJ8aetCMJyUY+nS8bjSn2U/q1SueDPAgSuaaHqgjpPr3DQ3JNEDa30WwlOOLS2+3WHNa5zvG
5EKsPwRuBuRgHJlKfp0GfBv+LD+xffRAG7SLU/kGZxBCBNRnBOlTWlrqNWu3vmgkupHZa0Dsrf9j
OslJlVOaZgcJqaTfi/injWwq3HZAVa1Qt3vbDn5NH7gaP6qQtZHQMY6S8kzqTkDKl05MTAlGY+J0
nFhxCJFolYAPmaKU9TJtcwn7BX/y+VoGVTSv82B4wZJftjABFN8ik98RpRMV/uWT8DYRoWdHZP19
d14g4GL1m5nOl71P1Y1wxsgxPw6t74Cn1IboI3x/+sjezI89diuf+EAp9T8vjMzn+oQyjFoQRV8e
sKU/5np0VkgLmSUmtg62fipZsbQ09RYFdpJZuz7wuoXcblt3AfMYByfwpWJVrR3L2HThKx4Mbwd7
ZA2w9Ty1qZ7wra0qxqx/OeYYN+C9illZN7DKMTEPA8PwcgjeiHluba7j773oso7ZZxHNco05bnUf
O09J0xMYAV4L2v761b9usPwPBaUzGO7fFML1hn5bXy8MPcgUKCtIOvV6Jd0e5r8PRIPhapG5wwEp
Hq8X1/BTYK1wO3kDDKpz2dDir0WYeXrx4u/DESJeyNkaYbCL/jCegj0jUOmJAWtl9MkAqfKmlEgs
/7zziReTb9lo/LbrmiN8WcpGU/B6ldUoUrIGYGGd9Qe9tYemcJWFNvfJhBIJ5IUUqeS7oA9Zyw4f
P7fXPErDIKegXIPvieW3Rkv+AeQMmGuVjhqYfjFFpN+XyEKvhCSvb5i8RwZ9Je7Tvaeh8Qx9eZxz
gZFyJ0LhLSyKGMKf2R+gZiJSZHLT3YYIBW8aCaSRTv4dtDNA1EA2/Aarv+WDMKHOWrKgRu8aHU3m
svWRspIIW8PLoAe0Lp8Y7f5MFtJw796diUSsN+GqBMP368NmVJOanaabLqsGpuiU8ELXlYtmSYMf
e3j1lgmD4GPkCrsl1J/L8mHzGmK6t4H7FFlbs6S5DkAygVxEbYJOmPHDgQYKBBJl85b6Iv7SoLoN
FgtZAasx2GNO1xHGfN6dwNJrKlCzowpPEUVT6e1wyvnnYmRCiSN1UBmee+bBEf1polj/1Ku81kKd
jRnlSAY6FIQoJH85AaydHrRGtCtjuAfTp4LlHb/5OW0iVAIvp8OtF+V8/F0+8Cnmc10LICcFvi83
mc6AJXxWCt2wRXeBP8Zkp9epgLb3C3b/45RX4O8yRt5u2MDBaDgXi5ylL/ewc9XPnxWF0cXrl5o6
2Jqvo0+/vF3D4YaHXhduz0sc0GW8mQlpNLykUoHS/xppijEo73HdxgEhPG0sml1p9tCzl2Xl3VRn
OGKG/PfUHWXBlTDVcHdJphR8PNuPXwbM7NeDaf6Du1JagrwuxmWP2Hu8HfTCZQRh+75l0hO0X80Z
g4psumumJwYNin1Fp4tVI7ypNkQWkhQ2HLZNTbVecqwbCgrTu/fh1LG7PfVzDsbjdbQuHQWZavxt
rNgVYRl5BLpUq66Fu3nH+d/qUGZDCEONf2xntD28LFSOTDzBrb99yn6tk+LOpyTiYabryZmsoYO2
1AnBoMDZt0yq3nkWtZsZp33PDZL3L1+GssJ74634rhZpsVcgmzcS9y662rhv2ocOdSwJto/tMaUJ
v17Hh1TO5DtDsNNNyPzl81sMzwTsI+7YQki8ExNAABF2B5GC38TMMhNydA4QjoXUXUco1hMU9l8Y
USl+VjQ+klMVqojU4LlusQP1HYNxP7mELUiNg/YEVCnbQcRDo00UslK7KpRvTvag75EuEzigAE0m
HgKHuB7P3VCk6dLWPF3JfaBJwX4+BefSG9lNXzdZn4llvZjERKQbrOhYqN82L5vlghFRumbeIWyp
/CyeB8aktGPQODxNZ2Wrb/VOs8NKpBSBvp4VZYvil298E0WGsJR+Ilso5Ok2FYNZ56Rbmu8ulq7e
oWSBnv1Ed9giCqSFBI9UJAjB2Nga904muYPLUYtUI9atAOeHMdOaMPmdGCtgPmD6nzc7MVxdVQKd
wIsfM1NeWdlS0HbuRsFDXASSrecvu/agalKbuVD2AN5zWO/BeygmKxsGIHegy3q79snVXmL5VjjN
HlcAcGWkR74TYdI21FkQsYln/nb8Lj9bp70T2VO0vbhxCLWyDjhIUMQbmbbM23F0vPHRLWkjLwtY
G8NjS/VJoK1brTYnmaP3GvmkK8l7cMoK8v/O+32xYAiml2leWXauqzmI3RqsmswzAMtq1mv7jBkl
XX+W6zTbAKouVAiRoYWSo1PudHL8hbbq/fNVVnGb7fkfa3WZAqoFs3RslXMIbOs+jIofsyuwdOLg
nX5/uEqXw2J+bZ5DVHXZZVPLrBNoIuPwEtggQvyrINPG3oUFCYVyDOyipp8DR0o1duTLWZJoNwq6
RfpFU4VN7fwFmFE1dD7usIMqh4MzU9s6wRpYh2c+aMeqkQdjDE9hYlG5TeJuaEAYymhgXolHMkW/
Cxm7SC84pJeWJMr3XaWf6zHegyAODuNIaWVppJQyTvBx/YXDhxygwLD3PGMOv2hyGzgE2xUTwXcc
fQ1/jDWy+EGvxqptcZUuAH5R6o5QX7cTtUiXmdzVKuuZz+inJ21APgQtYARbVlEHnoUkmS3ikJFE
DH97OzD5ZnEb72Dj4sy1QFPMm0MOm2huo9CFbDDMFQJyrVbYzk4wrZn/n76d2KEIJREHpgazgvxE
KzfoLlCaH0kRr0kz0j+EFW8bITVxofMFDQCN4PNkZ2/ZRifjufFnbcmViZeB26S/St50mLiyupDC
EvS5ERiB1qsvkMXN8QvJSrLCS64XPKzE7S2Cuga6lk4pYNL21XWb217bQyYTN+Lhz9ESSf5ty4Wc
1fFSENS2ONozfwjM0Oo5Dukj2vgtk73FVPay8ZMlSyglPbO+vtItKqDaXlH2fPgYyz05xYW+uWNb
wVoc4eUFfzoDHhkiR2HFjaorNkjI8Wqwn0IQ5TRp+ZDgTsNKrd1gpQXCtsjAvFxTTyh6GBz/Dm0n
lIiI44e8WKVrw9df8LX1JD/3mrHVD3my6fP811mtpLN8POqpbPxrHeNQ/wyLKhu5sK8f4iFE+We7
y/OnWq9oBUfMGLpKrBRZSsDqAfv1y8w3x/4/9wF8PhN90eQbMYzMw/oZY3dNJzmv0k64dAjNFnkF
//x9r6v0LxaNeAOfDc5NB5WRDMgBJWyMgu8BlT8F5+4gXm3pkG7wt5vCzQPRWej9azXw2egLzGkS
ixf0+4kJHt+WqfQKs2B607HRHdbVGc4FKYRHQ7W7u2Ns99V0rt31mqQJinvHDzOQliueTc6Hl+dC
Eezqy8HVxCpZWOg6OmYmR907EN3BAUcTePSf4WVUomPaeZiAU3ZIqs5x7hCfbvlMbYaLiIiutln3
WBiRc00c8HbyTOmji7BKHdetMABkVZ9brgdBmDtmlEFS3DVLEPOoKa0GOAFNBUdeE/aj2nBlLnWN
wiDFv8KnIQnVc4bBj7tqLt9Y2wUvN2GD6107q0Nnl8xXg/4U6ENGZ1dfm6DUlnwgHBKmT69YrVJ4
5XuigkuDXtESUxxFVj3P8LsispMIeKkflymvc1dFjNpSCEm20UZNyJYWillwsFOmyAHs1TI8uT4W
vUecG2zev3tHMLGbnXYC6n3mpOgJsyQ/Duosy5z1OPLfRQPESsa5GtbuLoGVeutx0QBt6f17oxI9
ak7PHMg5lOtevqzeHcW2uS6Oqsv7H3wUEoUwsPY7VJer6CW++wTol2AuAYf3xZ2pw91zK+58Mu/u
T4ETwd/oJx3maj2WFtJwUf9kJwS/rNdwa/t+Si2ZQXKULtrEXi4p9Obxs7FcDZqe51YEz373oTve
p5RDfK+VAGLTABpGl21C5UgLZaQzHhFckkBSVkPmdf68IHHjALdAlinSwhH0gU/nsHZggZRys+Jp
k4DUOq1GyET4T59nYEE0u9Y2UqYWZ6Ayk/w2SOSYyLz6GHrciCE8zkCupcAlGW9WiogVI72FEHxF
8SuQqLFf9PbSAFzHu6vokTZkK16XEjfNS5kV5zmvDuv2+epeSq1NdSorB3nTVI+2V/YZky94RXz0
5+BdHE12aqbICCk/iWjabFsJ4JiyYMTPqH7OJN2hjEgaexXuN2JYefxsMgtdUS51VMQvk/o2T4aB
ZNgp/3zti/kd2ofZeICJMurMIehArxmyIiIZXpZsv1dbEwimxSGgOImIAEwHLK5Oz7PAVJrsMtGu
S7yz/veZHEsnx/fs3FWv+Budh8ohVEZqV1Dh849y66KUolBR7jZ/LQSpnmYBHO1AdB63NbwKFOko
CPWJWjd15LmamzKDSJnXgu5VlCwiqTU+4UUgEU08bc3ILd3jwpKx5R+YuzUuQijDqK3xRe7qEMlz
ie0x7iLd96LwKqT7DloUe6HDNAJLV5ia2KDH/qNP0vAo2QExjE2ansVPfYRAn53Pns5GouPeCZ4U
ZxR0WWF0f9Td8NNsczFF6rObx6sMn6UqvvI4q9iFsw9fGejjuWMEH+csOzI0EN9KJz4K4AsFJR/q
6IGH26Hoz/sqhjnIT6no7XRqyeIZ6vhI1Pubo+LnFNvupPxzigXmkGndGwhK+asgRz3H++nTKA0C
sZt9BxpalQYWkhKUcf7Kcz4EkUfSAohnF+mIK5ks8kRMks4MSz+VBT49RENe8olbE84rhKPFDA9X
YS6IIS9mkF+G7hIvVaER5MxAvdoFtJXQV9zaX10KZqbKtelMTNo959UvGsFnat3xhbRVz71Ap2D+
3zYDZTBXrpPehKnXk/hsLOkaVBYNKDH3Uc8Cb9ewYzbbnpa1hPFSp5aOxNwgdwJEfrGsb6lTK0JT
045YaOHLvbmorUHd7nvAU7uz2W0O31wnPFnQTWBOMz2U48HgYtERMwwm8AW01DtFXir/ixGzs8kW
TCm3ZF6Z0rDNx2vvIaVZi99osk+dnDHaXZ8ZNclve44628oPuRq9E7AAWBanXzn0YUYmq8OS+FEK
AIzZssFPo6E0M4aKFMfIIlgSU5AwXhVQgA7ycfihfn7B97Xe02L/SXte0E8DFTMlg4MIgRQKanwE
VP7zSTunHPNA9/Katsn15qVukbOQn/CGhWIdmH8lxoazcut4YPQExiUCwDvsrPGmuvPf3qYsUUE5
KFOA3ZEPY0zWvclceSpqTbY5AZ2AIWURpj57MkzqcTEHGBp0f4vOzD9ce52IwJ/OR1YKSFJH/fTC
1io0BkoSKKLBSWyT0ulKdCxbkeclx3it1SLaprBdZEe5triLTWypYuMwLqgDWrCQ7uxQt54JRaIH
a08mTVvCdJpc8mftsklSq35RP5gJa+peultbTuwsjmm/jlGgbJR0rKPQ0eUA0zeno1aHA2ZIBEl0
4LbEpEpjHfl+l3zW1jGUisEDH108s1NBctSV0NY1WMBhGJ4t7HMtpWIy4CalOvOi4MF6fgn5DV/7
TrJsE3ki/2s+124OjerG8hC2yGEqdWPpvH/hiEeDSz6cHMsfIEfgDVWsK33fA02GFqzUC/DhhYpE
23U7ruFh7/Q2czZO0ECnsakMPDhDXYLLUA1rIUiLdGfptxTxxkwQgQxOrDfDXTe9tIJoHJZc2bmQ
HzTy8oK+2HCkG+Dl2j+KK5rb8a6h+1bNA6SnjbXEwEdjKmrmgwYFtRK7uS0pqv8ef+hwJNiP4rcS
nwn1HW2iaKagL/9lQYpVlhzhEfVTBfBioyFaV/FtgBtk7aYJnlpsbe/x/0gW5exJs8Jis9LqjuNu
H2thQKS4drfgTgq06Ymdt7in42Dtrm9c39DNGlkq9jxuSir2mTVn75KKEXtaKV5PYeMndQgDrcCu
wXDvAvLJnuZcwkw3oxV16TWaYlYB9frnG3Mfb5QOQw6jiBkzioNpIixvE9pVo4fRtZnAGF6XH9om
vS4X76HMbwoOzV7XbA6l0vSBLD5qm5S3yRUoCG602zSkkRdfEQT/0oKyTMtFEUL6XOkhW7E8UzAR
I3fEAVEPUCKsnrj8ktF6MhUtLaKdxWub5+aeGS91kfdD4u6Hh1FLaS8E7SOmYGJHxgvtdqAwzZyJ
LXe7MpcQTKXw0Oe7oO0Bgx3FgRLd3AY/bgsp7xNHB85XFoS5bo4Zn9FDwYF1onGbP0JAoTjsyfUe
JUyIJsnR3pc2UmdtSIepT3cqSyyRZ0LpdKaP+T/l3ngWo2XhhdPSVirPFn+i6/PdzE8O7LgpvxA5
LU16P0NOv+/xagNleMc0qtXrzWMPOr5Em7+xufkfQP5LYAj80gSF3MotBoX6J/vswCuBkEe06vvD
V9+4DKXJEf/51qT2hj/xJmx1B6FhWe5yJGoE4Q+M2sBk/etteAyp92L7C0MWmlpPPlL4HbIGJ09C
kdMnNiTtK9EzYA3oIRJz60ESQZcERvephh84IkEJx8Wmsq9tpDKm0D6HbLYWU6lMqg8pgH22FSJC
nG+++iUhPW2Ys86BAZWnZjvZai4+vlB15cLfKTV2ZDJjf2NcXZ1S85CXGjWb9sAZtKEXrKnRqz+Y
T3Vc1kGcERIn1sljlKIuWOGHxLuoDiA1PV1DPHX8P+/ddS7tfyyK1rmPP5TbsTmLqjf4kw8aOPgu
vU7d4GVmREave6zV6T4ExrhQRPrWB8ikXTzr/0Vvuyzp6sqP8tvOswiEPC9gSlHc3YjppaJQ+Art
9/qgPW1MM3iD87oCOB1NBd7YoktS5tlSQBgUIiqzHOD4QIt+fobAaxcQDTOdcBbjWK3Ip55ouGZp
wobFP7jJ0CUOL/WRDunR5I7BMvmqFaVH2ZMNdvOibwuLI/08O74ugrig20D1ACErMobT9O4riGqw
jDPDl262p5OxcUQV2bJ3hjhuuX/V9IdWCotbhhIdNJ+yripJCzwvW/O8ENxPtlqUQKDUUrsQ99tC
RvRoRAHYNiqFW1KcDA6JKk2IpV+58aHc/3RPC2kDH/WKUm0xEOS1GRN+G6Qd6PeCSPwi7v+fN/WT
pHtcMPGUQxQ21zLMM+VqHGXmQo4cY7N/V/NgwpclDGH1moQSK4WjnjmxTX+PuufXwXx21H9DJzr8
01PBUPYUfUS6ODLj2cmgIrxtZX2ouyLYxim9XD4AFC9iFmqrtBpJPLMf/HXdBDcswjnmdDjdq5xk
qQ1Izli+cQp/RHjxL6v5oxCnR1JuiPkG+fFBNyrDTpbPl4QcbGXNgaxFFhERJYv6gxMbSHmRoYqI
7LNm949YD+Y0fLR7s5PQIVd+VL4o8gXszZyCze63UyrFy6UicDYINOcuQ5j0gdVoYqk9l2CkySJj
z6JSCLw5MNfTK3e7LslLiKZUu7tO8i53CS3+XaKJAIv2p8FSICLY1v4iN0CtIagLAhFvba/X07LV
dD8SsgIEh/HDsJcrFHpvF7d6AVoyr1vA4oaxccBk50ePqnMctPviVHhyyuIi4lQyudV3287CXw3v
sfDuoNCjo+HUybJzoU/d28Ezbg/7UGii81tAF+Lm9Lr0ChNRy9dvtV22TgGa1SGhLSxsZerhH1Uk
CRpWIOYr0MGFxwB8WlqsDNIQXWuQyimR8Ov+OZo3WjAq9kOjEaQr0MWvvU68OazHUJgy9Oz3jZ+f
wp4fXaAzTrmmWb4j+oAMhCVdbcZ+saEfED1pug3kaOVi+RV9lHwN8I/f7Zab7X385TDtU2kPtDA7
ZKJoCvwy0Zv6au0gMGXgBZnzFRkkrbSeh+nc3XDkLnfhQYTdLY9QW7IJQXqRjHTdLmVE9NfHioFT
t6JsWrWb3XMDmXfzVkrQZEgH8dWyPbREn9T0mjn9Ambd6LxuHkTzA4NC8ea+cs7foMvOU34+bDVT
eYoM2m/M4aW5AFxiL7+tUts9B3J6GQGAtY5AT6SChqLJBPCaUpe1D6jHEHy6In39iOhE01ap5ngF
v5mmxy5fcqkGzCD8xwY3+7v03a7RkHwgF3SH2vLdqCBopHYWHgU2QXVukfW+gRZ++eiwI1KfWyRg
aFwyUO8Qjgr8t7kg99Do5BCCgC/FCgQ2lLGcguogHUTNeAiOaKopNR6UgsTc/7pjjnZAZ7bX3Cuh
3Q2hzrAHDpnpQCmd93l58qY6IgEVzqhRmtU5SFM2CXiQvLUhP83Q+4pxtenWf7qHU2fvvIB6P1Wn
fS90i8ajKHO2LU+G2FtsfBDxCb99RNkHr7dF2Wm3gH4Wr4SDJkExnkEo9zaa1to7mRQ3t95g36vj
GxUr3FNW7/6G1606dnbwbAD+gmHspyqmjPKW1YGsIk0KW7Ps+rkuwzlbZ+emcklOwo9gK7+iVUqF
BkgjJ0MvX2fx4z/lbeP6lYzpWWVAuiUIQlCeATx1jYjPJKqezW9IEr2IQcPHcO5sAxI2T8A9BMRH
2mvpr0pt620Ux3LxEUW1qkR9wJVlMfAvJZmazxmhF8XShSfvgucmqOiBgsJF9cWkfrglw5OSkPKo
KlzmGYaSxfG19ZmhljPPCezP08JtY8LdFrRXdxBJyHJIKFimGEF8RZsJkvkfZR7vdE9qWszJvJya
hOjX6LcemA8UVF7Oe5Kf7P4/eJ1iGMCzYji8x3cdQ1J47I/TGrFFGO4hua4moTk7rl031DsS6b7m
LLQjy7W70/RgGSJFivArLTQrJ/m7saJdT5zpKnZdkSLFSB+e2s5DizRpor82meivXpRWqtp634im
kW2lQw2mbPOgpsEuk9yJwmHpCeh6DCZKIGndANf9n3807lzfO4UQBFiytxSTG1ofbeMfUlq/wkhX
i0NhK03AVPoWIpTFBpwDHsWgTGOBEbvbLEwQzI6rx9n9TyYn3F1yzr5ueC4FhHij4nOuPG+DSZP0
q6rmWrdjC7dgdL+Atur1OaPGjZ4n9rOEO0QzUiMF/wUikafJ9RKYoSwgodbbri6L2llxn8ve+G+u
gIEfDa1TzLuydB01JLSMn4pCz8SX7Tc/3HHBcdbj2MoiLypzok8aISnCwUmb13kvulg1B4tfLiy3
FllQvY8Li/mfUKg8S0JRdFGbxLIKBEck09oQ/d82L3KKJ+wtgzux5Nj4W3tN+ClGs6a0BB26f6Jz
M9sxxKbEZhPoO8wJZ/E+IoQnlhdoJ+8j58LieW5EupjeLtli13MCXbYOlmbWxHeXN4mHbNkFfsJq
k30O0pENE86qGo7YHgKLgN9+/THtgS5seroFAhKaxht1JBF2mGpaZOMMou8K8En9mc2P5mAReqek
umx/VmQ8/RQ3zR/fUXdpe4PRbl2uZVKQNtLEXDEWrcgf7S9ZkXJdZPid4F3/dmMmXnUVzRK1kg2Z
BlPgeTj5S3qyd5q3H3Lbb+0rizZioSiJOyDNHEGQsyBS5Fk1CHZnNll9AsrXCmL0+eu+bksFQ18D
HCsxEp46bGvLhSQIJ0gQEFqo7u3F9gQBcf16wyM6C+TAV2b+kUke4OA7a0m6cdsenzlDlbhYsshp
fyONCrLaRzoX4r+d2dj836AvZAuVJWFHuEdoY4QSRNe/CE7BDyECJ9cf5+0sbLP4Dz5T9zBfei/n
zauJ//dUhHxfy38Kz4dmcz4WvZCu52I/liPlr0HzKeheGf1mvPntrVV6ziAZK7GjQZIsDOhOC0bG
ru6QG9efDk9PA1va6HdGxMnGE3YVwX1X4VIVrfh00P/M8jNX+GR0oZ3OBx2BpKQylwkQzSrw33nu
ESBPHZfphh1bA1CImsxDo8luPAaLuXcGa2q/iZJEL7zyv3rRk96ufCRvssgizMDw1hCHs7sM+tbV
BPmCtwypu+EOtzjocfoF6cXPyB8BDae3+0fQMzQ5yHtemWzSz2xvYgsv4P+voOiFftaB5zdkh5b+
SRkB90jnA8DYqu78TSnxqWJlNZCWpqGsHP3r2dwwbA2GURiAWQokX7WzV6m4FpZTYB400XOmVVTb
PZgyQsulYPpwyrovBfOTmwS5wTyVfQi1kKt2cOi+WC6LXyVaCvOULlzXCH3fTo53svH5zIQxqnqV
yXRdrEHgCB/yarmMubYguiI+J9425LTsvrdVAsDJFrxD9k4Ky7I54h1zGjcTp19xtszJ5pzToQqt
iuzxPIPIKfblPLl60mNdEqnLU9b5vZLX+1vHpxEtaAEIiEp89ccOXU3kk9XiLomeuaAsnOb/qhEh
xZt9/pt/qHqAWza58/0ocNUdnTlSUA+p/n3QWYsl8iWL1i6bWvVm4QVRElymLa3MUb7Rht9+KT5j
bkwCpRixXcTcdf1XeDLPSSeYR2DKPpKG6C7a4puo5A9diq+nI7f6Rm01o6ITisOY/H64cjnxRBFI
8VAMnz6ZzkRYHTxR579r6Vj9ZghgF8iPi9zkrhsGZAso8/Y0jPUfA1NHLgOz7r0SjsEkic2K+PkQ
I4xgDcSGKA68bmIUCqeTE+taKb2xpGno55sRHOnkdYd4ecNU85JVwgQTd9233PK/NgFPPlhZD5sM
0eot61MaxDFlGh2ChfzatWJRcx5QgUrJ69shSOGgAkX6yqwhBp0fqGfwzF21TwzYJ8iWUXOGM8We
WFqOUw2Je+zXxAW9RJ37ixtHuaRc1GNcKUCFUxRLcaHiFNmjKVko4KlEWUIcTM6xMMTJlKv6kiNq
Rvl32VAIs9yEuIbnIdFgSiymElInIbYa/y+AlK+k28G7s0zNnMoyjNr4nkksHnn7xXW/r0lF/oD8
FjeZZQDkxgquJA8sO4kmUaItV85gm4stYDfBIwiYX8+lMdfuL4kg5pBr61ECmG8Bd0EiYYW860Hx
KThG9f2VpbmaTngjfs4hDGQTHUINfkicAE5pKqcSicNuA/bmU9NTNT5dfMVnobk9/zh6C/0syFWQ
196ihFUEjKtkmyMh/q17PLAuCZ8CYtpibCAIYI8d+FAj6+DnxXP5v0gLuXPBa2c5ifiGg85hhQLa
ainLR117MskvzX6rb1pm9q5B33JbC1jeO3Gq3WDa5HpQWEgmbVc3KBYJ1xg7UXVB4baDOL2GTnmq
FGZ5Rla8GzMZuADh+hHsmqQf2QDdkXpTkXyHMyWpI3CGbrSAEnhH1mYygfL761jLDz4Zqu8+uOK9
NVCzVoYYLe86HUr+PfECDn+L92IBKcqx7mO7HJjWjgwO9rq+OaQjYyEY6iOjolHcC67gGCp3ybwY
GKOKMysnOJ954vqZ3BowD/sJyxuhPEPxU9B+6b9eaWeELQo0upGHhf5Do8ETej4eABp/TPISYXy3
ZbHc9sO3Oo+DmaZk+JVhBqeJbMsXrFh4GRKFwM8NSkQSIiE/TmTIHhoW6+HRi5mHeATyaT7cbjXU
Xztr2UunicAhHWXx6wtiMXqLh20jKWEW4B8TZ8rEFVePZukyL44abQ/CFOMcAPjoZNbX3vEKgymL
sPeNasFr1f9xMT/8CyX4XxZ8PIoEH77pO9PvRVJRRqeQTxNZ2zhE+/Axfq3oqomohxxypnrdhXuU
xtYUcvLp0t3QcU0JRp1u5G28BgFfJ3Tf5y9CoFMfn4Gkpr2RGQUh5DPSDNYXBlC8WAc7WnYxFzh8
o2jYyDir5q39C24tYj1g8xWcC8/hWSrlmA91cTg1FekjUJdpB3yzeCpro4v4In17eT7zjSUobn3O
iFb8nn6akfBtCVU2UNSGa6ONDXg++ucgc6PDLvMML6892pYeOnzKuj5gLguoMCQdifTMQZiXySUR
y1DgwxraYPhI0ubek4Ru9waHXBh6lhbGiL6dwTUtG85glJVFIbw3bdxxQoa80DbDUzWly6peqD+y
FD/99O07+D8JLCCKw10Z7EHR2NmONVnhtpUOgh02Inv0ppN2/Cd5rc07tTs567X9HoI7w/Rsj6RY
bQFMeFmqbhsqdn1/j21MQ8XcC3q0ToadGU8EKwKwUY3PTbCy9B24ims+iQweVpZUznSfstagGOYF
QtS81wWnIM+BLXUCa0VzV3rlwtPXVkvZpVgcXyOedkDwORVVm0OPlCiEMKv5y44LoAPspdFzgp+J
ai9HN0Zln40WEvtb9lM119iSIrAjpTVHYYUVvQ54AwsAXbZUyY5nwDboMm7upZZjdJcQAR6uK+0i
nAmxjubz+GgHkTenDtilmRjBxmUxidXrq0m/gDGeqZcWhcWu+Sq/wjp3Y/+6sdq2Dvviu3q3zVow
3F76pE6ujTgg1ZPcNIcXCVQMsPVN6Bnaa2RbJ+flhvOZhisVaY5yWWoHZr27RAS3UiCAPlmAPGYv
58v2MXyRMNnA9Sbbl89twFWX/lgg9ud5TcaRq+KMD5Abkq7B51NUYMn+ZHx8g7B/LlRXPhfup/fl
1wG3PGMzZYmkALGVQuNHqyx+Oo2akSFX6PoDhx5SzncHNvTMySPAjnkxMxgXuDX/z7OV4PEcZ82p
Z8g+/zQagRo2pWPqaKqdnYLH5ZxeGALM1yIkG2M7eU+pKXdRzdfuHQJng4D4ORf2oBjuKVbdc9+L
TKC8ZSvI6eXFSyyaQLhCF5zVMpdDMYYcjW5n4s5ZOkWv/4fXZV7xVjqTcTc2TIuvIUEsJCaxjV1L
V3E6xiLlznktRufbcZtfaqG3xt68S7+icli9yfJb6ZRaolyReyeWjC/dLFKWTwMinmhMXFWJlHTC
peiGiNZQllQtL4rewhYiODA6xZJLSdqt9OJTMfE/RQfPk9RDtAM8/J9EX2CbIBwHYe/yac7/vKrC
AVc7Kynft1ZxqbLsJzwpJ26bX1RASu28LDUB5fCTGsHnbXKGFCH5miounS49QoN9ljJvgvVR5laG
Uh9WUKsJoj9VP7gZQkMi2V10eWrJx3d7Q7Ft+20aVKemioXnsFPAYdTuaOt+CBG3QZGtj/WztbRC
cHuGe9CGP7439RFF3kHAcgYVA19vOMdKBtuKZfrLyT4sM3hpoZsQsofjjGGsf9bNWZ0GUNxBMpbl
gftfbiQ4v18n4ACJ3vSxMv9tYLQodZv4Wcej6x9yWV0xwwRD+QadpeqyflGbSYhvpi+r+9ewvl2A
VZoqY3bg6SmAHBZhThN83d4MT4s0fKsvdY9RJ0F1oVYVV2dAKV1Rd5p/o11JHqy7MyN2yq5tNuY1
RDrXDBsoIQO5ak+tDQDWqEeMCLjsK6GpF6aV5g04ny9oi17mDzh3SK1PGG93BLTPJYzpJfbCao4x
Xz2WxDl1V04/p7juB5Nppvv03tXIhI+3IClnGvjbBEXeVk+4pLsNHUG41TXwQtswYZz6S1uJobsk
AwbnN+p9biHEn9mZyJ7BHox/IgzCNkXGPCWIGRkLPEdbVC6EjEMOMc42t5cn1jbBaCTwQ8IVKsHC
NuEIbc0P9UobNNdup0zf5MWNqCoPlnRS3q4awGjDC5sTtGmmfI+mshCReNRWiy5P9qMWbZV6Rfuq
XSYXEyjSUL4n1CPX94vT3fRcnSJZX2u5akuK9nwSrLqsKfJ+PiDeVaFZ0rMCy7d/i/668Wu4z/g+
3z6FKU8dQcyeru9j/iZqRmxzJGVqzNMYmx2OYzgSMX0G0Y8K9tVQhIhv5yRTI1FmqQg8fMDk0CWV
pvLhEOUtIRvQWE04fOYyjZx9Nm9XmVmPkCvFLAyfpnkXBLsrTeyi+zTCPjd+luZcEmryTPbCPbGw
+oaBF4fdBiaI9SDFmeU8NnIUzsVZOPyeC7HQgz66K5gnP9osv8kuqz4Q3FGBXjryHHIZcTGfszwN
rBxAcNnjCtGvNI3XTlJZ08ybZlid1v+vQ7sgSG7fzb4zRTUyl4VHYMubQIAoEqoMcsHcB2Ve0cqI
FRCwKd54A1imURpA48u87i6z/PYWATjYIyyVxQRpyPY2H6xVTkfzXbj9cVjk7iPmiKfOY+oMQHf8
M3n2NXaMc/hOkRmrn4++V1Oswu2aZ6cT7S6dhc+3kY042rE23zrpplbmdJgA13VZTm96KqKF6Aaf
5/M1Odd5aYPszyt+cEGRJfJ+N+h4k87XOL6IHKsvzmOAgMHCOhyAIdVProgG5qXCaorxkVqr1vow
uzKOeqwb7rbbwswkyYHgWFk/9sCAGmu5bNyb3Hp+ME5S+/ntgOT1u9GqyCIGM/INU3cmXIdyRh8p
H+0cpi1MLkAw0Qzf3ODfF1Bz5fbD1SUbXFeiPBErYXswesAMnJKsFdUUENqUZXrl1ilwUhPyVi6u
H3UogoyKjJ3bMFIwWsvc6qXjybXXd2tggvvWcXLXlWi/pa/gvtR+3VVnrbBq5kd6Ea6zOJR/4Zfu
AmYMRaNp2FeucosZQP/QQimEF3H3pkGfWkSClPg4AvxmvNq8uwNlmNPWXqXG8FobSBPi8WfUiCBj
Y0jTWEhFAMrlMl+WKOx6fQYSQGgCmbKvNk887GdbZFy0D/caiT+k4fc8rxhKH8O3rubMrIQiRzJ7
qKtLJ48O35HhjAE52t+d8q4G+/V1ftgjFQfP2U4nnMn/Ip4YePPPmAu9oTsq2qcOueb/ARDmjNrd
U1mhM/Ejda6J6khUAan33gZDh+XxCHolZM7+7QqeIVZz4i59p2HHzTzXddG/0jnJuHmjf9q6MlW1
ubSy8u6g1G61XRXeBgO/TAT+CmP2Q0xM7wBlffDfNnaijVNeeL8FNaO6l5GXEEZY/2cB/ncV/HOc
Ko69n48pEfuxY1HcpkDGdsyIaJVkRVoLa/HhXuquVnUA+6emHGkJlGRS1iXLuQkpxO4KA2tvV418
7lAbgVnIszSg9j9hbTAFIo9ptrxZsRhNPnOFzshmFYRoWeTtmoST8hP/c+R8pMoNQ7BzjY4qxgWl
MYziXX0JH8tbIvPcTFEUxHjvcF27YVgr4wpuLT+gibMcU13HfGodL7m0SoTOKnrWXvCvbAnlxNKk
OQTXWkvHQBWcaLeOfux84RcG0YB2OGP7zSj3lqAX/oJB1lfnTKeL1re44OwxhNp8+6NxAxtK6A5C
/Gv7lRv1/ZMXtXTZvxGzA8aqs0VwTlM07+gDrT5e5ATm9m+V12uVfTgAM5zHanZxOE7TpYfIfHOA
fJxyxpcNeIJHBgopP8DVUb5LeJ7Tw/6rPs+CesulXXxivV1hvxL7Jv7loLdcfPugdd3GOypUuayi
xiA/MsUCbs//wgHbboJ1FtkC9TkYbWBJN0UxfbYlQbVCmP509jE1wgFa6wtwyMRKEzypL7F5hwmO
OmG5POOX5ttEaRF7Zn9wlV7U5gFCLSfhU+eVzg08ZXLrMTZJxyy4TT99l7+zF8h2Cn7DvVfRzRDe
pHgaexNzU8PP950kMlsrq0Etv77zmNjSM5dIbJgAf9cQS2ifgcjVW/5G3+Zblq/eYKYC34bdlm4v
CIYeICBq9tNJz8LO40JmQFJBzczIgi+o4Hal0HUpWKEMrAFeBr2v6Uwwco3+/TwHlV7AIfQecT1+
UlGGxINaF3PyAVPxJN/gQhlwf3xiqdqjpyTA6ey/JcSFhobYc3wKaYNMlVfgEJ458YGZNUzc4089
hXhLGCPiP9bxGNjIoT9HDh8UxFfWn6Z5xuKqEbBW0ie7voHcy2Hby7JJHWS0CWDE4QqlUn8dd4Ir
k1OQlGJhB8AypNj9XQj+KMoiiB5k3s/qA6vI2lA6HNpPLRAb1wuOr/vYkwotkksylsUg/KsCAyFC
/o/Vnri4avkCih80CZpU7Hp1mtqGyufuu0IrxUROLXkiegEUPerBnYZEgnc3bfc6FkhqwheY7o1Y
oPqgqMwIpydeC37+KGipH1cmRl9YBQLZuY8ZDGoRRSfBPDWiT4N2CaXxF+joaiSUNeSzWtg9N3FW
9gWSf8JRdYV9lO0zhCfJQJl3oFVwzWLKiGJ6wafDHjf8w9Dqy24PHQe+Nil90h5ccc5i+dBtStYO
Wn9lI72ac3a6IbpKQHMKZ2DtG5+8P27w18EKs9zk2H1dxyTWsF9AoTh4JyT3tyN+vnYMM2g7aWoN
HQVljZFInCx5y/oh4n5LD49CLbRwZ/8sWtMESGi4FJnN0hgFE+c3fLbfhxKP60U7sZK36/eihw0k
XKJZp15c1gvbJBk89kpsM25dc3enQyhJ4ysXTYh2HEfxW6bqsrYVdosvIOxaSUXCfz0fLXDYZC+9
A4esQfqB5F/JylnSDAG0/XB4g4X8H8khchdytm5193IcwrZfx03wMsYPTPBKKeNPEoP8p1vR58Eg
pMiJgPkweqst+z8MB+4ESwi1ildsOFt737vRshgM2u+PK4EN/+bmvMkVwV5z+d+DbEFDmsHPoiE5
BPETyjAIa1idM3tSXD8Q01HWLKnEUZ4209JXrNfxIZVkiHjbPjHRYxtIYplgRe8xpjWMPy0ODMU9
d0ZGw8MkjiaAFnHz9oSmpcNKoYx2q4JnUfly5cOcgzcCD5Nn+4RBcHWYQ8Pf7WjqxUgzuoHRATb6
T4clSRD+Q3LD8B2+iqGTOxg38NoELdG/4/k4nGjA5i0qN4X9SAdjF/fb6AH6fqs1ooVjqP0QMs05
eyv7Zp6Oq6UdID6rL85npHvuIKc+KFTBw57H76dV1LU6BGgcMxjW33ipLxt3CBIZoBUR/Y0kC1+r
+UbuRyfP0ykvh//+N0IoYeqIpIw3yqtJWYRGtGBcOLYr+X/yPVLvBlxFxi4kbdBNtFJG6NcV4+F0
gDAYhUATuMwqOU6wvoFdP7yEpHzDtEzGBxnf2zCzNdcfIEEjaBbjbBqPIduLUzQIq2G6AVGg726i
phbm7yJ2FdfCBVbsXpBag+b46znRX3k+jHH69paXQ+i0V3MySMedi89vlT4xOV0GeCx+mHxxhVfM
U4cRNXlbSNoYcV3m5bemwdWy8WQ4Yv/jhdpvobMgiNBAjnoalqEmclrOwOn7O8M7aG6WjNpqlC1D
rKjNTODwNGdDwlMB4h742P5QGV+XzO42Xjh6BiNiAQ8IuNefCy2kQlaxaJVy5jW5L1ynVHPCv/0S
aUyZ85eNOFf0Khp+L8ChEc4wpB+4Xh7Dq34VA28h2O046KWG8hZNJZFYQtmVYUOZXeQkOCDJqiMv
QSP/hkO4AQaROz6FiTs/gReODufmhN6H8bz81vQuqD2qXaaNiJzkmzkJaHGDtKopkHp1JUYxgNYu
FbYK93ES9sCv5YA5YDfv80ta6fpbOyUtLLv+v0E1GH34ufUS2SCE13o7QxsEZ1C7k3JdxSFEiE3N
DtacZh9fNsx2kdUqo3b6AWWqK+wAD6CIi4+EfNPE4PEHc7GjblvWH0TfloxnxgB7P6q42SpkCwDy
0eAfHsXElezzSQDhetLs9MkzxGpZgWisM7oP1JnBDd/lihl9u8a7qS+mYvwhrpksK1xDRH9bv864
IvOiyFRdRjVo5OShUZmRXqeu6cCftGsFaT6mqJ/8fh4vzBOcsrdUkkv55Jr60r57vK7+9uDczkuA
RZbI/ptNgwjRrDraXYFDaQQ4KnMuE2AAh3spwXEW6SB51lDyQcfRZ1oG1jrPVqJRH/wANy1qh9mi
f3zhb46dmdjlSL0Bf0TnWJhHdCc+Hb+inysJLnoeKEgAZaYgfIRNLkVvCewGdwOHzDj9vS5UzNzg
VpF1gGuYE//8IdJRGcFuGzcJDnVrUf2LsFtgAf94VFOKj/s3DEenue8rDsb9Gdx2KbQUnoOq5KVX
Quys4axEwCpqKI8Yap759/FW8BQ1R6IJs7DOOfEITlBHizJM+I8QWQRUEeen1DYaVA/xGDXL/6LL
xxUp9vWRt/21eTJpoTju6uc/e9zq9dgVZuxQObX24lW0rWcnbohwm9Xn2LDGko5K/di16dbu3oX7
riJD8bvzNkOcAhQFkNFQB6KD5ddbegHoncsB4zLK+KTiZ79X8QkV1A0ILPOP2shi7WX9yP+4MHgA
JEUGHqjjiEcGvPva8pBknNsp2JWAiFMiXP3Y4nfnprgtejHPbAKNsG4ttjYCPAXYgC3Fw/3Au50m
3mPT/gyR/N2wkkj2cIxajjN7Rvy3z5757I5A7QBCvWm+J6yLjB5th6N/EtZ1AhDPRb3hIfPM9BOh
0auwOAe1x0x/BD7avQS9n5adSPFDjXjGUS2HMqzeE9Q8LX1r3W/eGSElak2qbxIvh7UmF+suPm0Q
uUklcjRYkNm4O+QD6kDB22Li7zgpgcBjn0ajKViO8U4x34l4sMttBmFAIH3K+H0kD6Nwf4ZHb8az
MQ2jd7PD4X7+g6MoKSb5RpP9czWNjYatzjeRXMISwmtKuA494Wqfhxfz8ZjXsWl+WipjpvhNIvIR
QfyDahhnbm1Ong/mc4iHOjZooZiop+VtAryrD6NELIn9foxXQW9TBF7McBbVR/1Za4EXQg4259bi
1U0V9gmet9KN1xrKaL6r3/cJclULqC9rPVjxO8l0DAvtGqX4wp0OAtLUJvKzaSUG79kPTX9H6eTf
udFP3GZxms4xEh2+6EqkDq0juBPtvAD7F2IFHpACIj6hFf+4ar7IVLdlPzpMug/Tpo7UulHFAG7s
neW12b8jPhVXFeoJhcxzHH+PFB/P2C6O4mDNikAAPdFRwYXYfuC/jxD3vecTA3fvcq5Op/sOh/og
JRe/4qGXS/WU8CSrIeGo2g9nQbXjiuDMYmknarENvqCtjSgxOiZx8ymuB6LOAgYOzss7rvHwk4Y5
lObkL6lrY0PeDVgfIkTshqOYdCGZV2sBR5JOVCJUyb1PCcpeePnDzc8ujpfHd5VEdQ2k/ALlAIjQ
SqU7UapsviFr+q/zvK+dn2FqbtcHKTyuJuzZVmsfJntByaWXh973wsf8GJmzGuWdtreegxWYKY2w
dWvS/LTVHJGskO2zaUdeuZlw1FjYGvKWearGrOwF0nkUAjqXlRlW3fqkfjkPyUtSqYE3QMr1755/
tQW99juTa+oQ0s2RSRs72fnk2OvdjUw5djIRfjpZuQ6qmy1d2s3dFNXvvqMBiJSO6iT4QuX2ONJd
4tPjlOvb3MI7Fb+Jnt/mtQ/jJnuKboIy+xKr1GErJyl1zD3d/e8IiAYACxYDBGysf6m06iMEETqK
U5nz/u1PXaKxFV/9qTSju+WXAzOs5O+G/fDN3e/rZbKiiD5aH9j8ZR/YdiTm8AGCZ89uSt32AkEU
VptiWtr4cR/hh3JUsNvsSO+xdfPetvyQYYXfQ+0OuCKwuyDZpeg3yorSICqQQXdOsZYWlsPIsqlR
ncpyB69h7GuNlRM4zlC3WPt4SQOoU8fb+ko36ZACFtEchIiNGlJLIQKp6BZBQX7emWZqtRGYxdSz
oYftN3UOpDtluYiuqWXQp72rV8SttnrZDoKRhsjKC2uM9XDjPWrlNNjUbc5Ja5G9I4rwJB/bKYAa
rNsxFtaSJ/3YvXRkEWhuM7eUCxS8Y2C/W73Qc7IDd+CbUR3kvu4DbjvtTuxDd8Oasb0jNQOPCxBm
bKTB/5mzEt7q7w3TRfk5fp/6DI9vd/UcdyNCcSCq8IAWe6LhjLZZFJ1r+xlhHIPop7G130RflCXQ
eQr1wq2KCY335trCLmulrfAzvURSL6AGSyND5H166k4IU+raKn44gzgrCF3geA4c6grNj1vGkpXw
9S8JJgq1kOuRoyIc++RHmskUSeP/Ousa3+ngJJ/4ANk48X8YymYX8L4KRFYyMRe8WNP+WK1BSuBK
oJJAIlT8p0esx7gfrGFPhdFC6iquwArZCRGFipsPs5ida23rWXnIcmSw26a9afhRDGnNV9+GSMMo
EwJa6dwC18N9h7Zq6gpl4lXQxXgg+zvS5mr86BYf4e47RVcBXMqQKmqLsaxm9634+2CxbELbEfao
QYba3sLdQkJvfsPkUhIKaDUgfsVNBCaCyjD0dC/5sG5/ZoFmudpdr/96eOXWFo5rowjRBiDaVk/7
daVTp0PMK+3DDrOCQq3qvlG6uq8rBPrn1KSbPRI5M5WsmiQ3Z2X1zBGrgKGs9f+AFyJrXF6nVFmq
9evAOovaOjAHSzxjQ1o8zC+qBA4zp0GpO+/JTGUFBDSSsPTArJQEVSsvXl5BA4muQ33ICD0O1ZMC
bNvm0nIBhlS5reFrAEESSWfcLc6XD2JPMIDr5OwZ+gk5Lu7MGpsRZwckAXv8RKAigz4OV0Iq6e7K
QAyo2RG3205nFi96KZCIbri5tJM24TNKYqm/jysMoPdAHFBfe03nsXtBY/AJxJc1yemDTrlLUdik
wqyuelscNbdzqVmK8nHVSaZrLN7JkRXASr0rTus6KxXoRFPirp9O1k71L80DxhngRts/Fzf4rpgg
8TdFoo4rKrgHXoexgdxFq7RyhWrStf/1KizJg3AOxHkgu4u2XWWCgIQOOmSf078XudIgJsW1t0sf
1ZIw0h3QuRTj/H68mM5OLUeCrdn+qLekic/y6JEJwz7weOnf6lh7Uj6K1WC1FL0kUkJtiatFESOM
+Lp/LKv9bFKztdaK97S0jzYeVu6nKPB581lnVFsZMQ9kwROzLjh9hNjkMuY6vCVK78I4QL3WtKfU
2AP49yUA8VxpU+JPsk3c3qt4UPdzG8ue2I2cGEnqVjpo6M8BbWx49aJJeVQXKysyFL26luwE3sI9
ZtONlYZbrVcNScT1Iq/3B+Ml8yk3wOY3Mk0Y7RSn4pmJClaBxXLm8qPh3dhy96qca+XVYlhXQpg9
5MLkpYHO7hV5lRprvqdnvTaXe3Hvg7rXhJmCkPiBsgiuO63MWjqIS4E/svWa3C4sLi659zzA8Kds
2qzVRBS2dNQd5qJ4ssF5NtuuR9RsV+2XK+v1ZAktq1+zaq0OSiNEc2JYvTrLZ8NESZdS/v8fqH9J
9Nh2oCsDlsWe5ZTVb5g1IuaIMRSzztL+euhOJJyIItTxP3aojch1jqYyuHopKTnocDtuis8aKiBD
uzZYlbbKuYbCvhdwG8cjCT8BS0Nalr9ATB986xhxexsWcmb9P8YcwBlB968QrlTNmKiMF2iUVOMo
A+x0Q5obGxetoy80uLn3FzpyI+xbb9uYkLhny++/swVK1h+Jn3SqBWXTA6Ufq7RiURdT4dQi7eJB
/YVkYA5Hiav1yf0zeW43QmhkcpHaBc25jA56geNqsfftwSxdZSGbBk5SoTeQkqsT+RfTg9UpV9Ys
4eEdR92JYbA3WLntobh6sUr6gRkNhqvIPgsT9klaAmhXHIYnTdGH7Q3Ha+86YmRfQwBaCkMWnmdU
VCdcXeJZXO25yRXRrZHxcTm/8ckWYc/LH41gAkQ7qa8Uhv4J7CBGCnO6sBwWlpzz1bJXb8z3DdKi
YUTgCZ/mXkQSd4HawTUtCOqwf7IP02NQn9sPBgahjyGzza43mftG/WY47Y6KcP29feAX6Mau2dzM
EfbELKzxBGm+mwiMRai65mKDgkADSgpfQFjOc6yBvfoAYEKHG51HipJ3Cw4ahW9xdL5JTFDRFvpp
6a4kH4WhsQwxdGn6+qVdtxe1MPwsjVWxAiPzfP2aprRBo81VpWJnnljBDltFzAES6RGtttB4PGWk
+xiHlv0pMsgxzng5jgfgl3vLaZ+72gf4GIZU1nOWB2JpUSW++aJjFtoiEWf0GJlExAd1UZZ914e7
Vhy7k4VJADhrQo9AxJwVaFLI8DBKUWWGhoOJt3/NUDMQy0NURP9RdaS9HUeUUvwTlTR/35fWEZS2
Sc9JFSKqg2OZoXiZ+koozO8xf2kJiyFAEt9aNJsOvNJzlOfA/XLKL+FeGL5TP3AKANazVDnC0Mcn
qqjbGErMBFO7OfMJDsCOP2LFNdTJE+J1MTgI41b9UjscrPQRxQ1ktOgiyXpA0/CGe3aIpJtwe1Q3
w6wZl+6Tx9tFCBBB+ytby1cqPYN1An/JPfJs6nGQ+Xgcj2zgEChXLkorZKB2UUo8huxXs2hXZJVZ
UZJnoezqUSVKkzkqbwKhaYA9raiVWBmB+DzhorgxewJ1FjAu8GmPWknI0onkYa3OxomPxA5UQGVH
d/C35RtzO7Dgk6ObQdfqqyxlxNM0Cwmz2YQqjv/VaehpUg/lBFzS0q/T/i4gBO7sNEHbpqSwdLON
Ii7+Xf5Z1129MCkGj1PvjTUsPh4UIAvNZrrQrA//G+hrJf6EuyPaCDUlf9CNx8Ow90e146YDQbXO
FZO/BluEFCXKu89JNAwNWQZJVOQ+eAwrFyOVmuOm8a9mjDnwE4sl/u6JxAP/tT/8qfPnxI9eNpmp
qIQgyUPNXnN7zhu3625oO4ZtqpY/lqKWpjkNb//ZOYq2cxZhvVSunfSZfRM5EmmjO3n4YziNAxIK
PYXUhEYOsggNYtjW1XYRMnuO/oGiSxs/5/PPkLgrvOfbJ8ulquchqQ8vZirxzCoCy0Zvt4DFY+J/
rkE5gBms34nZO2Rk5ZWqshpu5kQsDhFaOTopFLzmLA+tR3Wt2HHW4TZY86nE85uE9hBzLYWZTvSH
Wd9nAhFUMQMLElfiFRH+FRYnynJXBXRyH4TO+oO4A+2C1drRqcWlmSwL/pxnIKHD3rRvmAaWtF9y
ur1aE7KyE1WPkSnZ+icXx61sTYJukKgCy1NS9q5WlVct2K+j9yDqS8+qPj5qcDzjGlvn0o4D3Wt2
bOn3PStefnMAYtXbZGSA9y5F2QbjV+ugW4Kc3PMa48LHU+tvY/9TtcQ/E50b2pmFgWWYiKnZDkMq
UF83q57cBxurlJYFLEthoUNBJn/5IxH/4QopE0mcZvSeeeUfCSz4FfHNRiQ5xd4l0uIWFNBgsg0c
UCYoCfGkPgSsSE52XYbIVitMbUqLgzjZHnWu3LVD6SQJ8Ncaz4RxQUNcIYvqCV7p2J06uUJgkMHb
JskqdtFkm6aCNvQzYe6ermO/vhk6Qfy3HLn8psLxZJz5aKFrVG4uimVTTkUN2rW5HZcLWudahGQ3
35NFSIaAgz1G7cttkqhBhu3bz+ew5NPrMBrWx4dWc5xj5Q52poq8F55wpkY/nvSytTmsHw/D/xGR
0IOCIECrk8xD9w8/QiVrAFQEE2y1hdsiADhkSI8rdLY1uIvWJ+zG5XCjJc5y0jWmZiqEOZNWmaaS
lb1LJq5ZIDOyZ/M5q/E9mNh3M8/oDY1u3qaSzTQ4twamUl47uDrCsEzOgU+GPQUWb63yROU+TXbB
VphrvLR/2SiskbjwcmhaK9+p8pv3OuxBxVW7iHzKi57vxYyqXgCP4fSq4Qugc0qtu1u+/4Fj1PO7
sYJdt13JdiFlPI84RM1pQ9OVqxlaVqKmlFXLNapk0TQXM0hEJnCOFoBZJdsVB4jX2Vj74p5+0TkY
2qwcgSCdTGLKoOqbHOga5giU9af8fW9M9Kkied8WHkt03ItqYFRO8hGgR4pc6lLFgquBVDr1WEry
cqG6MFb9F4EILk6OoJZhOwzBQL0+SVGCi3oS6rVZuH70M1cD9IdKuV7+pPt111/AO8ffONgzggtT
NjRIHaz5mXmRM3+bJlnLeBHSx7v7hMKqo0eUspn3gbD6E3xsomvMju3uHdvU5hFqIe5sHFBzsDNl
WMwbElAhaTAQS0lxhBa+uThshxOcbIKdDH3FN6lV0Qfut+XtTC5WEN9lZdR413d6V39ww5NaHXDr
GQ/iJqus1fz2uVU/kaBkn2SdF4VbChJ+fduk65D/tX9LW2LQnDM3XRIrPuq98xxUF+vblUdEEG9x
rgrd68ZOKHTAE7bOimQtO+dLgkMKkyWNQi6nGdEtlCNvWJDAsseD2gIW0suEMca4h6PNZoapxdB6
E4odg2Du8kYLdN6dKwTCzJpBo6NTgMo8hpP5Ig0O580/2rLGz0mys+Wo0jHb5k+XdpERfjP88Ye7
UBm0O88p0NMovuOzkPNUim8fW9oh4FP1uxqltAzO6ARojiK1kHZxuWi02f97bkD44lh0Q9StzOzt
+sCIXrdhXUbBgjCj7sy2O2bdQaHpuHiRIEqqVwplZlLIybOCdy3IhoExUy56X6qHrlfWKsKV2HOb
j6NQUMn3arRHYqdOIf6J5BIAyXv2wMlI89zuE56P5mb2Wujq5PXj4l4FIrlnnQL5/RZVb4Ce9mBc
5t6FP0/+B1YiHo6CIwEyaK1+EFAmqkQxvR93Kx5Qs160I2GZvj8sR7Jg9U65XbaM98YvRCgBxTqu
hhllobwMLpg+dqkMf5/gTbRoXDrhgFmGKgd5R/8BHiEoytn6h7YCYheNxneaEOQ6fGX7ogeNEncw
APlUm6LIhOJC/w/0QgE6o2NvnsHjXKkBafjVaxrd3Rhypmxi4ovrKpHwiPvksO6adzJIcT2dzknV
XqtmJ7Wu3CiSEGKXLAtRvlUiuuHS2r6V1lv9BOTrVJGCcdEo16Q/pA/komsDmC/s98gcb7FUMtTA
Vj6JGtuupqf8oejt0pYONY7bD+8yuS2DKEz6+QpoL/17Ii8Z/MipSbm1J9JDD+v2fMyRA/iNoPAU
nTDg/FSj5GWg8UASSonNIOdGv26yK96us62eos9c6q12i5ywOXyJ8A9hCHEiIDmUzRXT6uUL9rYP
+qQjd0JBWJ9hOecfk6n/qUjMqqE1frqF204hVkOy92GuP1+I1pHJXazDueK8s+3N4QJ+IcPednIp
zR8wmh3l9ccs07xVmANLoGKujEXRzEyVZwwZ5Al5VBtosTFdWjf6rwRFh1Ye7uRgJCGkj0yHMspr
bSSDAnL5uO/bb6SVXJNO8Qe3mkX0pIiInDhPDskp4l4714fV6/Vn5+bU5XFHFxNAprXIrq5nKxl8
JyiLvIjNyWQqocN/Jf2GUAiW5M+E9wHK+cWxKMLUdfFaAlo09rlPLKLTBr+W+inW9yZ/8VA9y0Gk
CIV7sv+FxA33uyWM6eyU/JZ2fn73s87C92lrQKO/uC2+zm3rlQH8f7KYrhTMFnm0G7CFM+qbWrlr
VyJjzJDxdYKNJ4oPuIVVixaOVZbH4CFx64TYipJ7Jwb/GSNosj3JExivuypLv1W+Q7R/e9NTzybi
qW+DpbFEinxMznIk6RuJAOKElqqWWNFTRnpy+vddT0waAVzm+4mJfCNlftVfryFLsWspguVKdlFT
Xb97pDqOh/5qfW1jdChUFqqPvvrngFMLjwQj/ARu9TQm/3DekZ9MYVFK8KJ7OgP0T8TJlg3J9odD
XdGtgl7vpfQ+xbT+dyI7fk4BSoJcBF4k6NILdwv2+SGPbCVFS75V3pAUsCi7f72aQ2CBRd3ICp20
CCxzXXkj8jVC2ViQ8mnflANGxwN60+m3iQvjTaeWaADNoWDTtGeKBujqqXCIdndHVzJLTAT9Jkit
pA7N4L1pZ1WSZSXCZl4mA9zbFelQoRboJ7M4IJCek7l+9iRUHeyCx44NB8aJnSa8qEaJ3e0VGJX9
q+4/jGSQWIHx1bTgdANU9ZKdEe7jWeItrBmwD8EkJ508/1FxPT2zuTPupqjbIVj4EWKJHmCwJzXP
6Dd8/pEq+2U3AgeCmnh1Aaia6pLPBg8WVm61+Kh5TvGNJN2kchMsWX3nJ8DcBvm7+Nd2QfiwLN3s
C2cjWoarWRCFHilmdF2eyeQK3QLoNpbcrWpmtz5U93qggzmKvgS0Z/XecfygEkRkL5vX693WqcMu
7Mpr/S3XExIO0DdPr7FIMdsZjdYqJjDQLIset82BTI5NYqq1fkU8CocgkMBbRwne8z8133ZjsMqQ
y5rhroEWo6JfpdfQ6HMab48K5JyMrIzgH6IKbWjsvVXJd2NBfEMa62sNjeJm4FQj8ioCaxfcTofv
H4kDOYC3eXQR4zlB643sTFOFgkp/3L2r8eT7c6lVOSHUYMEy03Tq8DO38cdKe1K/gU0fgBcGQgqD
BYRExC0vK2oOXX1Xv1iPMsscETk3/yDh5DmdpZf9SsIQGgWKTZ+R3F8LnGzglXZl7LlGPBmYo74k
1VkoaGagxrmFMSDcoZHIRLUPF0qdBQxy4MM/HGhM9gtKpFOfEhuDFeOcD1WcNa4euLANvYIKD2fn
Bgo1f43y+nSiYCUw1ZHtYueZAhdoEMf3a1rSz+6nvMQ/85e/eSc+5lwnD3/Dpp6XASCwa1mF2gVM
Sn9nMIB5OL59vlq60pc9WFbcYNOzbEfOGtruuGnhMaaX/lfxqx34+OMJn50KN9tTWn7BOara7ETV
fhBM8YFihbBoW4AGPyrvjPbnv9WbuKgSmxefnAWaz+9GU6BLXKV9wNCmGzwqme+LHsp4ohaY1XLN
9xI+MNxmyLCiMAciZwDzgxBejKHzNNhS/+AdY0l6Oo9juVA0mpGrs7HIhTDNPyzAIbku9kFeGTJR
HyNh/cN+Qw7wZFix7ReWkfTt+UBd/+z1FAmUUzdZZdjnDLaQmifr6rsO2ZwYQZQCq4kyq29l/Tp8
lyi4flerPEpgy9cm0itpHUqsDE3e0nEyv534SZ0Gfhv70wwMnwbmT8puJRc24FsnN7saQY0lCVAP
UA++FSn+FyBDeL9HaDlcn7mE880xITkZzl8vN73GsUvziYSoQpzWIiz8g5E+05GFlReKd2EI23ZG
CJ+wTNxOhhrcOKQj1lpEa4Z/N2BB00JyWxW3YtwotTYTQpl+iiMjXd5h17V/HD7QKbUrZr5SxQSq
QRluug2GJwNObc440cLADvIMxBpmhf5EbWEMzB0GvgX8GdDZhxJHZdTjCJmO/4TrBuk8dArnTI8H
VaWCnOjrZMGxMeTaoyFGht1UhkMvUoKuQtphycEC0T443mKHhbYNGw2s8Hj2OPCt7Fe4DJz+GnMZ
4UW2LSTzlo0LTL91umDmrtfHLWlXhqqwgwWPSCHCoDSTK4kbh7DBCUEmBC8zbZRRN7VCB0Ljm3Wy
BnE/TqchIZ2fmXZr2OV5qm/cw6ydxdiuGzYnGxawBAOzwA2eUJLPzYHdodGRz4c6H02GDyUs6d+E
qNcREcp/Umdse22jfOC5hKUDdhLuaazG9JjaVI9NI6Xj7D1wDLBEHqBSTxohd2KNsjuIFqPcZ72D
MqhHDAnlun92Gvyaa2GlqIpmp7xjkDC0afPfav2K8D3noX9M4nVha9RfOaD/BilhELTV9K8j2qPX
25wVDgVC9BEASHv2MHT99/iLNt1ZMNXUdgv8N+FFLMpPkC7f17in0VTW4YfYNKFKXmrmriMD1y8E
HV6MTwyHcaTlpGB5U+pnTKjjJG13kK78PrwvL6KzutZnCtpfHSVNaEhSzjItC7cWlPiKXmPVLrC8
59ghZ5NGxq1ET4qwbO5svNji239aTOAJw1cAoQawfJegrMHT6PDHcohW28+GUVBNhOnnq1BgKCuY
98tAWXqpoOuG4NQAH0gBZTUmlQCuYCCS36S00YxBL89gDwlV+549nLUuQbNWyLNzcaUfQzf8vA1S
kYXp30FcaCsTDwzQJrjvDWjTW/mRYIQvkE6GoWUiF9QvZ4vN+N7DV2mbLzXxrNjmTZ4eo1hB50mi
/X3tQQOQTPrDWSYOeAMbIKMQZjlg05x8UXmColJKSi423sIiNbUkneZ8JM05uDY4UH++xfvIGl0n
BFZQ4cIQjAK4UmEqkJg7jK4ogMUQcFsPt45Jv1cHn1+zCUe50L971SJit68hdotgJlt/aF77tb8s
GNlkFdyaD1PCuY4BzdqjQhB4Dh5PERA7HSiUXJX9xtSoK8DptrUvAKxXDf2sh4k1P5g5iXnvP+j0
XLmm8C5wUZWADQL2tAnStEQQjQZK1l+Feca0XbsiJLMhrGeGBr9rGKR+c4pr3Gq9crCONOL+2Nuv
g6YfS0rR6KjRX/s1W3CpxiG0LxzQl1kcqiRxuGVbXZwQ/BNVED0Vp5RIJppUSQNl9LdPze1pbhiB
rv/hacP5H0KKA0WCvXt9beNZWtIa7mWc0H+s2WjfXseMSm9c0MX3wdeUr+jTO5MiAx4rIyOxkbiz
4nkUTjiU87gIcIHFa+U/gYDuGWlxQzA//8YZ6B9isXsDuH5Ua5dhr/lUTJngZzdGSIGTTsdBsiEL
afJuAv074YedMLaVeK564e9WeOcFtkeMBdmh0HOKhJHig8bCCIrwMqB2hvMnK8s0cT3QK0Lff/4U
vSm8wBXm3QvsPqdNMt4Fm6j1fIcUbE3XmxzkbGnvvSghtx2EgFf4ezrgdkoiQ+1am7KcQI1D1IIM
s5Re0hVyC2QCq0crpk6I+J8HPLaFX8zD5mCJyHwPDIsZLOihq62EGpGzHqxiyhiA5V4qS2qS6znu
rFkCBNeAwvBXy1w0uSdusYaxeWFbOXShCmylO72HYBM2ExckUKywjrKREIrVu0sXi9crzq0oKtAD
HEELgP4JjVF9YLgkKjuyqo2j97tO+R6xh+3vtCKQ1y3vqCKwbVq3FDP8HOhGd2DNFFaZwOlliDVC
asOkXgrSEZzQqG99zcPb9SUqhnSK5XXiAZWsI70aP+VnGvp+rMwNtPXMYvqeFsYmh3K6ksy7tGou
JLfmnbBh4A9hkdux6sjUayS8vLEss0xx9WkqK+UFCHJ3BPWD8X6xkTVYbdO1EeyJyA+YoJ1WmEbX
phN2VTEHYHqljODhhMWVZ7aB2DRQYDUfwwrq72vk/mJeLTW0crqySE4p3ZT16Ddu7lVfIqg2nwsH
hihjQZWWoGu+MxhNCz+aDfxkz2O2iDtBxPL4DlzYawl0kfFij4X88IZy+J2knoTRxfYZf/AsiC83
9zP93ngJmAW6n6Qm4/ok1qeWT0y/SXKpF3kk+btYK6e5NrW4dZetyUtHlRFTIr7IzQviULOPd53j
BZzBz49/tvGkePUXJTHwr6kEsI1OxEjILvCLqe1sBef/34XdidPjYvFEQ7qRaEnoon4H+An2KRKN
APej+vqvbwqeRCZ8WDL0ZC4IasVOa4vDpapBgZLpIPSy4ajm1jAQlSJe+5PgwHJn+z3II62wXthn
8/piVPVdhtgO7OFdNk4x3tcbHv8J55eC/UffJOs54jqxHEYshAr6tuVR+ljT9SNXCnxwDk2872Ft
NoM31Ry4/JjEJz2yQw9r2cYEtVmo5sV7FIu9kzgD2LMX6z+9t3mV5aIci/jxf8ObCTM+J4ueWrpd
dcrt4V0yIF7+h1yzLIA2z7OlfZnJWpORzjI5Df/gneJaxjS7hL+HQco5VmMGZZuXW0V5hgxffY58
16E9LY4CgHKQmMZ+r6ioSo+81Iz8gtkhhWlk9b07ZyUnTqqLLVhmLpdOimz1/+U5tcVBTqk702A0
4OIYA8e67qW7EFfFdQ6p1+2jChF0eZgJQ+QXFh6P/UgLba6Om0zlRPBJDLko3GBL6n1W/I22eWSs
+urcA9UsCsqSHTU8oqQp++6e1XUy+TVySw9klPEja4a0oRnUCRz6gu9KNPuvBRz8IJSYzkWGwI+e
mKRmnz89wKxI3u7gtQOvWe6g2bY/fUjSByH6xqOhwd/FUFj734zjRmUuayjPSvNUJ/foJizjchmC
QN5mybVymuXbxGiSRbRvSgqb/CqgMBI/TiQLHiIu3gBRky+wc8FeQioYAD3xjhZIHfWnTxOOq9i8
/CZoxnnQjp6Jsho9Db58StYr0JDWhvhIsyzkJUEYCFQFg/88HMtd+1YjW8ZuVfIylahEIUeOnTPm
xiWNRv9GcxuCfrK1vPgVdIlbZJWl+5uLqGhALGVdDmFOIyFecXyQMuVYiglpJj/mK7Tk6zglyWaR
xq1hyYKh8knup3YVjm0WEM6qdEfkhSpXSsER5k4uvNKV/2NvWIPHm//faKllqZnIQOfneVWeyii/
0OmPFx3JareKLMM/1N1xU1c+aZkJY7crZyVNpNytHecjRyn1bzrFa5qKkpb53ufjcU4FJO9Wpmqo
XqtcTnSGxKeLN5/ua5IWoP2oLUc5VWo1BILnwwocZi/CJFwooyXkPED6vYU64Bb6FvJzlq6KZUdH
XXU51osvFk2bkzujCpZbHcJvwsHnGxC5sk+bDqhlCIVCETy2OJM6DpBXAm9jqWTowEnlzGo7XER8
PiUNYcO0zUvJ6Omai6RG4vd+NssLkFMKr0DAd2lF6lUn71eXTLpE8MgbhklOzWMlz9kJw/Ei76MD
SXhBACHKYVs/yZqkVavEUtAQXQwtMSwsZijAfhHVeezS5z/vrZTFdygKHVK/tls9Kn3B1K47MLyC
GefludALt7CckUdZgCvFIJgqA6hvceJv3lGB/1Ps5ZYFN46hz1G8k97RzwgOa5LSPQDm3OmBOAbl
Rtjc5OeLqaU/JeOkC9Ms+iSF1eP13Zod3g09J4mif9i+EXPGd/pafpO3RZ4ZxnCM9BlNvr0urvSL
JoKj0PYDO52fITk87spWhQKMLITruv5i4TFaxl4wDaO6emuOIpiGcwCw6Unyl3PKds2aYDQUCRc1
3iJUPdXZFvz+WkkmSw60QwZzPLpLxtKX9cf/nL4TM2z7q3vOuD5K240MGJXG11SckUixTpc+uktC
tMjmqL2muCKrKjugRQ+WNbWkQ+JOEz2IssInvDKwGEiujhe64SUtG9cdTRliP1C7Lfz+BoB1eN+t
VeAeLR9pUNG90eK9z6dHBX65Hcj4+icktTRifrzcZuXrGYIXgoYJfjEsEPFjvVyfK3bbh8zoaYOC
Gv6Dz4JQL8UmNthx9SetZA+xRIybPdFV2oafE491Tzwa6ruC2yKpGkbQ9DcKfXjr8NQWKPJ0KmJA
sQDK1OkX0zkQDdmMahfGQ3Zl2rs4J0XNjh4JTqAiNzMahkwBeN+VSkt7i/x/V+95vvz2Li6kWSx0
9oontv/kuqud1aJwTPZqH+W6RcDgGU7wqiNOb5rXNzqjk8tO5dsZd88IEvkCmszFONnaIXiarGpz
PR6K1Btz2W1bXuce38WGPvuL+6qozXtG8xNErCaBGDxZOSAR/iRC6G0+nysdWfx9mwUj38YQw2rT
GUpQoJ4wbRxP4FCe5xkcJBnGmeNctHadFGTv7yTBoI6fc2+a9L/TreFwOX8nl1t2p+BCse4q5+MO
HW+nqEn7X6/NmalEfNI940bzKrly6aP/CpCjHsYiDKDcuHE0+jScN7vDTEXXDz3WsNiSKloWeGfA
wZm2gEVMxFJG1EzunbWb8E+csp/U3oLf70luJSW1Mnog5iTlV10m84DSDP2+jbBArx0vUuyvKsRE
vz3TDFt50B9mu18BQSywFpgLJ2hhS5/DHhak84xkTLznMhYl6V0woDzAWEeUi2N6cfIBKtolzXNZ
VPxSX1a4zuDOOK4okBV5Nx00rtBMXiISz6iIDxgItYBeU1+lSP/lLECgH2Ia4PZLwOj/s1zr240Q
5gk8JbpldPE/VsDqIyOMQUHqgeOWW/M+lR1Vvguweq5ITRBll2tbNwjBnQyYyX2IQHGuppJdPwQa
g4lY/6ySZiZpBIsKqWVsc2I47hpYvXQJvfQQsgCA6jFQIWdSWJavNL6EIQHASdfFTzz9/pKJE9w1
VqvIXI49Ni7OmYKU1oP2t7IaL1Exl7e2pAhVWn8cLGP+8P3SZpVfhW84p1mqmN7orkYQXa7U10IE
Sz2ywoM1FGIz/NeKmwNG0Mm80AD8WxM5OTvEF4kSPp/6tm6wmYPxPxzckFN95fd6V9uppPETCBQ/
T/F/+ScHtf55EmclKwEQ6IbkCeSYMthrmxoyq9MnD5uOV+OYSmKDXi291jGRMPFL8gSPB44hDSvL
uv0KN9E3Lw54GZ2x13FYLBJWdpaBIS8SiRZ4uT+k7Vx3c8NaJzR7s2f+5eVOD8p0eiMKLG4kZTUl
rYzRiGYdIur7fLSVJ7qoGpC0BrVl7Pe/dCEl7jQWs+R1fqxefeHLfC29gQ0/xmvwFMMQRI2OZk39
QfhIkW6bq/TXqFbJ26HJsy9BO8+rsYaS0kbAfVRjBGyyBYvAhF2q1aj9qE9GJeqXT8ik3h8cObor
S3Vf6WGLc6OSC2u1BQAiGd5CwVqEaZUC1w9lF9fBnCwqHWU3uKFQSUpwLrKKsfy3wbTG7/6bZ4q4
vTcOEbcTzh4Q1Shid+c23ydjF51iIrCG/Qb6Kalcxohng1RceKbWpfhZz2X2RZtuZjRG85ZyvHuR
jWVBhZ6ua5VjTzATAZxYNI+IYm5AO9+PJrNWN+VpHn8HfL043J8u7X77x7smrzuWLtedETm3QOVf
hckmD7+v1skF61pPboMxjKJ1NgyL3w0nxCNN55CS3Oqwlf/bKeHn1t/+QHmdqAQF0CO61+HujOL1
3uAlJjiAQnvHQX5GZqHEd80yZmV0NZawwMTGiI7lhMfuDLnm8laH70amHUUsXwFd4T/xLirmXl5D
PbFIpRv4rdl6WoXdgVnp+gfhhxfZRHhZWt/PrO//n5Mu/AqCgUdHHpH045RHD1IusopBUaGAl5QY
s4LPlzjasQAHH9+70bLyKrR4giiI+sufKx72c5NR8wHJ1+Rn7whANCjhPhlsaDvGmtKfX5RtfPDG
ZrEJU83CvvoRGZtIcEgKhTq+rGWjELa4D6h+hrG/vpog39LJ1ZgaehUvm2uyKKBAM2A26uGC3ZwK
l/YkPeS5pPPJ2D4W7xCr+HaVjVSb5h7/gk3T1MHxmAjHaOBD3A0LLpGbYGO/I0THRMxbyO+SiOFp
aGEwwLUGCw66PJPj+M4/GrlC6uxMg7e2Uu001sqnV1Tlybh46cX09IQx9ifJsH5wqZqz5UvDGNwg
ChYG2rEiSXSEf8wzdoUxUuSHivvhioQ7e0gvnv9KC96oj08KJIrS6WGdbc44h+6OO6Jf+vZ1fjIJ
47J1jc7UuIzOM9JyDhcM8XaCsHHtJsSm4eqfigFKY5rqDo0tMOBr2JlZPg1fRTS9c676a7thBrEP
muUzmEeQ+dUeB3qiIXuCMPHVHYltFkkCORLkTJHm3lYhAT2JiMOmKdhJCCdGbPfbbCKOMT+uMppb
GzqE9QlTE1sJ4MchuGpj5fTc4LtubJxSc+xEsb/RZamNlmmKvyL1cAnefoQD4lHfcYXiGKbM2xeB
WH4qo0RSM0gB64c3is4Vn226VXh1jJHMMjnzx0haaCepbHfBaU3vC/t/9VNS85t7J7noutCN4AYk
tAqeGItFo/nMSHlM+mFzrHaiVq5n3bwoVpzJ4CUwXUA23qMDX81F+J0uOUPVNtPAztLiTA8sTESG
Rpgk/3Np82AFv1uDZNHKZljCfWhgmDOzYlybuNEnL5Tbve0fyGyNrdzH0Rn/7E3UbaxFZrweSzwA
7oHDFDA3mdFEhNFFuJFgXTa+OH49exIhlUHHmGo/H9Rm4Aul5QlLSmywvZOBV0vi6NsWfrIdubAP
hPy+J13UPT5kw7QtKsPjnPzU4TyyMnsaJE0XMJ1rGQSiq0C9wZGMa6WFQt2gvMFon/KZz0qSIR7S
DbF0XIyk0F0TTv2GhOGFiH8upZmDSSmrdAOx32OuEpFqgutEWZM/L9hR7n9RRwuYGRKYCZwrLLov
YKs7o2CtZOfFHHRZvC39mclhf9e8gKPYKVbBEeKfD5i7VO2FrL3bRNb3bV+xTd+y3IwbNa+y7AUV
O+i89lkC0RqOY0HxC16BdbU9VdZTpQRY6wmzT+Dfepc7bOZYP4c7J4cCnhDtiByZQutZKMh+KCTe
dZYUOrvLTn31DM66ke0rUpdJ0wO10ZnLXapWCp2s94gvy4r/CWbWQGkhhGhSAua5IkYMpSYkVbkw
kq7DN4zkujjoH1TQVppZH6dqFYwAVHGEaha+rJs2PMhqgDQyai2jzgfxGNqEzozi8Y2AXcxHI16f
X1Jf8EoiCQcWa9ndJ+xkWb/vXgMQ4geE8heqp7SdrlLNGn97T6xbf520dliP28h8melWw4Yd6gLQ
HmRfi+KlAFYBRCLj2QhGu8UZ17MyZND3utqyChQi0KYCn1z7NYYND24zUIZYXQhpc58H+0uYRCqL
MryjmrOkOPDfzwfWpL/A+Vzf99kbnFJgHkHmwnAQn5wYvUCYKei+RJOE1+fAgKfKRGoC4Aj26y3L
X29t296Zd5Hg37eruiUtDP2itGo3cPAcaX9ufV8GWYmz5EmuufQ8y2uARZjxg4WPZv5gIEv8ZXPF
39TgxSBZ+eD+NnTB5/h31yCRFSbB/kpYMX1UqV/Gy+HrKVQ/5ZgyJv0e+iomLuH7psxkGswufciv
Xj7k1OyhaIBneAHu1lVrz03MSAag53eB4fcCKl33/rrGynXVb63m6NUuK6Z+3YwqXRR0hUFBqbMj
mMxX7rurcSXJhjt8lepIu8/r9f93lDGgENpMcUj3ybc04h4qeQkDlsJwRMyU8W1U99JTIDO7YWcY
OAHcS8jWd2iFlI4f1AFyINKxu+8StUQ4vyUT83YMgaZDiZvpy6PUk76Y5PZ3Br9k8u3BHkdGyko1
qp9BvYiH9f/r7gwSPMNbbY880dg+DJ5JnabFj05T/AUr9B0/RqUyEGFsWYz3lV/2hxrB8BwXUegW
lDCfNOh/GXj7+OqBrSQkYNyZIcMxDZB+GNJuYuvvNZz0PgKxOP2fP1QL7dfRJPkTgEuXR7t+fD64
b4RQMYjIrUGIA6q4O21o/08HDb1OaiUvyiNPHV6BRUuc15QJP8kcbEzlpqO/Xipn+Uiu4LMKwnRZ
jdagjeyEWXvrOKIFsyRSW9F2tdcAlJvNbIoQ5jG9JJz+ZLY6NMyynbvYz2gF5hYvdTX1uMYCDJ1h
0C1wUFQHFuhgV1youdnQGsNnZHd6fGGI7KIvfsYHNM1ScrP57RswkIuLDfrlFVa1a0Q2S4Ioy2Y/
Kf8zA5QyHfym4H5vmNgcDHWNe3gtoCsx9QOWcdsRRA2YXyFOqToD18Y5jj+HoHbolNhar9qGqzSd
0d9XXU3TYK7z2Hv1Tj3uT0m021R6YpiIwBiUAGQa0WGPjLce70LIo+g0grK8I8ODmP5DzIQhFDTj
967uapjZEa2BXMCTxSCHavRDj7MD4x+KG02yXwo4aXr1oNDtj0d3eJR0OAnPLM9lq7OpUlgKPyg8
qKbYp1dL++q3jYoJ7aVA87BpD+8kEyzkWW+l5+IssMxvWQjSth1yeExYIvrQQLrRl2xYdyDZveEI
tlU38GQFT3OH+BAIUVdqekJmNRth6k2V0eEeKjUGoZe5LFFbPTdO/GJUI4xyRzejzHRuNloeyewU
gafDR+dFKDc9FunKVQJr8RrNoi537UnBMlJYLWVChSVcCaaCEqHVLd6U8iWusMA17wXN/KTdRMKW
lFE7dGSb8yOKpq/R1LTSvQtN9MjiqDjXzH5xvwy3yCqpy47QJmXRU5U8nZqntnm4CoX1Pgi7SO3M
5z4GkYGzmpDJDCuS2NiFsVwoVyXbRpFYeVhyXJ3gLn7/TKuQcjOKC5jVR8LL5EKCzEnvHNFtWrdd
Yzr1+bO2oKlqd4oPHgFnVz8pth4MvrpVvLBbEojHZ05W2HqoGDwBumv2JVU2u0sPAPNSKyp7maXC
c2AYypQeeK4sq7Iwr19fC1W8U7tBjB0LUlUJWOYHGj7LebBQCMLFGnH2lnT03toLXI4vLH0yEPo6
rJVjX8sljbQFGGaS3hkXRKoPRe5V/e/TpK+xX6wiEuSrJt4T/S54V+zw9t4pHsyfNde4NGURMOml
+Oy7YkwBfqHnQSv+lP957nHRw+b6tAd88v/oXwcGtPJDu1+0A5+A7gVPU8/XpiDVCydolq1rhdJe
S49BLXXMXB1hBHf1ZhKIKKixQDEx7JUD2qiK1rlEZ54aNXGfstr9/kTLqpHKTH4Hk6Jt2J5wLjr7
ASELCvRwmK+M2+GL9hKmZZMCGIfiPl+SgXDhQNQAKuYSGegzoQgx9WSmQweOb58paOiDbI5EnLvq
PZhcZzy2jXbzhpkNQXInN6vqA90IJ2xBPdRGPhl/HDtrEYnzXMl6Ees1Ro4w+LFbxdrm0QaxKO+M
mjC6kf4yBNF2aM4FZuSczEdnnKosC2Z2MgC3yV5ooHyxpqc6yQM1l/YV2cH3xKIDWm2KIM1gFDsu
sy7JZEFE8M8WOjE4BKrdpVztzMWG+3D1Elm8Rg61jCN/aJzRrwT2XWPLWsWx+U2eAcT7nUTpeUYx
/pT1OE4eYUXFp6FXBrnji59XmLqhSwas2jpC6BKs620a50P0nTcK/3+XHEiP8s0SzIOvdP3wbfM4
gKrRb6wr7bVRpT4DW4NAdGJbPySd1CAHzEa9rFcDK8JXCfWDkOQntQSh1Ad+jHHD8LjVQvKfw3nl
ojicp2WgZTiVHBQgmdOU4mTYo7SkCl+LStgcvldch1o4avVjsBXkrcPm7YIGB0ngbyDXb1FMSx0Z
hROrUjdhg+F6kVwhql2f/K/M8bEqMlBsPaVAN9xFvXPsbuEC8y6vZ4ITX8xhVXvAqPcdLuL9XTv/
HccZKwZ7nDDRJQd+cg83HJOj6rbzOIstwuSu3hSv7unRFNVc4XZ/xOJJW4dftfUGefhZ7JbV8JyA
4IttAYn5qrGXuR33oJceUS4z8vku1y38ZBAH/hU/E15RzRVFyCeaOiSCzHgdkoxani1mje7ZMaoN
XTHDA1p22R2uBY2QiQVTcNc5unWjdaGCzM27/ozSpV+IjzvZxXNSUL3UAjfT+1JBtc60GJ9H7QCq
zk6Up5RGGhfQguCZxS0YfGcUwyRQDEhscggMSnbu3IfJF6l2sSEhb+zrHFr+bLllsyGtwKlUc5dE
JwohmQ2TSR45YxQQqVsqNJz9Jx/xEIK4ftHaxguM1X4f5qgVPJqsrJgjTOZ9PVBG9vBYwE/N+u9T
QnurXHXjiFjHzlrXpD9vwy2Tnf1nxl7hBv33aWSazFDvXy/15FSAEgFdvMPTuAJd+v8JGzG7RqYf
1aIXPoIwWVvNnzeMwXOQQToDt8fbhGVtQ2by/grunYP5vpmzZA8iTC2uh/W6dEXRWFpPGPpsyVVx
BgXkpKkSSRVtTMESTbCSirUiTGUIgjemsbejBCx1PX6xu0nknaYNebSpxpgSodiwuRwutPoGR+Xf
pU/p0FpcWpHaRBn+xt8IShoENGp2c9ocPY1AzjhSStXHLq0m0htvky00RzimshM35DHxQpVcQ3bR
+i8tOjmvPLMvhw5vUD/7ZeTeRw8RK0aq33vcUxjd+ms/JfUGLVB05t3ywIpqyD2m33qWGl9HluJy
hCoF42KSxjVzItBSU+uYdfbpBVQWqY9NelvpH3HC0gA+pceh905rJkH6fU2Zt4e7KIzGSkCwE3id
QzmU7zOpMjsGuZdpO5JeHnblOWNbmIOKXDH42ByTdaT+emciWWiT9hfHnEl6eS0Ryx3mpQB/NmwA
YX8E5ietA9FYZ2+OxJYtXahaWI/TSM4txq15sCiLC2ZBVa4NSfupiwVYD7DBOdtIHP6EkWs4LOdi
6OslI+yreL8AVBOJXtbICOv8862waDGub8CCroZFww8z/whCu0A7OxpdihuGqd2UDnDvJEzaSNQF
rY1pPN5DCHl/fFyWSSMuhcGWMbWceZgm5/OsNceOmElz4RFSghBDqUhtfaoR9CrddDiouj7QgEGO
UCoigBp25ZosoFQQL16eJZsB8o+eY8h4oauqS3mfU50kDSG5nD6SnLxE28fXokgBD/DgdK/UBM4v
X0MupCLs/ONZWYo57EUZrIk5i9jawgoDYnuEBcdDVxbVLnMkDlOqNTQ/ah936DE88m9wZTSWWId8
NNl1xs/I1VE1ogW+CFNemcTdix5LVKtnlAF/rSWiMAD/7ztsNHWpYo97n39rGWYY5zZs5PnCtPLy
l5EYNPPfCPxO6AMXZRVrbp2JRRELF+DgM6eU6bKvEYp9r2JVpmuqEtFhbauZplY9uSrwnQ40VBdQ
CuzzeTnV5VP+AoV08uWiCy5xxR5M3NjbAwlKxosgijxsJEo7QjeWE9IVTmYLOlyPitWKnBosEBJj
Ipe/610cIrHgS6YPypq2KqyA9iXie7R4SADVJrVRyswTFcrtDeq6BJwSY8oOmigDt3bjD16K5oF1
S9WzTQlliHHBKsUdtXs63KIhEbxcmUKmSWfleks3NgS1zz+jX2JomJdwOXb2CBcMLCijaKqphf4y
Fx/ioyBLjUyqNGiDUsttDFsz78485r/CCtS3AG8YimBMXHwwyuIAn6C5CEKe6MAiWBcdYwxaxwcJ
gc/VbjkXm0PYGjBDwohG/qlgQZVnke/mvXKKiouyRMDqb9CWycHomZG7KoGy2g1rTQwbYau9OLbf
/3PYy0JcmNq5aqDIDY//Kz9JWa1y8ikCgjoy2A8Bu6iKjUIWAr08BSO6M0UxYSFR2eTxrdoZVM4v
k9kMS/U9pFKZHgOx96Bc94rQJ0+mhFdU3du4/i+FrTAnNqXFheszr6IT3UybsMFhNGbJizGzdJcU
ht7pGd98toJf+0WiGs+8GL1kSeH5b58luc21Lpw/i3Job9iM7K80TlbkGzGMqvUoGAyu4dxu+pne
pBePTr2IxDn0p+aJ1G3k1ZwMgnnulmwMN1IbR3hAx9+M8p2LgLriTlTDB43TzsBm7f+MLD8wFCxY
rcVMlezw3dGDo41y4+W8viHSj5u0aoZpKOiM0sp6wV52Uq/SyqNyf9zeuI1QGQiR3btFaOJ4RtGQ
gGQqI6HSL5wvnYt6co/wNiwXjaxAmfS8gjNJBzadgOcM8Rj8mDRUFasYRai0kp9J5CMmwykuxurW
CeqohrVPttKubG+NTJIpcBr+/quigIFNDQGmjOridPgICdCCBEVcvKLvbUTWAghc3KZ17MlGG60C
PamGb+Kkih4QaRCQyWaApJZc1gSMMK7LG5c9BRlDisAc0SO1usQsKcr11ls6hikavCS2JPW0IXEx
DamoKy7/FXVRU1r4akBEb4A+qgULkzA+TaxhanK8w9SVyjbZ1T3dQGErE9aYIQFn/SaWo8PCa/Kd
qzRbmuwOVrsq9k4m4QYZUry7SKLHFFjQec7wuYNxXPmsgOMk5pwT+71PjxX3MrK6KeWx7UpPa5es
zV1ettcS72UApskc6NKw8oeUV4okdhm1FaaWHgmI9spzwdFBH2uBErt9loAFgULFLrCLDgaCQOGn
md21NkXbQA5MpPGCM0ohWP+kyI+BGQjfNi2ndVx/7NnnJlrUlwGeQ6S3GXDUJc8kC5VOe/y+66KP
tGX3qiMbC4ZMdyfTxz0Dtr7QHcxVL/Z3iA85+hgYl4uVG1BJxO3iWjeRDD1sablVQGCOG9MTw/EP
uT3egZqREft+2coZTCF3RvEZR41Zqbfy2T63jYI4gW2EaMqLKLWm5waYeFgfRjXbrM2Jlem3qN62
eDJ+Gk1NUT1da+xzXzBbO/d4jA/9pcHQio3D0xIUYOBIRbr9BOKCKlwT5nPBtUH9HTuJbXHLMCmL
ct0AKgWBdiNSE1ZuEeWQjv5hs+AcOcyDCWuR4+zkWiatTrir16ld6hj/haflb9aaQvo64FcEdhsw
wuilYCYz44GV+e1WuRLLTO8U403DZ2Qfdic6Rgni1iRRqXLTc/5HbihOP5ZhjxeFHKUHDF6xHJU8
wfIkqC7cTaaqyLFwcRYdViQ5hB5ZdjWx9oOskV0HClarI8W2CAK3qA/mtmftPpLCgZ9MkYISPYA8
5NS2VTtKvHeqDd/qb5js/aW79HacYkfblloFzDp3xYGAWDyk7kYVRSC1zu2tZJmeKRX9eer+wXn2
xIxI4xUwdVDolkQgjiFDjG/IrCV//KcoGOAUIStvm+rDnr01rhGFBGeHdkRUpLQ1j3+MVhhEc9yB
UcFpyVOFPTdtwghrGT3UODaIx9o4mGGsYTW6WQ/2QMFsjPaSPVrWt/hWgpDLZM+dhsI0ZI8898qC
C46Ld4OoDCOq7ASL1c1MItzESbWgeY/Ip2DwJYU+HA+glmAkNPo30LqBwwdqHcAQ5n5K9pKGJAwL
SRpcRTDzUPopE0/HWJFVv2AlqwAyECnx0MbaCEe+B9JDWX0YGVxR2Ha7oR7ON5mFmSBUDXuPi6Sv
5yb9uWMdTWlfxMq4bjeYOcX7/aLETEQ0VfrePaRRnbBfxJdBZh8kRE2DZyy2kd3DfZezOqoDm1W9
TygGyv/DtIZQerLL1zQdjFRg/PxjYS473WP2dCHoSYXiYxGlnmKIDuLBOiBXJOcy9GH06eT76IDo
6rGuXsgCRXYO5zEBnXlpA4TvQktUncPPfeM7aB/zEFtgtzGt8vtLFHX5GbmXqF6MojzLTng7Ov7j
GZLTI/Gpu0270KIitpmOnteqMN0A5r7S3rHswc5h3QXj0nE2jKXPjNv0D2KW9gxzt9NCC8h7+vSt
IhEtDvA3z6fqNI7pdDO0Gx53+m1V3Z+fmBJxzBX8oELx1sFFjg+KlANDyGGZYf9iY6St7vP1Aw2F
j23x+FAS6KIwYhYKycj0sCPXt3j5+P7e3s4HWyx6JteoRW+y/imBBIhNlG6K2tsmOw5csDrATNY9
EgwV/VmsQlUowwa5/q8JoBwO+i+9qtFhOomDWPQk3dqYv/OYtJmFm8VS17Dw3jFfBJiXPzlLMAsn
aWywuW66UHqalbqwOR1shAnU2gtSMbPkcPOH0SuVwEQL6DtabkzbgJPG0HrTymO3uuDjiXpwbr7k
F9DWD55eDro/l7dDzHxXxADlDyPR1iTWbmSVen2zldjCKwro6k/vJ7yjxiZ/sscoJ6cPbaswSQCo
4+TIVJGflGUYOmDHKyTXzMO6iSFmVTrLkeMvlrFasbXgicmkJ2E1zFNfPL0I5vvjrLQyI0cFDdiV
lRG2qA8/m+g2+TbgKQ35yVsg8CVuBN8AxZnTtkh6gckDipusypmRM4AE3k/b6g0BQ44SpZRRTJKB
I1rxqbIw8znToSAQGK7t1ywqhxxW4rtvdCHlM1P9SB/yha0YsCIonIHegHqkwXx/OpqO+cb6ufR2
O94Bsa0hmqTKnjO5qqPyaWBnrnAHCigDihGT3SJmYx57qVEvIgHiJCaNcqubXqaoVMy/hUtZvJcW
rikj6RPZYwKRrwtkTS516vXKkfbyFtHGf3l60S5QJGqZw8uQs4ou89JhclT2Ilfh0jQJam68kb+v
AZra962TScX1r8qQFRONtd6BTA0/jjmYQqOwiq+6PIkl+gQwy5fLzKNlVBc+24KAOfCUrq1UqVhL
A3RaruqaxUy448ZfmtT/hDB1CiFhq6Rp+fe4vIZdDE0fJvtHyzKu1QY+gkEpSdzjgJBH6Nr4Fsnl
0Pk8PlL3HyfMGTfUKNQRAHK3mblWBgb4nUeQ1MF9MEjYLFjY9nY8HP860wrVGaUod2ZUAUBnUgJl
0P7kSWwRsmRviqZpsu5rJS85LTkRBANM5auHvFrhguKIAXkNOc61BAy9XM4l71V6h9oK9pBWBN7C
f2Z9gKGgt4my2oY2WP2K+5cf1dpO7eyYVefQ/C5ZKGfnxgFsv7pOHDhSwDrK+FDLbc6OhKwq0q4K
qYCkZopWGJMl5U09fZPUzfwj5vxlSWekWbt/pd/Br07maahyAxdIRD4sfd0bqyft1Oyren3JQDws
B0i7xU355gCcABCP75upH6pj7+92xq09wgpe1Q6Eg2zIR+Qgg5ueQ90kU75/JBogBdrn9X0GP/Rv
BXRdWYmkxuaqvn+ArB/nEiFYQT/oatN5EGLqrnTPDW4HaVP3maJC4lrFgCLtOQNyvqmeELPo7R2G
/0rKSZq/DOvRqNMhabZzYr6cpna4NQrdKW/H9ZxoVmjnQVMhcs5ofrWnm+TlxKLn9ZJ2Fjlj8C0b
WgHeN30VOnDp0dVRqSQS6qjpE2ecfsgFM5I7clKDSZOP9uR82ZsOZXq4jep8dvtJqUIiNqJIrJIm
FJTnlxvueqk4yXqUC2zqw9MfOhfpN0OcqN9EuSOFoqTaXEbNF9ohfLWrYXnVS8cX7oh1MS3+4NIz
zp4Al1YNiz5Fzvhb8qdtTo6z16ADrqwmXp1R0Vq49rgR5natKVHC5qHuZ7w5EFJRtP/Rme7wSjUz
vX+u3T23qEJELpMaCabcKhB3iMQZkvI4bKG8QdNgIWNfnIZkNkW+DKNEW4qF+8dlGKa4HQ7DJcCj
8qlvnsW/hI8xEvFSVRwInwQsX8tQMW150ONw7Io21V1InmeYQE9IorW2aZuDdQ/C9ifi1Nr5Kz8b
OSAeRnKXQA8+Y9eLc+HEEE0TfV7nhj7vzJacgPi43exGqweBDeFJ+An691xhyxNEKQtqCU893eIR
AohM23i8er/vYw03/zj0uD4twgVK1Jizg6OHTq/lzOX0m9cK0onWt1zrww3GuJghbEWYVmEFK2f1
p57/FYV32tXFPjqXXev2jo+WgBJHt5RRZzPg6UUCks8lU4DmhWU14jToPzYXBzzJyUNeoxE23IQ/
Kq6CdD5Fd5LrWSC6APXUm1yLUkZov4K/cPxEsumQpAw7gk1LQPXOq75xTs29V1yyBTlRBb87rxCX
xWNxUv8bdf//JoUEK3D9aBsNYqf4s6dGeCe8U+nMnxVntCzyHXUCAbt22KYcsGaluf9R5EJIAoaE
jxUlLa6xWw0iyiyYezTlMctcRmcO6Lj4VdbOWXBiG8johv4Tag8Sd7QTcE+4MHrAh1/pDzk7GFHF
cyv3NyuvbcoKjlF6KsU6gpFY8Re2E8j/U0qOxaN+9TBsoucaOfhI0r8nA4ox5yGh5JxB6tPdUm4P
kcOHTbDgpQbVfcTrWP3RFNI1VXmGpmpjBJMa0Rx7UYepaCOkmZHXaHPo3/fzCRYSRxVypFHCLV8o
ZNuHQJ3RKs0EADy225eEU4NyWbGOIuwbZnF7c5nuiLN3Q9lDt1j0l0DVnZD61Am4xtdNca5EjkYS
it9ni8Jw5Iuvs+c+MwmfZZLVpppL7EVDSUoSr35SOSzdJUCJHYYf9BzCpuf4hjm/XoJc7zyE8pAD
tMfNbZJ1Y6h1mUq5+Dm1mB/ysv+SePWxvvC9BW+8mLCsOcN4mVXtxZmCTqkn6JBdeaqcjuVKcF1s
eaSXJ6Ix6LEJeLOuIz/aOHcZK6E6Ey4crOmWKPeRBQNhsekp9qU2OPesdgC0koXdQ4U/IHjfIeiB
2ogzSGhtdza5N/ltVmI1lE3jwmF7G99pt/c+2bvM0Ex+H5H7LXOxswcZieEC9ovCR9A0UaZI6mWJ
JBUZwubk+gNfwMW6cTD2uDX1sKTcVhM+qmN+s+Yulov1HSO/L9x0T5A+K/Leiz+EYnejFqRtnSC5
njhv+sgpwyOBpjwx2QWEwMZDTAwjp27uKKaL/X/k+XRiff4AT45KNu5qEHmaMB81c9I1tml523vU
8FzgmunvtWTxJ7BAhK8KnnVjvPDWjbNQwDENUP2iRf064/7i9JpCqL8OITS4eCemkMKtcZKvCjzp
AD5SIBxaDuJc8kmLX09tA1N3elrflRq7p7IcqQxiRi8N2MicyEi3e1azxnashIOVfDhtf3GQxbQH
rVcxkS3ruEZK7Pt3mDgvFS9jRjbpnfwhF9I6g7WUrxLzF7NOCikTVarTKAO6RdbLblP3Wk4Nf5xw
zH1s9SR27XghkNskCEBVcoBniRCcEuA203I5ShmJqCAklCD1dUcnIT732ZrVH23U3bd2b1qQHNTb
qt+OCVn3k6tpBL9HoclwxRUN+wY4iBJlwYPo8d8/0slsdbZyK3oLDf32lZgp3tajNNwuzRXq77ex
ua0Tmhe5mfOzxAbbWCkYGqNoxXeZ+B7zQfQF6VSKGdC1yPGuQlUdGNyzqMCJgWRnlhBRdJE43WF/
gFmupGkKqOBMBnQNrLNrEJrczicWxUxToYAW33yPM0GnZenGwBIohd2hAcTXI/+e7OGFyRZ8IBwp
wo3qd3vRCG3K2b/xXw2K12nDWFWmgyXdcSmoXJ4rYMp/SxH8nrmv1EaABkcAfEo28/e/MD7yBNdh
aHqsqOYxg1un5IbcsCNr7u6j7BPLZWPYfqbUJ8UX9wtwK1eRUz/HMkQaXuEjdeSdcEDnFbpUXtvv
66QrKGPSYVvyT+7Qtv3EJ2FYAfD6VaHT3Eo1ZJIAIc73iQxsjQfCcQ4kJ2A+sJ0gM17HOgt0Va4u
zTui6pjkbiHZZ+OUiqVv+TX0b3SxV/b/RVoCaE90pJYiZE0FW2X8X64vdFAyI37Yr43+O/Xro/ZK
XpFf9RHLLLUSWVdBOflmfxD8D6FXDnmUERg2BWiVb6DANp3WEbl/HFeZB/IXKEqGU5ky4wK/Kiwt
8yN9sqc2cJZ40s4aTDtMWZ+XvcAJPS6H9YDiPwh4Jm5mlDx9RmSauoewOYDlJILlTSrKPPYczEXp
5j3VGskMyk0HAjWFKKvJzhRySkFaiuDCorWAOtoxPGkmIoANxEIdWf18cEjtopgBYrAcBAoXbUTS
m2koKSynSXHPDqxygkNavYXvm+QlVlhmM6X3bTMfDcjFc2O9qk1l7uPkTbUQQQci701egWf6mhHi
qHUq6HHtRibmJN1Xm6I29QX+uVElBIv7tp/9NUlg27/2kzHBBMA/tQbJ0d+b/lBYPRC2p2Oj610z
grCO9LHf0L1Acx3B+s90BoZK78T2yi6Awhl/wT5P1sPsRndYb8ZYGDhlICI0BkmLH3Cv09kP3d7n
Rrdc5wWJiDvJeF+oVyEj+uFTV2nS0g0Ff14zEPXgOzuXBcobPilTyTx2UGvL0T9kzAfVc3hij2aU
a2TcXe5z5Txy7JxB+pigYVCiA7h6vGy0zCy0A95PaH4tzkwOKG35s23fDADvEBdEW9/F3IBUpC5o
yW8roND1k+b5PhyRtJL80+b2gHIZtnrIyz/vXjV5JWLlNjnJJmjdYijX85KlMa63plQN+OAEdvHW
OCr56ebwjtV40D5vzaDcOxNECO7bPzEuTOC9uqGPnbdaWLIdJYZTSZ/9KJi8BM+8MGgkeGXKQyYo
k6Eg00GQfDfMnKoEYs/Hfq7E7feye64syqEi0Uxif2Y2GaZIhjPovGz4eIl77I/flEPTRJbJVkH0
eyjAIBqvuiuOjdsfdSzPGWh2beWljyb9AhQETqQ1vjI5sRStZ5F/zL5l3UiiJCCiDiZr+IPw5fZ5
wJTg+Q2uVlI+Cc7wttbNd3iUZRM9Tqlj7qQtk0WLgHW9RSHcHZLGjhumLGd5LpmkojI4XChCuelf
46Vv8TRz1yMHg0JQJx9nAFzqDRt/2/yPTifFFeH8GrUryrs6R2UOfttEZKwdcRNe4Z2vvyJl+hmm
W42Y9z9b7b64rfYhGHlbykZiLcyuHpJBxJyGpdav4i0RC6oBTrspVy79SbTUHePXlNUtJcg6IPPo
EuXSeVSRlCIsH+YHZfskuwpWjThtZ0AFStTj3uVvV+Azp5xQvKkdCynlUgekbQWNDj7zZoX8rSEe
Rv5j0pbdjvHCkh59xA9J/caI3IEFT4rBs25rf8q/daoHUO9nZbm3D27t+7cWaPB6wK0ydH9GcMdN
2kxDDsJxHdO9vFVtviU/GWUtnD6sUIzETaEk+TMw4+sovRyqlvqU7T4Rf40If97FJJleJyJvPHS5
6YfXIy+eAN9EVL28w9PSI2SeuOTRfFeD/NGPf4mIhAUIcuoTytQLzwfPAw6j6Sw/IRN1Q60HeNY+
QJC5CRZjXyVefNBJcs7HvIo/7HrCws+6hjnQkZicMegH34rsjJxzLN030iw8fzzds3DXz+xFM59Z
HR/ervFuSD2cRJgqeS3MnmnWN9F9zIQuRtnvArO9Bwvf4o7iC3SbBa+t5bgV/4vGwnRAZTpWSfT7
sfriD4P8U1nVtE7OpKZ8MwKHA5rOdCEljbRmb9fY6XPuafGUYLCEGbDaalmCvoGt2tYcUjk6dJRm
542ebCQ7CHH8+VG8rYvxo7fU10lRZB6XlpjujBEb/+BuXF2PQnF4iTKHcZ/ZLeGcbazs2TwMJGkB
GQGGjpJN84izoPkAnIg9wFI77Dp8koaTl771e9AdoU3n7RiANqs4DL0TK6zmCIqtFRRMOFLC/t3f
LKedqXSc0TPkpbGEJ1G/juMHBhsARPp44brTZdIQAk83lU+iG2yePu+akyeny/igd2kGLpO/SOiR
/WqcWi+HHRdUkg2xAsq44i8qu/ud3o12Q3RPM4Ew7Fs2uIPJVuvYihxZHhYaWhpxf01GRNTSXiwp
azz9s+Wk+1OBY1klz1ZRR7m+9RU9odf1bc26EdAjohukdRR9g67JGu9bHNjMGlVgR5JKWwF/+86y
AmDqfgaq4TeYDFpERxzCys7ySuwByTOoWvHuHdfCJeXvhZhfkGEDWmZf3/lxFlGZ/Lf/RPCXLZVL
OT/M4gEw0iIrv47cIyERMKX0UUj/q/Y48X9HlMHwR4Yrr7ek9Ng8z8P6GbJSstVOYG1FEyTb5ueE
zm465Jz8PDTMahNvW6TeB9nXqJXwv7nWHYEn0rgNUZTXhUWLEIyNQ0p2JGJn9eJlJKPSAFWzc8Ds
8LYUNKU09st4v7NbUdaet2fIJuar9lQ23dzWf43aqb9ZGs8hQ1o5NoGlaSSGLriy1PlhVY9vltSI
qwGfbbm4NgVKVjHRdxm3du6wPKEaIjYi2QSpacWsgoShI4XqfXh9bN0sN7Msn3OiAAoh5ytNZsbq
UhQPP7Fq0pGgEYHunv0wveG62JPJL50MDKCyBW9SYOjA1rZpisttZwYxRdcjW9gCoA7xG0Y17+Ek
rpcPM56VPxqunV0vcj5zMQLfDkyhPWZD9tEYbE2SGhLn5bZSeiHfM071DY5q8mjDv5InvHLJ05ma
GPtvgHxeHyvMSfi60F3AqolBxReNnwvC7nTa5tD7UpgZ+4cJQn857GTWE7gK/5/JZHWFELdxXJ3k
bH31AyVMd8AoyC6X/KhkSXWDyQnkzynO/ZS+Pdtn3Dd/PdSeEoaDRQO6SL+6xPCuzK9A7bBe0tZN
qloDgwRiqaN23MfsRRq1/Vs4dSR4S6POTzFCkqCEh2w/8kjZRTm1D8hWKNZphmFaZOZrbRvkdgCn
BKB+5s+8qWfS5EAXHXZrKB1jkCso/JTK3tNtePhIGUXL9V6Rox3uvrZJoDI7TbiiU+JaRe1+IHnU
3affy0HNzHT64mM6lYQigqKZah4qSwUlbTUeBm36Jac1j0fI5dE7li67DMHLcV9x0t0uoE5M0x87
No9zk/4Zee8ss8pJ4K8uH2k9RC/WQ5CsSZC58W+gzCoSz9rA3h5IKUcZetTg5mCh1iGMwhZRA10S
I9I2wKMj9GWkzItlO2hh6wt0Y+/UGMPNJ/85vojUz9/tmzk91D5lRMY6wjLu0cSukDvBDR9sq57h
46tMP/q85g/f3ELybJGA0vFCqIIH7ZY3aW8wV529B1OX9RDM4xZl0UERuipq/jBx6duY3BnvpdSU
rJqEw9IutCwrjLz7QoLKDgMza46IQM/l/pcouZqNUIwtIDbmvdiv+zUSV6vFuworvwfgIpPoEBz8
arJRUuwmNHAI7/LhMncQCJZ6TzTwWzn9VcZWjG/r7BViuBu9SbaaKzRG+QWLEDCcdDWvbe582E+P
lcAGD0I1PbeiRV7GZeVREGfZedNT1JDkAc3MH/D7lFPY0gBEMWTa9UaxJ2zsLgz2/HVpbL70ZS4h
UzEqVKSfjDWIrxCcRyhSiW0WdlsRSxKKuh0sCxViAN4EfAP16Mxv91av+OmvcLiPTHa4R627/WfD
12b87HllmUrvG6FlWNNMKDgRVWQ6K0g2QGN/tXsc0Mg2GopW/jWRFFOnMGdGbzrczuwPDOAJ+JwX
g9EamfXZuLKma0Waob6fovbfgkv0tKpIvYfhCDz9AUgYXzwQVQFRq8k93OlD9T7U4p/vCgM5bl9M
A05YFniVDYJucNKmVBVwnGYHeAR1t5uOAPSJSQqL1KFdJN9IXqJgHfS1MjbCDJppnGY9punKxHQL
5Q0gfzWswX3ADxUYMMnAjhHrWu6PMDQsV7X9kuDfTbbbWB9pue2eqrzIg4qXdrzx2AomWO9RQ7RT
kyR0/qizB7rT0WwUUdPeKRbwruG3MzuUqgDSnosFDbhVRuoAbtCn5SaKjLlbwgir1HPpzaXu0A99
pCUwUWVz1lDTCq22lTLuYY4aaEDQChypRy/eYRWAAGr0bV5fX4zR+dPLdCecKC/cZU3/QZjNCN38
JCwpyAnDKndgRmksxCW/Nx+dr/nmEbpBkjR1MxkzQvMm0ywak/0dtau4rEaREbPi//D82WUw1xuP
ULm8WNaWXz7YtesNoU5pHlLpfWZfXM3QtyH92S/fwUv2H/R3gGFjD65SZHYspKHx3OFuA5lQtPVm
Wdz3TG6xfkxg9C/qwsJDm1El+wUShB0sEPYuHNnO8MGjSE5ZoECcqQarHKK0bBm1hXxDs6s8lJ94
YFL52IrLReHD6TIoYowKu4IRrEo3As28L3sg6jZsswHVoEjGhDm9Au2FVaw9lAiKoiI2xKHcp92H
QPxb9Ixy/A6vB+Wfc9Y/4vlcW+dsHarijLPR1qg0vdEXYcjQcdFFO13sncwExlpzIIXxAOEo9FMA
jrstUCUsarfsBuv0jL2+NSDyzlZEIPEi/l5R8HBN5rW8lhDzP6JW9b//Ep0rH3d67yldEw1lGRaR
6JAOmVmfG45sDoRHi5g2THjGkYjS3GaOWiUinH+d3VXT4PmUFdAaiz6fZvjG5616t31lHmLBDgZL
5PYo8Vkaxqo7gSKw7l880AS2dApYQxC2GUIpwuXktINKtBoutDkkj6BmkYwb1WTz/8RQDFnPQVk9
B4RZYdwKtx0vNjd5L8h7/2Xca81wnw9DfbH/+gPVQeRm6LSc7nXWu8rHwaA8eelgWkdWV5d+/URn
nJkJJxL9Z+1Uf8yxInmj+C6Z5WTTfewj4Lr6crmcbZGMeYEJUW1nm32OLVLeK2vnf4PMMEo0NdBV
iJ1rbwwaowlYZ2fRTjr+ma1441Zev4tO2emSJnV/Sc60iwOdoYjIsQhqNz72t4GDz3ynldnZm/45
RrzrA9VVwkJNHZ0lvy1odNUBqUh1sd+e33QnFprR5WKqIxF1u38134AROrxBElV6rSfWfgGgHqUp
PnPE2L1zO9XePVSynd9iXreoSVDWYddEtSZqkPlUEMt1lbuPcj/UC/wnRx3nu+IWvCMsYOsarw30
K4DeGXjOjcaiz1reu/g/uSS7bbac6M1+WizL637ZNKzsUcew6zFjI5cNZwQftqrGIH0xYaS33v9m
w3kxH3KRLTCzy+7gh09UyzeCRxskIklgxcJYTWu+FHc50v2f+QGpB4ouFoPorY/GR2yV0D9HM1Uk
8LrgGmc4Mf4u//vdzx7oN+lPR+moaxjGRynGy0tLeDmRXBHpZu3+Art3gcBYEgK16Cujjpm8Vwmi
JH/HDpWhbCtNwSP31BOYlEYeMbWvE+nSE1yja6GUbtZr/FNlXX3Fn6PMzMs8PYgQoKGoi7iGxA6T
U9qr+yI8V0JmHuudEwEDBpl14xPudwLmDY4ESXzjsy/HwoIW0wlk76FHMOAN392lygNza2pFkDJO
U4KnkQJWWX+tVWCZZ8Yspx/vXFentEth07S43V7BYnNL7nCQrESyx62dPX0NdbROGGi8pk/qWOWY
ILcDJQH2+KlA9YkvLhfagWaspiiAsi4b/rgj6+Yk9KpfwoLfXTaKDbJpDYyMYoyxZDt8VHrn/nnE
ngvJdhw/ZPBzhwCLfVEti1/p4y9d7nxzItypOgzZpfVxtVRXoKbHZH6Esb3qW17vFJAnlswZHRn2
x+MUwMkiPv4HN+aki+A0ZW0Zk0frhX/Ero45I/33oNioXga4++yWydwlurFDCWc1+hOy1qd18+pg
lTknVtE1cmZ4/xWpjGQ8pHfOZhHil7bRJeJ/e1P4S9nlGC8kE+QkFn2Dw+r0wSg2B7u/mjK1T13b
js96W3PBUTYbii1mbvnc0VRIX7r+OTK44kTCvUctfnBqZjSySU6LLYiJVCkf4nU0xpUq7hLdHHAr
IPJOgibmA/L8rCJdKv3G9Uq9XXLzNXm9rYAl875VYEhRfp8RB2tycP42kIEgpMSYdkIq3LYUBdco
n7oakaJy7DdeutXr9uceUlJb9SIQnmaJ2rMuJJ7L/Qgr+yRSbAFGzj8hG1p+ECV7M2N5DgeTAV7J
BfYXwOVX6fzIOliq7eEbRXSdDQ3JbPBBY+YxhUxg3vb/2vOn1ZLtlpXVdMuGLr3zb40ZFBp1LimW
8fUHUGJsacc06gw8D1aPoI03eibC7xeGhPW+fv2yzKEw05FmYBWiHt9567RPnZnt+mWV/XeGx78U
NvOVKR6vGsW7VNze0NLJvMPmD8wjvd1YAZcYWjJQT/hZyS38zcAAiwyqBeO4+IY84ILYEHf5rkI3
EH21tqDyXDROktOv9Cf0kcWw4sxY1wLfBtDqCQIw2EOn4B+aM1pFrrZVJVmG3b0Dqt8WNv6R7TJN
pm/aTijxYgdknUBB+cPU7Fo1HUuAafnAygyR5UsjSwMsz2gZuW7GksjQUYTdP3N8IU5IbkHfoKM4
KxlLZA0A5NSuqVLkhi0OR8gZp8q+5D5D1QM4abcHEAWnoLcsKsBfjS+dSHPQ1G5OfNdgvIb2fDvM
6018j2UVJnKLOZMcUAS/w/rwri0c/VZSoSK3Q8o/kWAyWMvwsJNuFlDwNSOgi9Wwc2EdEFtLnAgj
Eu7ZxLVxZY6fQsJsg2WgGn482tA8YiNhzQqdD2NBbm0IXLGge7CdbmmC16MUj4QofE1SHO8MWSiM
TptVguUK2HV3ssScmRMe5qa+ez3Avygkj8bI5RXkP+KoESlwSwlkEl4cOmf7+S3Kk4QbQEi/SbkT
DteUd3abqB3fBY+v6vW8we2/HzkHmBJheaKqUmVzZMOm7CUN39/wgaLj7eAqZqSjCTV5hGi4I5S4
5xAJXKB5iAOeuIHkBxcBt3mv6KGm+EFlTCI9SuGoJj5vikT7r3lmFxwFP9x6fTH10pzpgV2reocC
ytAyjyTSqXzEyv6WC0zo5m2fH0vuunyy+uvelTr00ftVz3mUlCH82G+Z+NnK+t4zLYNLN7USO2wf
wYcXHBto9kJwHToyORT/xNl8k8L7bhRDqEf3rgzwgjJHX1rJL6gqDkLyAwhPH6vFDb6q2+QGph7I
GFk2I2KdUhQlfc4H59GEhQp/HNEwkNOb1aEMx/RKgHfswdfYIvWPMfGXrtv/aAQNMtOSjE43bLKk
S7bEWaMSuyU4qLI7QYpGCHfH5D2sr2plBDGZIgG3RZkgZY6opkbLpN0Vj9N9z9EQ8OpQIGem4c+x
7mFuMpnaIveq/MuhGy+wFLzRi9qHXCuWQtpt+FLRz1ahnV1b8Q88AhCJ4dPxeD+eEqr420b13VoW
Mn9NOmD5uh96yvOBPgZpiOm6KxivWqdqL/GIhAUQbkkuSwcMfcH3sd+IpmYWoCivuMRC6FHiYKpl
aRZxnDUsgEAau8hYmEGMqI7YXMWE61DnnYBsX7XSa0Remt3mF6Rh9m4gcKWy7rfo9dPSYfSYuamj
0lTccycbaRosox0imfs1A70MrT8N9ggKZaAezmHCxuqPOWZwHGvHd0T4vHVGYLHfqCI0NP9ekPUc
8JXp4M8wmjvNhtYaFRKyE4Sdb9/eQ6/vIwtJ9RY56nMDQ35aFxQ7Z1O8QFBCQ41IRzzyuCWuzhrK
LJrlLPM/XcKLAQprDqXQ+qqQYSgj8wztdKCEmRgg6N5UF2CCMfleOPYyURHDveXBELOoe72ZRJp7
sXGBqcLiI6QFKPj6gSxDF1LRPXABi1PRBDrBRtr4kwt0urN91Y76gCs2kDSn5gHHxsgvze65Xsfy
WLhpI8CvA+a6BkpJcp01pRAZs41tuSsqmoA5eH5iFj0Y6NndQ3e2VNC0eqhdumBIahdk2u+ecDj2
uMgyEgYUen94rqHQP6vMHx4uRScisj/IwU90U8Op1MEVGJET8r+v69EjF/9Xb4BWJHOuZSo5B+in
Ew5LZY41o6SuofgGa1r7xwUZKgn4c3wKD7V+IHltX1K0VNnwNJJyW0gUjmtgTcxrxRc1ZSstV55B
cYj/m3y7F1TAruKwJMeQtBP9YAPDA9ldRFEX9qyDZj1c6Fjc9oV9TrPkgMCuP9UJFWprJW5dAFY3
PNfENcXVFZm7zvE4VVkaKYoGaNf9FBRi+vQ8lww62Vjfnf4MbeGl49Q72k1iVyiJxJPAFrpFPklV
ioNQpoNHPQCS43nFEDb5djInsoFZb+PyNfTkxdEDuZfCziDhqH64Muqr7WwN8noSK4yE/boQ64Kn
N3pD5hHoLhg1HFy0OxpEPjrI2qJ8KM/wmTGGY26xQ+MEmBnhySUuL52dYQFHoeb287xuH+sagajw
Asg5OXXlDdFn5+dWnYEi/G5wjcFazHTAB3wPX1O0wAzqEO9P92faszyREs/OVOxUqbAbA/grHkeN
7IbK02Iyo3iPKtwMXKjMUj3o5lSn8kZ/uqQJndsWNfxV5s34lAcG0JPQTjir1lciBknvMWCI7cw7
n9Nby0RqFaRsEhDf2qmgOLKmxbtj1TbB5lySBuLOzo6bOJCfSzKXAzk//n6yY4XKPmUrhXJA2yh+
kWBNnlYgM7qg5MlXFMUQCAmveJ3B3Diccohx8JiEqizF3TN2qAsr62y/vzP9mUKx1D9D1xeMxTch
kt9RET+Ya1q94C26FnBZ4dlymYvk3AaftaXZW01f9JBqV44KhqCLa7eZ0LzYf4CzxxUmDnPkqcTQ
YZ7J+IqtCxZrGDY1ieoTjeTJcVVHO2+6DoONcUxRuNylk2yhENafgbCJxyyE8xaDKhmBi02Jgz83
VxgWyU2T+ZJWiK9ou2RI4VF6wIIluApNuC4UESnOYXphrQybCs1Q5sftfg/Jg1FechFf3Duw5BjX
crK619l5ScEzLsY8Oz468sLM6RV2WBIHoRGdi5y7hDrlvhyhSq2RV1SjMxmQt2G35M2NPPfoMeT2
aifbhtAlmMmdiYrV82204DeMLhl5mw2S5Vj9HGkb+qDsVL0cElApxordBIM+smy5s4FwHD7422IL
AjfpNgJ1fKe68ye9wbenQFQUhfbliD0XBc+0yNLZiysae83pFG0LgF1B/Oga7OcDAt+wj7O40wmY
of7z6gfdk7lkoFJh6GSqsrqvFxc6Qw2auikebO2AByRvCsGOrzIdMETFDlkAAXVgHxf+waCUaiz8
6cBEH3R5MR87nfZhyYgOJgWRTIpn+bbO1b8uUObc9ZATe0XB9YdTao0QknL6EHkTpmYz6NCoqpc4
IBC+gZ1qkBfJ0edjE9EFyCEL9Hh/ib2V+5Ex5anfd3FZaG2Ee4ZFS0inHp70XwjwBJ7zcwUW2rQ8
slVqtKUUOOjyMTgjP2+OrDfSVoWsq4X/OpA5oWuhLZxC25nQ5Kza1Cer/kP3yrXdL0awdauXPX5k
OYUP0FjrqAhMhRl/IQu0muttWIEBbpZ3DnXpGVhQzGJ1uPlXMh97qDuW81OgZS5cU1GKmBJPMfk2
YkYPHnoDn89E1EXTupQdf1yt7PzVciLkgpijm0uKBWQntx+uSop9CTBs4sonCv9WoWBX3dy9bDSE
d7hceYyJNkU3ttBr0mFT4Bu+uYfk1zQ+S6G31/lYJ6PA4UdwgVy4vT6qitvBm6oDY9vUd3RjJxda
cG1Nnbpv2d4h2LzJC24NVoegUy0vr5TqiUO/J8jPYBR4LbBe+Ji4rwzU+KcHsDFxlcwtgN9jnRX+
QpkfKJWYn0WYGi0eJpA3G/zhg7EcOIXO5hwH+RmVoFxZvTX2T3J6rIET/W4uqTn7b9UyPx7NtBQb
/ItkSTSMxcaPmjSVQ0BkBlMRKuzOez9bwm2ZG1o2YmiH5tIl4GKc765UWFF+kBZwLqSap5htSK7x
92YGIY4MhKOvVNxGOAJiKx1cXDnlt4FTqIN79OveAPF4+yFSsWd2UbQGwoQyaydrswpp9EaKiMI1
VrYOVyPJvgb5NQKVZ8Ll1LoJlJlYN8kdduNkkN5c0+D0//QYqKF0gQndfQZUHL56sJt6girx6GnS
PFa97U0UBI3rYkm25R+Ksa1cVh/mMfa57ai5m1lVR8E7w41DEyfziU4maf78760pziJRNm8PUlr3
G6JfKLfcvx/yNX5jvcgY3lJRx5vytQHsenAoZa8jxuBo20w6CXnCG61vt0HUhz1YxWB6mWRBZiBp
XiXm4yWg+uyGuo4dUhZ9eGhCiOZdxuoW4GSox48CKwYkNBRaFXvvz8MFDJqr4rMnkaa/ojjKU5AU
wJNvWB30HNUItV0akZK6iTfOu1twTFhii3Pa+/VEHmgNVHzHjeNDUHkCArbbMacXuyWv5gGDYHo9
BJGq13NfgGSkglaVamUs0T5Y6X4wlBEmoCOJF/OPbj6NAPioh+CvvX+1Drq5ogCVaVGQ0dB/aUmC
0jwT2DehBQtwk6bdH46uMTEl3VVfsGiMa8JrJs8YMJH/ArD6tfPlpLTcj6rKkJtwBqLcEV3jFNPV
OEg6n1pqsSVkHoOZPWAkTwV3x2sT7v7eP+NKgWxpcgVeH2z/RIpGyocsRO5NFUBA62EghxKQ1JVW
+gJ687DHjt5QhheqqO6Hl+3CgKitaroovTL4qJxBtPC8j1zyFqj8Oy/J7iCMP/WsuhOjoTDXM6mx
4JQvpZCY5sYiFrxyCBGHgCI17rhz8ahtWzCvBcE1KJAQLqQm8tu8IsfnCgvyv9uqb/I7BDhuknDb
ByQHXHOPkhOcnTJQ3+igeX4o7gkqVAsB7/hKn6oCucbIuA6l5KznOmeYyALiZniW2scd+9OmI0Eq
drMObqaugN0UWdsYny9gevCubDtp4Raf+psDWojaLIi5xSKtY7bT5CKuCD/ftxY64EfZf1T2e/d5
DtiNZADaekgEii+IH5VeS39Aiqu8kYfEHxYfuCxGeRod8KPXM5ScHStTMhHmmGgo5+FVf79hOp5l
0lUqGnfXpKW4iHSqD3Rfxc6mLHSaLp+wE0+gk7AFPggmcwxNkuSfbcOTS04GOOaRmZoi8Je5Mmlk
SneNbRqdCYkCS8mG0P8pFMt2Yh6Ayvp0GkQ5r1uP/r41KB84w7rCZEgEtl/wJ65CdBocGquYdUw6
8c9gSZlt6BIy81xAmyfdxWMHwYiLOrDXQ+sz7n3GrmQNcdSWeli7cRIbmlKZp7wxVo3z9M7GeWJe
5ASqY9S5WwfS1RU8qRJd8NxdAsrlVaj7IJ6jqBEV/ZrwkcRH/sN2bbpdxEDlBt5+qKymeOslx4iq
o3YGF6ocWU++HvV+AWBsVpEwLctPdy4A3E8KrkbkFR8IcaYjEsSWZMSFuyFbo13aYdC7rF4jgqi8
yBUkaODbRh6nW66bMqhLQGIS825uXAlZntYFJIZ/eQBQJwNBW64zZnkrFCnHCMMNWcdoK98YMkFQ
A2MGbNeHoQtJxMuBOUIhcKh3x/mB/iPReRMj437/gJssCNSvsAlRuD+PLNPhT4f/9v0dFgtlIYcW
UcSbapdPeN1LCfjUOzhq4wwqoaW+i0nBG1EpxH7ufZpLsQZK8/Bj26r5w4cSAXC0v4s+ChtyUDF2
pcPlUYVMJUyxUR7UBnpgp4J4v6MpoAUZr0bXtV1Vcnap3gT5qCRCRrJRc0h6NHcQWaV3p6PTwNgH
WpSREWC0r086M1iqRcDG4tonwsbWq6CIcpJdTSnhMIOFhIuK0zbRHwvn+PuniE82LlhnsuCrNHrA
nWi1swf33LZwUMs9epTs3z2NMcNKRMUA/P2r3hkjuNHfJ00RDpstyHvdIQfZAPlCKrpz7uljaMJo
1x6B2vR+gyunmNGe6hbac5BwZw4w0dxwVBzpswabPOm3JaJQlR4k+aOAamMaOF7wwIU44tMOg6+C
TT1QIXUE42h+mH3OjYuswBHxI3g+GHGnPLCd/rcTkDn3lBhbIL9TKxXNjfVRCrOuB7f/H4tm6WsU
z+lvjNZtp8mW67S3IZA5dwigQyaKhwcofs4cy6dkCb+vUjhl11pyphVhHqfB6eic/d2l12Pqt9mE
PlQ17+xZpsDmDMQn6Y8GOtrWKAE2EztkWJj7gRYeQZL63NsLLCoGtFtonAxjAr042smaDOtHQUS6
bLtl6PljaZmY9358qVgdpryg6bo1s7NWWVcX+RezkFE8BQZ2BZ7anYIBYDlZ3jR9fI2c37l59HIw
pJghND1dHj+Tvk1azMDyZw9PBXzzdLqp7MssXcwzXLaJUlZ0zL6plV82jAHWEp5mgRZMoSl+rAbr
XBejy9RvXL7ZNySSmpcza1oCQt1FbbvWhXwtuQFBxzpooA62q0UvN6JqUz7KJWXcZ0bloNWiR+/w
phtOYq7XdOZv0/bYTVFv8OEWoo5MZjFbDx1YISblr05wyXyghxHaJTrZHjDGjlQbVlDqswLbj2Sn
j9xuLKMJNP6qkWVDItGBmWDHZQDFLB/yisfDwgojt3YyKHjUu0rty9wbajVy5NHDx7VulEQxQK0S
KW/RXOOu177nskGeJiZn40vMbTIknFWDsf44+Ngc5/7Bjr5dYKGq+cb1hI5Gj2v9/6kcANq0yl+z
8E1FNbIqArdMC1YxnaHtTSh0XwQTst6qTQL91bpwhRoOPKRBJRc3cZFCaqe5jfMhdsF8VU6hyIp7
Obvb6pz8dqnCVWLXU6E2o81e0StJX08LCUlmbJHYktHBcfDXzwg7B+x3ipfc3wteVVyMH57E4tmh
Tlsmb11ileNxn+BLPEThPKDd1+qS3ye/qn5N9Dn/uH8zR0IWOWeBIedZGdiSToGKTVkRW5NGl4me
Puis8L3gEvtx9L0YVE90bGLychV2QC3RbRpSL0mimAaMNS6RNQsWd5P1JMWMwCl412Nyq5ttnBHd
j8drLA0krpTDoOQHeo+25OTAVgAmNVnJSeknUs2m1dljbCf6Ln4zu+yrVicmeFPJ7aJ2o7jfhcE2
+HIIm6VM7jJMUK64kyWWoQW5TD10MvEUvH1obSbuAk66UlZHte+CMsNjUWTxahX/aNjX7211ZqZ1
s4lz2ReZ2S1oz4IFgfIZoITdUe/u5Z5sbUvvtRKRWw9HFUt1IZLntq3dGlX/EYogri4RlVamvf5x
mt5GjLefkOM3Sye3yed3PCOyNNYyzjWikUMpx1S95w2v2zgOziN1ebgizvrMrqutvUPZvRyWs206
N+UYZEoz+GpVp3wtycd2avUgxNZrqaitK1Up6M3VTCrDbeuXy/VEpIroVoWp0AePlm+1ark+5i7L
cLYgzalsmOirzhh9yrCtAVlBPvCxL9J9EksauaNtAS/uANWB/FkyT03rX0FXPovyRaIoccaUZObO
j+7aIOaM12Zm9f+VTvxgMoqzmOGn9lET6oxfHlIu1HC3zjK7chjZYdEOYrHXRBzUGMNDDBJIp23s
maXEqAKSN3KC5IG8J42Tymp1rOlCCA5+P3HbTFZBFu74CWpQH/BJiejW/hEUxX17Hsh/LS5bDFzV
eEN/LkkI9U+uAFBw95O9YmktXmSML2UZyVvVnMGizTb4ydaZTUX/7ggwZMldcXI3NPEJZVkvkhdz
7MUKb+kLSaTuM0roNyuDq/BuKJlPjy4pSfMbsRnce6M5ZvBVb+DXoohSU0WBgSKEyy2e4YKiTnS9
kCAvr7IjGAEALK0i8CnZAw9flAPSkus47lLtW/UdxW12D0PMdNWrRLedwIxqBOslKOl9gSprcCeb
BUWEQfSk3HNsvGTUKY9CZKpg/wiAyr6pWXu9bREBtNx+i6nHeiscyB3ZhPke3Dq049dOS/G5QYrW
Jm19tctLD51HvmcBO29wJesKqG3RWNw1ZL3kDga72Iz/ua8E3rh6FO5+iQjjg42BHW44II4hin7L
0nPVNmB68JeEHoebHhTl3eAgt70skP9/GGkAai3m9u8DwxjAF9wmtGA3iKuwD03rNtmkHKCj8TfK
yKlYT1jHCvHO5mlfmp1pwhyTBoZG/LlRxDh934W95GKX+YhQaYqCky2tnb7NG6bFiJa+mn4l6fdQ
/KiECSY9hog3CSPQ4CFg060BS9soSyNAv85R/GYp2RajhQ0LQC2X65iowvQtbZgGIawjvvzbT2tL
Jyn+e1yIrpJLeyIUn3MZFMiPWMzGgVo6GlNR1ED7Vbk5rewwBxuXzQzpGdY2hUz7pKBGq4+8g/e8
8U/HEioclKeOiEXzpoO6dXBK3b9TE/FfqxhfUHtK+A6ij47GPxrTqC8CUx0wWnmLLiDExyjzXd3z
+Xp1IpyR+lbqn0+qfFxXMIQZWINN0bE+aH+l0QQelUkDepxNYobH37reRdDv9op5oGfnB4rseCgD
k0zSppqYsJ0No75kG2aF+bMHsRYjdwH9+6UzIm3NY+5KGxZaOZ+IXehsMSMuK2Pz9pDVMayqUVr0
eF7l05Aq63LHzGRuM3uMyfavzpYI1HQM5ub+oZwJTedBvWBg3+rw072kky9GQObTjCwLmasKfNHi
g6dHOtXtTzNtyD1eaC+e6oegSGFdjl/Qeuf9rj5QcOX1W03FFC9y9rUzlTcDcJLKS2ZqEW42HH17
Ck2MOvXUR/fd+IUwa+wJ3CtIfEFazFmhduxpAPUhPMWEEA8OSDPV/njrBI/8gN+Z+IRIZybOWVon
p0GxoyCuTjzFR2AesbsK4xu0V62B5ipeGvEFQV4msRB7tTvXCPykl5/UAbu5TK5EK51tvFmAYH2K
UeICazOFAHGoUHxYuVlrsebAE5PzzUChbpLcQeDi56MhrW3tBatOQJRGFdKepdTH+B/9QxXH/Xo6
D9h2qYxzUKVfYapC1Hv5XxPgN2m5eTn6wKzaqSCGmJk/jC6bGmn0DJScCMIamqUOqTMv2ISm0q0I
U8iGnBwZfj+60JHOYsOC4vb3eLbNvSkn1SxeniVqNDwVHTFWu2eKUxB0IytJOlZkCOJkvmnvAlyd
pG2jb/KraS1EvKbkGLQvulCiKR4SdhE0ezWpB8r4Y7XappN6ONPIlK+G6EYVNdtCZvayhIce1sU1
CeFtmtoE/Md3wb9jUb1UwTgbpSnO3bHKxIt14iFDo48+Vh0/w4LKN2mMF5b/scEJMwSmve8RaabQ
zz5c7nyTmcGMSmAzjpNYoog34iV5C6RCIFTG4WKJDXX+uyyeVa/9iyyGL9xATX8YZ8+kAwIpoux2
RGcqsuQXSS/8FHre8T6dPJ6WJZhUwxwYSJWLR0r+IK8DEpzu7+EytSWiCLL3fdiUZFbLNK1U7kdE
upZq04eonXwo8kmCXzKAbTBgy4kWvPIs5nyHY5iqHIjdov0J4H+0G5xF90O3o0a59wTAtq0WTFK6
jL7SWBU8sBl5QWE9Lg4RckrnkQuZHOKLa6huVVVy0FEvUN/JfQvhN6oxt5VrZ42SZWe1tPlBtaKV
BCkLE6F4S33a/YM3meo/s/VheT0uIJMoF7P1pqI7NwvYbPnLFYeHYURZmWLP9JOiN6ruXDVeVUTR
LLknIo69WrbGVT++UT85dbaSBFZxv6T+V4B5gVbfwX7T/0AD/RjvxzFbndvbs1YSsmWho4fpA4bu
DwXx75xFHnfuItsdWIZK2t5ccpRrlTSmFDJ0XWaLQuoyDp2Tz/7ZzNapSt4TlaANQ7eZyenfBWSl
CJfB6IBOv4DW19FRqZk3wxAkYGcHm/OLBlyWV07hn7ZFFUQemfeM5BKGPhwXSwrq1w7ereaBZX/P
vCyfnqGJhZL0fDkLtT+o24OyxGW670VL7FgQA3lbVGthUOqxyLlAjYUirlY9CUUOkEA7XlFlfSnQ
JmuZYSQaPg6yTPOiS8WvRTKtAf9BvkzSN/uWfvTHPZDyLxo5k6tDOXxofU40geE4kIlQaQ9dHnOZ
xrANHJLw4GpRo9QXJQuJei3vOkppOYNixLJ5PrMk6yCSBraC+W6Xrom5QrQJSvZ7875YtsrxiRDU
BTzUW9ZGn+4JxBOgFed2oGK2EIfvDXwMTtpu7R0EmMchwaSb/cKm7x2V2GL1QYgqEEtj78gkE/Mo
rWor0XbFyhYuFtLTTnp5Rl8hTGR5I1VZQGcJd1j/cgJj1bc/CNaFC3cz69Jt0oghwUUpdq1Qe7vi
uYmYoqLQv95gh9oJaC4FH4tqXfgvUEavDRtrAcdlmVCkmDf4vXbLH+WqPz49IwVcZ+DWTWBvHt6P
BhTGZ/YUE9txqXlp+rkV3uc8UHrceSxyCrPVpTXCCeizGTAikEdaGVilEcWt9LK/I7XT++ZV0sVK
dLMMTMw0PN3FsiCTttNcNi9SKcOE7rrwDAvr7vELGXjlzwWbr8ws0EUDBgE4p8d+FiTj8kZxw78V
erADvRc3gIaxkrrtL88CbYOUbMPChhKNsTJ3Zg6spTYCBe46Sl4Hy/sN1mbbdE3s7MNILVxsZqqr
iKsyjrbQDfUXvmxWhqFDkVmZeSVtHssRxhJ2gM7Pn5MM4ngTQf/3rJXt0o2XYISmNPQsPVeeSR0P
RwcMoetIlEWFZPvZQpigbPpQ3bI6JdaW0mzQRnNze4WnnDs7kxOFJbPXdZmIYbo8IhNc0bIPo1Zc
8/HgM+NUu5p1Gge7nKHAc7wPfB+szUAyDxVcAh8QplTr4MSU94okjt+F60KPaUwPKSpn9ELVanns
24yUBt93oxIVt8EC1kmx2XeA7XVh4P36ZxNSZGrEbhjD4PS87D7f0Kf8QS76QCh5KIY78+mItEUA
TZ4aBTscVUBQOZuH+InCAQnlm/P1Eplmv+rRo4/AAWbd2a3Sc2s6emOX1sDHITXwZNYuvg/yk7Ih
CubPEhp2hrT0ZVtcW1Q37a4DqGzVQiE+4L7+eUPCPGFBpJEUnZSWr5GnqowhGUnscm79gwK5YlPl
jmH20cYuZk6GIrLD/JF9PQfE7luE1/2DM+GGRPFmFJ/kVkeheFA00QO6D6WXXhuBDBM1HxI40rgt
Jq/7sIezbKqc38Y+drVtpt8W9bOFJqnsU3fLokQxLhuO/iF/AaTfpSafSQdJ0gJ3w5Qf6xGTDPhF
2U9JfPJTDGrUwwesFJKsMjKApwEHIIZaw3JA+rGH5EocN7fJ27BT8865X9EaLqNzD3jyNy6Yzw4c
ai6sXIVODLoPTYff+sxrQJXAx3b178VHYHtWak3GVABH2TXrhiXAB3pp9YdP37O96Cv3jfyYDi/A
W9k4M7LdFvFJMYB2Ez6bpDbuWd1bzOJfJi5saRy5DqlXLH7ys9k667/Ah6WqRTcQfQpC/U3lapyi
bvgHnlViIcBvsO2DkdGwVJFQQlx2eCL1wJxq0vPArF8d9N/zrDzeNocXsAt751sBG16/ZCaLdf4d
jzRozvY9Jma9jwEu0UGqDo/hHKNsKAzsRYDWdhtskCXTy+AtvuGaO6jNwiZ9owRaTlkC1w7c4qkG
2Sy1scadFNWRrzeiwV0TnGqzicXo5rJO8wBR/Rdohj6ecoNixk00H0VhU903I1ZOXduiIqzyK/tY
vMr+m4fUvfCscDtrOgrcW7/9Wpe2iSaeVKqWdUh7muiVkd/kUGMJPh03sP2l8bdV5HGVoQE9AiFj
ijCquWUruyB3dYnDWZ6xy/HJnOq5XO9XTsKwepRuCG5ecqB+LCohSb2L+U3qZyggOlkfWLcABS5/
Wk74Snmqurw+iFfC94WtIpvJB/ANIEjL2lOF32oJRul798QUUly44lEwX+x7IBiFTRPpTtzVdNLb
2Y7qXn+OZ1N9iep0w5vyVGrkmlR71ZV4se+E5xiMh8S850BVqYOlFPg1rHSI1xkDQIyu8bcL7g9G
vznzcqkjseKzz+wGqzYyOOCiBU4q9vnmVda9NbD6CC+wKRzyMw6vUocYohtrqZyvMsRIbc/Z9Ev+
m8OeCZBxbolsQB+Vrt5mlozD3yJ5z+Qh6sY9CbKipK8iwOOy+72W2RjAGzk7NxuXa7YDZEL+etEl
5w+NvKcDsxWFHy4PitoLpe7BY9TvlYGLMMI9vv8NvMPqLz48Hl/4PPdUQG+unWQw4cFs1BBnuG3X
hDmKcH7MGyHVl3PX9RcwvDGz1NYJ1NzLeXrIuGrOzPOn7Sb8Bzmsi/MBXHHy8qesK6+yKucLTXiy
ejScp80g6wAp4rzHXMhSBaiHMvcEQCCp4uUFm4vQKVtciOic2SP8D3AqfXvPWCSJzwKYHUQv2OSL
pyZ0SdIKH7m1Mg8pnxtaJkJSHZkfCZMA48b4taDqmsownr+vpHfuBsZHvhgmuD3TItly2bBFb+Nq
l+3/ftpfVlb/Uy6ARcncZdlqr8do4d1iCx7aOM7ZIHnnlYM3ShgVqpJ/fsLa6yIDcZNhKjBDslyU
sM9Caj0HM6pjJQ71QfszHQHa7/vEz0QEEpXKJnlvUgLUneT0MX22iSKjYTjpc9jco6P0fJPi6MTv
Hx5X1NCYcsP+afWChHfnY7xkUfRmVAO+TbL1+x07CK8ZfyXIBAM4xhi1gSMywFXm4Sn6pK8pnFwD
ARm/Km+KStkaMoUn+X+ogW1kz0wTJPieOO6lN4xHqMpEmN1Y3CWwD0F9/vq+SvaCF3k7MRTV82ZL
VC2NewWckQdnvV9cPK/Pzkh7M+pJv3KgcWvdl8EhBuQjNrHFDcavf4PhDEKUHgHkItCeaM2ZaRJu
Bzq9vRfRLJXh22Hg+RD6eOdIW019ttVCcsn2LhE2OxdyuGaFsBzUwbUpP3k2OZtIAALgOFKrVN4n
upPsTmxs4RYfRlPrKqpI61GNjwAbUUaf+iSNCO9F9xlnaA5ANUl5b+J/InN0aECmF8CV8wB96gOK
Zw9AlY8X23ZZplTHe5gq6JR8oLSlM7Ob06hbQ/fDvuEdH47UgvnUJBMiMBzmqSyAZbc+8Cs7GBiE
hAK1eVr2C3eMMgyiZ7qTZlAX8RwcUvp33FzygXtHL51IKB8mjxknqeBlgcbJdxfHKvDs6IMtcxyu
+mf4p8fvOLxHsH9ZLfV7gOtq4slWircDkbm5jBsw3aDzDbgt7Ey0dzOdkA4fnAYPuJ5D9Mn4ZbLC
Um7AENoUK64t0Zi3pOXa4jzL7HtW+JB9fKEBZ3kFZVd2iJ2YdQFy1EinSNX6n9ZiMYl4oqzBjGwx
1VckRXasZ20tHz19wSrePVGQGYyEX7OBiymUZQlgNGHtXb5zRyayzLkW/LuoxnfvW/6eF1satyxd
yhBO42gyMHcYWAfJmflPrSGVlyijjhM+t44P9OHFOwxAZd+KXIHF/h2dLyzVEUjcrmr6Hnc/Xxdd
tPzSzKnpjg4kdyRTmcGSLWh4fmSmNriLExyABM7M+UZcEo/io/c7tBAyC7JMKQ1rlMq8/Dniyjml
Q4e16hyccsVpcgHKGnwjhYYI9TO8YkL6eP1oI3qTotGZZkWZmru+kMHDlv0p+VY7fDkxyzhrZ1P9
KV3uHwzI334JETYkDpi46EMDsm+dAdmchZdg15oCzHy98CMTluSEn9nbDFvDZXmvmBYQWrCHBYcc
rZ5v0zxTNiwvLtrVNpbOXlvMQWngR3XupzbsVV3CnJPGRzcjndsLRe9CgRG/mUnuN7UKJowFywf0
orQQ9EtenD8EUwe+onCpeWa1nVTtN0EKE8DsJb3UI4/xzXQK6njoQsADMa2kRFBcV43J0BVUV1HV
KDRHe8WWLmQLSayXdTE4HkS0g3buySm7kToF02eoUX299iA1UzMMQUpY+DEc0ghkOsPGTsOY5hfk
8vKeVKj5MolDkXwgVztPWqUg1qFFhAjKVwaFPJ925T3aTLYwJv0DrTJ1kIo7iYjAh2dn3pfrP3w8
traDGORFseWrVzTRe6tyzOx5cEOJtz+Dl5nyrPeTVWdbvnbGLGRGYAFC8sEeUam9jZ4TilbOnxgB
8D+J3zFP4Asi3sl/LydhuzYI4dMMOBzb9FgDYKK2W/P59clog1aYyC3C+M0eW2DUgIOX41tzXU68
c7FGinXc9FCIdtUez3VzzZeHve9WC5R4YchRHsZHg0RtYKpYy+Ck+D5loIkXR2nypHRaw8VyDF5k
epL6AtrlVm1PWdPhHsU6mTv+qohuzBh8m3cLxAHrlK4alEAZiTZIsUQqD7xpZyn8tJf+W0d1FVOK
5/GiA88aF/QyDDyyO5R2bTeM4nSrsgSukzlSSm+sVnWjC8C3mMvyNG+8gfvg3HZlaXilUsj4iXp8
Z8J9rY8NCpIShx5/Oee2MNqUnbuX4hpTUE3VRXAP9oDMffNmxBPtU59+myj8bf99lNVAtQ+0ppXW
qKcH/UJ/yxt0D5dtMXiR0//2UScH26BOh/BAWe9BBNUQ53LWCoQr8HzN/Ggmy49z8c+6S6Luv9nX
bREehr44ki3Ox6VF8KQTuEhhUqrgcmX5b5udp0gYyBYpjfIs07WfRu6nrflQZnYBod2JlDLfGkt5
3Ebz/VNqxbSMllUpboSaxXRsjp6vX0WACSRDh7SnV8b+bQrsJo2Atl0XfAEYePQ3zgOc0P3ft5tn
pKIDp3iZBRP7qUgBx/4EXnYagXGC0xIs7QcC0U9dEUIyqyVr7YWbvoSAJ2/iUyML1jk/PjCB9hhL
xwAdLB7Es6BOBLjsOF7jZHeI4OgPbbJXEvYIZvfdcKA0f2eR3tzM3s+oCfF5xd4z/Y8c/sZE5O0H
tIlQ2mv+IMPkLU7cJOTT/Gwo3Cgu7hZg6wRWy1p+xHwLZagJrSDKX5yaH1qaJ4Sh1vcoWxG2a9zE
cGNg5tehZBNEsVIhEucu46aNOdzaQ1ycjxb1+T3rih98x/qOiJM5HoRsfU46sGIXPHuxIKi+ZNbD
OCUvzyb/MRgmpXRoZ9HtRuE/E9fjQ1kyF1BEEx1opr/gRViy3Y1Y+fqVLYmkr2ZwI/WiumzwgVhP
1ruPQDPlN3AZJPmpVT2coN1IW/KUpVc3bJjCgxDfIWgjkhIif6SSdybCakuTZ1UZ0KC9GOaOjAWw
ROj0LAQPNkj7WaMAg1XE7A4U8pXoicyThZIrajNlJQlJLRBOOgHeB/mcm8IBrDnmxGHBwx7IZ76h
6W7CeAe77kwJOO/zqCOswSk4yhuni8RpfMF87fPvzusOcAP34e8wl7lt2UmjHVA1GS0mg0xbAYEs
eVzuaLvo0xk15TALem+ajx9YdebDGvl3Po/8V4appXpjfAQWW9g8wB/Tn5sIrJphze2OGoFqQDqP
VI1CzHIigJYpH7YkXNxoTOIlayRDG6SYfObqXIJhjAqkU9gOI30FvXXfeMBqX6S3LboCYMLPnZnD
3aAf31GxpDXIWRI0S638vVibhBZXXi0g/j3Mg7GiC2SOadk6FifYxyrpzXI4yp0HbjaqM+QdB8BL
lDsG8MUsQG91q2sf5vE8MXFjC9ot9I8UKlAibClhMMme1w0J21d+4FcO9jO9a9rB2KEyFhb5A/WV
nHCysOM258JbGvxW1BNLvy46oGa6F1gTr5xFj0Fa8jnnG+1UjrsrBJtSL6WXCfIAXZfjKviDpvYM
6mP7Nz0P1GBa5+PSlEAyZEmgpbvQ0DQPkTTOm8iTCsGdE2wgl22Glic0Nt8O67VwsFd9lQJ4fl1L
ijam/MHzUw9s+8lQWrVrNmgARTwILmG5AxVxHZeLaCSRoMYkK6w7+AlvxsgLrAxvyTflTZ26EvjE
LW6rvmx/6LGHI4hO9VYALbknyW5CS/aL3nmstRb/kixrgARwTvN/StP9vWf7SHu8op9rdkF7jbWY
bTlcAC+68d+aS52KdA7apM1j0avjvYTiB4WzTfP+cBK2Va4tcmoJ/whCqQmxOkB4jhBL3Z60184+
6lEeTz9on9py5dQT6SM++zbAe8tAWOiFNzMjX9TpbHcwKu7+MKp5Nn7wjCZxNjhIYHOsImVZQ640
Y9edoF8Sc7UE7d1ABTrU3xBmPDe1ZUsPujrN7q4YkeAR6TK2nkH0RaLp9DYOUUQS2AQLKaWlxk0Y
MRakZA2asVI213nWtFfa1N64n5lNHKg6UOROq/ENH6i9/aSRmFd9FlFNxM8TNR9sAdUtuBFRJR6T
N7G7SuNWR52sVgB5Z7vQadhcC4Siiju7gH9iQhpoFr3ElynTVGCGeRpqaqsLtCJVcToDBwaMA5FG
8tmYzTpyuhefan509HXqaQaFyWiIhLsVLxJ5UHj6dM5R+yYn12IAVQertszfckUkfc6doIBz3ogU
FXfcZX5iyjHgsy7BR5G67aAmHcGVq7Jb+UCCXXlcO8bKwlesfiIZBeP8lmX4T8mTChrHzzXHB1yZ
1sRG3/7Z1fgrRrEAl7ErLYQp/jYJIm1jNEVnawgw/nLfB9yic8O2V8A9EPCYptlSTCTla2q7y7Gi
cHm8EQHXj5J04qMOTdaeAVYJ2xgcgTXDKVs8CQIJlssXiUG1b8CyWKrIqIm+Wg20E0J2vP0e56Dw
Kza8ET4+hzkQkRhyk01diWvwCIxPosbMHelkUTDCxX7qxHSQcj3BVKqkvu1Azno3TWRkNR2Th/xp
p+FLsZms6E2BST8Cy3nTcUhod9rVtBCSn1X5HS3XYQKJUwrTWo3iPeZmNO0NAD+wWgBMK7aOFaJg
m5kk1Sjl9isd/FNHgV82XtrBQB1+aMflMLqc3LILNiqS5EGCbY6ngAkdBlSEck+JDsHZOc1HAlLW
b3Xu10No5QVp6Eu/keYrdDDyLeKQfvSmCXo5eRTfbm0wMAlCxpVLgSuwCRkK0imy9yFH2RTL++nP
OUgbmU4PU7/F09A67S17SKx5kFBjkKvfFtxOJYqDp5t3/+7O3MCJjnESFTJwrBwM13Rwr2xgNKgz
MPv4/7myYeycvTRc2lVdxzs2uFwEyUP5t62eWX3oiMJ58F4tj3csheiT519s7flPQhw+OPhLJ7Es
ozYw2SyzstkCEQQBqBnTQLoEbrkxQAkxV9oPpC2KhibJKBFPTKxhQqNkNcPlu+xBFkFuxARcPXhH
FR9NwE+sucPzJwSBPelFgqw4NI63sKyophHnxSPJHRt0m5z62tKJCYUi3hQMCAh4w9FKILvCcEQf
ZK98Sy+7IkE0HKNdGzq/x7mbvhAKtUOj1b9BGowKfQ44JJWBJztDLogs6XUSHFNhQ+3bXIqI6Nqd
iK1rmC4Yb7IspL4RvJBUPwomWlZGfCAvpvYQQR1sxFc5AxCl5y/sqBwkX7Jx1EjeOD4B6yB4yh4m
LgqNv/vPda4PaJw1LemSd83fnws99NQqSu/zJkWg7JdafRNAdar1h/JSLVS2d6xnYXJsAE1rW2i5
vPrEu/aDU308Jd74f9djgh3Txo/uyEpXLwxPtzhEcuLuEcm4D+hs/o3f86sCcS/MMKDkaI+hG3Zv
faWglFyYxqgLh+GbFa2eMU+HK4Bkq+p5OMTk518JG4Z0dwr8ztwoH46GAVB5MDyDTBkMlbY0NLW5
7WOzgW4fcEtjhX4rBjw3uKlZc4oZvSz1Jlymy+oMUzamD1KNhEZdiqjLmoq8u16ZiovWLMRwrlTB
/nJsOnBmTBkHk/4a/8EsRQm/yVyba4ZUT6KotmyXAw6Qn9vtZ/hA81ocvfWorXFM/Mp2Pd+CIISw
jhhvD2sw9oKpC/UoMyzYelc9U+dwzzOMmWfdfGU67Y7rjIo5LcZZDekG95vQ0wYxbkxOg0SmucQn
lEJ4NHAXJQxhfGqUf81J1bSj0Bgx+RpdKGlHYGEDDupJBgqBZiaL9nxjOQ5cGiFujwQjF8CPNShg
5sMvJVzhE6SYat2J8CkOegVg29+BMDD+tx044aS+u+rKvramrgo5jbBjkVKJBYXBVo85mcrDKAwQ
KieTZl8f611nShkdnpSe6VA3kLjyGFYQeXb1c/CpX9dQTwdsdXZbH7sdeC8OLG/nnoHD+EjHKi3h
jbCimvpdy9Zibh2j11X1sYg2KClGGneN3CkgBiXca+7550/HEXcTNys8RwProeIU7t+GRCfwPS7E
X0LbpX03DqJLdsD/4aGHDFV5f8ricXrb1bLClbfS6Dn9CCWHxmYd6L2GBfgfTxFCM7ONUvL5s934
+DDnyFE3G3263wa/Z+muZem/GS3EOyRs3HNr7MDhw9ylMLT2ztKK28VCnK3ErYRkFoRDW6zRdEjW
JqvCeuY7lhSNeYgxC0W7CGKVzdwE7MdwszCiCho0nU4Dv+eWEkz0WDOEtQDGMHCP6yZA8kTwq/Pc
L6IrASW7S85Ea/xYOt5oT+o+xnORTbsaEA3KVoi2TiPwy5DpqeMopivIotnMIevshh93J2W7QttW
x6LYatVOuTIAkEP+k/a9BVOZWMAhxCVbOA7RDBvhCOT/ZD+wS8xqRfJWDqeDuZoeB2+ZOhHBEUsA
bKB/nyI9JSzKhr3eDeOET58pneDiNWAn4kPglXM0arOm262xXQEAiUhEBFQSi31o6tKk1LJ/4UPN
VeAhiZrA5WoswxPn/vaqQ//aFJ/gPIDb4lKpTmnQInIsYueZ0LXba+M4wH3qVDc/hBxZ7oHzebTh
fq7S60NHtBJfnftVWAqITGTiaEWUGpj9BWy7T5If/phk6ekq8n/MR5Vb7tEto69G5BGf03jsDzRX
0KUUtsG96FMCbjTT1wzMnuS0WZxSxIFzeEK/xco1/fBbUKEIji2xr2ztWbx5UCOm2uSNYOUYWGi9
6s+0WQj0Sw2f7I2hz8my1iCRv4V9H0xZpoZdYVpvvj3DxSQJWesWF4WwiMhDXAEWI9bR19fjit1i
ZVTqZV1SScc6Y+i2Ia7aRK+5j2WRkpzfd79CUI/Z69jJo/eKQO5H1pE0Sal6Pf1+21eWIz/Glagp
FHUqoZiD5uHXQ1AqcbJWrNa5mN42ADJeOuUERwYhQGs1ELrjcr6fryDRuH1UmTKMjy49TQjx0A8x
CWrWlhu3+rJo4RlUQRWoN+Xz002cdreSeJE7lWsiVSl1yuO2NOqHEAExiiYKByyqGBxpeqEgiJT7
RCw2eM2ObT/UFKQAzEHVSH7jBJsWuaso8vUSn2DhVg81b1bltqp837fZzAsEoHO+UvBSR94mqtIk
+e9xws3xUP8fo824SvS7PloQwJFmEMTsx5ilSQnuMgBf770lYj4JrL5K2fpXpTvbWhWbevSNuqfK
lQN6I0tcW4UmA7RMvjO6bGwyDBBimV346V/NMGF76Qvra0Oe5ZYEglVmGeuZuBzVjcLozJSG80zX
FPEWOpI256jaBzo3wHbqDC3YCzWLrPkezo2vfUiymTPGsU77V0/bnSwakHffx+WSttiigUC8lg0l
4dnJ72oo/widjTZsqKq+NuYFXEtzJxbaPAiToan8DK16ALJCwTDK2joBZ08gaI/FxcZK5Rp769vz
8EaB7kngNVYprX3hys6rG70A2+SzRNlS3npOFssNmDicckkhh2hl6rF5iVtls9LupO8xjxiSKS/1
BGCI0OeHui8uXEI3aRtQvR4DBt3HnqVo/fGJIAqihfgEC3vFDFXR0UhoQzdP3ZmM5Q6zzbHY2zV3
X7PSaBBOpNbcvtEOTRe2tccbFtVJ7fPWdH5b0vi4Hli3vGNcKRUbp2XNrKc9C+OVGqM84S9E0bu9
smOwtY41jdtXWbnRwBD7jDFiOOB46jO3fpx4xPvEBD1okGFjNrc/epkadTUsK0YSE0k/tGWZUsYr
+lfaDI1McCiWQZvqvAkIOFQmKCJIVHA8br00DKJqW2j096CiRVa07Ux3MiegndHV/eJ9g5QJU7z3
264i2G5m0Wq/9sh5OzXiUARZfA+ihxZ0P2lJFsu/Bcu1uDrjiKxLUbjaZae6LIICLanJUl7uxan3
yhcuV26XWc9E6GvEudnGbNn/iboUKrYw9TkqNBrs9s23ezlCjnemOzoVg10q2Fyv20AN2nUVoqjl
XqMuNWYe+/x2cCFWfYLSecdeu+BgsPHptRIMgNXBbyemEuMyO31GU5r1yV/4aKv0EnWR6/O6C/Wy
UhMCJsRneK36jTTeEr9sJqWUu5j+op0UxgnoWBN6jVsGRf5JOXbUEaR6jI5RuonJm/DYxwp5RUY1
9/0PB+a4YvbsxuAwsF9/P2RlmCdIzSrKBtt+e0p2JAZ96VAPfesv7XSXQ+7DJJb7OV7Zm8Gorls8
Ndhyz93RCg2cHMKzq04DFo9WWVNLEQG9wDkGnOnjTPVg1QHX6vtoyy/6eVPrpeZ7LfPG0et5g1QF
r4EgfsAG9SZQM0DHMg8twtwElrUEx3BlsdHiWEphA1QirGgQAZog7reRklN3XIBaheHFuw6o5nCW
BPlK9Lk/qAjg4ZeeK90aaicueixCnl/s+SPGt74ky5+eZrATSmAf30fOpNKdhLfl7LkJ6dolTTaC
XIxMXwpzDXtQdHjR3xr774k97PGcecACqs3V9JdyTKRw8mvrvLGNy3wdPV7NvKtXnv61zQKBug1U
5MkyFJcbTNGoRtar2YbgsF8uOpACP5U/S5qjSTTb++Yu62aRTegEw+8JQJ+WU/TD7ysPLrUkoLKy
wZWtUUSeU0af0LzU39iLs/YmexHVUMm6GDCfsb8fV9lqFOsn3nUAzzVSW3OPhOn/7BgiHiZXGsgO
xQiVaBQ50Dwx6GlY5qLVfp7OVIeVd8xSVVCTC+QmUWyVtmFSw+erwGi2UfShPVjfoSB3+PeQB91v
8zxySW4RcVu3HLa9Pu0oHXPOqmbIh8RGAyDuTaNeT/pPuj8eS6l0+yK2EDUKOI5bl7SYnRS8UVNB
qy6Bjc70GtZHy98EFKHd/XHCDsZcMmR6Ennz925kEiOkfhroax75xRwMRbCsWc7IcCJjPAGgTqjy
bJUfj4qAGLrdiBG0ljCDuoZIcONWjp5a+55bjSLhKhq0CBYu93q/UNLu57SjNDARHf1ZtXFutfaR
2JGXnLn1pw1O5IityrVRAXc4up81myQ+/0FQ9sKDvO3FJes3iWIZwYApH59MZtbJMV2bLDhb/WCH
9OUYzrImlkyXQmn7salbSVEk4f54jlgshiXLmGYMMNGW4FWGYVgdKM8RE/dw+uTqoPRthkpwFGok
djccg2YYTEAjsNlrb8NGY5PW/+/+zsG4x/hjZnLFolg+mA/fRhHw8FtROVfqHpcrMQ9LZH3Kc3mP
lbjP0WMdBoTWzT5uWgJrUXlAiWa83YmQAkt+Vn+OoXxCueY5kUt8bBKTx3+X+QQwG2ki1RabFzI0
90cgChS/27X4vZKieCI3QTqwpOLjEskJWp5yoQrHVbS1HDpDkFRliFOgQlN9CnrnftzP6NZRxiZy
B+i7R08bi5hFScOooMeHHn+WfxJBMLZOW9jVQ/rIS1fpHCZa2SVgJCsio1GhTzKDSK+J7/DLVSfH
IvdX/nobOf4izMIVM2YxYRnKOT4cZMRA52HLf4V59WwSQtAyfUrFH6ToPe3QIisgMKTY69ZWaW1s
8c/yfZahjG7diXjEe7c5G/5TaosSDM+BAdqvOsCxpZUv0vQDAva054g3pMj+yMXxoUmr/bVfVFmE
A4XpeuVtmkDqwzrXdaGGQXJSnziZWsHngH5ioJXx5A+OH65BR+t0P4tKg+BhzkqVvdAFopzxoJyc
zO0g7YTwdId+UwfQHJ2BJklJgZXBlYxAb+WIuZ5NkGDPMdRQ+F5Ffi7JF+3OipjU95nN60ojQMcX
vsOYlOAN79KF8M4mDwLxEvNqTKK2/u5sQTMkh8eTAKlsVzA0s7xl5C7o7iS9st0ljboj313MCJvF
PxUTJZOC8e20qmVq31zby8lQpwiFyGNxZdxekZ8eOFEtTyP41tYch5FsRQlaJrmkIEbfjkyj+YAN
QZ0CGB9+/ZgbtYly2yCvJI2I4CgFOnP49DbdHG+EJYuZNcuI9wTdZiG9wHeJCac8O5xdOOrdnoK8
13b5LNWwz9aFqHH01aihh/vGrIdQAEAqO5n+wXOk+xcYPom39SigwarEzR089DUQ1BNXQhk4YN5A
Hb8cj3dPJEpFdrH3RaT0Xkf15znvtsCcf+qzgRKM9UsGegykmln78AeTM/ThPVJ8M8QldeMrssBr
zBQmHrfreXmzTWQLotQjnwvhO7FoVJOCAmYbJmKWn00HXb7e9c2snq4SYxCSNpoMUVpHNG0WEGVZ
7tE2cXb7SG+X3kTQJtfAC17yOfHDnjyPl2Vv2iW5fWapE3F8wGU/aOdUzkrVloNiG54Q0Cx2pD0P
sJB1IIrRBpixd+k3eNFrvFx4bgPPvvYC/ZGLBfDFU9SnzABHkBs18ES1CJl7nb3UrllM7Dtobbu5
/Ib5/LlLLHVWoPrVSG5gdEiGVeOss0U3jUH76nUNBhH1s/XbdKYEQvIuYGMZcbRVyoUOQRXktXdq
K5hAZAyST7stwH6Y8mH/gJZkZUqAOede5mmt23vz7uaRXJLKm+Y/kTCm2ql1u8v+FICG9kJ95AWN
5WtNguEZffQEfet9YEFYAsLTPcQvsghBDiOGElXYcWdrF/2LPx21Ril8tElHCwn4GqmicCJiGeQy
OyXX3PGFEYASPFyETg8WVJenhA/NAIDuNHfdAe3jE66hOIFrI7j5pcM+a1aQEsdC9dur8K5C1drK
0jU6kmDdwEb4MH3W7n1Tc9RLHniiidd2WotOFS+X1FXF3yDxoadcc45KcvnZWATKkYRztzRFgI9H
NErZKghp6UwX5ieBy4WCKNnEUihy5FX2g3vkeyd8AhXI+UXMQzlzYiklicAoeGD8+xTbzKA02UKZ
ojranBUKjTaLR2lNWRbwKWJh8GJX/iKLGw9roeg/eI4UXO+9mRythUIRX9XLPrtugZag7O6K4rE9
m9YtBoOVDUKSjz8eGWsf330IOqlmgilyfLTjd2HuoDfcoWSmZKuf6vt5YqXdalNdjzP2iYhjUHoG
D0JrjixSYVwXzMFIFSKqHxABAElgLqNKelLOwLr2WX06eJUcEpZYgoyd9Y/vUzklmuLojMVmg7P0
1mgKr0bO+nu3cRyd72S8mEFUbYuMyQcAaNi3Wlt0jlhtJgb3ng9RbMHui1Hhtk4hvIXSUCF0FFV4
+uCcY242RkahZa+3MLEpUJMg6YHv6pTQqaxtHlETH/3n2wqxpLCF+MU8sJhkOh2qG3kS85J1lE2U
ZRhJVuaCmfk+LRWoPjLrA4W3OW3imjK1bl5WeAJOVJ2FJvzr6WZMwGzRzxExAuITMEI3lfaRz17f
NhXEYd5CVOVjJJ4Yb2fqCgVRlCLUJBE1j+A8N7S4E+Er7xSPQrQ+yFjtGcElCokzahYk5KXe7NDk
2+/uWXpLcqzVCks4wPfg1c1oBKy608eUCsA6Mz6/SBc+Hu+o367OFgxvtmtgV3gBDah7Lwrww2LO
aOPJY3e2XGbtcJphNFum/3rfyYzWnxUoKTVaMCnPI96E1SUZJ0rM1bJly9C8n6khL1zG43vverR5
QkZbqurCSuM0c9Dv/JRGNbmhhWM2SWHJ8+sYbfuAEuVS1kjzrs/+LKP8vn4aqUZ4IFMdE8e6AqdJ
vOUn0LbifQOw9gP3mi+zn3KJXKNM0X8ecehUn34gLTaQLiHHQim4xuafjyVIyH3hdpt085h11+0f
vKUlDAAKE6wiwL4LGpUqX8EIo2uNSyUTBZY6X0d/0B1+OGgjOcAJo2OGKbL5jYhrxp05g5Htl9sD
j5QBx7oh3O6HhTMr5TXO7Y2WmlAffddvYl1NImKfxEZXswoDgz2TNl21s6WHUR0vFRuBKETQC44B
JI5QD7QiUHBD9i2Yw1KmrTuSskqXh7Q/75F4M1uUxI3KYwY+dVKK2Mgl3mKt7QuMdsY2pmuL1uos
UCDx3a6KDG6tGveHHpIFc0dyjrwJK7i6yV2YQ2mloJy7I60qZc6OaSI5bFAc4kNQzz7/8Q53J9Wv
L/6OeP9ciuru1zJrez0citrW3d9JXMXsvoP4qUsOKBuFcW+w4m0hWRBaUGXPY+WuQfjYvwR/xZPa
N0Q0+ly0j87pGJA70la4RUllDqGJLyGkZ4ezGkn9HscQHtFHLeLfdXCdW/WeTsUC+giwXOKh3G0N
Iib+UXc4GC18mYSvqVLmi1XUZbxuQAZetOhQ7gmo/amlTWmcw3IvsnjoS93lBDpvFQuxzvHAimJy
MREGqXVgDQpiesofysZUe3icVKqWgBKM8s9GfuKuRB3I77jcAaJlQ7NPFa9EK2MyFhvEgj23PYib
aK1AWnD+p8K+kHNbF3gUPGrtDsmpYxCIlU8BAIk7B61c7MdkEq7RQoHmWkUm2yHQmwO9RWnR2P0z
qgXEjnsUfjr92vuJn/YOpy5RZ6TDNyCqcNSmxYc2bXEc105l0KK3vPlWEm7fkg5nPysOOMh+gEc8
C67PvmIPk9a7JUi9a98W9SXQ+dDMqm/NpsK3vW0biZserJZYWeladcXeoM4nUXr+3CZSZBsvEeZj
YDJRmIdtIewNnEhfGOm2Chk9oGsqy5ny/byoGLwqbj+t3fEzB5W+dt8thaQIr70R1gY2ys8UVFN7
5VelzDCB4xEzTdDNLmXUACiX/Ugy4zLcdH9w3BWTqBeQuKqqYUf2sAQxNgdsyyvtYWIaGcKYdtFT
9mn8iX8PmAGfO/3BfbzXJYDWr8uvDa+IoDWVCCE1Kbif0s2ftA2pa1ZGLnve7CU1Krk6QF6Gscmi
eWnAdRD4yKaJQglRlMxOIMqN6c4FCt+deHB+TXUe/eZCfTcdGnyNuCAHpATtg9EqEIeCRxLa2O5L
d5DIW0HtgTdLyEemw1TdgznPLw5Ks6uspHyGvD//XXt36mfjIZkTgM9Unt17qpOZpyXY2V9ubezO
vFPpMO6Z49+dCnvyrsU8IDDRi2yRYHBstZUHl9v2wj3k/GcdLmoGIV4YTgdR+CVA/WhnSHm6EM/F
wrZ8KBkojbcTvVVvP34im6ddDz+20XYohiN5YKDye+x6Vy37nn99/4/CzGa01pthVfrlA5rWQ8JR
S6XRTIkAaxh4oXGkcoXfZHI5WE0Z+/aJn9IrMkfEgGgHIKqGddFm1uTo6KPZJ7zlZm8mti6do79T
ZWGUyZpo12AUDGBfxm0KOm5pDWPBkBu03czHh9y+GnOiSnzKYxTvS0pVAZ4QxV7MPn3RaejIFCcv
3FjzJpCv6pGd10uyUfRzyCw5tHf6wWoUsJP/GT0iYvYUAVFck/YlDnlVNMT5fbIi69j9ILrPXVSu
lZEG/p2YMJlGkyQxQrW3WGixrrSplTeC5roKoaZ8CTA0hnGZvEe6xGtqQyxUCIfdmMUTbyfZ6CEC
+hctzLrQKDi3dIhwv41Suc4ubigYvo0QWwpedk7Cdps+sZv5lQgqltgt6HDDbU68JrnQeQS0VRob
mA+Dfg1/q8KpQkK5cLeNR4nSgia4mDslDEvSEIUFsSCyl38kED2xxIbEpnPuXCrq79/x4ghc1xCW
kU8sQhp0T1+GOaqHvwPGOPGWmxEbZktcMq1TfpQu5TKVwfnDoTjWw9MlU0mggD6QCpaiJ1clZFbR
cOICN4V0b8C+DqaB3BuHe872kpttZGeeJ6T3pzotIWSNdBLKLXFelQb8Q6NlCMR0Ra5ke83qfxIj
6T9H+FXGsPyBWgiwQdrIC/9abvZ17QUVfnV5QIH9UpdHbBfJKcc36jJm1UCk6tDC28ASwggiA8Bm
ffGkfQn75fsP20frIi9aEV1WYFO7BY7Z/9MzrNieH+EpgWHpMgQ0Qh+LNVJi6nGgZiCFlkmI9PN5
TSLSs+Ee1sLzMTZsBp9yfjxtjpqoVHzgPy1anD3Uxpztr1G2Hvfh58uXqZxJzy+pVnEEUfweOjdA
uwGdJ/QD8XHLfCUeSOwXJcWyRIcWTIBcg76W6bOi9rigJGCR12ehQXGDVcJSWaeVi4pQ7fmRo0jM
Rz4uIdMajWm2zhP86I9uMpPPcOxdKoLJ4lfxlY3Fm7YczKdyHhM4Tqcy92eiBE+vKsbTbBBRpUMR
JXngbOyASf5xxFzxVgFnEH+0SpYMAPAM2aPzCUWA6a9qRx0HDphUOI2ENBaEc9d4TITmsFfQ71/u
FosyxtfKVc+LF7OQR+Q+5TwAD5K4Eq9nZNs5ohfbjAh4UG0/c6zC09ZhUIMveN1KOMcUfkEr0FP1
/mnVGeXfG6X3wV3vfg/JjyOVPd1Ev2z5eiEIubcP+yq3XiGw7v7YBX2AQlHR53U62qhdx8ik+7Lw
tSGIWDKdqsQ9yzcJcb4VhejrlbW/UrK2cOzSTtDj7tJwESCWPHlPunNxESxbxt4wGX4SFclDcNQm
8ggQEWz1SpSAus7oOPhWblHyiiv8AObaN4CiEYGChl+NZ3sJtegzqRNa/ZsPD4ot6ZFv58SHyYcz
ATO/qFkAMfowypXm1xUpF+CBwS3fn9YUBxlm7vtQk4ZNFlFJY6RA+uCPAwV4328BUWsR0GJ2m1mQ
R4wZqS7WK1VlTLWTeiJWlJHb0DlJ96h7QFtVHfh2k//xJymRIWCp4fgJ9U2wQQR55wKRQFY2Bn99
0Lg0Vh4Uz8PSzcravIfMTpHfPUNRXsG6B3u5CwrCAak9IKfICxC2u68I573Z+ffsbF5KUKBbmqP2
gQ8mx9S0I//uTfNDVPMhpY5IJRLfFpsPJHWAQWaXEdaajZv0S9O2gxw3r/sYkTQSumQuNRDZpaqI
Xk5A97UKq+gbQuNljMdWXAVdfahgroZ8sJfA+1Y+cGUEHbUcBnKPsk1SrMkp5csudIe2pYql357m
cTl+V2iQ6cUBCQT7976dAd26dsjBqOCMjv4FSQQAxPWRgTMt9dcA3xIlwmImo+XxH82EHxwD065+
DzpDMTuX2fCm8rcvVIj01ZTjV4XRtrfGNNlV0NosyV/c7hX1roeHXCN+ZXaqaz/igdn1ODBD/iMQ
sO/saXQB1zFe6LZMmrg2kz/RuRFQwwLyFlzuxQk0H0K59BdkYkApWGG3rg4hugfeTA9dzVSej10F
kB+yoCjyddRpFR/gJXKxKJoqHgZ5ht9dynatL6iZNjSl9gm6xcT4d+QGj/JYGqjOYV/6JAK8biRk
5bD9DmuDy0VNziZIg53PrYkZQuU9IkBZqnJoc1z5hqdh5BZLQ0HKoCeG/FiYP27jIm4y/U+stHy3
3+yY33xJaB1BY9y70Rx8GrMyn12ALLhWXnGBm/fhS/DigDCRw0SUK81En252IvajUiSsN+pkXyR8
5X4TgSWAeLO43QULdx6fNX8big8a+qI2M5KNcB94Ju/5qQAB2eeHVXaz+vNdv02TcFgCBZudhkUh
88WUOv0pdHbGZQ+EsTJfXqMvGix0Q9Jak+lBwycW9zx8kVB/cg8ym6VuNzsOsZvg1eIlc4pMrR4Z
mhsf+eD77Ff2Fzot8ksa6pWdNcXsfV9EwW53bB5IH9+NHU+5qQ1K87FxDvV1AnMbctazQCV87IgJ
RVuskk2mlGtfSn4pO/ocye35yAZf/GYZY7nQEswbWOR1orKaQko8OlOSTjupP+AU81LcGQ37oy9+
YKVkpNjnH/5XM9WM+DX4P0qgfARpPMaslNnPDnnju5CI/fuC65qQ/7GLSVl7ugHV/e47gcbP+d0i
QSjwlF2nxyXlOmIIVYE2UgGjmGhl1uFYLkxFTfZp5kFt2RsA4uJuKJTvViXFmJ1p7yh2j6Yhbbfv
qx4uLrMzeZu3P38iGsscWvTLlD7UOPkyvnwQOm0CH4rHLIaxOyKpLL93zDcF/E3KOrDWOj4FRBHp
AVJHVqSafPti5Bm9BPU1lSvG7fhbhi6kuMfreqMmpZJkfj6YKfHknNR9cocBYZDMWClHM4X1wjyP
bclrk5B6by+RxXnPitQtqdDnQVIWAo9iCF/OvNXz2N/mMHK/t4Ep2cHoC80e2ZlPHxZUk+msQ9rO
FON4K+s1czhVhsb9CprmWq5GrHsG+T2cvIljH6AgaILsYXPoireZ8zW/LXebBRSmcHIUQW+Cvwr2
OfdVmUdW3/7e9BsbYuoVjO+RcRUUCbwNX27l7/U9biDYfjWNS6LilDNzKF0DzXPCwo0HxVzdEYFT
HAaXvhBM/V2O10kN/eFhUI+bUU6Oo4Q41B4bM7p/NwR4Vmuoj5ELBHrnUVaXIl+lrRF/sosq1K+T
njbqWJRpuLd48RGkGsNyjhG1PZY/gX7eT18oqaQeFH77wG0LPdhhtgYLxj8kxhYKdbQ1wTR3ReAc
e6WXAFKdPHw0DmBRHIn/8zyWFrVrTyanyCN8MPwJBxiTAB4jzqycJfHzLtCYI/Yjpff8C/S1cqOO
h23SM5F7fIrFFFSrHmy28kSWzemNcM4Shwo73LPnBiZzNzzlBs6oSvJY/aJAqOlAT5/tJQNq+zm0
jMWrDeMRSJuKPqJqf8Fqy5FYLFerN/bJc/vhleM/d6mpkK2Q75cjMl+CwgHwZuBwcgXikTVh5VuF
aETigsXNj9wLDZdw614Io+J8QOMU0TGf5LV3PdT8mgkxUl7yGumXzOy9Bepz8EiuQ55QtWuOMu//
0RII7bQfpcBKxUySpY3PMoOfTZfkPQ+2ahZGEg+gFyGGYYzrh/PA2j2kQS7I/JL8Y5DzpYvpH1vg
S+mycIn4SPDxfvvto7343/RYI/1nz/07EPrf5nTJdVQPZK/ag9DdLZkQbo8ccwBy5yIPl8rgydV4
ewxhNMeqjOHndGKJII1yhpggNC6w+k8Qzsrw8WEUxgGCf2IMNDiQF4MKgZXH1XgoVHfOtJAGMGmi
iVid8ksa9MooI8nW94rsZ8Zw3idYdrtPU24GaFBs4TI2c3ExKfh7hVcuytQtvJsb5ZROlCtJgYv2
FsrtUUE2+V2C9Cat79hQJAY+znqlqXWzocLleqb+hQJNclfCga1S2T2WxC6EOMpJaixgDFsilJ5k
TTfvh+dNkVM4R6Lpc+mfrmLXX9PTsG97qGJe/RTMS4xAXTQSQHjvDJruEyi21/c/0l7rK6bpURvZ
tFU8lC4kCQUUO5s4SYSAgf+d9TU4VL8FpyotJft6Ygj2s0vt1bxGsidfOYfMB+gaGXBhNi38yscl
xF45kB0d+P9lAJ9GX/h5Xmjqm0r/WxnNjwoCw8aIrrzaML7qEHyskS4UktbII3Hxn3DCZO/pkivZ
fpSYH3CA6l51/IDokSH6E2x+6jOMgJDT7yPPIK73TQAiIFnNfAHnlo3RpdLkPB+Cs0oemHOd0mS3
2BL8xw+QdqWfIvG5AxXeSye/U6K/epxbPjE2i9CpAGeQdTCyL2SE5idpc5SMQBlYIwXc7iTS7YZw
LrOa7BHP5yvAoEwetVL3vUrCsdEp8vaSoENaC31Jlz2ee/Bl+HChm0y+0AYlECidItZ2R3lLmP2x
Md0nbsuSHuNrxfA0zu4fB3FB8k+oY4KV/g7qtulzD3SGhaccDu9Qu9pth32mOxLEliwCjlRVUIDC
F/ovAAOUfXP/BDaLHeDnmpW1cjEFAQQ2/MFOEdaC9OcWL9S1JDmbIxY1akxuVFXTpw4LUM5hL+2i
xCg8tDcSBQnJtXKfeYCIdpUM3RkPlN2YwtpcNPspDxjAgMsHyykCKF+UpV/JBUZAfgXl5efnHC8u
MJCHq8oBsru1QR1x9zis8bFBJZOghuvykVaGEaq1qsHEMaWF2Y6nblHRwgMjYM+aPImsTaWt4Dbw
Lk3lx7l3HbU49VTeMfFPCoXw+fAOTqzPYDVg4WrHkr0dByPOq0tHLIsuFKjXyDB262Oui7nub2df
RzS1jdIuAqAmwP9DEVCW/yY0DsNQ+aqyMxJuwEhUMv91kVDt914ce+Xq0FN9hyDHzEhOYKekDwkc
ksmWdoiwjfw+M19MtYzhKdkD/xM8hwFynrCi5NsXeSrnUx45F9uR98fMSmDFRurkIUREYMzjfiHa
bq2h+oyY77+vyRwRYKRpYt6BNRC91wZUYH+Pf2paruF3p0Oe/ZKMfnYdEB/sJcBKwevz1YjHw4ac
a1bt9qoGx5XDJ9oCdCQsC1c3VhjLUbA3b0qh6aDAqIOWs634Ybw+9+QZK466ubucz9heWxX39g5F
C931ijaF2d3w5LDLzmkyrgOKeIDzOr/81rpz3ptI4u94SGuUjI0SpmkxuriQstpbamUxrzJ2Zzim
lWSlt9qWGicfjSVWmt2cn/8NbIUXC+uvPOg6y8+QEgXWirE/D+r3qv/K11p2/pIetR8i8qasWm5S
9a94hQ8Ok+Fx6Ne3REyshb8hPCXpdvcQga5CfKoxwc7f85SUPB9N6eMqczI7k2u73lEHeRwF4DKD
kWCV2H63crsZ80Z+IJZrXVH2UQvIAOk3TfPM46GKvUZV3TcpmNnqB1MHQ61b1Y2ghcnqpOjzpahj
yYa5ldncLASV9PiJkPEbInVtnv21phd78ODcpAIuGeptqpuT1+FpEdfUexCQatKMVJDk7GaYrcso
MpswXQGIAmTstrIMJ8SB1JjsDlTtpKyxLSdcpmEMY3DkQUI029/1Zwy+imE6V27j85djnVXKa+BS
9eBjx9HVHvW1mUW17vvI7dtbyTDfVX1yzOfSb50ukzW3TnuuEWGBvCsxtgeZuyDTnCrkZIGPSc6L
nADmVKy0isiu8Ccj9Tcjsk8iGlpZEsVUfj2Qtg0JWzgWpioOv2grvf5lNHqT0ZoIo6gd282T6wzF
Dm/z8GEI03eieGLKOLrqNcUE3dZxLAl8kBQDtCERj5Bdr+o7/Mtg2220OuQOzny7/kxndMrIG83R
tsaZdHCBz95zakneRG+CNQ5WDXTbWMaPQehSqjYB8vhUj7OXGxJdlnqsMvgXcOEX5v2fo4sQTD9X
/CSG717zjPYUM93AedysD/kyxKGSWgobR9GY7QyBpsFgYdjpZiKvi9u58rnAueZURZ85SpYJdVAX
KuhR8J60Io1jwYhAWemhz+y+NCddOEaHygNqR5xRksAWH6YFPbGvGgdYrRuvxLcbSfQEvKkmyMFC
gZahtwjB3DpJRWKjqm7ySk0IpSBzODJ9M7S9tsmfXNL8xkIemRozKwm67HPGQSyKaVmQzK89T9Ld
PkUaP408p7P+27RiPwteRxsVR9p4XPbiMJ+KIrHtInY9jxYyNMGddZRZBSlPkNnjt3YUl0rJ3npi
Y1jG31lDR2kh3ohz0TSNT3eBbuHyo+stTp5ri/2XJ/J1qNUEOEBU4/jNDuZZtPXUhn+OitS0gJSZ
BSsm+a6Qg5ltmB5f4pk3GtkX5XgrEp5hcxuWfoklrSPy0rBmMvCqTSs4rzfCsjRTK/AXf7n9e+yr
sOgm6MMP77TPg17USc5Wt3PwkZ8zdHeaGZJ+PXNfpvbH69LQv+CsBs+it178/b0sxKoVCSRPTmbp
xrMsQtOsj7NrwYawnM6hLmNhGBX1ocppk4e66lG91QjyxzmWGK9rAPJmJXLQgR5FqnVaiAkRvSp6
Z26i4PKitd7spjAGozmRPPLDxQZF2lLwspj90EfaU3rDeIrH5pGCC5BdwBL43Hz2Y5/vZB4tE5ge
9TTJOm1r7HpnRDlDf+OVaiPkgWKr2qGJ+O4xbrh96yvlovVTs5PeyYz6eOEeYd5pCaS6JBk8jBbR
S5D0UoBhkYMcfK0G7vFZgEcMGR/S/if+DEkZDnRqQweCga9HWNvFw9BfmaurxYWEmjcdIitp9/Lh
ogMd2siThiiUjio9uH6/70vBWfyIbG3Xg9AbeNwqld923D1uC9VYaCrSZmEo3+30otQ5ycNcb9nU
EFxy1iNU3if86rv7DBaoJWHJc1tly4gXBX4OMQ1GGjF1k1kntWFVw9HyGcVAdblxZykSSBQHmOtT
Lw2wUY1pszFpHh4OO3xyPWxFc2kYndqFXUqHt0Nuva25UpmxNWElyXTxP7NJHqttlt70FwJn4b+I
tlFZwJVHl8Xm99CHKzqsaOQ3c57ABmbsamlaLZpaGrLXW52uDaPUlEWqLfhCVqnBQpIg2kyvE90Z
vCRXhc23h2gjxAv49t3l84yf8CaX7pTEWFnr886IH44pUsIeXQgC2Ld3vzig2khfLkrdOfuXC5di
dHL1KAc4VD9yD9fiAot9uBk8Ava/lIt1Lz1/bq0VDBtuxeQD/f/waOD1H0LRfwD7FgiUGVJRtoNh
ATwPOTWCFIrPOg02rO4Is7EFn8hp2HvsrMbsLQ1oKkJEXEqz7+hBU1ZEOcj7dkVOjpxb0Z/HITux
B7FpO5Lt5bfn3m6ck+AXl/gp8qpze3XEyMk+ok1UJ+Y1pmdPBkBdLdGc0KoyPZJF53ZT2iwQbHIO
cs5eGPqCqwxJ5Yyay2KNPRmrlz245vWlovfQ9ODBypQo4ppspd+qlQ3NdGCOwxLOxHr7KcEECgUt
QoXtOZVeGnwG0kG5q9mX6eL0qUhWbc2VUGWuYnyEvAiO0jgTnFEMOW2o34l6YfTA09MV8kihiSZz
tYrvkeiIqv8shS0fNEtOEwMKORJbJ8c7FCMogtbGLOWwdjoUCUaLxqjuR10br4VR4qtOgOeZIf7K
slERzJMmjHyTwyIemecgjiN7R+YUimWj8vWbpCdrnc+Bd2rGgSwGmBC+FNOR2LCwE38sqD7pE2nm
+kVTUPNtSxT1o3b3KYAv3smMdpLmFHIGOX7h6o0zVBSggWeetqULirQpkXsdxDigL6F8EgGLBmPa
re0xWgK33gXsEUzytZi2NjXMRsZwhzZKcPNbJv+AIU1/U2BhckyIlSbs6aQpCDAc9bfXOwcMPllu
OV+IqXkPSKcibjAXAvNLOYctD759YyrG39TLMx1JKs3XSYfCUUplc7dibgAwUBITHFL0GwBfESMG
8/iVN1t8AoG/1Hqvwf33g+obXeMMgOL2nO3ojYevs/dGSegjl3Ptns+MaCaQ1+eS4MMNkdUFUyOg
34JqFQSGywJQlKzvRapIpM+97KmN3m4VvpSXJU0rm+64JWFMy4zXA8cwX8wronwv637rmDWkpPQX
nsOmOtpywlhEKKbhG+Iqz1yt72zZuvTiTVIx6Y6HOfoi6ycEWta3AYqA3RqTh+fevqFllDX9tGrA
2aL37fZQjIl6KIrSR2eREx2EIhMVRf8CiPLGV+yUX1kLZW4zpOL9qNlvCVhbLiBvvqdaLkA18Ubv
5S09jW5Jg+0LwArfZ0GXuhHzGB9yocKik3QEOyhUu9kJBF7Lvd9qsy6vFc6nHelOTkBTjN0KovFT
33D6TYTnA22CV6YcFLQB16A7BEt2NEz+wYZ82iuJgfha66A2XcFiO4tq3MKwUTCp+Te3IqEWnQZL
BUX01da7yO0NCCS6da9n2TWfVjNkc37gZ+oIjDUj3875ywW4w7eUzquduM6R4gl+hG3FjXJt4Uc7
sn6Hosx/WoJAhBhfcXX3XbItKTN6AJhL2rUCwqoiyF+fj5m5IKzOOTOi+M0XNcr3MxtEOPscFW/r
zLxno+1zWLSmfJGpqixbkGETtKT9n73IlLds1cdbi1HG0/gxQ1C2jCe9yvP+0gRncYmE/joE8xpJ
q7dHlTaII30MJEIAV5w4MPD6OeXzdQQ/Y9QR56RkAoslbKweJu03BJvxZ/6Lj3Cdi5MnKX1V8Psv
v9N+E2CE8r0vXtOiJ9nzr68vWl2Gx0AGrfooCs+AdVxySeb/zxHgxjHwq+zPfnyyQgClnIP74bkG
iFWwahAxHwr8a7rMOstkMmUs+0+KTP/snwXZRDGNsblRUnhcYqQZUkASnvfYNHT/vca5F8TDevAr
0v9cXuXWRStaW1Y15ZxYYsYl18CJzeR25jgFo1L443iKJU25YMIl/qW/8vfY6tXSn/5aUq6Z7k4K
7dvli0yC8Jyyc/WCmoXnj7G31sa7JNbXugHhfY7+vxavx99A3bNzFLJhkMgnojafuuvoc5PYHIW8
KdqAz2v6bW8S3o2IWahlk+auzrWuN16oat1A7UBzRatO93tog7h7RIc8z3l3HYmtzz4hOl2oUHWv
UpmgxKEjc/qn/oSnAu15yztqRFzmsLOIf3SK1dS5BoJDqWA/nAe2fCbWL0c7sc7aHBT5rGzUjpaj
m2lWkeW7Yq4wx5eOjNlGJAog/8OIj/XFouZqeXRcie8Ntq0utFEalssS2Xl2MD4r4ipz4/Ip0m1e
2M5jscaPSqqW5S/w7hjssfjitKW1o/bHji0pq/r2FEGJ0u5RI8tt2kP5rHiUsDZlavbtemPPyUPD
q90TmW5jPF+J6Iz3L3DFUewnFmMYPSqI0QDL/W3GbpMJiyA8iGeNzStfSwv8UNwcNank4ZK88QHm
Hic0WnrpGUGHtKKvxkwRQJCm/EZbYQRblG+OV+6tmaOhPR/nX2pwYFHeM65d0q9AGo5Wn3sjf8pq
yd+SGv/scaGcB2F8rZ6Cazo5elmOHFgnBTjfniTf9UgCYBo9vZLZ1LHYeCB6T36JeYiBg6ZJo9Hq
1AR09iyI9mPQ9aEaqPQsEaDPLdRRvMoi3Yh9Hw53Yf8x2Xb+XU9SC523S6WFOlBySRFym3ym9m2u
E/21SSDxg8SQEFri5a1daDTt8iFln0yczkVShFOKifn+at+Wk26xJQsTT8XgS5Mdx36jsuGGXJy5
8ArJwB8VaLQ2JeOsgesTY99BV0ZYiHu0e4VbdkqQi6st6RL6BB+8IgMdO5yroLK/SQxCwnFW7/BQ
11gKeFbqEf84Xk6jLCHvIouOdf/3iwzsmJPIssgB4yL8UllDss2JutWUphN3Tc21g8d6b/OEYk+l
l1IhH5lzoXy5jd8Abf+mHzQW1LXMwfCuj+z28Wds/pOZVnlk7hfvc1ZMRbF3c1J0seFBnGoGzkS1
u7sHcHtUa7wY36zQM17QbgzFfbGkQSk08QcvcF57h2bi+OYO7iUHhe2LQEKT4wQvc7a/Ou+D9bU+
ehdiVBZHFtt96gWQzTx8DTwTXNvosMc5h8RBVFVmTAIDHP9vWDnkkS6qgUawMzUkUo088bD4/A00
sIvZEDA0mcvOWyU0zGzZf4OFe+0IPwHhPlHeAQ5lSJ0ct9y6XOEGvhn+K9BCFr4i+G06b0Y/78xl
e6YH5IW/RGDYIoA06+fPr5DYMGqy+jQO1p1r+xjm3o7uDNXe/YMLdgNaESkNqqNHat+BiMZ128tL
h8XQGAFLTpU60ffqKGQ6rmdKswqvFuOSP5O7t19PEM3sjkCzFclTkXt0RtbIA2Ml6mK5/T0NvpLC
PSVW6At8pvuzzshWtXK0MMdH8rCQIiEfWQUpt2BuUEObjPvKcX47b8GFZ+JBtNnk8/R6tUEy6U9A
zKDOnfYS5s3PHERPfoPQPrM7qDw+3529fwGNOOjntlJ1ZvaYKGWhAQ90wPe8q/ztmyKsRmuvANR6
i2MC7LBXnhuW5wor1wb2mkZ6aN1As4T5JvXYI8ZbwNjtCshvqZZSdfLJZgWsUhBqW/C7XDelKR7l
RFBm21H0Exl4OFsPb6aozS3Oy9EJIKUterDfww2OWhUpk6thYjJ0fTJUvI81miJTy+MVSrGRJaf+
JIOsDMyxAZJjvEFERJ8r2rOEDkou6BAwgPP8bBZCacXBBHFh/RvR5oOrm4D52UOput0Z8wHH2/Fq
MaI9fRFNWpc6dQUNmxDXj6cTa1TOS4Dn3jnostCEJ27xTsPeKDEBjsYYhJ9ATgE0uEcKz07jB8dx
5NCswIq5R5GjJsIq4TxwLtZgZem0myZKu5x+PXpefHUM2N8P55PxGD1zqXB0x4UbtQEUYFhw9Rd2
buIEQWu9+aVnuY4hjvivEsVCT73gZf8wm5rbpuiSFCx9Zc+HkDpbPZdVfqI7haaZ+aozXFuvSMHb
ZoBTGVWpp0gqj2jid0jhw8aqS0qML+JAKbzPfhiYWquZBwz4wpmIrktmHkupKAVAooHRmld0Y5fk
O1kdfWi6jvuO4DIoIZvDBxfSw0hEOW/jeJ6HH8Ya9xuMFZraoBXGi4PpjX2/lqncF5vEfRurKdU+
vbo7j44Ljc3M6y1Sgs7CkKo/vB3K5vkGwc2Rprh9/kAKqABQlTQYgKwBfl4lzhFaBL4K+BYnYmgr
xDnace2LNWyuvpEh12HwDnwpFYEOySiVoW1oTTGKWL3ifUjIv8sg5yZNzYCGEdbAaS7fhY8AH59P
//j+Lloo2v755beSDicUxP1X6NaYpKfzeGjGYIuHJuudZfrXYPLXk20DPKReHJ/F5GYoEkUZRSEI
5lS5LwolXc3lsWqXEruXtp2pcviaWmfEvjAt898XgPAzh3DgDWCPxBs6zxerQBQzIxbiXw/7YSEw
b+i0GDL2c7/BUdJKsp8utVO0HV4NCinyp9thamqxpc0bJ9DSa2G4xplkBlDtORXk9XBfE9CMEeYy
CnXd74lu2XMRH7V+5nm/d+5bUWi3v4JL2EMhcrtku9EDebAD7dyNhfXiCEUJ4xjX9Ln/m3MH06Jl
n2SDf+qv7QSG1Q840RSa08Uo6P3/VQgTl9ynKibkPNyZmMf3Unck27YF/J3kgFbFX/Hc54sF3+gt
YF2hFePNZ8jemoLAjovi9njghUMTOmbl+sQmF10xDg77hGUxrkzd8n7kgyOJWSkO4L5UoIOYFZ+w
eEBBemPK56Ya8InnmeU2h39DevEHVnh+rYKFhP387liJSmvKMd1xn8vpCzhJgZkqPcTKdrdS1/yc
XMVC3p5+3JDgcR8dokuij1LaEFPuPm8agldgDZn6rD5MrfeH0BHL5ZHMoNPPUFxwm5ikMVC+hqtt
5Lq3m59SzwWITdNDZ2Z+vPV2YSffsoJFH1FQYKVSdcXx6Hg8nftFhkC8QfLIatspm7CXM5rweLRm
2BQUGiDxApLlOrNTIALj12RGfOG5zdC7ft9+4bc2MpIJPBR7mhy/wGUPqs9kAZAh1GJ5KwWY/6Em
Qh1+3JeZrnQIoAn7IntgvL8UIilCRw6g5WkbGHMOlHRpOrwWnUFeq4Llhv9F/HEf7BfqwtNXPE1w
Ta1VrSTVMlA0m+ebwYoegoYR1N3236tEg6b+qUBKnmZ5X1JDRTQQ8glBJcRG9s4+pHeTRgsIfxvS
/QiPfDwmjIdV2R+s8A9obxAcernoLYBb9deMF/e/0qReZtx95HFfIsuGluln/g+/m8OQSh5n/dYg
KG+xKWRqz442c2pjJEIcV9+MDTx9qBFXce4lUgXxE8ysc1yn4XKlCC7ozw8LzR07UPK13xU+lBcQ
p4Q76X/QlUo5lEt0iBm2DAhvnKxZTFLs7u9jbjAicnWKKw8Ed93lUCxHs4EJ1pnfQqHEkzMSPH24
V+ltqFAEYZ+AiweOG9Wt3spJxsCaKPsicDgATKoVW8Ei9Nfy0bOvgnbSkB4OzNjE09mR83R0U610
S4O730vasMRBICo8taU1zFYyh+VSNsZ173OqU93gcwKtQZUh5nUZ08sx0FN0we/vRyv6EVYZFOkU
bq9JT9bKP8ahnq07PbkqtfNfkntKcUi59tUUoY1M9StIq1Qj82SGtGUwiW3uFm0xzyvs1lcBdIK2
l/N3sn+ZKEoXVNoJNvJ0k9fNyP1tojj0fswfYtn3ESGKUdSbxI0PE+Oj6WkvEhy90LPjrqL2tBaC
uAbHCq3P6qW6JacLUPCZtVf4xDXKVI6g0QtofPZ/eO/qryQubHcY5sQ0AuHC7zMU5MUvgVjW9gpe
wAEwHQGNX3lBLwIbRPIKpPf3J7BXmopcRythikarRjmcRc+M/VbsplSDPHGEaySYLQOQMyONoEJk
ONIqxfnArkkNEHyUQesV5JPls3XgtyWmScy1JZWSD9Kv7YbjHQWMG9It6jFjLvmFTApXl0uUVL20
mXbSR0/NOH295FKR/09A/kjP7fcnVkzJWzPt+K2Dq3ifko+OzN+mWp68o6LJKR5RecCJLwQ6usLZ
jfoSensmmge8exHEGdi36uB4JR0mYQ3temuKdufKYclkBRU+W/yEemMeU4Rgq5z8aKbWHb1xPQwv
oRrlE1io0EnNYFr92T31ypsm3o5bLyI+ookXqnFiQUScm3YTO9aP+e8JJijOA3xLPgh1/YiHLO9e
/sAWoUfdNEb6c/Q7kYULR5BXnu1wAfMHHioE0tQU8/gCkeokfYqIWyQHzKce86H//NdkExkejDp9
CyaQKMdyRs6J9xT2HRjqJeIFDdr02iq1EDiTwdu4cC/aWHYwwHvW9dqfP/uzMth04gdp7Ut4s2c3
mAXyMW3h912uUIqYTrWhKuL9OU4RKn+cUrZPRYQ5lyZB14nW2C3bOta28LXexeX9FLmKh0nwdtDn
ul/J8QQGrio5Imefj2luQDA5Yub85l835z1vSic6i+9Q44FFrvwL1ufgCXAya2IVDypl1A+CrR7T
+fCMiVpJMiZv5nJ5It2uCzcl/I+P/KCgsL8ArFdqDpYoXIY19upxjF5/MX4Pia8JZTNSXeev4Uo4
lPAJn72pz57VxzIEv4GdNeqoa0kpYMxQQ4Dl24+1y1Fsk4wtjbiKrbPDV6cz1dJwRSNcyiYAAniY
GMwx0t5sOffN1svORpHERxeqyPGmrXTk5pwN2RJg0JCYaXlxkTU4t8e4nfPA3zirJsiX9pcQg3lh
aZdRgOFdtOjhGafB/I4mQ4Vh6s8xFDc7UbXUPTM+NM/BKhgRxmCYE5qK2izUUXwt/uRO2wipHRal
JbHvWhdH3lHAUkl4+QEY1kD96BtTdgi/tBMtZUMg8jzNeJGXwLinrLPLgftvxXy/X4if0Pm+KTD0
eT8RNpFh9T7ME6cA+ak29892x6IOrOxHk15+lu/svglAE+COJHbJDZRmF8c9j5L7xCk/f85Q91Mf
xWkX5qKQn9RltfETqh76amigJo9GEE2uDgmxd5wBKTindaF9Z/PwqYY5r7CDKOsZDrZwj+S2MgQq
WEESzrAIf3DecnVa/Rs5+1gI0SB9FDIkS7xpNWHWccKbiwKeGsFN/B8uxaxCmdNGPB6iKKoRhBYN
rX377rjyfxu/+wawKIH3/U9SkWxyZHspVzlBXTYYXGRwUrsHfZAhBPwEkfgyUZosqV9CmL9lNk2o
/mRrEc3EKUrarji0kXq8qYjSNI6oJkXFsKy00Ae+tT8XACSheJ8C23zFYP43hOTz7+92pSP4a/bC
BQs0q1zSh3BCcgrVKJ/dXqUUSrf8hzq4aTVz2TUJHGCSavZYBhb7FW/3iW0pNMiEwqgCXoihrzLv
D+nWvQTlfvHhWWosJ5UdMYUQyGvDAHv7D1N1R9V/+L6LPH/SHBtphO7NzO5wKkug+aj4Ijus2io5
0akwch2tLOPMJkIxhdJA6No+N1ZCZ4M7bWMVybDsOSQ8HngHbQBLD333ih04ISm35xlOvnhB7RK2
PejkAK5U/+8CGhDIPs/B9yHURDwYWGaxrz7F4P26g4wc73C7rSrG7N9pJruI0b9biCRgcXAawmv4
QChS7YSG4gPTXfMfF1lSeGvfZ3frnVe3kLtcHLmco9BRmKzyw0Y/NyN+0JZpmxYIo3vS87KHSgNp
T81tyJ+wUxUpFXw31nXyKGH9Td/YBC07wvXMXlnAd/dwfhGXD9fkcaME3rCEabm14nbHdxuWyhm5
e1MVEL0RNjj2ZXn0+al0d6ZIpqzk6/KPFZPdmlS1Jq6W3cbJVXj718Ct43l95//RcRVsbRboUR0G
4EcL980tlf7ekpHkkj3z32t/EI8faDVInf4pSbQqj5JsthHE1ZlCfkVznO42lUSygD2fuaAsAHW/
TJ0f7ygyJplGGjjN4xo5tF04bjXubLy2p3mfEgk3DIP4fAq//T/CpvxwXK7pDR869KT8fjxTy1F3
e8qApMGMLqb3qJ0Nki2pOrXGXEncJVETuU7HA6U7/ws76C4c6JH7MGSRXjamG7XAqnrE89vph3ka
wH8gGZcD9J7B/eGLMlGgQd01bYzE3Ztxyx82zIicRMLBlcFETsZcLYa52EbW2qnioILABcgVa1Q4
AeXr1QvaPOFu7oRgSmTkKmKJTR1fUdUkJBHK9P00wr5ALRDtGX/GpOi9Ui60jMjts3a7sysqnDbV
IU0IyvmkKQZ1M80VkODhIk1CbqRotHx592jNKofcxBaErU5YCg7TzQKxsVJ8E2wu38EEk3IZ2Ms7
uDNU/VHOLaZOcJmN05hdzfJh5+sx9O/13X7sy26tdTqhPkAGXQ4Zlpdvfgz3LAV8bFWN49SKOqjP
1YvShHFZLGoIr03Xk/g88Baz4+vo8P+1vIVgvd59ODWYahgs1+z/wn/i2aM9y8vc+HZBHoBQPXtK
xcRX8BOf7wOMuW7lPtSeTU3Ibpe9yWFH9WONh1aaVnxdzLyYFpU8spLLvPNAp7e+YtYpWYghyjyG
LIQfwsC7WaKxM4K5pUDqEIa9hTMrnFiUQS6R+OxmqxyyMGPMjxwHHP7wFdz/TC/w53hHpFGHfdhR
+MU7z0v9c5J76M86BX7a3eVtNl9IHBZLcXa7Skl3PTGLqsBA9pYxSb5X5PvTPSN66ac+ZK90feSu
tDcib3eZW8Qy+huYkXo/5k2pYKmP0GWVDAr4DbMY1fh7q4Zi/HHhn5wWg5oarBOe+Z4EP/FbNo+W
YrzxfHWZWTkb0DiBBFzxIiOMocq0hqExpXilQ1irUb4p2ZsYh8gZtLxjDmaqC/M9a9yi2sDdfKT1
s+mVvXaZgaF9yF9sbEn43sjS2WLhyAYvaSunoiPD1mMGcw20PLmubGYIH691HMvO/M5KhbfqrSxC
SunTMNgANdwf/MBUY1PMRsNWSBeyTsGAT/5G30z5pZRGpQ8hYN83NlQATsWjOHb4NxKYmqJmXfAW
hXjUa7xJHcV5WwfmCzEP2Kp0VCt6TcEVafQYfG8hO3A/wrx6RpWLlzV5ftJutPxCu9zvRiSKNnw1
ICoRBmFhvtsdnbbdOcqK2LLYyQt5oDfEp6kRGQnMeST/kiV7olOZ8Dxlq59rvorV0ZaFd95qjLQB
fJtSuiP5+Lo0plTukyhCremjNvSJW3KkIWgWZX1ZdfO4AMX3YLWrQF4RAxRpHkCk3W+qJw0YA7PQ
cDBAT8drBT2nRTsbOBxmopt07SG00y+rgAb9H6ycjTLdAT2cOLJpK4hERrz5ap84PaOJcUxEHMb0
3Ldqu8s0fCFOBZGW7QQSirRjmDnZi5ZOTQfq1J2C9/WVIu8yDoQWNk/I8IWEWG0fJQI6lH1OSmel
7+hLXjVxxGNjoZyNZnJHxiEBdvfgFW9oL6aLUIFAC3zxmLS40kC18O/U7wt6Zh+cI3BYnOIwOTrQ
5cbjVgSxYS+s1X8KDWHIYrqbYXGb7E7dfKbqYgtJyFk8UKmLj9d14meXrziLsFvsHN2pDlw66ypg
I9h4hk1xNLYyKx3JXRNQcPBUMW7yZEeWvffQLGoAIcjNWSahAjH8mY977POEooI6ByoWuS7lYtoU
wxme+SHyZ4Z60uvISy6hf1pNi1KVS8ACpv6qmtypGn7jrM0nj26i2EbOshMNEdEMpxHJgLulSHo5
PxsLHF86v8j35FniQQJ1LAujkpQjtN28bnsPNjw2j81aFolyGcSQoGRW4S8U2Mjbn9H3R8+pm1lb
wNZ4HEyjGplEXMtaCC1ZDCjkCajF5aQYOoC3BK7DQhRCQ0xshw6kAaAJaKtGzWBroRxGdIqTVOO6
gsX4IKpwD7rOkHOKjibPEzkP6KSZU0x7KIQp73Yc6wdz18r0fXqiBaqC6DUffyyWEhloycGLjR11
sHstjXcBnu+9IltioAZGMN0viH+kfsekLB2MbDSJGxSAnDWC8FitAtKTJ3XlBcXMsbnD476zwm3p
3VzcQxED0ebElbz0eQ8C4epjVr1JiNb8veFXjN+tb5+18ur3itqCjIoVqCISBABAY3zHN0QKO1sv
HfmqPlQrSZXBXddwxWWp4FCvyXpSvOGHFJlp1k3PYHhFyfG8tkke0AEDAufAXlAGlek39gn3FgVC
5EiRqj08vU1xO2y8s8mM/p3BydLDMIYuJVjw+0Pd5NKZsmVrNW0oPmuwj0Fu2DsX/aUtpv210XYL
5n/O3+YX1eqba5QteeIMaklOJvOJ/nVcCotDoimxPnlkcckgUfKbo+Rtgwa42oXg9oOk+BfTw7Cm
/AwYNJu9YSLLtetsutzfJ3tuxLhGTfVyLff//r3wkDFuy5ZR/+pv969hPkuHi1d5enpv3IEZhv9E
RoxPn+xx03RiYxOqXaavOQYEI2DTZQnDO/P27eakAuv4MIQNohhVopsxXdSVUCOjawO+8YrakCPD
Fkjg7R5qrTScIRo665MXaCeigShh3PPIziqk1sqtQTz8oq1/arx+8ZSelU4KRR9jRBz9h8l5Wivx
4iPdjhDocm8BCkZB4HhzdizSCYsP/TUot0CU7a0h4IwuGJDd/uPDzwYBrCq+Nz+66HIrr943+qkP
0/QFxu4TwS+HApGWi3Zub4+ilZdTheuM3Ql13UZeV58L8lTEHc1dQS9eSopJyawDmb5A89y0kuZB
gw1ezxdmv+mi0yDkhPWOaWID+m65yKxdtyZmfzv3fD6UWW779lNswkHUX6hJJ31ANEJBzByIDq4u
4rCmqRlXZOnmMimg9TkFXp3ODUgDeSiMSlTZpd5Co0PrAIrM3oUHK8Gh8oJXl6S+S9WQJo1AFd54
OdaE/IChZpJjP+Akd8O5HEFpJITBJqhbw+fvEMhtXtc7pScm/xN49oUxpAfHcV2ezjpIGaphTn5u
OEHLk4YSDAUnfBLqyCcSyFahI5USwQ3impMt2xKaMGoU+OhkI9cCYEdWCRKN5Rbl9n0JzHvjcbsx
7++YrL1zXxCCqwDhhE4/jFIcv1cuPkTWQ2LRWKNF84F/LvuYuYFvyPTJh7pnyt86OKu+qjW8tAJc
d79JmiqinZPHTLlAWS41H+GjChfl1pT+1wPAfWiWjM4mvbQUhTaBW/7jk09b4zKI7w5rru8qEkHE
CdIrZECBttvYKOKN65Aa9K2C+uUbFbvEkpG+wnSmiZ7e//XAvaUAPd9GIWmXXozZcLgftazibasY
unAyVGJL3p1js0ZciMWmPrcrwqNaGiwhJqfl+0gt7XeGbtzq82JCofbZeB9YxcccyzM9VxC/ptHN
jpRUJ9T4cM4NJy4LSnyOl0UCmV+A3HT25vP9YpnuWlz3H+uoyalKCpWfGiDrFx3LIM9U/Kdj6qkT
tPQBHY2Z7ehNg2zM5IZYNFdOyNe1NgvWZjDdnLfGynx+tVIdpCz0c4Asz2Ixslw0OuiKWrXKgKa9
Gk0BHOsOROCi2u4NNTQOq54Qj2IZx8D4thYMSiTTuw9euD+pAFznSFIukNl/O7t4hsZNwROPmJN6
c4oPOv/lO+w4/oDYeDLK+Xx/Fszy2ODGqUrDqTsHd2XRdez9qorPvPAvSMZqJ+qSfKGNF7N/6mAB
mMJucWiCJRYQx6Z1NuuR6OtFiLyhko3WOXvkXwkVq66mliG6/FL+b5UuCa68kxzXHQ2tlbyQebBR
LZu1GvBDAf0vb4AUY1ybBPRNgbrCUykb7VVA1OLyW/n1SP10EE/Nb7k5ZDxnnPhpl9Bxpw0kNmBi
rALA0mosGLOrxSQ9vh4c7PZ6mJo/yggInnI8Bc8tEwfUaiMkBKfTOIuX9f6nvtQ0YPV+yDGQY6QS
JiQfdW5s2No4teX82nlfxVKosXOSwy+MSzPDboLqfDVlfFlK+7u49CIXFoFlA39vZlb0qTgWzBfw
dBc6j7id4iG1T3XvEgynK6b/sDIc7jyyPISHGbtJPxOFUH+DlaU46lkRB7diK3WGhwNLQODp7klG
aFGH2PyuowBMlIZ8CEz/V20sMT+AhBmT9L7JtqevamMkvqqm6idn7u6CHa61MHnoR2GNF995vu5A
SwMTSdX7UWzR3xab6CIkw+NSB1ZBu47kSUJxUSkCYb90Cu0BdLLU2z+mHMXu/XqyG3k2QC2QRGN5
snGjJlTT990KhuFU2pfJpNxIn474f8SGzag73uekRKdud4xVdkF+VYZ6vXEKM9iV0nRLR+qtYuOn
282ckd8bVWyCZqo5JJtE2OzWD2r57tPKEftspwwEwLJ9l3jhfSi3ls6CYmugUHvDBPT+oZFHio/l
tUKQkR0qI2LO0P00CHyHbsBv57QqALx6sNyZhWHNTCknFpgBzhI7TTUjGrE3OcW+e0gSLVJqHUDn
QlM3/NH6+wpqwWCrp3Fe3b5UuiukCtgQSBEV4aWKN2MHGvp669bdY1j29Nh36aOm0gLcH5kKAT7K
E7xIp0p16X9LUHLUJuNO+eKZMs7U5Bn6QmOARWsMHhZhPE9bWBY9wjkiAYoSHrFDjo9mKzGXkVnq
0hCR+1DpakFPDGzJaaH9Kz1A3IdK1KHDhtykagbCKkeHCnBRCSRCQ22wf5i5cL8iBMPkNbZn9h6p
j93HCoyzj4NOvQKr55ij3drcUrjxlLLTGGaPaopjUwbWXRfXXrW9hbGd7++i2Onmz5luhvtw5l87
eMa92dczqqOhLKyKTdkb0hC5pwlFAb8RAiAGwyhJor2F3xjcuenZ5k6fVP2qvtHR+Ju3N2xG4c4t
312TyASlnwXI9rMiv3IYfUe6ZJy4IiosfDN8Q1c6ka0khIu4NCNCa8BROi/cTSfndoxfZKkKZBd5
IUGyLZQU6cmTBWTcETq+aRTLJDAmecnRMArC5nMS8EMpU/QBDNIS4dfnXUzHwLJbKfvEV1uxtSt9
8f9oKtZcpM3MfPPC8FPvWppUpsodHjHWRLDhY++03aTwCdJJs35KZbLmhAnbmNx+jcTtkr3JQXsN
bVfVx1lWyMR599ypVNXHSM7OBh2hz15xRgeKtvGOJQ36f8IFjljE8cZMTuPGqHvzUG4V/CmpvW+z
yCUpr82CgdciKuPCbQSgELk7R5viGgmry+xN+CqA2da+gJhheiw6oJXLOfp+7bM0SPA2qMolvPqm
exa2uC1zPTLvIWCre1I/B+vsUygF0uf3PMhVtxJ/7imBO/mJt0heJ5z+N378Ag3eWJnJu9nCXoY7
9J+wE3rASlcdALzwWPZXcyQl5DO58OQTp2hoXPlKNNDVIzaCWI2vMag4kXNnYcO/kMvpH3luxkDg
HRzDwKzcUdOYahkJeMEIHjJCCNYQr/v7an+LY/kIHt4MRZ2WtUlbrhWoLKj7oIv0gwEBgb33b4KV
MoDXfwWGvekI8MURaHExu0fu5rZtXff1na7wV0sXV7RLi15f4GqG9YxyIsCG9SG7SPJfo1WfGsE4
BxSvaeXsf7FH3dRIH8wWcjFjkgxBP80ZYmkuLY3fcbGYe3iB6AnKHVFsJIIdcWaReia/hIe47iZy
dobwM1RwIZceLM7ata5Pa3mzMxi2igd3w4XsEL5upldUAvArFSo8r2yYa8ROgZl/5y8w/TCZCPlk
KbW4r1OaWEkxYRsVyZmunI+VeISH29KBpJMeAkqw4nYumLGVeY3X1YEmolCBly6Lf0I1b0yuYS3N
jXRcQHB1GY8sqKnJ+p/BCu59wK/ynuiw41UTYGXSc8U6sgy6dOKtchQsLo5rNuuJRk95Sj7bDc3X
Gejq4o1U2CQMRuX/Zx2EGLsyG/1sx5AiwdCWpE446/+j9pQyRpnmxDtJ+iNBuFS5vWeiME/YaAlE
JAHFQ6dJR7oPCMso2pV9lGq6a9VTQ0LH0/ofTK+NPZERFhhqwKSrk6zpXj80h45rDm2MAPrD2bKM
u48VDmG53o01QyWe6+g7tuQlhGUUmTcKNkmrqsD/GLDhyXGe3oRDzXcsVxYx+VkeXPRpaDZrJrtV
w0ITQT9QZBsP2aOG4NVSc9b5B867sWBt+uKxcHDZ5I3yIPbhwL6Wck61V9M5zRUu7HIMQnfYpncK
ZGEqcc+7zqvOSzLZvFUcAVWbkAuV3/uaSUthMu0RqCHiiDtCKHUlwAGbbHIUwuWBfyRZH35I1G8x
25WaKWKhCJv1ef546uunw+bLhJhLO5+FC6CVGN/rreypflgewj1u+F8SRd5GJ9FtklE9aYmlbbMo
NkkIMKCNts86fYS1dq8zy5YGJpvf3gw11/ZIr5QgGNpAXGmWhf5iM32c9LKJQ4+z4OgprbcMQ8PC
5VcZEZ7FojwVzCiZPpugYLaxONvxy9ux9RasmB1XxL5ZEy7eHx6A6cxgU6iV3uGqK1h4Wuspfa2w
DCXtqIg6xq9KXruXloA7ujjBuksd941eUePhTeF9rRYaa9kAiUe4355iKLd6SFJMw68L8NnxArGa
KGS3005X/4XZcLSsl7VS8uPwY5Oj34KK478OG0dmlXjRXsyz2YfUkSYwWaWLH5nCN2bNoCY2fVGh
4o0PQevhbUe5DVtI3WOJN2jshS6rsLzowJy/SCKRd9IgOju5y22WtUK8hwc/awPcK/0d1BlQqpHR
jb0G9Xrdt8J78v0e92CnLBQBd3eLPNBD7LLzLIOc95u5C8K+rbDsEVzSzWIFOHgQF3svLV+FhJwr
wTdzgWJwpgUdkinz/PZk2107N7NE//OhlKrEQneT6Ng8M5pinUugU0P3x017Jkb2as+K5ZS38K6N
AO2Fu0UYk10cEwySc9UjaUEBqn7TREfJZj6ea38duZAQaqrlzz2lhOeoYdkBVtubzPHE+o99nx3I
gpBc05IWIAQL3A4qMnxPK6ogyzEgalAhzbBCHS/YN9XAqq3AdR19SZ5bO5GO2gElpmlUSndt9UaS
nWIxn70wX3+R7lBZTtnxq0TaFEb/IKjhRASs53yfZx54u/pWjxbn7dQ6iK58NE5dA0eriSphJvIw
boLvx4VIRFN2QP8wa0dB6BLrVm6ur3t/ubZsFVi27Cf6cMjRVjxVcL3Omt5URE8wKrj/9qRDSuzr
rUg2Hey7RKpmkak8jYLUOkz7SiHoeSrqcFEf9jYLDXqRnINfNJN0rN5NWRluTaYM/fxovfTpebB7
aOOLaiWEoI6XwgrYSRzO5P2T0/TWhKxkpzdIkxhcwHKOh9VMSmoYNYxQTBV7glze3tG0hX4T7Jql
Y3n9FEuaC8VE4XXbVv92bdeHXT4RqjhfIySKGLIrsWMWkbyiki8IIzlpYuxA2rwU4awNss1xg1+f
TxSGEt6jzKtifM5fIhVkcnnnrnAqzuhc9NTWgeUjXbYqwAEFgolQ7uBSb1WDr/48NTTLeXT8xK05
+ffyxuX2w/n5+Ia0Sl9B8RR+dccUGrcp+xeentf/OqaYVvA4EAjW85amsFNPAC7T6XfYhhFp5BFX
Hr4L7SJT90gw8MwL0hkhXWtzOmbZqAnh1Lr9mfETcj5kuLY2tEaVbyOJy/SWDy3ltd285zDOZGBG
E4RTrf+ugEAUIUDRoVrIloEUAkQ/+k3jLpF3LXJrQ/UvOwS8riXAPokmUcSQiemFk88tnroz0WuH
Ehxw2JORm8NOZlb7QQeJPPPz0ATFhH2nM+918bYVquwrjwwCyuz/bFkhSjNg3cGfe6MAicqtCVi6
2RzVHhDaERCIIc7VCNmiu9Gaw8DFsWcl0qVzvf1toPNV+QkwnL3WRC9964YqajitU6UVODFTJwji
rnE3IlhjPMgC4pOdux7pbLYGiS9U4PNgJYuPJrMjq4vqf0BmgTS/uIUnyE9SP0hsItKHnd+vdi61
YCSidjDY84GXT/50FK+mhjExJ59aBJ0JzwpByWnjiVD7Y/7+GR93u/CFIoKCPnM+30HWb3JPNkym
k9bQ0f2GGS0acJ9GLPbrx9894d7wk5nFhbIBqpBzW2Zn38oULX+arNkA9YYqSNQeb2KFKXcpReCk
JWYf9b98n6BBmCg9SMYiKIpMc/b9p+A/t4dYc3pqVZ998n5XfM8b+9VwAWpWnEOKiodcsY8Spvi6
s90fsBwXQ9pVPERMbRMJn2NJ896+NrMRFeFOpyg8WSWhKeb+XR6aPWj6tuvYHW58WXboP9h3SedM
Yu29CO2q/AtF5HR5qegBPbI79dU6ylk7MHMlsZqIY92NX69ecINribqsFOfzHJ6BAWY3s+1id/Jc
RmYP+UNqFdjuokpXOCBXYRjFWRONIDc/fUF7gTZ7k7dDITzcCq9yMDoV9qpv2McitR1vVNwekLVG
oyXdNOt23ZMyfKRJKH84JQNwnqtxTxSzGydVhSKkhowiwtBEjRbQQELWxF1KxEXze16FlVUBqhA2
zp/OpI4Y4RWwjXgGttI2LhD6OgA0Mi+4JP+Cqi5fO53iVHn3C2JQYWvXCD3XEcFtfkb3/vO+5WmU
JwsX7Sdf4nK04+YHJkVGrdcrqWeMbVEFrdnkiDWLAT/A+5dhkfKfoVJpRkvD+Qc0sxIWyh2/8N7e
e9EfDkkbAg6xPYOtZcNfdHqno/UDkDlb5j4Qw9o/3lq2I1J0MPQVL6n7pWYNdC+AXBNLiJNaPklN
mHK3kUZR8oL+bOQlLdmYmSQlEAly0Hrl8ltXMGPDekSwlMPS4dXfILoOu/N649vUcFoAlQFSJYLt
ZxZKXavpeEaMxlxsX8I6aQvguK6hnxCxuHW2JtgTQVxHqu2TmiRl4PAJTFmXiGJOm31r4FT2K+XZ
32dL7zQGvQd2mcDfYkptKTUVvfE385ZjzXia540c3oRvRijOoi1N4MGe9odvGrJl+GPB/ingJfDz
ExhgA4Gg296b7CJ65oA1KBXVFinXV8U/sbD0BJv1tqcN26gfYB4R249TWNvBZW2tTO/q6/kh/vOJ
hrjY99loF4XBrQeCOVB91yCaGrgC1sohvQgD4XGxZbjeYtaHuAv8Kvnpa7mcJMz8HjZu/0XlG/Jy
NTiY4gammyeamgQ1xFsyxnPNzVIbK2xrV2yHW3+hhGRwiPGaUWiDHp7racdkmZ/ANdCpslQp0Ubc
7Qr3vVOuqMJaetACQbB8phL4UsvdTI/0bIkSHmFrCH4R/KIDlcSqMDw6bUaWeBikUPd1HUngCmWe
1aXx+hBAloaqRIk8qpi5VjeSE3tQCj7CkMeIK5ML2ZIX0HhjOpFFpy3mkKGwCbu5731ve4N389+r
mVksuzHhCX7gO8CI160Q7JO2P1c6ecPjQSpvbZQ57pki/Wm9yWfgf50OltgCs2UNyx0dL1C/WeID
p7as3ME0CpzQSggAe7fO3yF6VdWPi4P+8wi9bvk0ZzwbMfuHjKi7/SJWfzJaEVfGabiywecdVbn3
cAS+QUqnqkQpZy9uDgNrkzhMiYlvsSWl7MtiEoJQWbd4+60Ltj7pcKWdm8xANu93Is4r0/OYdQuV
c07uvnDzW2niCORZjUgkhgOP+4z8zpC3xwxaRO/IBAl9m4zXzboK8D8d2XOuOffSV/t016QcG4tN
5dBVcO+NbOg1r792rk5i/8Tqunmu1wrIzGMxbY92aFl0EcshYaRF7A9wpxOrIu0ThwrAMPPK4kt7
DMdB7OmJoYBOLxh9u0u70PVc7x824VCjb8Rg3AcyueC3u1hrfU6OB2BAKNi7eN+eaaDZbxnAkCAX
uH+WlpPtA9Omv0tpRsrwlNZ+nRSgQevH8eMI2cM6Fx5doqCNzkROmf1cNxux+FhKFWJuUHCi9JN/
8FsQm+4mZjR9Z73OIdTe2AxFZ0Xl1lNa6azBjNCxOj+LuEpZZ661GN4wxOowAOi552TYQJ0fk1LQ
gQMYrW/tkJe46+kwWkEConHhJdkB5JA9nQOIHDcVmB3FlyNFB7kWs161qN6ibWtrTF3ED4JHcR1f
GX1mC0HYcMpRX66XAOoLsag628GlvxIlm7A7NkkqAaUZwQDRoWDTj/P1l+qvgP0jCVC9CnF0asr1
BR6N+twEA5wA/Bg3pYaQeW8nKRdjaR5cOO/kGOlGnWkT46f2D6Vk8PrhfC4vAhzC2ImYfBa/dgQg
qxI0WOxX8/w/0Lzvs1vtsWun7m4Yv9cD0AktbYXS/CHfxn4anJHhh6OAxXaGBA7FHbzwyL2DOhVa
T50HFLYTn3Mq7//6qdJbvwa6KYDk2ZWRcDLOFiuiXqIvlhdjMX6j/Oq8uzoAbvnNzPysex//y0ke
hFi/mZnY1u3EBFJUYKffjv7+rVmJ0fG23An5H1Mii6mue82QEXm2FE7IlJI+maQ2R6Z3oaVjKFVr
l6HDTwo1DpSlhgipTYrxY9w5Xx304s1wkcuWKBoFkf2Uj3cmW/44I9AF/MSA9TflaaG4lD96Jj7i
H8KGdblwH8Sy0zzzCT8JTlxQRRpjF1oXtjoeBSHzu4tmccW7uGtFw3fjtXPld/HwLBHO5cWfjcH4
/pbF0j+xCFMDMkm/zPoUHErTE7+jS/c6ewzIbQrSqQWMtJkBy7x12xCRFHQG1ziurelznJbPLM8y
dA2czMjWJvDDV1BxvnvzmFiBJVWKfZItMC9p05FQlaezYGAGwTrsmeifWWP4osqWM4ppOFi7Tz3h
GQvazqoCkcZE5Ivr2VQU491k6EWU6qxJ67J0nbnyluYgNaKD/DTExux7L+CZdqD3BmIcOlmyoIYe
larJKuRv8yO5LLGoFXPP5W/NL5apX4lVMbBrjBNSappP/Ccbgk2rb4CiXF+aemTkTVbi52j9J4IA
Qdz+yUeG7qcLtPXqtGEVvi1G0dmd9MXxs+vOwkJDC35vP49eUeSjp2KBKyDq7rqQ6By7NwQEnowF
EIx/T4pVeZrFIdiUm//acMl9ECGV05VS1zEq1A9XK/TEFqCn2R8keMqvA8PqAhV39viMLNqF920P
NqACJmmZcMovJrHyzPn5jdLjNMJCQ8MwpxeXxRKuROPvzhKkx3dOzrLsP/dUeiQp0Yrs++Pu/fnG
Zk71ODUHtd2eFS0hKAHXqw2moIC5kXOvfwD/XY4be1FqN37b1/9hrsMWDFG49U2dSa1S7lNxr3km
dNxOIZ0Xz5Of8l63quwHrIefSvY2v20ixt1VZonppd5SM/hbZNCLtAdLH+l9JlVOUXiImeXGd8Rj
XLtjIeEzqnoyMzPRpUbPy/dSrQEOI/n93MBvozSCq1y7U8iVcc4umKoUzaFTogwP16Ps4g+8xGGw
Ep2zDauE7Ew8OutPkjhavW/kQuYQ58Nw4cmrSC2yrhKRRZmN2K321q2L6w7CI5U7IikKV2TvCPm2
9eA9niavxEI0jSVm/Z9GTGSqvpEno3wpmsWBzBNML3lhjGTHUFsb8ub3F0q27aByiZ9MiWmwI/F0
SzGtwAH0DlMZnj1hZs6lqpQTFu+Mrdc/YdmE4NnZklOIPYWQT3ofZXpQR4LgadoeVDtaqtxvSvOh
3V69JGizNDBYmTpgtLBu0SWWSPglQcyULCz7niXdwegteLWIbfZCm+LcSnwFy5B4GmznKLA1KLBq
BaCfRva2vzDFDOzX+e1XwQJQyA4l6zLabPNruRYuAjW7AQ+wxRbug8cOYibE1ZNEgYfI2QbyvwJt
Ah8XFln6eVORNuh4CGymcP4dTasJfRAinmgvTHy1flVlAZRNaLHubXpPraraSpGSCr6YwxMO0Um9
5/kid/Mu3amYaXFtBxkEx5FCc0GNSx6NBB0sQs+NNwma5QUf7lAIiRYarQWDWFdk+bG1miEo+NQI
y3jxApuHpWRzkNHZm3svJ2zPrEjNu12Py5yKb3fOI4LZEiSOKWiOPpQ2pwz0+KYmvVK7HHPk+yR4
MbYfLp3nmqoBHLM/YOb7rBgBF34RzY8h4oivgdxxcOPWjfo4u/TkqP9m3s7ChudGUEBfmQDDf158
9C6FOUz54afoFzpW/dwYVRKCKzXf6QBmNoe1GIiNSoTXRs8RdeGXINa2un+uXYGm+Oh766Cr1qmb
c3ddrldgnPPS7Ajhb5YUlvlKSKcevGJv5SgMg7HQJJRNL7YT42dyJkAxg9ZsxYO5O0ylzuYTcpXF
Ymk4d1w5uhj5nP6mheiy773fm76rSg7dF0Gz8wy0k2IzJv0ezUOgQYDwk87GWgUKsFseG5EKyiDQ
q6oWo8CUGbh9CaOGlGG19tlHtVakHGbOYYzNeE6crGaJSBP74yOekIt1Fiod7imWillMB/8Yv1kf
fsMRMX21KmrWNE/SEqcz14/vWnk3MnYH4jhkJQKCs9Nswdp6ltLYfuMhVRmRTzwrBsQOZFoyx+Cy
WQElcXbZgF3PdhgPdgFuDtt2/JF1RSxBIw7yn3blWJ/GSsATOlZE6RdhCmaD1pkNhbsQS0bsqNfn
T0u8qFc8GuVInBzjteObO5SqY5M6RIYtbKI8XsBF5vPbihHpFspKynSHrW8qnfRvU1dY0pIyFXca
UHVdi69B0m/64ZwtQKHpCTrkp33sMzxLPC6rS5aI/VL7SnCNaREK1RtmjlLgEo2Vu+eC9XH5NCap
dvx14bcEO/eCyaGRdHmrqqgYNav5mD+Ob/mlGpq5bwRqPJWRoCSOrriYz2l9Cb2L+/vbnc5h5PKP
VvoPMFBhB2qVGKJl+pnePgLMw5pp7Nrn39Psan/ab22kywHuwePTS9L84CTxjYjfF0tZgqoBEHie
A/QEWjEjK+iLEfipKoL/RY+ttgdXgVZMf/Fnn+OED/EyZyPiP442c6iDJtnqIjcJZ36j8WbZ2ulb
7A9n/oEbSJoRso2AhQa0HjN1ETrgfgaLOhKWIPdfGLF6lFiEWaBDkVkyx5UPC7td2XJf9RCrOfrD
G4lNCsfCid1nK4aSjIdTxjl5gYguGYN6yYRmUUho0Em2kEyT3iLG27ODKBcKFEQRDFaVGk6mqBqu
6KbFsxmO5fLrv6sBIxb62SeR3A27TYmElE4xB5n9ZgN7/P+TvClOUOgXY+Eh6DCcI09xoKnhdK15
pI3ESKYAeCMf0FoUcx6WAS2JQ3Vuqii3On5EjUt4yQIGyUeeZsXEqA93k36OqYZWKjb4weDvQzfv
gOkI3C+xfTYyufe4a2XsSoK/hLiTP1EYdycLJnm9VBf9/YTYLWdHhc8sHZIQOg3IoLK1ZMWJmEGu
9qjEovHxZ7cV7Qme742qmw30D0GSWJf6+ZfoTPviaOrz2VkLBdHUhcRlz9xmlwocvphBKLpucJk6
fh+m0yDJeyA+43hm6YehqGsSDGmuUwixviHi/VCES9cpguheffzxeicGQ8bmYUagimiJ5kJFNFzf
+wE87hq6aazz5eBZhcYkE8QKbWK+omCYMg1wpFmUHO+ny3pLa3rwzeiOVTtBaIflz0FuD28kYx8j
nwj/dB3HksQ56g2baBOo/Wt7mAsCSigV2/Ht7g2yw4GcymE6Griiy4Tl9GqvBKz7n3ia1ijiy8VU
5zcYRDqupWF6MwBNbk+snPCMZ2zlp2Zn4/rQGECwn6AzyhSHe0gh5SHijajsay+We7Jelg+B2gwi
pXj1kNvAlRwlnA4hroM2NRlBWxSEM/CPZALKoUNS8G6Hhcuqy9eKhaR7avKjxKEBEMEjYB+XG3NJ
mIngOi8JKB2zzZ986V23y3oQodrGxSuBIC3vxRHQ+VqDz3HCrz3Jx80B4qetZT2kViXnyLI+HmQ8
fkRSmSbp/LZKHvF2lR/NNvjZ4sex8alKKaF0CDRLnIilLHyq8p5tFt1yd7OQSHktRbpomxphJIuC
18OE+dYxSNW37WVGBp9gXEqaQte3QyBUG3I4oBboYT5xPQP7aTY+yaxHoCTwaraWFbD9t+nq136X
9i7EPs8TMSrxJ/r/ZX4Wy8pc8aDXOAf5KRVEBoh+rT9l5boRMzrx20se3CKzoUDAw/Ptab86Vs5K
uF2ukk8a3nHigI8OMHAivfE/6p051wJFo0Kd//r5hrTUcRRlY0RYsEtFsdyAFYJROVrhMkBTF7OQ
wU+F+BawS+Wh+CJ1Vnhg9UpAz7HDy/GQlz4xBIZFgdQq9Tsklp8U/Im/fD50DuTFb3/wKyOFnZpy
B6iZqK2UCweR/+RAnqDQhGHEawj5fsXCod2n8/bjL2qXtUZ9FONWnF0phPX9o4CGr884KLvx3GJ5
kQsMpbf64Vn8Mc53oLXEMaLBXzTrocFT3h0eW6DfnSflBNslH8dMtAGeHQ24en1ciOEUlXNWDElK
SLK6bMlfV1FCcHf4u5NHa5q5kAexwBWT0zKyLqVCTatVXIDan+000x137kKj7viPnrPtTAIeRmU1
AO3Nv94k5WBs/MKxUtmR2l2a6Lraob2Uuv+vHLJG8w4yIAt7MZVRjeB1+x1ntaTk0HfgX2uaP/4e
82J5c9mLfMF2zxT/RTY6BV3Zf0d+iW7W7egsh4+f5lAAKK1hLSOJ0a8Z6gcG+CFckkboBoWXwaCs
OnGLUk1liDoGtmcR/2rMIIiUb/IjWHYae+x5s1x5ovH1RfvzgeSa24CApZGdS/f+ZCwwDS/FpG2w
/0m/KfGijs3VXlUXIhj0dfqgOfO5O6qnqTGs0NoWHUubA028qd1b0ChVNkycElUIHNGJtYTiI2Um
ac1alLAMR5mZeTDIvESsNkKX47V8XUWCWLVhy3zIvL/EX4rEX4ZsGFEAW0I9GDN8cCLFNhFrDruE
8he2psLS9wZ+rFnFd8V+3YPApO9klGGqRcKn70J+vN+FGV43th52ylP9heFc5xfRZ8OsyhvURV/8
tbesulRD6KlSUlReh0V573vtPrqjfBv+sqyb2m348zI/mh02egR4j1hmEKBeJi1ZKv+uEiVS0q94
XF66tlYATU2M2olkkpCVVk53He3AfVC6slNyjMtTsTTOynaTBQ0k5vOthHoD3WAl57tBxo+dR7I1
8239ET9JxlEkUMsOHbNMyZvFfndQySnfm4GbP0MZ5xBifFE+QvmTCGdQACAywzklw20BwgFliS08
IpX7i/wMSTDcG1lKsAXmQe3+GrgbkqMWas7P46lU46IlDUJJYlVZFIs5+uJtiEhpUz3dJnrD4ddn
J9UK/fk0yz11e0SqR/TUDWANDWMvYlxhBE+gBxwHditTsi4FbI+h9TddyHtZnaCSp5hvRq962Ocf
Vn7aYKxwqsxg6SbjkwBRPirxK7IvPjZbNkyoo4l87A9xmoY+XF3rx7rDVKc3lpE2r/wdnA38UfZ2
wGn4jE9A5BcsLM1oEZf7pDZPb9A/+siRAd/fTIVQMpMxJMBYsMXE5y5djfx2x9mdYDuHID7zVRa8
IW5lZQdhRpgrmK8zqvJZHr4mqD23sUDFWhayhFKfNXyXXqRsFTKqYH9GLlSdikKQGB9TV2NzT+jR
qfG1Zq/GUthAU7ussKno8fU/1bINsCal5kUmZlBGeBv+ayDY0ErBo4JEBheHM4StjNEM93jreFQv
zy5I5aYWDJhJ5mYOvTDCyE11W0dr5k2+O4QBSd7NF3CW132Hn8ld9GHihQLtXahsweVFVm/IQ8wH
zheVC3Gu15PVil7fpDWPJ1qJTm6Tm/Wn3IjGN1MbW3r/SY3Euu+jAYUJ9r91Llvs4wQ7knJhvJoY
sT0s/sdoUPAYH2X6kNV3T+N7pkzN8oaPGW4/eaQ/ezw5vyF4rh803z2hiNhk8hjKtFsZZoJT23WS
leeCGegOgXklPoWo0FGcq2CDWfinvGmqebxiQDr4yP4nxMuMglUG+pVlUrmsE2HzV0tjQkUP+0m8
qyVAqp2AEySotm0bO9Ph4EhuIhcsKmgHephgBY0+13WKB4H4fKPfkTLboYwDvJKVG1t4mKeB0i0r
1JyNUFKFLwUhTF5GCx6NfEhrYRUF4F4uezn2S9M0VwuUC9SlK1jF71rUdKmCZKaJYLs3UyQFbqaR
EZJXgu2aHFTXFrgjOZrget8KCCq1BzgmYH4L6fwGHYV9LVTm3BN4eobTRp4q7qcpZCLwpy7K/c5B
MQ+2+zJbF/aFlNddzdL6Q2AAvKj5whimeavKqt9dyPVANSCr39m8xHTLzRQJoegcvVOnwVb7QAED
nhPFO/ulNVk5L0Us2XFZe3sTld9aanpNy223D9hPeh3qOmuzahcdyydGyInzHl1E5I4qOTe3CgVa
ELYEb1Q8yMB83qO2Cal4rF950k6+p33LbjM2Hqh3y1XSxOq4aN2am8n/B++/QeKg2yhwIDoqwcpe
9pziL0VQ1tUDpNOHTA8egOQ7Ls5T52XIqyCQ+2ccU8Uxh7+Wcoptuol1d+00oGXS3JMhx8sEKo63
IlhQiR7xxGk4FwpobWjYqPths+x9cXEor34RJMg65flYKvJDgVBLzJr/Oj6Esv1RPApOOZeYqxUd
vJ4FktM7mmeThazWD3dqdhjq9F0nI9nBPEDrqgz3isl+f8XzRVraNbfbanS0r9DyTbVMBbWpp38N
JwMPY6Qn/K73/4+39ztcUVE4sLozLlQMfAg8cJ8Jer8hU3cSeke9Cmk0ozmZXMf/t5w5A9a8FmNb
DNnJgoX3yUfwXSB7jR2o4IVLIO9plZEv9SUquhXH4F51jlv0d6nisBMBo/Ob966K3ntJTdlL2IwN
qMxldduJO/62Bm2TjB8iz3ZQYlQEAbDsr39mFw7dG33huwOaXcTSIM5GmmzxLP7U+mUD3LzyVyBP
QkfdPsknurIR5mIFeBHxXts911XV58uORzu2pc9uKN8p5V8EXRoUPtuwQCwqJlzBHj6tj1pHJHNF
yTJFQJiona92QMizkA7o3aZhDNTaHzLp11+dN7NKSaV2U0yxEk6uvpxgeIGESOHbmdFBv5/llauQ
IZ/CH5x3tNXWXugi8xR7YdMX+Ak4tFrBXuz2b1VHs1mhd/cx4F+RF+QH1ocu4GJw9+/PL2pNQIER
ip3SpLLbhadG5V3j/pwoCY/S5lbte43VWdh/llrZ3Kjb9k/82gzJLDFf69ONlXA8j5Hic3pWT5/8
8Sjtir1lb62XduI1PSYwzvg2lXl6hF9Jh/Bptr9+g1qd6sqF1W2pThW/uMP8nGzBlxwktC0v93fC
1fxOJ53l9H21OXtLu2VFsiai2qdnBLAemDLLMatG5HJtUG9ndW7IC9PVmCa4kCpLseP1sYZaHk5t
yPcbotrzVy6kx7co6sH9vKzDy6ktjJAgomyjy19SlzxiIXQEwRZGqIhDe1kb0LqWHfvhIaLNmGIA
fx0Op97eTKzgpz7abiEeQZZC+khn4ZHKtKtFKOCP4euE7fPTi0V0qMZGNi1fffEFIiWxHxjaXyQX
0OK1AtK1BhqJOGtmZxJZbg7QtyqHAJlls4ch2hwMubWqtLNP2mIl3vVb38ZJJpHmDjO0komZbwaP
Nf4ZRnzLs9kjFZ2ESKykICyPxpG2D4bTQBDHTSlU2Y1gwgeqGfu606Le6rhGvbTWUWrHURbtOlaL
sFK+YTODG9Od8VZWOFpLz8i0xyBh6dme3vua5MfMNsq3rD2As89qRRSI0fxWzpVN0ZGzdkGy6bsy
qLxXjEqK6P0eNFc4KaX/a11Jwp2yQ7rgbJ9OKo+H0PR0lbuJUyFkRQTKvmjBiLSsuCsYVhgAZ2O0
PA0D0C21oiS9aKGr1VO/SkXZmjqoYqKVpAnOlGcDZV+MDfZTcJhvsmzuyrQVTnt8vxHjngzFKJKj
Y/U5oZrrRs+iSjrLDOJZ1k8AK31Z3EkX6g+5GVVHqQJovZjtGVuvkrDhCJSX0ejVwc8JRAxTkc8W
s9bb6219MT+wfvpo8JkcACP+2NFl764k6mAwaTVNI5a3ltD6GJ6DQF1wdwCN4PpAIuo8lyipp4ZS
lhvlZqDVwfyPQuxktpnl5eVPFaUTJkDEEpSgScU0hZWMiC2JWrVxKUEgo8y5hns4PQgzsCgRk+Sr
iV8BBtcx2oF0fCxbie49DGSqIftD+uBY0F+sttePa6m/so4BBP0jHglqdhmBhSBCHd8n7NiKT8uY
uFMALctF5bOqfUACOXc0BK1a4VSCbR0WlUcf/6oMIVyO9QGA2DuXzO8ab2jW0qE7FVBzhL5xJ3pd
juVNvAso70ED1+TPukCAUUL9vsWBqxDIK7dlQ3F8r3gBkqLmS77vjmpSDirWs0KNcG94/mEMdLKE
IZygQddrK61qBjSTTkrTWXCpgGQmrf6rELqU9UpDsmxURpv7fyBTwtMWp+ZDz3fnnvrxPQH0y2Zj
Z4g+JFd3NmtL+VfO8xMdSMf3mRZe0cVnTEolD0oYQd/XePpwjYUEm9kNMnAGbwkNsymEO9kbSjIY
iwKY9BgvIoHu40b6Kx65eY1jBvLtR9pnWkJAoQtZ+MYCStlv9adE/aC/2J09abfwkD7aON0uTQjC
LxO1jVq6PKMesHEqanhYPA1T1z35mX6LXBe1haHJsugzL4Z9bsSUdCJ1A13stTLr/eEpSbAnLux2
vcXFUMHVUQyTjnm75qI/0Vixd/HokOEcp5e6rf/u9bXPioBnNRylPT2015Ajw8sRvBwiooGL7wtq
KDLUuSpJAFAcmImwTMy6hDBMbQSTiI2yCQV+6cqDsrSOCSCHTrKmzBPXNHFBw5RUZ9pu8cJrZVtI
8Zy/AKFz1O1q5vqhOSWOVENH3pDBObaXL31ujcvoEKcKoj3I3bi/GmRQOMQdPgWKHOtPSg2TTdbq
2wuFPoH4/ejx/mucEy5q5Y0g75j5c9GU972DTJI6t3qO2Tdkqa/oRk/2oDH330t43ugHP1wCoaho
JtIbJhYXAvU6OqPSImGftnPTgiIJhxGE2QY9DLRPc9I8v1imI5luTgnucQiqymAevuEolsCdhPEd
3dS2rN8Ip6f/DXqhfTJmCt+12BCTgqKj9J3alPHCsRKdNBn1tlCWiqnUKK+142cAA72DNn2jTDEe
kkE5KPtz5MZRX9quJ7zMCsRh9lpvmSViHjMVX+QT/9vl9B0Dp9tIIKW+1eM3gBbYq4MwqNPxmnOG
iUCwzuFDSr0EaDSmUI4hKScfgibSzTNhZgYTGcIsPtvWv7pzMK0Rjs8iyFdYq8kb//49s74eiWvw
91TgQ950oIEJ3pMQmGJaEO0Ej86VhLAdwrr2aUWwFDnH7FSeDxcSc93LrB6fkzJqlyQa4TvcxtSg
7AuvmynnQz0FINp/oS9B7J/vXFmcVciNjhpzzwma6qVamKUkvVlogt5DV0IP5h/2rgcfn9poquM/
dPtesCa2xNnSb2e4zIT9yV3VeJWf+gHSC97yqPRMg4poPSVO45WHDkqD5OLyVN23gI+/PgNKtzWh
1M0wk92eC+XCH7fXhJ2BFvXrZBesF7DTGLGX/D3qpa8PcwAne5nUOhaamJodwTSd7eMf86oyyDUB
y+kWHXioAQFf9yXQ7r+KaHjNhWSlz1HtzBzRIN22CLGyzEs5fY82x0V4T6s1K24El6ismuv5qYEX
FsqOsgFRWqxZb971Vty2DFR7a8+93gdm4F3DU2waH1HBfd8ooAD9Glf3DK1tpfuxTT0xVI3NekbL
f/4VlX5/KLI+PMVDa4MSjPW5xlIS9Zy5UIDy7GeX05xlHBuxorpN5IkP3tSIbtx9xcnAgn45P+XF
yHgr1PErVtvhrwo8gqYKQ8yKzTR6yBSasrkrkFirDOotzfOM9GMqf94KcKFTIfoZV9c2Qnl4RluU
GW+HE+QgQJGxUZLM9hyUo0J7hjClDuWG3+zo8MAm13bFhJEZ0pu/uuYPjcgUFGd8vrmoPIdfwlPH
bGzwmCidQzGkTzgI+iC+2mEEGFjfk6z+eEuIV/mxCbhM6imAlhSeTm0/xUwNkc70NyB/hLbiSsSp
+h4naxsUAEW7TkpH6nNdeJpyjrHsoZfjeJrfHPW47WyXDRY9XVrghlN+rK7P1xQuQoJja5HG0/Ac
Dy9zveddLp3/SHaVFEnmtV9NY3g2rE/Fm/6Fx9p9ECMIk4mqcvDR8FfTZgEamq5LRyR1DDnHTJ3k
1AkvSpnDWM3TfFeT4hdm8sYIYGEhUGLRKkpTMytXQVPtdqzo873l4QywhJS3AhTK8QHcCRMTGaj0
IrzzyFCX0JI6zkA/Qrop5MCIDMFImv59i4GJBA1ael58hTXyqydLJaK8D1xp+O4E/STN1zAvdbzk
J3NRAlYVyg7K7fIOZ4+/RurFnlsh21Cjc1tWeaJGTW1GtjQCaCOWUK9QbJw4kTZDSeEFFbi8YFmZ
D74ruEgP4LLElvJXm+fFKQbucS6WCkRHIx9DRix6r0kGiFb/aU0xmQBOVlQ0Zj3CpN7B7YUoQ9Sl
blNKxUDHMOezAxcJBpvdyBNtgupLRELfRwtNNkaFdp5gTyUZbKntMSSlMQCZl0W0DXleb1epL43D
Ngiuy40Xm2AFEoWpNKphikIqoiMQ0XM+hqUV+HOxIMlWd/4K3BlkImrX/df/vUK2PO1iueU7JVAv
4LZqSDWO5+jrZXUTHJHCMZkzKaTYxk/LUs3LykWZAfEfYv7dXyvOXpMja3q1izTkDGwl7xDGUU1C
ooCUnlwQtK0WYudoKdt3/ttjOoNszCl3Ogdiw7jRP2JuVOGS1vbjMeEa5/rneo+zHk2MQhzrgDs5
dJUxG6PQGeNYwsbNqAIn7t5fUnkG5p88+pKHTyk7G+rjeCMPvJN6t15lJeGaFpsu3yHQTe5q4zHu
efR13yrH2CC5/LaY9JeRz9BPDFXqFX6RvBK28OE+KWTRyMy0msKIlWdhI93Il+xjqfxETFynn7Pg
RZrDXQSrkyap9yvLL+Gp1cNpABbqLDmauudSLukNQlP3cwSHmGdv1Rr/rEbFWImrSMVR6s14xpT/
A+oZ/hnoG45WLHBCoVJd9zDBuFBDJmZd9YPHhnO5Y/dcXdEy273/BL5VE5utSLALt/LT4t16Xfk8
yXQpZgkpQPAUSJpYb80wwcUJceTWK1NpoV/tXfjeBqrrLMJSnX9Kc1O8BSQW8p5WhAylLHXFWG37
I3hxppP9D3okC/9titxOmd4wPGOYypeNNA2YGxmTa9IMrGtm0EAv4zxaHNlytqzCZ6JQcL9jxXFR
KEaraFIzCjcNVtM9tLRIwU/FBfdo9kg4GpC53d2K9pwDr3jYC/8zEbpptarTsWSzWcwM95m6OXlN
R82tQQy7aVWsvPOd/0bK+MAapzxYhbhZWc0wNkZTsMzetPLSBAJ1q5L/LQeNd0irIAq0dN6AXmRL
3QKHHyOtJrBBlAxAPfrDoli6cXVHY7T7BuJOh3vicAhFswcfVCpyabVkUdxfZdNdJaOERtcSid2L
WhcU0op1HJ05ulekxspsEZtvwZfqqZ04u1zFrzhBkb0H5Cy2NRGSjnubu9VBgBTEPOxNK6s0Ngut
KT+ZTLuFrlz4BDiWnjJW1cn+yuD09x2Mng1bufDodQIY/Tggz8Zg+1xWApHBQPITCTv74T2ZBEZI
sso+RpjPsVS0xb46UjE/4y5H8W9TrxhZIAC6TEdaujDY5WBL6JutUAh+Kiw+/MW0b6px8/YXHKly
XpRvy+SjzULo8hrr7c7+4D0cGufvZjKsx1zMc/nC2cuNfkDE8YTCgDIll0Vp3cbnZgYvYjABG7RQ
CAKAeJ5V6KwY6yJx2PNKw6z7WB9/ALXadDHPqiUvpeTn4NV6ZlIVFSyhRPijGhQP/7Rd54qXOH6g
7DOb/BPDYbK0cdNuzBKLVnw1sVrAjYNtpPN9grAsnw29citd5NHeeOzHntBYCiHov8ns0j3NoTGn
7nRgRuZbXHDBYwYoFl8txLn8IvnwUU3vQDSpDGzBmUgvyMSTbnG7udgw+taJ+NP6QHpzepPyUZKb
S3gwyGxgan+tTsGBrwZ09bJ/oNASgJk9x3S8mjTGJpHPuCqzJPyLvNBCkbujcMinh50w8xDcduIS
vxts5fJ8QwZUpUHlJ8HpLzQi8MnrkgSTL8A3E3xj8a5QaPiBYoKO11G7t5vJoOSpUvTyZT55cH2h
jH6JhB160sP9BnmFo2lU21Yrpw1ALMWPUUacRLwG98Xd6FQSxQgjYJ+Tj3BQ6cm0HU7jbAKDcMo/
HZUpoJruYlMOWSMJMVdC+Kvn02XJEtgB4+ApaAK3HWo0ynXix2T8AVX+5gOGB1csfO4uBnXlmNgV
mLxuPakeOOXtfY+Z3matxbMNgR+KKAJgLrVhVRUUVVV2tnmBR0M4YBte9fbF3KmhcdpLOBBAzGEZ
wx9yOTBIS4VuTUVCwbHPHRXXZzHP2vXNdLDnzb81wtgo0NwYWX2O14C+yPkiwLuKZiyRP8ioGM1b
7bqCbnz4IBT9NEuKDR/pDQkorTdLvOuhKAcR5Tc6wwA/xQmY5LmwFNcDpLHvaL76k8tnaLN+uS+R
fWsCcKqP+1jWqaG4l2UdBKS+tNzql2mZLs7ECkT1ysDB4NqjRvZ6m0VRNbbVf7DHZD24oCGWaMfs
N0YP1PIVAxEa8GGBPyij8ghHo8mOgs7IIIm85f0+p9Gw4Hdr8yLyzQK+57kQSV/BVJ1e3bcF4CrE
9MlAMpmeH/HVrWniPtVmO9uUsBHPQ9Tglgjf8iVsDkCdh0OsGrR2USCSF1TgCMsrtrbdhjQJ0sIH
wRnbc9Bpxacd4KzihbJgxShM7vhSzRWdVQHeD292rmLN9xYP3ujv9OLnAKu/nVuWxOxeIQC3gB32
UbQCvJcnDj6ZwKjrm5/xVuLNZBQrIXxuqpnTfj3ynZDZHS7f0V+2tyil773Vle9T8KEt/n4q2zdL
+cgQhAE1D2TPxT5UMUxbOuFoJD2LUU3gZwXMuqJJkKNEDsgbdQb2oxdRt2WL+3c/TFRl13/ZWG7s
6RnORCsZiKuozwv0i+53ZDoW8SZsU4F7uVQPRttYE1ySkeZToHpwsQh4NQ4MH9e56GXhkQnlQ52P
kJOin3lK/I6zlFfqLzGet6JO2M/d86HI2Q9gJb3GmDSU+ZyDQejgN98RecaYuzxfvEwZKaAGIfdR
TNsWV7h3mleBnaNYj3/wMK520m0s1bERZFtJLZMcNYq48ZGPO7H+MbaMjPo3SD9cI5RkZlqNljcX
yTfbhJEGT/2YyZnv5Jwn1pAzFFau2AJpKHX/tjp02CA233McqRIgjLjFKt6I/GfN1bi082/mcj0x
aqC/wWyPZ1APFfphJsHjfXmo90ezhXVb7W1iMTm6tcdeNMisYowHXIf5uQYqTRGGg7kkyiItl97D
mt6oZXwKw35LKHlyP6m+MIhBVoAerojmxRsb4aUEWnTzyWPku+6RLFfYm4J9wdjrJyGxFlOUO+iK
6g+s5FwDTeG7wBudVSsrIT2u4rpZPq12jRWanUbcfhnIwb7nkMoWR73OQor2x0AEEMqEZlfKwq4g
wYock8oetZ8wm89iFvo5SO9Z+Kc4bAyh0POb21jVk9RXJOowQKlRbigcNUhmxH/mvE0YI6CpgoRS
lymzvQ9JNbBpsZcxJGnny5ENYVALy+OaqjyWCzhPhCrcL7MgwSLX7Y0o5PUzt0jI6xCCC+yvwGvX
yOtTMpcpAHNivj5iHQ0/7LV4C+4ajuDAba3ApQ1JXr223vw97qut3aw/qvgPEAKZc7uPGnuz73kq
74fuBMphbRCZ9ZQscLEy8dOT7cz8t9kqUFumbu7il3IBCJAszb9FRhMYuCHRkmMgpJRrpBiPQ2QW
lmCMn8PgnlmOHVrrXPv1k8HqaNh6J2MEbeFuSxHa5TfpM4wX45ISxCFXSzDKekDBUGaPsooztQ2y
QwsEPGNuDI1zH9syeCvi/qRxbwrKoKdSCNffSN+fPxOewlhilbVCEAbLNg93AwdguojyDrdehUfZ
2Y/Gs0KDVfOBsDK1YTzhC5J2GNXg4PWBNMIC4XyIuvoLeu3jdX6Yb1FYc8nq26v/pnWrNlAMUEzG
UCg4B38HCYxqzUnlt8ml2pHL9tu6df/YZUS6PDZMW45F4wBGD3Xs+Q4MJJUseHpERV+beyyqyThv
JqUqu5j1KgWJEZOVOeD0Zcilt16ALRgDNEqIEewcEVy1Q6DSuu1zhskt7O1g9mUPtGER9TZfifQK
P908p3i+w5Svzt8cGzogKU1/K50njFkcVHYs/hBCFql7xEuOav51Gh1TbjPOpv1UDHqRUnzb5HfH
sezUQ6x0J+0fGK0uYAZGdtAKlc0EAindlxhgDL4Mlgpd0S13/witEotvdQ/ohbRB9U3mnD/DL+WO
1WccyX0l8h1/SakMK1EH3O2IvNX21r2ayllN1WamniVuGohdgP9P9W4nargUYOwhLRF/dSttUccV
j1kPlUMcoBkLBy3MV0e8XL+KBknKCRj3DhSO4p13UP0RWQbaIVqyrHB7Mtv7hayqtoPGg25ktT3a
YAJrYVd1uZmLX0yvWsQYAFAB8Y/5rabbf58zWFrKby/aPgWU3Z3v/QNEYj2AHM30a+wK77U3XZjF
zLw2WGPfzgveHguV+J9IF4f+kgbGagsH3V7EMiInbAPjLrGDx90lmdy9ozhhr3BD3OfMpaW51Tk9
qqlO06yVMWgEjhicHtBYlFFkriHb2rZI7O8q2nhCrpo1dEFxoSr/Ur8qV8S5nTvrLzWlKREX2S1v
1lZxUku4aK3JLyHIGhtT7ECAWqT5sRURaOehN/8TFWXkiQDRmTcWP/ZxA/eBp7tx1tujCXYNC5dK
2Xueh308FvcgPLT6b74eK7ccXQ9G0hJs3OkMQxc4kDGwjVtuoKJYsxd/ofbIOQe+ELbZLs/OxEJn
c8A4Q0bK1iT5mjt8bUxJLpK8QuOOv45xjnhO3gwOixQa3qsHUcJCetC8u0C4tSq8zAqkT4WVFT05
qTA/5FDCJfT6SABeLcP8T+kK2Jq8G/NW5EF/ZyP5xLOrUQaQ+atiDNtSDMWUKMvazmWdLZsLC388
pn5FYobe460+LYoRAIHcymxvLHtmR2O8TevCGikLVzsZtKn47lfk5cmf33CG6+d/kKsOZBNXtaWw
aLqZ9Tgfm6eXh4pbSJhyALitAis4+cqb8lzvf5rtBq7W62mhiKuW3s33niYVuD/8YoOHjy/sbJNj
mVSHCRdBy+I0KuGHeddeXlS8xTlhShFfacRjYi4k9tAZRFhmdrSWcQMtB477Uqei42DmqALs5iz9
QhANud99jEZXLFDF/64FLSyGbgom4PwMp09zzrNgLs5kMGTn16NI2pXCTKo/uWuZCU98hVWdFnoW
XNdoPmDYbYzq4t4RjzQpLaJvRJtAyI34gO8YtKHLMIF2aCqJsLwltzlzDcYXcjBitL2UMr3TYrWd
v59QBN2SDhHRrDZ6XDixhWUNDnAojq3LIpDjScwWZBCSH1wraj7eMhMSpm4vT/sxLddI5rRRey5f
9+yZAfoa73Arwr/xhyLfPjZq9M1yncjVGtqLvDUHX6d/BR/6onFLGeLqG4gu4SPcZmHcJFxFU25R
hzCnKaytmYuM20X5bLPL35FbmdyyrV/K1ocPqBktWYF1/+z2WJBCpLxfIgxWbmU/hqBqhvWRZ0eN
q3D142e+7le2bj5c24EyPivklSDSFvzqccHVZ3LeVkuUefgoc66qwe0oFpWsBmeZbjOYF8zBxEOT
pWDsqB4Twmr+oQ2ebwJZeq0+hRoCQ+RcCL7KIOhvPMrNZxwkYIRhgt7f4/G+xwMkMUu+XxqIiZjs
Abt/4Uf5lu2mMIPaFZKakmblcCVcwJMA20i6JJXIsIkAzW89bK/FzMntKXeZ77xivaEBjBug/D6k
R8Qn1gRMxuQt/4tmQGgxHG4a8uufBdGMeWj82YSAmsMf+gnYr0BJylH6EZd4Qi+LXvJHiGgG/yME
XZkZ9G87TKwzfp2rr3EdbyD8ARvAcgm1XswOGmABTWRcZNVgy5PEM5mvhOBw46EhFyzVx5Dm5dAx
RFUMV4hrBKPky4ebwbbyqYT9oxM27xNmz7qL/W83twbelF1JtFv06ZLSJQxzrOFZRMpP1ov1jYp7
zoaHG4ATLb91ZJeqGZrUh7xBALUDbZk4BdYvAYyVZ64dbB8RW8okH64OQPey4G+pylR9M0ndllHI
sU5KWkRtj7aLonXdUv5KMimPdyjhJ7Ew1fuO6dwSCr9IZwfSeF0uBeNee0YdzjnpY9XMXhkFjqHY
yUrbfCQORbDdX30l1zKk/JP1fPRVtY/vsSvvpNXA3MffH51GK5girO2+eG9PnVPIv/FoRtAZ1Ofi
x5xfEF/aayRN1OnsED9uAILXVztADeUaOawMPOYEaFfSSLc5cOpJQvc5Zh343yItEVhsJzZZ15Rh
z37iGzblJ3qPa72eKB02cMQkI8sHNTtcBeOqrhjT6PEDAQTp9RzzUWcikvdvNounbZz08wcunKIL
TYoe1v65BvrROapbjkW0IkG+B5LpKR6bxpMkFlQzoz5nO9nW6fZHdw8pM/dZA0IPcxInRJDktQzp
fe6oFVba9IcbgNG80pdT/n93/h6+AkvftCT+wP3auobp3inCJJ45YP5UepzwsY3h4DS+T39oXisl
DA64C+r9h92ZN1yJ1fKXLnBUrs+cRX6IVTb7BSUV0uczVR0rH/PPT/vnhT5spcWI6JH2q1ND0Z36
TBY3Pt4eggSmNaKdslVZGyvZhRixnR6ogym0OuGYAJlQUJu0PhYuQxTgBxAXwjjN9J5ECpad1c25
W7Lb2gPAsYvt0PwpAPn8xKqMoamxAZNpRFocAGBpRjv4fqdt2PXfE3Pdb5FOgbPJmpixTalnTirc
hOeYVwPiQTRjLGhfB93TkbVDHvqVHbrjiIdYjFZZk7uf96HVblzvjVZatAxW1q1AYw6f45F5rgco
fYQrS9MkkuItcYkjIglV9LtiWXtA91H8E56Tvad2kXp0gJuiO6atGdLfsbngl0DLZVGpUnO8NG5s
pJpD3k6s7VA1TI/+0o8/scJsnabMeR/S97K7zky/YG/wlUIcNFT/8inZfc7Qmfsb0Oi4YXFEB2ug
Lodfu/9GD81NkSv6a3ep3PAcpI6xg76XxczLhbCmTneFBMOVJ/Zdb7+q4OmeC5COb4zjRZPD8eTw
ECukHzYq6ZsB5sV5YlJx8ZlDliVD/l49rwRacNou9GwIJn0ESLS47n6bfj5dYas6HzrsPAd+IF8w
IQpMPkZmyY4DUGLhyL5V072wFoT31fmi7O9Z98Dgz5jcbuC+Pzkwqgcpt2NKDKaI62V9Ylv/Eqh6
ikBuRxFYn2QwsuY1ZxQNVFR49T0Sc5LvzHMwwXZyPcPFrnJJx0H2OquuK2ccJ7OFcQiMR356C0ap
UMFCJWFxI55qddhIDcbViy17uLPGQqGmsiMn3BpC2Twzpou+TaFaOBR07xpw2MfzywTEIlU1Zhef
DuVXiDGwiyNFduvnr0Y2Zy/f2arl/9HPE/XkU81iJK5cmANrN8WSjNEpTPcli6dB7CYxCzm5Fhdp
o8LT3gfBlUBJ+N/ZYBHW3bdYOvF1/9i0HeI9vXTYeXhDOT7xgnJqN9Y+rhFz/l4BysPgvFzI+8PB
HTqS0cdNQuZUEz16ZdKom6+YvUeJJQpO/oOjIOzuRG5SGR1S2wA3ci+PcRv16vm7iEDnbVsTnl0k
9KBY+C1FZ+O8g2liwQLk1ieWFELJXwqI8iW71TPLhJWsuNV1liu0oKtznlc6eaSA9Ug6Vb1sIbtc
G1A6Bx/izK/qejnqflJ8q5Blqd5oPFStb2XZMVW3jzO5k9SUVVC4CEZzqWaLtDO1a/buC/ndOAd3
2EBRKfV42LZ282SmNpJWTCdQmkSJAexCxaAbXiB5fN9vcUwKcNt02m3gPnuR7VvGU8oOwQhUwnL7
cUicqqGbFqS98u/Uw5XG1wVONJjYToRCqP6m0SyPIZCIP9q35MiFmSqEf7gtPaggC/9/jsBPdPzi
UfqsuESUEeaWEzPPJKW5YUjG2y4zOmKi6M454CXzjOF4XD5X2XH2M+Gp9lkM3bT2LKonqE7WUEtr
3nOoEFArECtXufAhDD0Dl0U4i9QQt7OhnvyD+AdWS+O82oQzGphrLsKanx+gVYGm9NvrxJQGILZX
KZQU5Hf3Z3d5hI2ZTCo/zdoTGg6jDKBEFAXhU98bm5EHhUHB0mTPpurOUlgDEpICoLmF7xYveKtH
vdcDI582fDM3mWoFoH7/kKzYLCDy/xIlNkYnMyuh1BQx/MOactGP2yGLCtsijsxFyXiP4rRiVirQ
ZSQTlAFw+YCcf9PnYZIirRTHlvP64JFK9x64ELZvMGCMzLEsnCowd6alx53O6g02T9QJQkmG9V7m
ddRTBVUMKcBkuMryJNd8//ewrPZo3b49fKFiKarl1IT8z1At78ZYBf8ugQDY9v39v3U6YaggIkN7
3K1BL1YtQAz0nm62dTOsRWnlhiztntbK+EYcR/MALToN9Hjbln+UhAdMSRbjiTklUMkTgu9Qq92+
cu+5WQqGO8d4TeOUtbWiOn4y8LTOv/TWtImdvLunBI3jvlrStzmOuqCDICuXx2SDZPYM+7+/E/CE
kq4JZ6dqjugZbC/ownD0W06DwSdiOupbIEFSRBTwNufHthObcB9KXd0WAI5CGjxjDLiPFAEJQQT+
YQ7TFqcV//Y+ZgVvZb2E3LibgzaisDizB5759WiJ4PQtAzw01021Dmrwqv7nsPjCh2h5TxW4d6qc
VsoGEuM+blwaJGMZqfUQJ0eaXwqRMrnZq0byTMMRVAszGovcafJcFGkDlRge/ToaFbIaQIivbz56
63b8vlQ9Wf3j52xfd2yFVhBLWKLQYPmb6+TVxJBvsyJhHIZ2q0P8tro6iAky1N1c6Jq8yqk5PW71
PUx0uR98l0RgRA/Qr8HKF5Ba+b3JlPA1gqyK61JBaipCqlVqq8lzWjQYL5eXwCWusIQX62MOWEaz
yO59KFN1s1RBYT3LrthEKlQ9EZQVsymYoxwfFU37Y1CcgQKkdftt6kac9TGaC1QjaXoLahzlH9Qm
WB7PyuK5WTeJODS6hR1yoR+LDGDquPTRK8WVEmGl0bdQOtZPlYPqh94EXOZ7CwF6IBvZmP5qWY4d
ZFnBN2SBYbfbfen6CVh3/Jc3dPIakgVvR5Avd68uL/PcKF1JeOGqF6YLGSEcK3cMzXqPqQofF/N8
+buvke2e6pom4HthoLX2v9zhsLMeEbn7/aE3BAsNGJRF8aULIBL3iyBdPhZP828J5ZJP3IGtRzUV
FCFXegct+5wV+u1+r1UbMSHC/8W2uxVdTMn70BBGJUr64Dmdk/Zo8gnqIHEPQEEF0n0nZD/W+Jgw
w1HLcBYg/J6aInK4LnwhlaWpAIZfCG2laIvdUrKgos7ZdkWOkxKtbJ4Ms9OKT8hXowNxiKbR5rZ2
cV/sLXPV01LsMnFXRVvXPLLYCVhFKbdgnWgL7xcHdlLRLXPU9vZTtzK/Y+bme+jbP5yLEPac6Hz5
w+PZH02oeD4jjthK82bn9hqcGLiIHQTx6ibNcV2wH1zer2UfpfHQAVaR2VaVFAr4v0zEb0+JnRk0
8erlXS4+V4WHJdsrjwRRXZGatXrshIIoGLErrLEbiykqn8vS9kfW01sGPll5ZUjWNw9Lw4xG+bGP
6lJocN3vQtTTYzjwLt1UJ9hpnbSwaQ2bPou/Bzf5WqtIP8TnEk5+MYWCunhccFaN7W02hFB6629w
SqeXpKMb09ptONP35Wf/Lw5cwnzzbgDFbc75omilnqMfSdHhKLfuU3EA27Q1rm2lkgd6pqiPMGy6
2641ALdXngwnJzlGC15x2v1D82Mk+kDXYnp+HBToJ5GFaTwzTEiAbr4bO0nEOZeMDhhKrUuU3Kxy
TDBiXorCUxuXMV8zLM0ES6Cb020/x5qkqnFr4/hhM38E7nqp8OYEcAJTzNY5Uky6oXmNeKb2BiPg
j7rBAFacvrt8ZuNU1dTa4vbT9ab2fXPI19r8vAct76cnEP86shNrqsjOLzlzKK9hzVjR0uyoLFID
QEABKmENW5aYMVuJkReF5TCzln/m1NJBL8goVxd6F+rvz0UAXfZMZwk45jsABwXOJj3i6sVFNJOu
GFpvIlm8HUrbA/AhSWEjr7LDaPfmWEk+VYwpq+wH+G4ydhHJxNTRGwV8gMQsVJYOMobUsup94LvX
3krYqmcGXGEC8puQOSVWNSkdk/KOy+3TMR32Da3S2eN4feOK/fz0THCV8rpN7/7i1JMBXPIe12M9
HzZcgdfn0W2EanqzdGbO8++9dGt61C4eUH+QEqBj9ug+SW8LCJEQxfBtReRpKx3e9LB2+t3XmANR
FBvDrKIBE+mREFQZjrnRtrGoOrIcAog0bdxmNp0A1PmpiY6wf1gjJWHLdJNqjHkvk46o1sjcbs82
U5GwALmRwv/e+lqI9lpo4w5chV0phJxtIrYPLVPqdsv5qCq1vQEhuoozzXzTEtH9a37Tb/qK/ZfE
CWcXSs9em/OoUGFcdtTpZ/ejlTcbjrP/QrddJDVflM2JffK4cToMe5MCasz9wh4jHBtH9BZTnuq5
Iv+4wP+m+LFrsnj010ZNLoZIDVqUF4m3e8IhxSjDdCXngnjQfznRBneumvyJxZC7c6UQpIrQuQuz
lFFmm2Tn7CWUC7o4ElDm3FwfbhjzwexsmOF4LIupNDVWdNVFsxSNPkpa6bW93ObD94wleWwJPWfy
svo9WMKUh4MrPS/kTDn9Z2NB1ofFCOajvn2JXLL+7w8qoZM7dxbU/5fUWqQwyYR0WhZ4Uk5lwCBV
f3oa70VnoUmaoF44eA50p+jpdtiZfrcqDrAKYFhGuNdZmHsEaYD1nxpUM+rq4DhMS/IhojDCZ99Y
PNsYIgJ/fw2vgB5aU+EzJxxdmOhnOXKY6cP2gHViAdrkhDFMcMasS0d2c4EkVtdXhQZDbMNHwXi5
zfZyo1AQASmmzWuvw7EI466BuIOOhbOXPCoPfPk7/qVvA2CpzEcrBThvW5cf2NWNArd/gnKoNMDx
3LaXNXRXtDDt6Qhr4SeXZKe/8gsaMmcEmZ37d9Nt/ykPXBFx+Wr6UedmGEPGXrU/3Y8fXOySL0ui
onv10gC5WwSPTt6M/qTNNuItjQEuWVjiybGQtWSde+Fghdnsn8yUpUbkwcLr7vVU1HWkz+wE4URH
iiDO1l7Acn4p07xo+3pNpK/HYHV5Mdkb6u021APYtqiZ05/+dw6mhU8WQazpYYWaug1Sbv+Yi0Wg
26iw8It9Cum2Xn7/QC9bOAhnDbujw9d3JmLRTCafl3rRSlBnD4S1XbGGJsojKpRVwpkbYVNTDO2m
hnkhehsG5G0vpqQd8InrhLSZErWWw68kNqSr8pv/tZd9l25xqPi/IaJSEryURkk7rjIrw1VFwu5a
HXLwf3I4MD1Ld5dpeNWW1rq2gTqC1NpUzR8EF/fwO+ITyoqGyXWlgMfkqjjglzV8kWDMK1db2zQJ
Lro/AAzAfhVh3hf3DFkylQUr+5z2rcKaDc+eXq9rHhNrUINLiqMF55JzkT15qeZ8Lw1B/3iYeyE/
PqUFRf22Z5zaK+hyaunvFzKkZBhx7/omZqrX/6Sq24+otduflcmZp2RckXOU+GqQlvSJ4Es1U6Hm
8Iquks9n/1VSuafomgN3qpMWHCuLl36MGCMfjpEhEADNhvKngfCKa7DM5AXQrK+SO2QqghK2d6Sc
Hmyc3gCk+/eVBcsM9JeBDs5lGmDLWzO8V+9wBwEmUu8m8cd8Qqe76A/+iVL9SirLexdGNhjfRukp
uS7++uwmiUjYn/5DdG08zO81S9czSQSLiG0E5eyw9IsHO7CSZ5No8O6GZm8VwFcVNRLjYoZ8IcPv
h0Zx5dUHAPmZPWH+aGaI+E631IOqs3XgWN5v9SX+wytCr6276DlirUH7azAlpcjqMU+BK9uftHvx
ftGmjsJ7lVrwdMsqR3pSYqHhZo6+z9W8rt7xuUSot8AG6Ap21vcL0IYPZhSaNUOBy4jGs1aKGkpA
7IWvLvb+q+JluMQl5jlnGSFY42PIZEFGHR+qjrat+zydFUMqsLQZdgQUG0z9d37sYBoqTENeo9WU
Z9xYLJdlBHqTI4X922tOoWSqrFNMTdxYJLbSFV2AEZytU0zi8MAEws+B2puugYJ1KOVK1IVh/sfe
1SeWzF1XYiIuP+DCQVTsOO7wEPAqaF5cZ1bm5P+Cqln2juKibtj9XHCIQEIK7IfbvcUcSutz62nK
mWmVhMRSKS6g6V+jdSiO9jFcOY3uhoi7Q8BbvnnRQbyAuNgOR7D15xHomPAabgjTtxuPfU7oMwcW
putJ8CBJeivsXp5PWCChmC9s+Fl06JJy7ovv6/uPEoaq6lSLTA8gPxu5NHpzM7WrajzxeadoSeNi
ASuOUn3rTjKdXAtIoMcF5E2wpGQpkMwp+/LKYiIHjOjV6QUBcVpKHIZaxfiEFOglSlS25+Js8hmc
5F0wjBin6aXruc5fS0fyDPwyH2n7mtPNoluvlHoiiWTJ5fTCT6cegJ78eCdni03n8iVXvHzJAqTi
ixWA9Art8RHtTXicmPsIwgtn7v9whUZKkSOcBb4G/lnx/AuZaFCKfOl2WJ6JMfKbtBtL6WK4Fmw2
p2Z9lialU2Q+XW7fJuRX8F5SABXytNbtDK3ha66tQGouBZ7XNOM4ws7bhvjUYfBijvy9JKBZyOEX
5Wgft6uVgcgniPtJxhAJRoSPilx2jj+/vezRWytc1Srt7PZU/5nWAxTVWk4L8evVtcFQ3M2BS2Ci
0JMjl0WPFWvwSbwiF2RbnejZJB8P8RRoPV5BxBDxydTZLGAZAnMTvdcUwNa6PY0lOLhz8bX+6UWv
aaMIZ7WWihXin8eUysXI/dwTcRwz5xQS8oNs9YI0gypFtQpxNFeztRHlBethJ9YHqka2t5XaZ9uC
saqF3TKcmv7JeootQzqZktbpnSc6GkJQUHSgxu/0iMxrP81D/uqTsesAFsN2RDigdbXeVX9hEkRU
MNBM5P8xygl3Lw163XN+JbifJhIG9qCdA3BzZNZ+2FSBIajG+91fGcJnFHGI+a/i2P8ufoR/1tLB
ZEs7swODuqbvq8uY+YE1/aCBZu52VrlimOJ2GgVnn1TAj2ztkUOubanaRS5zaME3jYTz6T6B0PYv
/Bv+rNld13eNeBifwSaJGEjuMw2JkvU00u+Pf1LlUgWMCiH6j8EGbVLbNUzP7HU+8WLuaO2pU18E
SNP3peYj5z0/77sfT3o3ffpqmUnqulRDpyl3SaDkZ/6vR991m43Cx8/fe5HktIsO9mev24x8gfbN
JHUR4MDNP2vbXMwfMXIHi19MWeerVnHIMtB9NnbbBwhpAhA9PBc68if3TWsvDx6gjs/8HeCjtgYS
8Lkt2605tFwtDdt+WvpEoSHp6X8Sh1UM/gCo0/KenznO7mLBzI06QOfmUTdc9Xdv69GayJ7nj7Yc
HR3iQSzo71VcGJh8dSw50dZS95Xnkuok467J+eTMf2T5K+w9o/UP2MJcSoOE3ubTSWXJpVOSYLqu
NKXPYde/Ly5uM1LsTFAj7NPC+Zo0X+bsS0N5hY3ytX7qLnhsr5mjlpjA/1G9y6mXaBAiDH4jtM5/
XNmrxkQ060+bWdHS6Zqh7+xFAGPPONCfvIvwg6vJs27l+8FMlTOCqeXXhrMdw5S+PX60mXnNK1J8
GXXIk+FVbW3VpW/2gIdnvMIw1qNX6HTaaJyn8Nn6MKEkQVIQAtG+fyUq3GNMUGJP2bm8dBA5Nspw
Zf2SBXY07uhCq8l7RxG3ULV/Js2bToWe+VBQW1mFr/UPI1U8I/SMmB8lk6Wq+eA2z4WqAZTKov/c
8MEpO+DSlOHnWSUcDmpbnp68Xyy9QoBaX2q7oX9w6yL3aIXy1Y1kS5z0ypsEenpVr7cm3tN90FM7
nlW6yJm8QLt7UhA18/YAzgrTJGMtb2nEJ0tYl4SRVIYP0JWoJ94VWqaiCXXK9MyMJm21R4BoacPI
74fva4Mdwd5kdG6QgG+NdhEpVOKPokXzQp+56euOAJaXIDT5QYAkA1MYB06LOq8hIbbSw5B5+jz1
0roIfwLqX8ic1jWuSODOGf1tZb3N7nAWLISsO/qJ9IZqZMVEweCI8jZvyPZaK7eGIRvcc94efyPy
wMVW5TjDSVZyPgCbD/dKi1K3g086D/Bt99+c+dwbXv7yfX2iebN0xq4lCYBMprcaul7ev4w6Ff66
LMs1yqlMuWB4cUlsk2kdmZ3Ki6OzM3cy/hOq+QgScfWM4iUbOjxmmk2Z/FsjDUB6OI9gbTM/V/6P
dE4jap1puovZmiw8KWOMv8DBrrpDuExyGHuHQFwUQP0yeNrw1IUjuhSZHZuMrkRWtAS6i1cl+uYX
Z45BjUhnEJ9fdkYavp8WwpysAvaxXf54bpFK9nqLbtM27ZEnAdfDJic2HS9VOsWaW4Wr7JHOmAt7
0/WJKIAO1Q9b43fBFBDslfdltOSKFxyoVQ2iYwxOMGpYGNckRQM87PHwTuNjqdWgo36tY3HJfJfi
iMz8t1lKupm+3xOID8skzOMnLDWhA+z+AGsVF6QJjQxqh/PizhqemDDYE9IVFehfPmEzFwCCR/+t
xhP3nS9PYqgG4T0DTPhSx8ED/UClif/1T3HidxbrQ9jnazdq9vi8ZABiA4Ov3kc5Kkp85PYcntZt
sGZmUeyPcbTRViB+836lGG8Hw8lMew4Q1zdgon3A1+vta0JPVZQUAlk9rJ5DGZF19WA1rsRD65Ge
oYHJmegMYnIrmmuZbUkogrLsG1Tb3hqmA/vQcVPcFT+zzL4PBH+OAIZyW6CvNq6qS3qojCQ4kMlh
NuEhDZE6t3qYNDW1rbZCYUnIKaS3arJwJRl5Q5s02aoB4S+R3l8+wzkx2DZ5xTeHlMG3/RtPWozW
exM1bU5nLyJPRvYnMF1vNdPJnS9FpYiZ9YvJsXUgQwoH+ZB61M3tJky+nqs1X58kh1ZrHC74JYKX
I1hGsAFTmc7vzs7WmQ1WgdqlUUdt3g6cdJC9X47GTJi37hqaCO+jdoYN1WeTbMRlImRkJBzCXrkD
C9e2HtpUo/hrZxTb1oLdmd8/ZcUihCdiIlZS3klWq1hQKIbWL9FKc/D43fUScEBKW0Zu6TzpqouN
IoztzDCmo8cwL1KkkAsL8dHcddflxILTLDP9dlBAD6qdC8mLfMRpdaes/kQ0gIIqUu35U3lwbF83
426zlqp5n4DZ2QBhD2BpO3B5V15VCoRUUScoUH9k63CfiZc8Vdk8xMakZ5gN8qkOryMWAdyNqWvD
Rpjq8hNjnIpFfG+QZYfe4svWuiJkn4tWvfYypJwPRxTlfaclGDOzVmKw9R+muvwqCLRICR/2rSs8
y3liQ3/P0Pp57kbHkZhD/VSv8w4o+nxIXxnuj1pIguzWpvF5AYDdJ5H5jNOdbsjynphFyPNf/DAg
lK864QcViLz38q8xOBvW9LkShDWb21tnLngXkgF8JSL45J8JGenJ3DzJLITyHpdKwISJd+nVJMl1
TRrxCaUc6/K0HwvUzfmTbirln0+gDTccMER2E7vpZq0lOiQfCNC9odPVZIMU+yzaCDQpa+OYqFU5
OjY6ICjgViMRQ/3FtwpLDHtqTbmpCzF9+aABuPMCk15/hDP7KUpBAH9hAbWTFKIbWSw0F0Y11kC1
7tVcb7PPOGULUMOhvig7hCcwegREp7we/P5GU9pWLE0ROYVcHTDpTt+AFU9QWzwhUsB26Hnj47dg
fdZGFGoCPSbaqGT+HgMTSbNjA43DaeM6HANQ3qMgISnX/7KUmYeK7K2XigAeOP2puWpP5u32+gtb
586HiOfzcB3R9rJbKK5KMS/1H1hua421O/mA698tSVbyq2RoHNWFpx591T63lyAZU0PTghVKyx0s
G/W8gYKGuvojiuGrDq0g1T9RpR90m9zaF/7bL3p6qu2JULbdfiFRbLZ6ITj5fa6WJRBMu3WJQc8v
hJwUMdn+6slE0KD4O1DKZII1ZAmldb7JH0ONHGFFHr+fntPpbTXacLeR/8PJmFcrqa0k5Ywl4VMu
1XuXtaMxV6zgl71ThWMnctDu/0n4WvowMlFHWvfrH32WUQX1M8/j1+8W+NB7lO5bXFH+lftWF2xo
IlIDoTf7GeRIS2oZuS63nfUpnoAbVQXp+TUsYMzTMhNc3n5XlHQTFao93PBfa/pNTxgjZSOrCUm9
CHLGsXy2qQNbd3YgYhR4CPbIFlK2D9ioMjJE9BkxBrxTmWghc0quymwjh/kKJZAEbG0yqgcdmJqq
3MZqmvwiOV4ajp69v2tUB2/yqn24h5n6TT5YQ/AYziqq7by1mwgrV8IsQPzKuOZ0DTTupWMJyWV7
aejHCDOJkcvjLuoa7AHhqAFcem4GxMOlP7ZICObc2yOVxsQNpnpYuRT5jwgPv7sGbYQDLKdmp0Yr
yesUcOoLueKZOKvbC1eElVHeOLLINrKUxbelaXzuzpWN7zKYo4fxetGRK+uyL4NQLplKNbcY1d6J
72hKXUrqid/ssFW0lNjwhX2EyISasVrvqG1ndmNN5W9gVX/1cQH2tHiH3+V9X5/HmQtmUqUYaIqa
qsoBVpIikSHkdPGl0jeseetDuHmc8fpW21Xvn8BSrS/vrnnOAh7JQ81BrX6BS/LDjf9CXgFKHiCY
YZTKk6SA6JvC1t0kA2EfNUk6OFCKG002l8GTRwiLFBLoNjBIEUT93x7FCq7Z1qXEsL0qT9oSf/u/
6WPZCh6p6pPvd9dxk3MOyBfa9phJPTf77YD/ZZqfDdDZn+UaLjS8QrUQIRK82jPF2iExI7JtR8H5
7tlThM72pFZDpAotiZOvQHTHnbCTlR5guU3VbD9dzNxPSerMdC9Xmluk+fGh/0HsgVzxX67YYoxQ
Boqn93pVVel6ZZlg49o336EtOALbz4e6IrXEXrpmoCFUYE0rc1KS94fVOzEstXGnSpysxKevm0Db
h9/5Rmg0QPGNFjaO0LyGc1tEa1IQXGwiCPKIErBd+t1sITuqUil+RAA/1bxz9RZsw1s/W7u+2CwA
acPE8qaKh8DKl20e8v2Xv7B6nMQZiZFbSBVvqtTB1hwh0ClYoSnYK/NaKWVwYOsbnzHIz+seVFc3
UEw5TDpF/DSRSmKVPIC3GgmxvJWGU6cVi1PtIzPHomaXFS7aMrFsVqFNst/Rn6dsHj1L/uJgl4x6
afEnXK94A7cqzTSLPl0KY/tWx9nAX8/GT7UDiXz55/WptTW49Uhz6y/Sr3WufuZRtW88cO6oY6JN
nLrhrDZ7JzpCKDQSDOy4qThUCzKM23vSzJWtztyMp/22KE5n5sGcah4SfcuF2+wSnPcTqyA80mHS
7YgtMHpjsSf6FjHQ8dqomHqbcHxiMrkaVWJtUoNctYEZrLAsbFxF5BPyhFi55UsSWPzKhA1OiB3H
B5hgQUQ+1znNwscWwplQ9Nt1REEmco/fBgGfP7I2X6LhaoJbme9xrQrcb+2yEvJcFMdJVUcH0C8i
bKKT+AgPxxBsNQ+ZRqPBDopdO1F/KYkxhvoPudLixfAOnYHCU7aAUWxR3/FGhi0qSh1G4bOt48dY
nWyIFO53LEgq6wg6M4/pkSl6s5vi9djQgUWtVwCtIZUNp+zsXEXHC2yqgYnaCOUi8fXOae2sY18u
yqPF9BqiXFnqyj50P4+Q6KTHoWo2IFTFwKprVBa8FO/lbuQDo5JHX66ULXzMCO2VKtrzujWdMTBr
J7WUDgiM/rfYmiWpZKfAAyG7wQlKenwMpdlji9EXNR/3KDiFbc+CXaQkkXid8qJfYT1MwZIfKUr+
qgU36RH15dO+ExWT9ACj4DuoKf1u1QMjp323x5nmc3UixazCaWx3mx8tv8tBlHqZC+z/gxjwDUlr
lsyfcFgIQUr16rJ3A9ac8lGALc97cqxiB/FMApwH927gwZi9dq8diiugpPNs7+N7KQAdmhSQToi7
wc+7uAmvo0N28mKYjEiw2VrYrz2ckKtF7RtYwr+InszBJ5TkF6mgdUtJ/VHYoNKwbL2K+hd3ZkZ9
vKMRXcs0DBzfxraNSpI00KSdEPWYgiuEw2sy5Og6Q2ATTnxBzRLzRgOPRUo9yuk04OVYBUP7aHJd
T9aIrYy24k6dhefWsB0Re7voK9j5LahmxxSnErgv6lTkfzd/1XziU5n6YFVzWCHACgcxsap6lX+S
AYVq1Q6xv+L+iEtz0YUxT/b9ujRDVZ+fP6vndsVxvfNTMpoEauegrpRMspWWKSfewDoomHNH+0pZ
a9xwPY2IWsxngwZIJlock1t6vZRjY5BEsb7lUfFZh13r6g/x2cjmlwiAGmyEIKKYFJ7IRx1xgrdB
OAuafs84+jrprzm+NnLp6W0+EXlVf5xSEx2sfsR/icdb0k8okutTgZ+Qi4NjDE/O+jEX9HY9hXET
L4TVoxa9bxgESkGeGahG2jAHayr1kp2Yv1Xsok1BxU6VV1z6IPVxr9JkG1bzwwR60qjxMyMiTdrM
ngxT/BAoPqClFnj4AWg/iEnXY5YeiYD6AnbI8eRuR20JroFnGm7qUNxCdyC8/eMxWI06Ee5wBPM8
LL5SbrQF8W6pU3u2yYVnozixVmf7NuYbTi09A2BM9DjcxyUDEnqcZRtkYXiUXduluQmoQlK8Busq
GDQ4niZw7Se+bCpY9F4iaCr4iI9VuSEWcUuBUXXJYfpsNCFEpTtlttm9Uepqg2q8JYxvdT8Tcv4P
VJC89RzfK1ZuHfAeFCT6dnI0kERDrdtoRmCfTg7RCaLRaUvs3jjkqwlNRptA2HKy1g3yTLcnQBzv
O7AHjE+WqTMdjqb42f9C3z36PvsOj7OlK2YVksNk68J1QaZhVvMLRdnSu9MogGXrNGhn5YhVS8qf
hgvsnociN+Zh3xvCE5vYuYc/85Dm0sVEOSnnM8YdnvcSTan6mt6iRAYUauFX0tHwOTcJq5CUDHzE
XRsc3+48pa7r2DwEEZQWRzxlf/OGVzsbYBFJuqXc/dlnaSfWHfvy4mZSCfobLBaxy2OE/1JD+aTV
heurFuznniAlfGl6H3UpNTIWay9YNa6En8ABBZ8ZFXqOO/mmmNv13vWFnzgIpx/hBYOCVGaDWe7Q
tTnIfNY3Vnw91sjut+JTIWG+Oo6/NdVTljQLlZlGcDghMg6IpRJBnXMCXCvNZDDeQgIjjrDxQlXK
t0D5yaotB78vc4FbGTqBAp66ejz71Vtv92+aMog5hDoJEiNsQoOIc7TGkZw+8ecZ0LsOGyKf03vv
fHFZTNaePb2J17xWAmZUf9YDQ2EdXhyC0xGou8EJOCsW85MAKkFSn58VsrEE7mGCLwpwGBpO1Krt
fMpsXtvx8mQeJtnCpOW8Fnc1bq9WrXEzHlswiD0ZtJhM6xhfimvooQem9k6bpSFDg3/hvaL6CnnT
RlHNwzhqh+NwN8KAkgrJKlXolm4ibn4cfyTvddpOLwV/cXH41ATT6rd4X+P6/Xua271hZSMCAvJR
oatHHruZ/p2OaoCN0s5h1PoBx10+0W7tME30nU3AukuVqEwuawCOaJ60aHUbhlRDhVfkr4+ri+Wt
1wVzS/VQBhzfdVogwSshthi4QFzMVhrqSjH423PqL7P+tSAQ3CyQInhlhmMEpBHsr59qgIBlhENg
shkO/KQgwMbhG/tyHABPY5QtkZvgIUiijPb2A5hMR1kvPfys7SOOeHLLQ2G3tEZqOjC+G7rPDg5W
uNg4xQXDlAkhJgEatlj3ac15iPyRgZXMWmGtF1x08wsVvxQwVAvzd7t98oH/tJpYl//HAcy/uaFo
ZmuclDDG9m2Zh5r8B5me9fvw0I8w9xRN1Qrbt8874+Bd4WkEoLsODBlm8rpd2xYdERqetmBTB+/X
zDWLqFw4ZEFpE5tBYrVXRCRTiyH0kJ2ebO3P+pEKrYLKyfLPzXsasWJHdNqWmfs6oH0qThVXmY9n
ST+a4cEig3qTHTqB6fAJUtGYTBRcKmoBzcWmajZvCjlAOnIR4hfLCpcnNH2h4reSuSfIZBwkj7sQ
6+h0BckcPCrl+Aa5ml3EDe2JZSH+chj4lix82otHoshNZdzsKMA24qheGqRciBI4/Fm+TGEBsLjj
qIQ7AMdOLk9BOPLxwrw1BqEMzNeGQEwG2V8J67Pujrw5OdDSXw4wnGE8t9qdXIJ5Whf0A0L1CQ8x
ZK2Vjidsl+gzzjoaIAJA52x+UByGc/9ypDxfW+I4ksWwHuXiqSxOCSRTy9QEyDM/5j1gButrqV0G
4A2TJvzQ5Vcvh0srwa3dsJnIFfBOZ6JPikTNKm8ZhpYiNc/PaW/cO1ZD/pYGqExpKr2NfR0alBxh
QAleBKJajhBXwmfXR8uxIBDcvbqY1ilByVcHjDhi0kBc8eAyfmu2puaZpbLez3S5hn7YPn/vnWEU
I5gznYC9drDDkaRPThuMki551aSO51oWLzU2qEKG7vVgu6VpH1W+eWbX4zBjVl14Lgl+LD+o3KS3
j68ebUnYmyiOoJj/PWMzGhcQ4oK7giRNGG333o6B7bDRk2fRpg1Bf/1bsA29oWYj27dzs8ri21de
tI/5pBDEDju0HlIZIC9AjKvhkvLLVy7Mvpl0ANdOiYotN4eBgIchocxnE1O/Jo7fKM7j94GvtIxW
5yJO4eIcCWj7dt7RYNExlvBJVSTBA7HBS8/IkwcSyzvGMNK2JVgQnPIPirpr9kYYiS5syedcA0u6
8Y/z750MyVQElQ7hP7Yty9v63Juv4U8wGt4O1gtsiHLRXKB1o7Bs97mOfLeYS0eGctEO1Alp82ko
LCM7hC+CWqe1VIv1fJH34gfQemOE65N0Y27HO58AJVFLltLuvVnKogzF76v/3mWBv1LLKo0qxYRI
RYWbG8NRyekacdpv1i0Sjg08y+PQakrwyq/6fJLY1cgbLm+j/nLKvp4UaYarJmpf9mDcwbXaLpXs
Ba2T8w3XUff7IqcZTHyFnWqQYwa90BO0SGWRqaSxZQPzZqD678EmfmatMgstDqUVCUXFWcj5iyOa
foz/CGPbysq6mpOxzw9IUYgfQn3x0w2gax7mVHj/rm2LlxhL59HqQhSw2Nmh8Z2e8Apo7oGblsMp
MSA107QSpWu6wUwN2slt9pu/utpBA9N2/xTFsDryAyeuEKvR5K+tbxe+A8fIHNopK3vR3s7S1CJL
S0oJW0ldVL6jglWqW1YrzBlfFdhHlRJSTqSvVWt+DuivfRlj6wBhuE0JTUeChEQHSS9E1aPOjDAY
wleKEkxc1nFn8oAC83HboK2Va8pQGGpUI4HNhz9HCSaocgmbVwAd7SyKniTn5Zq2/27myt4gDM0b
u8t9jqD6zgfVEL8A0erl9z/Hwx2sQPgpEdRwuENx29hbl6V4nshB1icmQKtWsc9qWbFgQ0UMTumU
hrcO1yzN/pPhqiAPziAn784yPV3gu/t6QKhzyHNoiM2KgqT03ajy1/rtoMg5nfWdtXIK4kV6F2u8
ayacHdy5cLeoBzGHEfmLdnALRp9xneWqBHoa1k6ppi83bpswd95AygT8TRhP18Fy9R8sCWm3iymh
lAHhAj+OWl7nX0upszosGOKLHkgORsXFXyu32z9UqFBzwNiMvkFO7f/2LkbmArngmaTrk9zc6+xe
G/5/dm1Dt0vmJogW0Rn+REzTBraiJ0RiEvefCv4QimZvnKv412qWaYhpcuYoy6G/JRkBNqLYl1Nk
JIf/XaVFh+EHVpcRLcLaY376JVXhtjUm3aYbBHu9q/UET3KSOb9BhKwsCnCdKTtQAWQQDwPHQ3cu
ylqxno1i+cqMLAmxvPCcqk89ZaF5zuO3ouUCUyQbRIs4XjromMSldho2o3gnbk02Wlx2msRLvReA
luvAEPulz0FUQs3f7E2Ejat2oL3gQmNV7yaXyDp1Ef66Aah16yK0dO+/YnpxRHJMy2SjfVWpeqoQ
yXUWncUihqcaFvGeNiSPInYXXH8ZgF3axBqQp6BOjx78ohU7Zm+/pbzcbAbOEagvFcqgzw+E68Li
qsdJXd7eDX5tizIuj/+KZ2CqEnxRNZ9kNZCXHH/2Bnu0xkc/ioV/FpqCF30ZzIdpVARDSaF5tiPg
+x3aEniHsJEv1xK7V55dSz2umhJNo1N7i4MWi45Q9h+pPjjuy3sRoSYfrceOzle5ta6FDmAbzpDV
tIc6VkAsPxeFmDkFnTxgzptpvqIcWDEp6nUU1thD06rMFXfyjK0bIy+7EwlhWMjBpwhdMF1nsvc3
u0LsVg8AtJnxoN0joOf/FsSfSgbNW9Aqizdxn38cwIx1XnGdr39WEua5INjlM4oexD9hkQgPHkkA
ftvKB7XIc7Tf8vnn1r22OA8/SgEzyKA4MBWgmWVuic2XiIUd3NpC0Iy4+NnyTw/ana1fYe6sD/lD
2ze+3UrWzgRKgh6wTcEdSKgdcKSc0ZDVEIc+nmJW4QoZXWvnhV/b2fLBaya5qYX11aTZGh37X/yg
t9+20Ff1gt+3K6ckCLgG2V9vaSvmfGc3LbFMFpAYYlgdxYqDiuB0mdeGUk+krxcvaLldOR8eWr1X
/S1IlWYLz1Nl0scnqVcZeUZG/F3bSGDyL/JAQQAKEkhmnscG11ca5KonG20wbmlROpeiLK3CBWIR
d/aJJYsOW25N1ypbMLL5iD8ehOQfhqtty1mtyoRdHBF1HwHDaR3na5Jz3avOuEAwcu/BSSYmWNmT
SdNJ47CgZtJrVsCWGvjxsRh8OMHsFNw/PXC4j0Vk7Rku/HCazQ8nmVWtzV/CgwLGTG0EOaa1G3YM
PEJ/zXIQCd/wnY4nd6pJZDu/oPvKAtQCAgl+r5hlkxADNjIFF54/VN8zNo5yZqOqDcJO61je3dZG
eUzXMn+SbGFvEd7lU6hr1KMD/F4zY7+wbHU90Tez/IIzt+SGkdpQjuCnck2hmybyxPNqV9/lTExr
lc2kXQ65hGdH2XWFDF8DQM5Yg28dr8d2tMTgUXrqS6b7HopcMLK19yQR5l6H6F9gNreBdNhq8bmn
PMSVo4pPfoxPfdJDLgXoiZ1LKf4h8DTCiQ4lB/9cupEnJQipW02W4ka2ncojlc4lobcrqDXzR4Ai
F1UNUy9Nd2vxC6+7yCStx+QQ81h+EnylyZN+HU0Xvx0RhwRhDZQ1BJ2cQJAkjAqJd16iO/B+gWni
thpg/VQUb6h5C1EWEgSmBsus4mIt+YbLZrkVs6I8krsHHMe9Vr0tIwr6D+8BCO1GC2gwqSWLruDp
0sVxB73yTGsHzr3sTDjk0eh7MKR7o2FY0BZByAgP+K2w5sqR2Sah9KWT7n0GVR4aZXSycZpdj12I
7cxGu7g84BWAZRTCq/K7goQVqtIdDJ9aLq/Upyw2kadMBfcgxEpm3kAHrdTl+KxTA03NaM3ox2Ij
yb+i2+1WMT1cKP6+zrjR0rGz9f7de8XNYtGkZaQI5Gt8BfE/sJJx58tFG8yrDblb54ply78kABHJ
8DQPYjPk1v1vlR8DxNc031twCMDnLRqkuMkhGKx9afUqNw2Um1qiTEQOy5AHIRHNCBez/ElNuBJI
nimVvA/TQSvyTgY7th7RtmUaJyQsQTZnqZ5OoVjQ11Nhol0rQGdXLlGA6bqpDV5MVsJnI8jXYJ9Z
Bv9LSMvEsnDKTK6Ckb4z51FefZHXHXc2LjuLR5svJ0i9dLYAVciq8msqsgxrvPqZZTKVK3Qu5mM6
oyXchUeV5EQZiD6qHjn7kja4MNQ1AWMtHULO1LibFFXVMaYmCzyfO7opCSyf8l0qv2YDaKJJ2NbR
boONs8sar29JQsfb9Tb9LDyrCy4Da4cmHIcCY8q4EJmY8NulKXMb47xGsAIqSXDPyeePwJLIeLDS
e/axU/Jb2z+VRisOjkZKkDlk/WnueUv0Py0znP8SU/ZXSrKNBqFLhKCGMdUrmDvAR5gSU+Sk4KCH
yfldH1Y0mLtbM07gvDVzCE+zRLUoP0TbPZ6/xzi3IJq6gEO/fNCztz8m5oTdns3gSaQjPpNkE8HH
RQpWXsbfg59pjlV7f6mYkJx/HH2XVk+hejCaGlo5NZMOv1gh0QeKF4BnCY843509/oAwyOTvW+7+
z+kGo7RLtXLAhsgeHiiKsbO8eqFp7K8oUDQ6fcklOrj58wJ6lAArVjdWJiI20QFmVEFp9nxQBHQM
lSfRMV6Bo/lFAPwoq8ynpcWGavTShe71N5dF2F8Kbo1K28weorGms2iW+2XUYXHiEvj9xSURZ97Q
NGfN0O/jiZNT0RyUkccbJOeDh8W6zdwfkQKV8BY2Du4B8QdY03QdsQUlPAfqPt6RoFFlI+5Pbce3
TebPdCPz7vxkVsQMpO1KzIp4ZKpR6b8/MKDtSsIeOKQdam++4Dpg7phVYVJcUdDRcUFa976rgLk8
57edM8Itychi8MNYYVLzNkT7xIIztA2jp4DFtpsAAQ6VgjoXMl+lL0/yw9kERJwK63SbzAt2hP/c
SdgJvEMW4uDSzS7r7FUCu9ejc8DwM979LUNesxjtNzu/0b5LgF/XHveLCsgUcG5qed9xmKSMIRn3
4xOkbYHp+cFEYz3UFs66tmUkigT2hwePDHlV4hmx740HN36mWGhG9pHv90u6lAyrqsHhwoOzBnzn
pBcE0dNlvk2mFti6XdmMQ84TemL426YuovToucug++Wjob5S980oBCQ4mf9JRuhMayWEl4EPQlnl
J9kJ4oE5L0V9h7w3xzRF+NnS34u94pJe9TBJVIQSLCftgrOZwnE/2ZHzRxQCvFElDixTiUY5hw77
wO1P6q4MdpHwtgpviEjaF7uusEbzVsqTSkAtIcivqECqdhSRAujoJELLVKdUDidra6Y0ZS3X5KlS
nagZmePthBEWbqjef0Fc1w0yaFPS8WYaG2lDL9pVpscIvmoikZXrSRFK2SQH8+C6ca/SO23XKok5
PK+I8dqybvRNp6ZO1KisecxZ6QPt7A4aHH3TUrXKKFGLpEx7JrUIpU5pgDNXk3jewqahHqh9/uA2
a1Ck95jlqQQU4GRdXZCmpVihoh6rkC6298tOVVqNaTv7d809ZgxocZWh9VGsYJFhmQmgM7d0x23X
ZxlzHx8noQokNCm9zQYHqJypQvvgJlGLU+misXdDMG5Zzy8nVs2dOjndS02nbk5hIMKpU4a9P0lg
TpTL6d2ZO+EWaMYxoDgBnwEbbbk03bM/ATyt9XyD3+VKvtwqDdfOfw8p/Pnn9N1PD1sqOIeXlbLb
l4Lu7nSBzvvRMZG0cgQCtcX5c68V+8gP3ORuIIJENNRiDSI3g8V18Huq9luIrqhmNKrNotHHzpRG
l+/+KaKOsIa32VFWNT1L5cIpNZys3XZ2eihGzXXRp/9dmJYv9aKS9YL1SBVMQhJgDHc3Lf+Jntyi
htWVe0PFPUHYwbF3xjFn/UK8TnBXecRqHoVYyIXcgp9NCj/NuR+3xRndQM6Caaz2DRPmxN793qXo
IyR7g3QHhJl/qSf0bXAw3P0NFrr6WXTjLBbV+zzYwv1FKKde2kUtdiRh/OlNYyEYZGpOk0BwlXFK
6CnYnjexb5m0YArCn+UlXC3KDClU9GRoYsBVNdgLDu5eD6Nf4uJi+j+QezvxhM6BdWvdBJ/FgzPk
d9002ct6zH/2H0UD6b0Ea2i/iDPSa5V81G+dgFMSm/h4cSWbrf2WLTwZJ/YJhhTQB9/CUNvEv0ku
yXDgnSjaKktGUaXVoqpQPh6xGI0U5ExJpjDGHWxNE5fWJ4+s9i+ahmg0ywO8oB40V4klrRkTqXr0
Z7uu6fEX9sOCSHNsUP1USvIO44Hsx0e1A7iwuLMD0tt65+/sEptrFzD5EgWHAC1UBSeDViTUMg52
TMfAZogQ6x/yOCAhu6CuR1DM18ePuVL00EBMcV3s7jOy3ZsdYSQLwsu4rf0HmFEWtPBh8If5u+ze
PO21wRbi3vljNjkdwYy9NKMnyBEM33kT87LwprdOtAxZyBsUndJQHnl+kWQw3Zp9fG3sDA9jMhx9
ZcRI5RyxJW8k9nwH7eKJTiohM+jnc11YyLldEqznlKx+1PRWOgiFDFGnh9HZTZNdVWuYYvbsbhvX
UZ3rY4kgETP5YzhuE0xhaFm25W48U9TlECFAi2OiMFKidv4TAqGxgqfiCGOcV4KknqMEGJ3YdboZ
HjrQDEL26uHjrYwPQns9bUpKnEgSmv0P77//bk4pkFOd2JLQOLNJFxc5x3h+QuiqJL2bvRRui67/
YGXlQrrjk1GHcfNPGInO4KlpmgpVJg+j7kHqUfl/uBFnswMCylE1Z+bZxK0u2LoKP08/YU4+uubF
/EOvGMpPQrjcJM6qqIMgZnXWg0abyCalIV3nfJ2F+HUWUhYamsnParqmsIKAC/N9tz45X12KKLa/
Fp083XM+cZ9Uih3P0XAVMFVeTDPnmN1Jytify3N0tc3FzTlY4lK3hV8+4hyy9BUBFBux6B0lpEtG
IwOVPeijuSQ6qkjdze2BsFldL220SfJCqDbj4ksRz/PtEYm5sJ4QFaQcAilgZQQ3rS+DrVEfOTs/
NQN5ecx+efSJsuLydTmTQNAM/3lrVw144YyiYi+SYeaAfBOO2E6eCFa3S4rjmcTtatkwe6gKNwk+
EVg2uQklbZ0vmYw09fP9XbWXjjZVBsXNoytQOSPvqS96pNNBiQM0DvzIY1ld5oOdjKccqZ64/Xed
fk5jMn30DNC/A/BShMC47HbyuSaPVmDiUG+rKIVXloR3MQtx98Vwr+dUhCsikxUVVsBBZ83oAZ1D
4zzmsHOH9SsgBKk/Ug44G2nstsC04brVn/WibU7Drx/QQxWTQXdUvh1uPgphYAbuxqY10hjRDYkK
It276M82SwZv7q+3Y8I5glBpuWYd7KIULPmBYU7tUsLfsE9YVMYTdBxOnJSpADb54iiSl0Xlxblb
8yaz7Hsw0H5CXWkhPiRhFReT1Y6w8Lhys8id627Tjcx38NJhW45pHyVQyoLg2iFrHDPoIySgx0E+
kizX8MDRAus+ysUmLHkvBG5wK93SjmFrPGnpFWwMOsJyp+48/5mbpGv5Q2y+9ojx1zT831TBeAPC
YJVz0xaWJ0zwlbSe2nsXKMbOOzWR90lf61xIgNhrO70GL9lXFcwPo/j6t4Ipin/bxhE0fs/iSXn2
XOd9Yx/dAcJjS2nymTkKdLBTdM1dUG5Q2W2FIsjR8FUIw5HhlAnJ+ILhK2tRczsAuBYpN0ZQeALz
Oc6T5k4CiUXiRaSyd5VmoaSiJnHyoYopVYBBCxOO6X7LsPEvnhB10vBjIMsjFRUv9lxl1+kN8606
7CdMLC22zmQe3sDqSfGaXn4+6C3mX4yASun6lBnm0esERrW6fmM3apZeUZTl8w8OXsP9mdht7LjO
31zrWO91dsvkdzwJmMg5xClppHL0XaP5KvfeIoQByM7VvsHAWu+yE+L4ovL2Up5f8b5/bwU42NrG
194grWIV+JDyPl0M56X39VUrTvILgvgna+Rxhn0OCj/yCEtEo6R2TumqVeOwTbZoOl78L21FH3Ib
mWGJh5SlBSe6C15od4lGyjCROUDaK9a5h0WI1SyjWKMojm0bqbCqhTBNvsG8+aeMRGQpMwTbny1t
ANjy521bgNxMx8zRxgyOLlGadWAZrogXzmU7sfwemnZT/eOV8dLEAX0PC1pVa2lAINkEfF8fE5WV
lqii7flI/h+J6/oArU+yguxcy8CbR4udsBTp10xEEwtik2IyIzP/tI/a2OlD6nXgHrt8ZkQvIwFf
dyLZvPBhwrcqEKuY0OlMfhC1aZPPMw5PW6L91hZs7ZQ5C3gwBxpCN3wcuXz81LODBZYXdGuchOEU
uDpsCCgZ7gv4ziz8UatBAAfqG7WUQXECDGfCtQge7MM/3PNfP3QK5UXGBnxMuKmwLK8MIuZEBMoh
eaU7uGXubZGuavHCMottAg6J9X1NYqijUySBxLMbNDTIJh10kJLMktCbs+3UFz5D1Gj3XUOvdsYC
qDObZzoIVuZPZXDAQyDmV7qA5gRnk7almXYgmDuDUc1iDo4KvJIfDsAHCFpIfwnd6Sp1euoQrUbe
JtYy56KLuiWJ/0PITeSocCa0lcFORaIfbs4VaXW3vlJETGQ8ZP8D4PfSATea6RpvOEA/FThQDaeF
ORI/J3RMdIoOHwYhfADq645IdmQdw2NoFpAZe3yWpI/YDnCWXvKVlW6J0iHAJEvF/iW/n4Ucn7Nm
ttdxm15yzxDear/KfDJ2qy02j0voXgkBsvaijxO1ji4NxtASSu1Yy8P3rDaNOJMujjW10l3N8z3I
5EtP7PPJSwocK0AUocfNZYc/MjQluJAAwM8qljBg4H/9/W1Xam8MLvx6IRwil5pn3gvcy7wnRoUq
R8dDx7e6lJ3op8iFB5u0HlsWpADJhoP29ajiavyKbeAoar+iq5PbLM5NlDE3K5JPyzTU9RXxS30j
01pEyiw6+kkGuiGJOvj3edERsYdALqYio+ZXaKEohZa+dMTgT/Q9hpoXbkWpxvQW26M9Z1MM/VKz
sh2BBFHy8Z1+riXG2RNihqP6Gq1Yj2QzDOeSZ/EwlTT9K0OsvLTYiuJ+ElA2fsRbU7Ud8LFFk4D/
LNTxIsecY8jiiuD5tgcosVV9eJyy/rpR7etgrhbrF6mmv3siR8f5bseiLL4UhSeHAS+7MpULMjj8
cIK7b8H+85zJF66TQcTfEzKsPQYeKmzCitnre8uTfmAMq6VHIjICbrgIwdeQdVfpd74nHf/GORix
gvqzFWJI4UgRNwozXsny6rtuZJNKFR2kst37Wx3BE8XqvkmUuIlUtd323imf/ikWBpBxgfzZbiCG
WJryyrKtcFwbkaVHObvbYtIvhjff3jR2/LBgX8uJMP+rXG+nd6li5z9Qe1DV9DOrDMva0ouGpRcL
JmyNRtuVjv92Fu5uy5mM7tDakSERs9ZVncY7UgKAUicQz8SL2ifKbNGu8u25zCyJG3PMQLjfGRA5
GSc2cZhkhlPe4HKJuq3jow15T8vXPKnfnVFboUPnpMEP0d/MQBQX+ge1lHga93NwNr0kF0n5llEu
x/XB56FzhanuL43zZ8m6vLgFZHU2BMR1a9j910Vn++z8wVHz2LRbzkcze+J3L9ZWP5miz2m4sVRM
2vSVrK4E0eQ7ermNBZFLuRGIvafx8QQgubrWiS00VRE4cpOttiTniizYncgd6fciXVIZOkDixxNV
ut3jTnryojathrmHwRkPaC9F8Gp5wz5Tv0iWa9rHhJngYE9KNsNqt1Pbr0TwLFMlziOJ21p9y2cQ
xlvUuueTV8HEBtOQMfhPlLsAYQLERly4IpeMyXVMdLv3CmZ2R7R513U4imvDx94eMUeVxXUWDgr2
Yp/VCcpIHgkBX4JntnoC4IvWLilTqnPDpe6W/TCGfNyJA20izZ+hVQ+5JoqabU180WavunzOoWu3
eGx7pEj6DNJ3jGcfp6jn5IFDsK0vDu4r6dfBboXOt/AyVRYcr9FBIpMs4sQCWy5R91PpWsCA3eqx
IMhsZQu/0PtErgZHkVTr5kae0DNQNBg+wJX70+4KTd/6fv4Nd6XKOnm6B8mtEB95TkfcgWAukvTZ
ENwkhwuhdHi42bTzRF06EInk6D/71npofee1lUlsMbNy5PCXvW2aYrq9k/LaBqeRzXo20nhApIty
J06/mT96Y1DYx2zDQWLTK5Ss6A/osInvcmzYD/pXpxM3a/J4QgG8k+SNy8Pqu+5gdCDE4lQX24PF
k6adhrt72AqDbMqk49QzHVfKN38h+1KPCXD3d0DOLavcygW0OZN2mdYDd+txlsHVsOZ8Dy1FO9bw
V4uDFlz2fxDXrTcok+3/oekCMX4AV+B+b34pGUcO05a49k4T+P9eARU2bgIRugvejZ10jrOfbTlW
jHaN7G9vghUqBfTZKGp0CCW0r617fovSz+hwES7ooqbuD9k+RrYzOBaJ6+CSQBFw2U01gEDNEN8y
KROkeQQElVAKOlwvQ4XgtjxlZWiHDhFzjMJ2fA89JAhXHveRciZ7Zlk4Pstp5sHIaF7Qiqu+hRb3
YI0RChV7y+1kzE/F/ZM0xVuYpgGyoi/MRw0se9zfc9+BGQJFb77IlQGUzPepgRlwPYSZvmlYyiq9
NuUZsi9MyiIyA0FVdlEy2mUtkq2tPUV87Hj0SWjDdqudQ9u5bt3/YKJ0U4Uyz9EQP04HidxWB+Qp
wbZ3XXoxmo+a5PwtoTnyjUoMwV77DomlzfxbzlpqxDzdu2o8TT3Z4p23tAmbK1OLVy6jdteaI2UW
mw0vIucufjo8Irh5HiB1l4kA9EeLvE87kSTJvkWpKMKy4pQzYYNj2Ab3epx3Z9JMLh+I/mNeiyeq
T0tuOwUVkmVjr5zTR2grE3w7lrf3MTpZSHuxlOASKUyCXOhe/sXDlPZnCzL9t2BEnN5OVQHaM+wB
yHssiXMQBc1E9o08eHLXWyMo8ri8XsIak16Yh0rbvhxpykrDqkXlUcWHJoI3xgKW+aHelbACQyfL
5tQfDxnrq1/o94WULZy5jLeWc1dfQpg/LcHJE1Z7vQ9/AHuS9Rxiks1fQLe5RppW2+mfwkw4Dc18
f/J/kQHdECUsDwidhAWz0GgztG/44dUdD0Ega7rOGgeuAnREgVaflIkTZmcYjrwz3LJNqgHWa7+Z
V/OdHS857DG4jsdNME2KX2vC8xfJ1bk1v/K7SygetsdSO0491jRn+uKDnLPB5UoElTO6Es0WAmqJ
6AcbGl8Dp7XuG7hw1InawVK/cUfeZ+FTyRSR8MXq1/POYUkoMpX5S5jWhptDWuNpcvXyMPPjPkUC
qtN7y9nDlMFCgwI/8Ly8LH43nwd/H6yxRJauTcILQiIYBdQQJLEENLrZkSEJNtmiSmV53ZgVLaQc
C+1+8X+U/89C3Pb0JQJvlUW3e2kgryvI0OSQz61xPmYLE7qrpjVV2+p4J9c7YdhE7eo5WGE+kLT7
L1C9Kx5y5lGJhrYwt5MrxMCBGfJUaID8UAEICo1YXxZzYORyku4mTnbYvjxqwyk7zSkLdDfqSXwy
GaWFHHKp+2bLAwrqD7TPgFcyOXCCl4IbBbbqbVrCyd08WRRPauRFQKY2BYdNnHGsdACm6m9hHzu/
Kt6XSWCvl1PhHVNtHK9RpeCrOSDwiJpwOIybkV7ZfRpby2EPFKDxLLEkDNIkfj9kevGIsB727J+9
eBIYkvZGx9M5n7z7mT/gEtzbFsllUEhrmxmX9jPk9i2KpOqO6yDL0b/8S/4zzteER9ODYL3l9FKz
YOVY6LsQ0e2V8QjxWTu/L0jz0w7HgLV4wPBpgXg1V0NQnxl9SCANJfOYcO1HZ8WjaBkTMzNL9w0F
HAnjv6ggbM3wuQ53FiwI6Y/Kx5UawbxAMuSd30qcjZYoSdtFKyfqVWMNZKQiwwxb8GPgiNT3pwEk
9OLAd1gcUM2dD5MY5KrgnQLIaPiNTueGS83qQuneTtDrOewcrZSp6NHXydF9ifPbm2GLQNDSWIDv
ls7jSQqpK6N7uJWAJfCnPOZiF3fr7YX58eAsc/FliJ3Ex9iDS9MQcu0Ef8XPtttI29WTf0NcOpnW
ExdLHs9Iog3HtYwZeVVHYekAJlfpttUE2zUjMElIiTflLIaIpAQyQK983KBBKL8fXQZ2DQ44YF4t
d8hVhU8Zw8a53vASVMz1UiGpWh1SNoKYWVaV2/9FIT/sDN6SK5ePi/CFXYIuWqRuxW4nN4FC2umR
vSMphYtsOgm56tSVvAUcfTitMfSCXMF3+UIkGxB7yXAn40Z9lF1aHnS/tkBx2dc+67WR0bFY+w+H
5MZm9P3F1IC7MHGPseyatUJV/9YbTDf8YHiY2Lc6rWwHTYKvhAFgGn+jJYWJYAHcXM4QPZpG+OCT
NFsJRw32IrzJU9VD2doze4dWh/ok416DxDPlcnxcMBlJujRQXRDmBTk7sG6iCVhxdPAjt2ubqyiN
FyOshMjVv/8CZO4pbdtnDsAbzYjHsD5YkmlbyLQzy7XJ7qjwYvNq3NhnH17N6U2v5NFmFlUZ44kl
sHshf8sk77t1L+wjjX3QvfTZq6zZJKr6CW7CXWc6QxL4lM0tNXymqkFtKT1ueoSo81qR0jIQUmu5
dpWyUJUrXY7DdJJPMETqMZhTavKpenjOtClyob+QtpscFy6PlYJCaEX2HrCG6IvWUFOQh6+Z0ZW6
EdaLyO7WSBVtiLFs6crwIeievSUfVYvRd46pF18qU5J2yxZcinQqJ1Ifj1ALEzbIrt8i6lwxGRo1
XcuTrm3AiwJ8YUxNrtldTH4GkHWvm+UTuDQ0hnWXSvcS9uLVHcwXiSjg6/JQ+s9MkU5knT4Fg/4C
D22JYkHCnv/dqjBRzM7tCZ+DM8JRKQ/GZioEHsUxDnMUDbXZlXLzv+8oIXf/lsdeHbrvohrCpR9e
QwR3tM+UadJkdsb+FyYyGqZMVALN0C0qIM7AjKQppkVZHxWrJH9YaBR+nCRR2g5wZlk1HydCT0xk
VlJ+wPPt5RlH6H5ID+LYghq3MNjXjKENjVjHy0DAB/pSevKQf/skkGzyr79WftHxNHWa+T/3zNG4
FKBzgSYQbCMSSkY+xELgWLSUj9Ahx8jRSg4vdXsBAfxudnM9lxDF1WKUSOs/YEAenhRTqL797+9f
7TNzy0kU2UkxQkx8CsA5tAYswgE1ETBf2oHVM6sPEHH12B4T7ggfNsWjwgXI8GGhRGqHCPLIJL+Y
nXZ2E/+9qi6LNvLY8p+EbB8b2+iKGka/w99WwYiTGkkcKtkQbCS2Dyo7eTGRbpc9CEtb/Rmo68W3
KhkAcjEYD4UZn6GwBJZMYwmUE1KTPCS34xnXZDv8LiJGz0LKaJq1LQdYNhuX2Qle4kN8KRnzBuPP
CbDj8NY+YWpf0tNoXHW2q/wVACgV/fv2symTo2GC5Id8uiQW8eETG5ai9Jx5xYWipdMaJ5mPetVy
6579h5L5gXZ2iCLNUmn8M+wSE6nZogFYJO9onZj6AjF4Lknf7Br5OpEmA2iXH4OKX5vTGAit5FD4
5al2j1M7u4Pu+lp4OItODDFHiqraDui5495UbQszf5GVTzri3fuVodmoBIStwOhd2T63yOU1MJM5
uWK6FQQKS3bXVUsa/rew8Ver8QKSUJxpJDjIyfS4Jlt5H/GLSJi/4BL6e6uSpDnmcdqMJ+UPsKAz
zqiHpBoy1zjV/4XTCi3drKD5AGBTVdghj7sJG8kHfV4kMZjVUdn5ZATOE6t32j8AnqFYaNA3ID2b
fp06t0EuelxMplmAyGcQMDBQ46zTHRplP0CQb1slAH386Zt8YXr91EbLrNRXX6yirFMU3YwM8sm3
Maj69wg5XeDZmd3tgC5OC27PNT+IpgxXJumiWzMCcCL4Hgr28ekMoOdgB6reRjoL/qzrSX05mUdj
8IL/av/FN92kxkowdSLy2ql1tdDwfxMa77/Fd1ZxxTQFPv25yQovEMgSy/I038/wZjaz9pnlsRnE
JnrQmajNCVM5iR4iq1XB0CE4Fu1Gn/mBodRlQ9O53Uj+lfBju/0AnaPAaMh5kM6JBsPiGTzZPJlV
JSEThuEVN6DOkAK9wJv2hOg+HQQSPTpMox3+lvTbP6N7j9WhPWgcUa5QmJvj9XFZZDIbLbNMN5Uc
fRUahGeT0H26sUyDeYG06yeTTn9R8wHuXc33E/PS/MtEBjHTkTws0fHXP56Vn043pHCHnMusauqn
YqJpt8bBJAPiP/MW1yVMlcpTqOMMIAmKC3srqdjkIlESViCn//TV23WtBpj0EnAkrfm8fcRcC8sm
mxrhxmR7jaCYeQvZlfKh0khdikbbQJGVyeMG4xUWNuys4sisgWabR04M0LSUrzzwXR1mYQf6954O
Vz1RSmMCLqVSgz/F8hjCQxGu1YDbuT0qiut6QL+AhfEGuPPw6HmFwAD9gtRAvvaX9qn+TkNeNfxD
G504yeeA80ykh7Oi2LL3Ld2dvfTdo4lYy+YxF86A1r0HheqOz5mVt+x3z8pIp617BptOBQMN8v6c
HDSJ4YZAQgy9Cyzh8TB8pLqNt5CTrqpKCU97r3rKI0kj5P3wdlUugHFBTtcNipXD/iKajleVNpu4
cTjhfUWljdshnpR0vNtsKcz4F/N/oRxFsxWEOSOWHBuMkddQ1P+eHddmUw4LJDDAvT80Oj1TUYt6
1ZckXVA1XMvmf/ooA9J3dAtV8OwjrD1B7CQZ0atZoMgEdVvwfFFiiukI3Yp3C575fY2qnypvZsFk
i2Cwgo1KzgjFSCAqSiZLI6UtbdTcwpk/AsTIDucH+0zSs79L3cqq76XCgPzb91j0pF6WYUW6B5XJ
Hehfh/BjX5c5GB48chwWwHxk7W2ifBHVf2tVqbFmKScPYw88Nq7IDXDnLHsZbzdycytzk5/TxUDc
ycCm+ns1wuUZvGgZfuy9knRcsviaIOr7AZyLoE7nwGwpGRxR26t0iFaSOz3nDRp9mXs7qDCTtdoS
M7sdjSHG3Cx5dohRLPatTCiSsN44lRE0DKIpUq6+Dv56lMlXoNjszC51U5FQvFr4lme2ESX+aqlr
k9SVEkdeCQ2Sddmz5JQ9T9n5P5viVMaQcucloYrXY4DpgYsG9+c9CtmTjyP2HsdHmBZBinj7qkRJ
JCuwk9pUkzBZKZJGIzJAhNZfh/7c86eM/t/ty4r6O0HGStmC3WlMxQeZS6KJn1oxwIJRpHM2nyTp
a8F/3pQfi5HStvOJPY2jN3Uej69zegHhbnmEyqE7y72xuM+BcBUqHgDYveYxBfHh3vIYzNVvT1/4
wNQ8XXmnZh3l7/c/Ib3tTP5kbzfCeoa1kXJoVlnBBdNGtnG2oh8T5eWj4/8ctl3MFGwKc/8kvznC
1lNWGasvfj1ZOLSbyHdYV43alXi42c3p2OPCQu8Q+gVjadLBhP78zPju6DujSZMqmTiun2y9RlO/
cRxizA6c8iMLJSVI++SfhGegKFkz9r31JhnSvAA0NoVuu+xUWVk/JKTqI1Fh+xbsPm6nkNcqQf2A
kSNHH2JCcnOWKYexIjKYw41MNbDXFCjU7cQsr0tLeekA6smuLvHdFGaq2zS39UESEYx0hCkzGBin
vrOC4CGkunPIi5w/CuTUb8EZUoz/wkXIN1FFQFWZ2V5zabLxmEm+kZ3A64UZUb52IozWpkWDVuDw
zE+hN7cEZZ1HnIQQ9XaVpAx92R7MBty/0yo2Wccmq7LckAmLY52t2Po2sRZt4XLXzdW4VMicXks+
rJUnPBFwIwkPr+/D8sXqq9OFHFU8gIm4ZIgZCOTx27Gej13McFjjZtm/l07mE5eFTQkPh3tLR27u
Pp6Nu1rz1PVAeGXaO3RFuvrXI1Y9mkKziTc9C/gpGLlPdHua/YcnKnCgMeaTalbWg9rv3cFhUfYM
ln3SXWRLhk0mDvu+IM1Vns/L0EkmEoyckllLwOrqSSBiYNjZSGUoNPFJTiHTta3IcxCM2QBD3vTS
pjej+zGN+Mm/JTVCnYgBU5hK3a/q0fzU9vXTBvhzfJKpsqtcKJuhL9Pe8L3EEBbNzd2g49lrTnFl
K6cL3PVFQpnEMJCVz7arZpfnVaqXI7hydkxILcMBlOLLVjeHM0u8MWKIWaTx0mROtC18Gc+/C1xb
3enqFuQyro2i5ooRYN6pg7+SDjLx3xk7m3OnAngvMXTl8BmECTpo3llX2wJMQhCh8TcmvUv+GaVI
uWXuRi8uVfDXslmXcNPh2Vlb0W6VtU0Ys9C7FOSIc1tFvxgGfcDdeYiZ7yX3LsiB6ao1kHZ40b1q
C2Uo97YGi5YG9PQgIl/qgAMsiH+VWgtocQUPJnVXLBYLE9R9dm8lQStfUsllNZf72zp7m6BpVjsz
OuAm71qi0orQErSwkHZ6nYKLzBU1ZRcSw6dgJVSPvVS+BFmOO2SMn8ciX4VVZRiR4y8R4A817Fh8
t6jyNq/cbsBDuTsux2+zuaTo2Xq54rTJpz0sJg1qoDBn9/32WYU2KFlEf4GQWap//WbVo/zS0Ebe
72qh/Khgv0p5TGDdQAaj6VltcXUu8SwXKMj0pd5Y0EDtceGO5ZkEAF2nbg5tnAUlA+CMCtwelObN
2kz6CnvMVpf6vzM68MN3D3eScu2dg/dMiZ10Kc4pxuP3HLfwFpOjtOzY/uIJJ7M+2JrNE2mNA8c4
6JJoFBkMUTGfI1g8Yx1oFrqbL96VO6TMAQPJKZ7uKfM3ylOO/f3ufvc270NefJlWLmRhKsaAY1Qp
gtshCwWw+YkGIOWkSWSEMZWxiUdXTbQZVl6H8fdiP4FpUU0WAlgVUzINSiCD0WejfrLP1ndkeZSs
o0H1Uu+s18Cl8UMXdI1uUQUN2BaUe9Q1B5I4VqmX1n1NqVFFyMfJZOlGVzfYtHVutEsc6oYi3AYD
ihvRUHHCQPhOkyb7LsC/A1ZBiUDXJQSMjCa9uZFSczAQSelFP9LToeYFmvMGtrh1lGvkBk5oTD95
F2Y3V1Ws3JEmP+0Qgs6cnlUInMD+lA95EjtSDjU4CZZJXDAeCRnOdnBAHS6yuZg/e7C4NEvjHStU
xCbitJdDFbiIHekut0yfmKU1kupe1IFrB92i8DIg0D6tLrz7nNjr0F4eT0dVu6s8hIa7CO4NBLIW
fZ5odQt38Uhz0Fpnnb7nks9JM/uKWwjG0tt1ghrjOF+5tGfsQzIv8DYo2PJTeGI9FkSbZFlKuvwK
49NJEpn8aGbpaNWgPdBy/hWI6hKgk8zOcaZnI5dLvc7YSRb9FCVMpJ8h9DOlr+7OAp72Wju+YKXi
OR0JLs+K0X4WelZQVl0UsSlWkstW152XY7J7pr7cK2WrEhNs8fNlQt75UvkXo2gFU7sbnZX5et7K
WcMjnMqbC8IyKdNfLJt+whu3GgY56DddCj9mdToGxEstp//E0g+8G9Dye4h2RIgVlFQ0yqRh3rZW
f3XyYeZJNWLnoduOSh0h9sBlwh9qfB5rpf4dAvSa+mUMP+mAvM463RLshO+WTQa1pJ7VYB/hggG0
0VmU0HyCTL2T5qE5mK5gstty8h+kq2Zoveoyn29Ui7IETl31+gYI4dlYU5Sp4NXDWqzaAvxw/GlZ
Fd8Ps9ar2+DsU2VDRI/NR4WjPGtXgu1TzE/avcSVbrFYUmbfrXX98+7hMFeeEtZWcRAYCbNg2HjJ
ZHIzVEffltg9rEvR8HULl1zvqi9wVhwG5OOEitsEom86Wd4fsfx03OuY2k3jKeUuiDX2VmBoElPS
Xm41Y91jea5moaL1Wyh+aVcVvkBKpOgQo327h+kXag7+a8oV/IfGCwWNYImFFLjSl5Bdg/vrrjCT
RcyFCjSpvo5JUQMNUdRjKmDFYzNPaQjX62n3ao/4Jn9DXwYMJz3WkoIALnzsnpjRxCWla7Bdb+NO
u8XVLDkljF7G6uXKJHXPplnyGc6YcKW1vzQEXTVXED+Rmqnu5HgjGJ1Ax43UMRCw+F1PKiQry2LC
jFDkT/EK2j3xmcGDGQhQaQUzI5yFPgU/76fagGkZYz1VysY3RXRjJBz+qd/g7LOayQCDaQvUJV2v
cjVMVB3Nc5ZFd6QSEX1zc3C4RGwz7pPtxRwP01qfHu6X/i3GJlL+SkrbdKqCjg+xDrZ2sE4K9V+z
4Dkkcltzc39DPVRAJjveg3/kD5cEoq53WjRxhEbY3MnVH+vqx8Z6poVQ5iWXwGzFWw4L2DW31NtC
BOHAPDA3ZkDPS39uXKSJqNwXD8wDAU0A56d99ASzasOYXSicoP9eD+naMKEM9ndf6Rdzg9uWP6Hk
JkSgjnfzicGvmJRsfASE0uQuoRDLiAokcL2LUV/kGJTpP55i5khyDnA/5s4Oy2y76TA3wpQf1L2z
gYXwCI+6pD78m6DZfXlv/eLu3Wl/r6nOPvBu47/l+VMgRSw58AxMnT+9uSg19UW7FcywjV5ji1uS
JBl091Sc84tYHIEnvDdxgX/0k2Bm3xcU2zwjBVDT8J0VwlIwa/29GZIVxthIjv42hcE6mR7tzme/
CRUo7Lw82YiUKM2OImu84J8qQrCdqYdUBiqNG34GGTSKNyEzZfHjmgf2z/crq/5pMW+5N/Kj3hOb
HtT+qWz2Pk0ZxWcrzMT6UvfColCDoZMUke9NUV15U6CwLoKgKro9BjeLZDBLzjeOfrFoDciBwAfB
4s5W2JSoU3NlqfzIvzhfQYcL5kDIzJMbp7bycQo+Wkj7Q8RaZCchNAaaGB471pYho4R+D5LLwcGG
EGzZiHBkUx5T2L681JYSoO2cCufE0pQQ5R9pyZtwd1JKkq24tSEd5kQ+aJQ+4z85BR2UqIb+qrmu
lMONTipKt4714wssSg0QIBEsQ5j5bUyggHnpCsUXJa3iybv/W724Zp/izSY9qF7VcaYZcvvGHyJQ
2sGtbyGrxDs3YSDWoHeOHXL5LgNG3YsCQmBHsE953sdtuBGIdqGwleqi1CHekDW5wvM6LULozK1O
xSN1REMNRVSwDFHrv5vdK39wpgmGMcnWXfj/szgX3XmzuCroUdr60XlSkx2qeTweeUArTVRi/Yx0
UOUmqS7tjJkZaE4XgiLFkJigLgb7Owan0nn3EXR5tbwv7Ab8YSZ2cVgLQHj1p5FOagcNwflYSCGr
sLoHZg4C44spCH9fzYHtxuvbPNuIrJrOitT8aE5fhgSLJ8INnruvG+jrkmQ48NfHT8XV/Dz+4Kng
qFDIWC1wXzPXWdzGS9rxxisjTnr571lxjFIdOdtaPbeT4D9oh+/OZtPS6QLZaXsPO4F62cfXNFVB
0rFGgxlUXyyrSK3nRSmt4fk5TZlGVM4b5ZSl8KuafbcpIiC0vixgLsOtFeCFsWFTXUTrn+S9g1L3
JP5QA6A3/9F5RpdJVzimMzKzB9O59mQAPes+OB3cD/gJqbuMBhVEXBTUyhcClGmK3EK+bEg2G+H7
n21NbSn224zttz2ZLAFZY7QMxmW8kpnLmkB68V5zcVDnVGVJawxxsQlhv3zYBw7GUkYLLFVzMWGU
FguT9LKxmH68/ReKCnLLaExUtWw+qAL9jmhTcub67dG+30cZHQV4ccHTLrcpMHnZRGF2IE70XWuc
UvPI94pa7ElTnTZbTy++U90OA/Z1jG2KXHiDfMexCdvcsyZ9iBpYbJmbJWv29yeqbySK3EdGoqpo
Q98ml0C1fEud/7FP/eZlbFlqu2oTJya7B4vnc/S8bXN5T0XO7k3nZ8DYACTB5N9rIGBlrXzbsAj/
4RDSgLElSO8o8z1K+KXuTOt5AkNhuO1hBYmnqYVF9DRZph8OZuPbKhK9eElp2mOouBnYIrTEUGqC
110efv4W56cFQYGB2aDh0r7wN3Lkdu9htp6j4n7mvHmTaDeSJe4YwyW1z3VSLdc4dhTuKhbdjc2R
naKvLzxJxV6Eorxc/DCz+OzAnXxdG7niTQrc8S5YFNd/9S753cZFX9661wS5VcO6kC056TI5eCKV
wAfijEwS/GaDpqGoXUCZWnKLuSZ/l9UrxarGujWt+nEmURYdU72waZdzSJDcGZ6czGMkcEXlFCRF
0eiPMRqTJiMjhBqzt3KYeSRy1ZvUQgiYbFMSiVXF0AHRoCcvP/Zd46QsOOQxLm2CEVb9HyrqXppg
ioPNkbqAXQrjZpLlGuCljRTKf8tq0ruDSo1EirYm/Nj1QnLXwFk3ygYTI+wvr25PEB1cxFMKBL9U
twR7nNrnfrNcjLxLeJppEomutSDvJ1x+00l9ZRJJndUX5Kxo8+GdvVrNmdxr0LnYDPv7r1dkoQOA
/lUqBIxO6Rh5iG4PIXg148anviguHogRG2JwJB0s3TDeTjHeU+OBydzmRgEVQGd4+sYXwmQ5//gb
drq6FEAxjxu9QI/D4TAlxA2atfb+7UloQwvjSF9sy/WhNmCrAvJVr6uO+vduhrc3PWwSJGxDUhhn
7o9XEjuqkMWtSLLTY6eAeu+DvoJPNqa5TJHEPVqishN+iTec0s1nrq94DvuipGvFBXgKksT85yle
rtc8EvlExHXbBZUE7fji6BflZ4uXWMJeH/SRgN88V1RjgYD/gfeT2sCY/OJPJi5yru5J99qnFAK8
aOgUFfLK6oLH8XOpC3VXJZmy4l87xD+ihoK0Zvn15taJcvpDet6ylhAzgmFW9Cti8FJ7Gj2EPG64
AQkeLh89ZuxKl3IhOzXXVGC2ZX9e3tqfT2MrqF5A0kF6rRIaTtpOBu6b3QkHrI+a/6f9+PAnOSJ3
hHgQ1TyyB70XJ2Pj7Xp1cy4J7kIwr8uOi2JzIA5vjbmRT2NhpoB1A4y13wZb+AEqsxlDjHyegju5
0009xz43CnMxY3VVAZJ8y+GERRszgFO4Zoi9JKNAZ+8Q1u3igTt5nRtZHLIWj75FsYgPY/hVJACj
jovjbRjyWiH1OOjOA0Uuvz7krlCs0qmkzp+Gnk2aCOvK0XneTa3yWZ5Z/YK01a7/TQdKg0x9HHl2
igvCioRjUVHddZzb0YWP0aVsJ80hnWCpVtHuqN13l2j2NMkSbb4rE0HKS3e7Kk23yhAIQKeWk3i7
L6Uf+4NvZdJMRwj9EhsRFvEkxRMdVm9+ojSQQHk5NztgGn+c+7PqjH37onKuvnKT7x7o6Qv4Isty
EctVXEx+xsGS0+hXSF+WVS2mFYH2aP77nVRzXHd2bfRhSxe7JZ59vPHszETtX+YCI5szPO20WoWP
5TFYtmFDZN/s1Cike5q3hJKSUc3Xh/UNSQADedAy6jzjZspOJvLfl55yU++5zFqqc1hKOa6zwp8B
xlFwyzV+vrwCFwf27T3b9h+qA6T4c/HUCnowFFPr+Q5VVxX2yqfYFWv6Zhenll0c/WLjkwv+U510
Ty2sH2FZkgZCpwwYEo+PJfNu7e2hbRI1GT1O2wghSt2YuWSUsr2x+ATp+s8Y2PfAltBkxAyMriEq
a9cllfZknHGU0TG/c2JH7kUsxJG51oDGplUET2gsOucSPsrWNWZct1MXvXt2UhrzIitkvQrMm1RJ
W1Zj5goDrKTfqRq3yvbC0UO2AgF4JpWgzytlu1FZTDmAqAJdNDPJH0wBkqw935K4WoVuBmq5LFSx
iuZqao/pY6vO6BoJ6RnkvE8kNBTgx9qjhKvv8YD1RmISKFKO/a+FJt2V4mssu/ahGNA3vnCQVc98
4OVQaPmJtTY876KGickfybjCT6jMwapy31Tl5OOEGj9fTDwsUKEyTjrDSftRFgJUulafFkHAVnYx
VpLnrwupf+Nn1xB3JAdrRHVNTNmhD6uWTl0w7E31Zb5U6lk80aiXzYxoOHEXQgJmSpbH019ppWNs
xJlNGIS/TltORz6l8KokGncakEKzb/gP2Uz1ulgv6tkHA+M1GA2MpLr1Qz85mJmanFXlKE+5/IcQ
GZCyIF1YwD6zwMxxxPRQUlrasSwG4Uft2PNFNlFqWJxOsKNzbmttfkQTaqOmihVRqwcRrzx4QyZ1
sAULHTsuwJiX5YYalis2NwMdVf36rVl++2yvGxXyI77xPtWTwCm9BocEeVfZtNu2zd7DLVoMn22O
Rh7RQIzquI4MXXx6WNHhS07G36tEl3IIvRVwPqoXJlybK5o0vV+XH1v8JUTADB5Rm+C08fX+KKlK
ZZDCnQmRgZBV6APCe4U7UP+lClR00N6EYbeHCyy2kyIlKQaBDrzEnnongOFwRdbliRYZynDUGHsR
M8B4/PR5Fxs1QA/oynWe1i2ZI33QoN6bQ4FBGbV7NHf4dQZhPfgJZ/IL0xMzUi4dHoTIC84EA+Sj
K8cxWnufuzV7VNcHWRmoY43LhpPKpPPOiGrzpQ6duL/B/ePGaY/GKf3KvVfNoUeZaOGY8YuVXxKc
NxxhGy8o1XU85d0EYvcZZowp5VM9USBVrG8ZK1jQwBVLIgGXySXzV84vxq2DYfFtqcSt6o8385JN
38onA/DjAaNwETYJMtQgYtn6O3EGj4OedjANsRat/DYNGmECIM8lboulm9OH7nPItDnJWUBTwGCj
HY3RirxGQNTqOACuwvhhjOzDtYzYRs6V6od1UmsxyuRlKigD45GYAMqAw92Tgs//GI0hZNlXMmwo
XITwpq0zkc7qpULztV3HOsteoPLC7atgHH+zugEgFRPi7wCPA+xA0BYF/U6p+iqjNYRw3MhwnisQ
WY4d/RqOoC8x7k2ijtCvpjgKHEPxJC3/SzptbvAKRvDlKbEPvYf8f34gjn+azuVkv9gV1q3Ru58C
eBDmwOP2zELJRY2iDui9fCgl8RWMMSiJJybAv8AM8de9UxSs3tcz/nDWVb56msyqQN9Kw84Iv+rw
LRvh9odKElU+jzko6axI88UThtbPFDvFI42uv/BErQXO3GIcy5M6jeFbIcNnq8yY5RLfM37saJHM
LEhXDkHL6Y/NzLJ1RZXzGb3o7RvIGPmtqq87Sabv74+ODnsfv7AGPitlMl1L3/mP9wdquleSWjMa
+sC3xa8rrkisgIHVd5e36dKhoOSmx7iVVWivci+D7k6z9VYTL1SmgUsrU6T4TI+0ZBQUms85IwTJ
D0+9XUtgpvAAcfBwmgqGyCeJly/IJIu7fZnQ7V3uzUy5hNvlaxHJ5PrMv49f2go1bfoWuyvwwL8I
KWhG9t+YZh8Gysa6b4MNu4p1HRK6R++5yCKK2gzYk6areJpQWOh9z9/3GefOtvlTcH6o2wjH0PHh
x/MuPAXGOoHQHLvzjQ/UjodqVIQlB+hpzWh/Z04BxTOWudbN8iulvP0bwFyvCvW0IhppyKj39X5l
R+8Ss1+RbODCPsJWeLeiqIg4tU2Ra9vOqRvnEPdUySfpAMrgHd0zHADHoX2D7uLKOxjekGyX+R7b
rBq7nRcjtMqCCo5cSHh9ZpE1wWdep3RleB8A7/JdNtL0qMp4czl3Feh6Y+RIu4j6q4F4eYMxV5vP
si5DD4F7uX2uLrOb/71DfnnjUC3owFNTWw9IvJM3Hm76tIta8B/wcYwGrmGR2phQclHH5ynkeZ6c
ZHyT5leWwdqhTjsHOjIiwpoSZzH0t6RLmgQPn0EbWLnTOZnJDk79h87eCG8XBsp28zNcr35FJx9d
aftD2X7oqK/zgA9llDjRar6t3Z2nrO1OxG6mHq/YAqOu4ZoN2CyUuXiV7nCZ16RJA1cSF5bGUAQJ
O6f3zeCEDi9u8Kk5Wi1rt6rDQst1XIlVywSQgq4+5eAVlvtbNrs+CVrqHgp71DCAlbyS+VULk2Dp
ku0dEDioh4RVnM8V0n+sfoMf2COW9OjzHPVeppRDau3VmyqbFZGlnWTZ1kvJP8fpDTC27gyZnac1
dxGGRyx3M95pz3MGESRLDlDqwG//vuqgFu/VoDb3EeKZzk0VWSfRaPo/9f9ve27CUaLtDA1O3tMF
rx8zmNbNMBah8BOVYkwVbIVydUEdGC3rRSvvshmryxRsJx4/avSrM47N/dhkmtl1p65aIBJ1f5DF
F0foS0o7Mm7Bm+ihWgZ4tSTB6tJBXp+s0TEfLdUhAj39tTkOdtFJnp2U/SgpUYH858vA1WSGbpMN
ab3J/DP/KzpJS5KCwdVW0FNyPsODF60qgI6TsqHFYG2L7h6hfr+bscJu5/7ZmZzrF/lbtDAUPcRx
1XSG5IBgryL4KNaDXSzb2+bE5QT5Xk+cbpVALOniS2pEPZTWPYdT9TllmHX8jpbIgafZhrfMTlBt
gHcOGJMMeioTUaQ57VT4UNiYjFJK9rhib9QnLi0hh0tK7bXkpe0tK9eFhK+4icuDW3Q7LbYpmwyu
o7GvvHCirns60jl43D8NMZ6sTipsrk877WwgJThfUNj9DSckPiF7TrEIxjnHSh5bbbGzBQ91JBgZ
XRTEHwHx1/HUohFbi0SpQHET3ENEYPFcFHUs1iXYJOGEzteKV1Kd62cpwzqepkMy1ArNBOReJHO7
sFIZZa1/SkeOJVPbS8Amkmx8Ct4F7iG30GSMdH7onjsHpneqewRXyOIxoQbmYrV9yZzsaa9efi1P
95SZ1YbbIt0nXQkxx3SkHSipd3Oy41O+YKaAaRNvqRXfXdt1wi3Al9Xct3qKicbJjhP6BjBT4kvc
hNsNUJHCtYZWloFnj/opbA8xpX5I8g2RxrvEuGCCh0Zm5zxFIcze//EFdG39Fvk44wabkvg/N1Kn
E4N/hLhV+KfKuD2Zi3LkHRe13P1W0/F8RFl7x/8E6/TCRuTT++sDsZh7hiC7/0/g98CRMneE+cR4
tH0qpxE0O+HuvT1boDv1TYhIqrMFW1MNNWWXOhN9iiNO/erRkJ3myEjn+Sm6384sZLnfgOgFxlF2
Bfun+67/lbxTmPmb4JmhPqRQSYJ00jpm0d+h874e3i1iQcvgdpeB1PxvSvy/G1KVhIq6/9e7O7/k
NiDrkutupLfKTzyH7C1hq4gTq+y2K5vltGx5sN7e7bb/VGGq42wHOaVhC3uVcw3nVGdruI0/cSfw
P237qG3zwSCW+5C34QE8nZeW0cfTL4aXzLL+Sw+20Wo3FPr/VytTQlfhbNxVPRmHqdNTPPNZoyS3
brPZEyu+mp6n7uuWKdoxrn4K4mxkyW69Jyo0tZ5SPzj2F6BrTLKmWajfUBfv7CHMf3jZ4g1+kLov
5S3RVlo4/0E/PiwOxfWTEkkaGqbKCKjJVPswvBv8CRT6wNQiFcIhHBqMyNq7NwfIWYHEW43vkwcn
OCMd1hYFKxEs8JL9n4XrQ3gMSJMIKdUp72Kx1OuNZ9xEdz0ZBNY6P7b11h+3OYEMU1OF4OaDAdcB
LzdMc6XWAvYE1hu9Y9AjhxUDgZIUAvQFrqYcduiFghtaQMgs999nGA139foHkfFD2D8rRDi3S1AW
C30FuCCc5NLSVFUBV2RLDMid4K4CnicgjeDyaj5zfX9bmBBqzuJAh0wOa8Yo8tUZ1Fd7pJ4lcG6T
8D66HYhPeq7oWLXbacevGsu0gfoLkJAr+7+Tt5GT9z0lxU5/nMoSxz1LwF9t2gQdcFwaZuJQOgOp
CIlS3nSt5M4+pWsqQsFTfnhWoZmQ3DGcsnBKX0fpnf7kLcBm5Es+nls86o8ZINZRxlbGvAZ1bGR8
kcCkSDrJYDVGeCUm0SM3KIh++5dFquNbcwd950XAVHgL7i82/A1nSCfTeAk5Lm39ZHuJzMiDmHoH
vtqeZat6aH5ykZTLNW47sHNVQoysf/Z5p0gLtYV8BfsoNdPBC8jPNffgAtOwRI0+8nEMs/NxK/M1
YmCY7S8X4cOAafANroJQQYQ3Fys6NyjS0HR74aCtWfEIw7A2ENK3d5b5DVsF1Lzc6BoDqYVew3fc
ggq6jtWlJSWeAm7BsfDpyPWsDVNnOGsm5s8BlgLs0ny6v7mBbN33kjQWUG2vmSAa4HbZivMMLTuQ
R13BlRvAarjoUHVRZQwId+mKG9xCc6y4ih7QL6BGc2f+mrCDx4B5WCZ/UwkbXMg37+xVl8bejz12
TtkraGNPG/7njH96KxDiX5Hx/KFg6/tAtDKVDLJ8Ri6MPEax13fYOuimaTjvdXy4U5q94Sp7wVgL
1beHP14SnvHWJpK73CDwCnArFm/uenvbh8A4aZ22V1kzJLhxUMaNYAhRJ+tucOyiqW0nC7DMC/IK
c270aNIMcw9mXm8JSV0cTum/GV4jxlnPQYYGUnLwaxMJzCQe8BAjSl7fRDmYjqoBM+Zw9W38HUL4
vv8wCcKMicRuAW3aAGGtKaN+d5TyWxp0U66CoBtY/gEYr2vkIr1DgvFW5mnS4NqDxE8wyqJ1F8EJ
J03is9Le86kUAy5aYlFsN682NBWLu3yMBn93cMYLjc5CsWuAcFwnCSraKomYGsUBa7l++Cn5mT1D
Bc+eewv9IkcRz7HcUNnk9XFaDW1FO6Uu9Og3T2sPoFQfc+Ss4CgvMHy6fnKVrgaHOgHWkCV1VYVS
LeINT9iIIpmmCDK8OxKQxOKlMaqFcbSpronFB8e6pQu1fyR2052jRYMjMHUxlyqQPvjTAG3BYzdm
HGFBPAag76nhzVoVrOvaqeghiJG5+jHH6Gb3/E2z1S3yUgWI9UgtjJCMLY//SUmDcLtNpnDIw3ua
a0VaL+d+rwlpBPU3eWTKaNDzKTOH9yUxD1GHl9mp9ATnC0XvwYgJyLPs9k5tvf5bivxCvISFqBsY
ZgZh4avUEPPoLGR8a0CJPvBvz5reTAl+lFV6yg9fg0c+hMOCDI9XMVKjacIKQdHj2sNLEPiCR2Cg
yaNTKWxDHYz6WNwrWCGR1ZNgpTCyijYfnBrcFX718S1uY8BZpzX8SO10eT6ovfJa8YmpgmZCiD5g
BExqtUVZPti4MdftWxw/EGS6SXq49UgZvSRBIDl+jwdE0zutQU43q/c/nknjLIEHfxwR419pG/S6
N80K7TjdEyIFcW4SY7vkdFTfEx+DzI5KfKYWRCDlloJntRWWo6Me6a8HmyWMQrNidYu4fyD9V1kd
bNeBIsGf9vPkmKNXAwJ0JaiRk1iNi1gV54GeeZiAEGaPuUq9OtaOfmTzfIzSUzwXpqXl7QdHN4sx
z9egLBHO8lJWrWCi1SLLzc/Y/QLBPhza7UF9ouqFNc4Vw/9YmQHqCCUaSQjwjoLvTcJky2ebA/JB
rKBczfmxcNaKVBrxJqceTRVFvdUL3U4JU+C2YvnH7a9sqweCva+HMaffXJO1KFiqs0bb0LcGVyoR
aQtvIdKN6SZiQcQHEXcZHzsGDX/4Cr6JFPwLPFZlezmdlP4In536Bl69h3X1FvztY5vdwVdH8M6d
E3CZtLprIuLfUPMiJ6mr+46K9vQlpXXkxzzL3MAUUPE4shRgHfOkADBFKjwuw12JFkkjg8xQ6uS0
LDATEqdNzFgxF7lwowSpC4oS0xHbJoxYS7KX7lDRbW2GwBhI3i4Aa3nbLYXB1fLqPStWGKAt8prd
jq+Ao3SW1KhdSH6+oDs9VAAHrKPfWOxGS3kNu/9G0QO6ueAiGdY5DuZphWeQ9a3MrxpuVRBll2NP
vKluWwSixbop9y2KLjPWKW069LCjZ3p86FaA36UNNbkalXcv7c8Bu7bjyTrirewC467lIaFF56Pq
JZvIyCiEtl/vF7rNlQXED2GQBemz7EUlH7AQka0TXCSwTMj3AWcieOiAnh5lBAFZXRlD2ez1id5j
llSigqT1Yad48Sk/x1J5tdFY53HdiM+6n/3P3jMmH7kLrDGPQbU/zFaqGeXJGjy32NNLmHOI6XkF
etLuGPBtZR8N6mwU5wmKWOf996ddJntuOkxGSD3+74D9XcoX6lKYlCzB6CsHBQdAvjr7KFVZlnxX
r633NyKfVHu6ubGFFfe5a6USKDIicA5SVOm/XL9euU514vxw56g1HMEDahuhFNPxtug0CZXcdwnv
zEiiBJ8Phji/8qnpBgWLcXXgQDhNmR0iMwIt7pvSD5iuvGhg+yGMIYI6c+TN2sh0W3KNNvJ4ejMC
YiKy8s7dYBclDu3odO8VnOGS+bg9V9+DjnnrsUJdrJ6vQTtO242BCIbVlUx/dtv8iLDuIH5J1kWw
jMX2UgLkRfd3M2hGT4a//dNr/eXjEzCMV16PzOPxpJ33vEifD+eUFqigZq2IxvLQFiIT101cjWfF
3wyi9Puw/L4wsh78b/zMfMT0eelYftU0uQPduFPjoNJEx0vVaoZQEvFKTf7gWcBclHmnPo77ZxGG
srGVufvYawDWy6Wy/et73QyGpCFuq9sujmywL2E2SIO+IsNhIF5dtEuj7JS+oBXvGbsW2nqNnNrx
fFQei6d+oFKwKHKvsydYSKD2cDxA+lGhwScVSwexNfLqpJdB5WMP7CSYsOANKYuR2FQ+GgsM29h5
8ijJfE95/Xc2xQidARUOBtNv9yYFvl2dsiw3JBsvh+9ICqmrGid6xw6D4KIdZ7WyBiQGAEWocA5o
tufT8svZe2MX+tg25722axRhlRES3fbcnlwiSQbWAXAUNJow0ITfddKmzbecYbobE93AeW2xRjEb
rn4zJniyBrogZNNn4015tjTqv5Q35r2/3z154cZM6CzCmQptsoiLa+fzWMMHnJNjZsPr+C7tjbYX
brY5Do0kzkkZWtvpLu7JfiAfACxpqqchpVkMfU7rrdomHkXTIcbpLha7x8klHJkF6LYh73LKNxb8
9IuK7dIyzHbJr3Zvn8vWfaUMl94e1Nq9MpK420rF/w51sCvGWHc4BfVxWwnLREKz/mP+ah167Z3u
H+O3Ybd+LGguxttUBpiAjDuZhWn6pWkGiHhMpoVZcYHSgTSUiyirPQUvoDKkQiW9oa/ptYko/O3n
OuLkLoXYPz+XrMpr0ka0F7cLl93XFu21mZqn9jt/E3EE++oZWnpDA1fAw/4LonW961jqsd2LFh4w
bF/r8tdCdf1fBkHlZtqjB8rwWac+63QIJ4D1TraYvybbxEXUjygwMtzKhuc7JfG6D0rwVa1BYtuP
q71E6sE4VJ7s8fYuzoJNuebYpmc4sfnhhV+dKb0puIzol4hBS3fJELdjFmG3SbdG2rdh1aIdfK0B
Ao6vtcgE6BwF651Lx4hfiI+9Gn8JX5JHfcEmN+LiayNFEXJvWYpKOK5okHjWL71xatyED+x90AfY
dN1LDMpEngygPB228/b0KGmrYcMjApgzQU9LjcPonLzLfiihVblnjhzqRfgsGr78yQZG1tPvwj0p
4U6yjNgNsTydwy/H/e3IyTv8GIyL5lBoCN20x3UvAI3e5KsD+A5HEizGik2gsqhbTfXz1AOX36pK
+Tc+3HdE1mz0hmOGkRg6TzLNbZZ33MNG7d/W5AXB+mHOXinatlgCiMUGylGpY1iapBYO/hH1ifYk
sRrP+PVmF95CNGOqlzwAgorXZ6jQfVniYQz1xyo8xV7017ymZilCYVnNLKe2JL+bq9tgNWXjXpin
5mOJzq2qfGOWUFHatdfFcKTB4b9wGqtdOt3kZ7Zt9ZNGU2QqW0pXFaDV+6nNsqpFHdfZXers0RqP
jWlc3H55cG/sCzjopElGVw4PPIEEyELMhUU/kEUGsPqGFCQOear4U1A6uc5axMXrQQKxLp9dXc4+
1YpZKsyuvGqK/hsWH2YUEywzC/2kQQBHD/m0jD1k98220qKkEQSOipykJlkOWdyr/3n1M75ipDWz
Lmgf92wZlEXS+tzt3d+djlfMC8u4u4tjUmXPchnlsdUWJqkeE2wPYt56H60a0Jt5ELDELG39etkb
zu2hHT/TSJQTl6UPNMqYJTJVqa31MGHgK/OhWf6yRGCWlSDsZZw3trQTxlCXP69RVpi4WeL5PoUm
FKz9qHzIpfTICYgM2y+Ux2PyU9PWYA+ikj4GVMyqe2Y9uYceggjUjaPdkkQqnNHL/vdvyzh9i2ni
mwOMzaLE85gWqwROVQr0GWXVJYXIMd3jYTueHtdselC+QnFUVgM+cbR+QsngLAN4qkQHKzvcBYsq
ckcpRY56oMz89ocCQKnOd3DNw9qjoBDX8VIcJlOSGA8bUFeb0mUqvjL0t0TCD38KbHsh5DSZAmWH
1R9iluqedJLvBwKRpI5XmcRk0vehmilznDPI+tjuLwVY7b0k6lXzXpHmT7iZNvn0M0LjiZ2/0C3O
3CeCdazS2QiEpH25mzLFio5HXGjXhQktImLAYO1HWykWGee2YuiA05rH/qrtV24YcwMk95uhGpbJ
he6Zgj/GFAlrPdVLLPlDk8t9BH6zCnI4oIXeqEsDtjb73QmOscVzt/6jUUER1WUEPTuereBGpoa+
7ZQQDkv+F1pNX7J94wdkaMyRi1avN9/IbQSrxDG/u41l2A4A9X36emFGzjEKtu95o5CgAuDy/aLA
G75kXlgtO9zp3w5m24XCOEl4LxkRUctz3i++66VhtslfwV2qPJceOs+M/dHj1iiIfay0zi+r0oBs
HNBkV+swSD9tvIt+GC6v8A9Qx4w667co20LB59UTT+zqtcuuObnnqCqUmd6TEsTBrPiWRxxBHkH6
/uAzVmvgX6franaPuEfjw0N7e52gj3yfBqqPJmlNXR26Lv2m/f1UvZWpRIR+/pYxeQNDaVQyHFBW
aYJG2aUrGvXR89IacO5duKHJlMzN+RgKq85Wh0KifoXLc6x+n/IAAP4pwVZ+cUczY81vrDqwYlHA
aQIOXxFPlNFKGXIPatZL6rVtApAog3yhhHGCtWhT/xEiDkOaw4ncuXhj+A02yrbYGM2kGvjBu5E8
S7k7jUplGi9U7UKgip8/kHBRr5lH0vQewQnWD6hb6Qgdxq5BJdRb5WiyQZz4z2YJrHnP3ql0SR7y
uIyk8yi0xMnIGeWIxY0TumvrI/hYPneCaCctH1n7bH/bwpIW1mKFb1tnkWtaDi9i6Y7SIFqjeELc
miWxVaWneouFmqo6CRYgj5s+mLNZ+kde/HnTVKhdPTOXwgotsrfJ+Z8OL5jHhdBsmNIqHQp2ULSs
duimt6TQfKODGuM3Pt7i7omh1wVdtuhRXiCIOA1kSsuMm5y7n2wmDpRHvalzGynim6suY3l7Z5mV
+DFgwlCam62ki0e/NCgR6/pKus1TfPasp6rMRabuV+dk4PCMSB5EHwxz3SbL6KqYxmYDjy6gOxNb
I7g1ks6k0VN4UnWYa+/6n0yOUbuGxd5VwHGAdJ+/AuqLI2ZlG9TVhu3T07znKJYriVys3AKSjYKB
LMmsBDTndSwK3I4DmQwNIzEIO0JHzx8u9Tsbego7vL3OVMd56CGZv4XLytC9oaT+4LLFeHLd23Ih
gMwP6d4jqw5CZsamwZ1irj3KbJjO1AK+Cp198QmyyfrdDowlQzcd3nQENYKC74/UMJlJDIGIXr1/
5c4zl4Yjk4W5lGIMWHpuWA825hl81qL0eZUk+mKDRCkfjIkHAKEtyyGNq6z6W5SqzSuDThQiikE0
ezSNa8raonNncV16q+0wv1WGm866u5eX5+SxxShmdExEGPW2SrxaJN68xz1+UC6iNDVWKpUoeicM
0YFXEdcc4DJnSsYo9wBz1WkgmlqmePHDFlaC7IAS39I8OnIB/mKGJouGdVhzUW/5Eagc6eoLWGZF
XkumqsTFs1uFOx8TszmQ9qA2eOShGc/GDyz5ZmEItWIfzMdoj+AthwXZE9xyBU7HR1Fcuq26RxH/
8jx/uajde4rNtVjM2wZFNJ0sDMeK67d33yrZDa5glDWphUp/T53nueeQDWx0Woo5chAZC6OSTLk5
yyQmyBPmTO5W2wr4gJ4dJ8Uf+uri+5QXlwmI+yRqYEB+hRpytaY7jBduEKar1W6Jb9ToS/tpOOZr
l4dthQ86FT8nVxcG7PDJeqSHqsusnm9B3DRWxAcH6ZxkUWVSaoUo4fSHNR4Ijl4shuqi6FWkr8Q0
eWuIivLTR3W/mKA4/aPki7ivjJRAE63b25CQgza9gocQT98m/50fANNoNc7NWuI/ENv0gCshtl2E
67OspTHI6L5sPOB/KMbguQGPMgMTV/afEGyhLT4NorflRkKHuztRzGiggJJtGF/Tcy0bETb+6HuE
e2yH8GX0pAHVZ5SX3V+T47F4eJqnTvl/fOFn9IynBNMZ3vGJTmEOHYJmpBYZoMirGBgP9ZBH6sCY
iX/77Q4w1iBXXJ/hznj/hvHX17qIH6OVuEvDLD2nXMuDtnFJAm8gUb57UDs6TQIyj2QZ/os6wQA+
du8LL0tLPo1U7mbALERJucmtTX65TOVUEElWx+C9vSNLkldxDFuQCw3A7gRusNf/BeG5eF4J2wy8
dt3VyjnEnNjvPiJL1jclzB9r7dGE8N0Y9nB8SVZK6knOS9ysP/dGQphG54XpV367Zizv6pM4okIE
pPvpPgH2QYjEmx4xQzokSXXILIHU2E9yQm4UNKbYUdpOzLxxnDlkcai4B490msSB9Xw6hsdJbH8/
0Js6p5T73IB3OEJCPd2As5lTCOuvqV5N7fyxmMB73qg0VuTkA/FxFvk7bqbHB67B0C1YFqYF6dtE
kTvnk2RxFMa6kfl2rdEsoec5MlyGeOmR4L6mM5ueK0PyQn0sMFUbZb7kHMEGn6/HgNczQx5nxDOe
3Sxh2jHpiThxX6T/roUKJZxzchGPt3WhTM1U9L+Rx8ftd5te4yHAKaBW9uNYJ1UjV/bXt6dAx9WG
9nQirqWO3qhBZQb44i2ioDU29jeIFAS3ppDfpsKFsKwaxDGpIipb09Jm8AM6D7aznY3IoYUPmdOX
DgsEmAHJKoVAm+GwR7cmUv333GovX8194KTtI2IjqQUgMWa4F9QsCWVb1Mxnz72KyILk+ccRtiDm
37nmBt7iTeJe+Lq18+VnPmSDKN6sls4OUTSpnzM+b/BVIOIHsBvGGJ89y8Gi1zQeCE2KSikVG+bI
H8bmmWjiKHYiFU416/b2EI5lh14p0Z+fORjCYHfULyl2DvcpRWOBWNJwRYh/H3ULIcPCEJtkWzUW
gjfco/Iq0MdLzTLBJhVPxzjyTnzP1wq+rfIGGi2ViJavWdPW8CaK0i05C0cCd6h4H14WDif07uNW
3wpO5BuEejARWT+57ofNBce95GWkDMl4DVxltutw/2ebAmlOylAYUa8tqwVtzzIlvMkMwYa8F1yX
Tj55m8bW6vfo8ex6XPOzW6srwzl4Vj04prJjv1wfTeMmKGpXjAs0QXEWCfvCZIVyR18MHxMG3lZy
KhAWM1VAUaUx1enkEMuaIJWGWXzYoH7SrvuHYiFvCAGFewD6klwBiSodmJbJTiChoOK8mIAryc11
7ZCzWmWLxfa3M5w27Jb70a0AGfMaIYrQIZOaPJutJPdAyLFvEBurss3yIkhKqjzjiN6yV0INcYMy
aH43vxs2DcDKyttssBF3lqut8bCBXm5eFH1rwEewOow1mejKZ+6v7yZQEAyyFWOZJUNJPUq91EtZ
FAGCAktfhBb9FvI+lyj9kFd93mD/R9NbMlm+YAv+yKYvjInIe+QsPWEol/MnPKZN7RCPPP/uqjSU
ChulMCatCSdA1OVlntwFabgD8LFVtOhVQZUCz+6YZkIXRTVZ3edASguQUwHkdK/vXts1stZgQjDl
0lI5A5MRMI81H57+56UUhb0HF2iin2vzOwtdlQlMTTXwL48Z9xmjnplXH2SqsyYqvmfa5wpOFhgB
SA/m3qiZ3nXKwmnphoq29rqXwq9OhmtGQNPMzLyyzHnUv/qageQl/a5ahBPxMD5qL+u/lwCy4Ipv
RuUcRiCl7+aHjom45c6LRjrgCH56bFA+kiPY0wJEdKJVNh/IBORZSaP3FjHa7ih01OYPk9QjElKV
7FNbWi0lhdCRb+4HajwTbgM6j7RTRX24z12cBqTR+MqzBtPEJ9uXVAdAKeiFOuA9iHF0S/4zVcRq
AzXZKAsCNnGzzuI0jHWO5veJxaamYvcvEHF6cekyieY1nIg6vhXruME68JyTCPRIlSeKzKxblOCE
PKXPo3d1uyldDAAzEP44z7hJqCvo4rtOchnU5S7Se5V0aLBJ3E4P2h61B/ViH6SL6O3A9mLXBE4h
ElaIEzGdol4A+yhBDbwN+HoyMiuljo8tcUq4nTyYCSQHRlg7F97c3VWjqroN7LFzB9EvjHFBtiTK
y4dSk5RUgLRQ87mSu9SxffuqSPGFR1w3H2ES+eeC1YmiJ7lkJIP3jNEXdjBu6N3i9ZsEwUxMEqpi
xf73LQIqfimRi7ee0ZMF7Dob/9XR0r1Pv5a/Yur7oXQMON2ZVxjz3DyycisaD4uvnMIfTQyf8SeX
bNSvSmZPe5KQT27YlIDRK65NPqXcRJpqyWhoXPtonxLvzIgULh7lIu7Bn/VsxNdUEhQQAte9233n
KAP+Q6mKmh8fBGmV9zcwqOZ7pCorDbQ8QhRY3WutRKAVgsL4S73y+R2d47wrjENCpVR9Xe4VCYPb
Qx/LHXPW4Y11yg4babg+CkC3yRLwyGPwDpJ2stYgu+HyPgr0nlDl2obt85bKBILOHeK3Q1Cq+VGw
m+pl8yigOjvCs4MHXrsmNa2CuA6OUd8mYuxrNjZwYD1cGShxKO8nMbcOiVV429fzc2YA/Oc8KGxt
QFP61iJrMdNMDcCRPPGjCIrKfw3ET04kP1BbrV+q/sve98/F8OFCI8WXluvSZn3knrpPhDiDYfVt
KNnW7y7KtNENjrsL+Sa6ol9Ot59rVJxPXdaoHAg6TgdGTub+8tzi9osinVRLDZMwNad4jxx0bYKx
detzySTZjKgkzD0lI1TqPJM6HmOq1rQ+J01Y3YQTQukFPdCyX1PkPllGSf+29ACUXk5Mq6BX/wJk
0K4fMIUlUj7cC3bD1k3Rn5xHBiji1HKVu2vq8tNhpuD+fvIKWEBnl9p0yTb7DS4i6zvLcHoFqgLf
MZD/eN0z8YNsUeAwEFvTGcFc1lS5l7jKrWV0asX2zRyKDLx8u+QAzfaoVcIeYRlQVuOtQe6vWks0
/57ULZtI7bJ+89INfoWsRfh76/egg7qDeYcxcOzIsK0CVdXRbs/AJPaEkFk92SH0rYcKMz9LQGM5
tcKHyO9mTMME3TF5wIMP9tF8OeHq8K2bCHgcHQ4s2sfIM3weXxdPUhBs3Cv1V0lteEuXb4IVKvyp
ivO+ce8FIGafn/rzYrUBcQ2cdDtomNvbpLvc5pjd6wEZVT6clYW4VXOwKRYsEhBRsJNUsbGTh6iz
iAmcFYEibSBQXoqI1oziZRi+MjFVvAxop73t537S0bMKIIbfCiCRN4mexcHfp1Oj/Xz1oghu1fzz
XJbHbZ5M3jXJQ26UHMfXI3ND5pddwcrH2B+y1KcT4quKqs77CO+v5volTQTCHJyDEJgxomtZWfaJ
QlmNd8v/btrgYI6FP0XqH2f3XnvQ6vDQLnDbe++E5zH9NqedrljoOjUlASBlKEihdkP6NzLU6cnn
/u8J/xYapImWkRzQKkNTsqgrBF/m6JLVuaea8CjNTGAWlIBNPMwnRFY5LuREDu3erylWmjHMJomJ
kkmGu34W2pM+GU07WUqR4sqaNFen37LUzR5esgPb0xBT2h8lJuQldQ2HhrDFd+TA6d4kqd2Eb5F3
VGvW0ZovwpXlRy0lhX6m/d1A9FQBqebAGTJBDNqguEQKaH/FOIHy0hkLtfL+CXxkCO9lCi0igrCQ
7RQTjJ7YhawiBxVTiLo9E9LL4SCOk+76IVwCue7aksExv3JTUsfQ0/Wo8kKHnf4mTNlIJ/pJ3JnR
ApxwuAgaqIHz/D2qLUzBLYNSl/ULL3gybDPzhp/JMbGxdRAbA0r7xZ0HPhU1r3J8F+T/yb/JSXLz
6Ak//9pkvLy4S/jr6dpvI46YxGgT2pS9dip7Pf5lmvKNn0uPRjOAUUCELmHRFzVuNL/P+cOZMqfP
p04YMvG+wPZGRnuEPaSUFORpxL/2+Pts9vOy0/NPozq+gM3jQlkkvkxB23rU8zBWlIizxA5WlRh9
aqIBkX6DDnZQBv2YQNne7kyPuBURQmKIUK1lKWaIRoe+Xu8fXfwGbMgZa2Lii4TP6ffIl3PmY2nU
O9RP+NPwhDGGLuc8rRaIJszbPnfrftmzoREtz8GCYT2IJFL6KDrlu6V4Za04kEcm0/i3rKTZKtOw
WRYYs8MxQasoz28X6q/FONJSkZngMyVuBDjSXO5mFpWspqfa+/LD34J3BPzWsIac4gTBbPICsSeo
KIzyU7/qoa3UMDhzyPJMdxiaoxeFKlzKWnMDBaalYSmc/mXUqbGC+L8RDw59frh7f9xc2Q/Wfee+
NcZrPSmEfw8EogWrW6tTpjLgZPnJh+8ZLUSAZWcwxtGh3KhersH0YAM8YrBxafzQMp6OSdUR1Rra
Gw9l9nEYWkBYDuqujAxhlmR6XV5X9x8F23vn1UvWKjnCtpettkiOcCi4nnGpZoCI3Vg58r5J+jKf
es7KeBEXEdcNrTp8v8SyAKRBQ9sUfBntJxRO0iFX3V99deN2ntleTRRQfDgutlVI1lDCg1/MOxSO
yA5uY6cf8PC7s5wVMZ47W5SoaE8nJ0BPWis985vycHiQoTsDzz3h6hu6GclHParVxYUOPfNkzGw3
aav3o0EJjvBes/AoQGW/iGp6bfh0xK9Hf4fth12VVH2kzh1Oe1EEckv7SKLAzumpfXvsUduU1fFS
Y0irGGCQXQlKpuKGgIN7iwppxyUX1NY9vlJcpPzbQTdU8ESjpA3fVZPfAXYzMe7JHKXDqaKQpcNm
d9H6hXH0iz5LX0QBshNd4qyGE4E9uD6wL4X6VntQdKygSK7ymYGaandkpSsStS52a7yLdii4/gnQ
Uz5F7pIc1pdRUzoKb5EISw7roNluuUxYOkvB+SKCvTA9Shlfki8MuQr2pB2tMQ41vboAG2qTA1GZ
iv3rII/XhyrIwWXIEz5POxLhQw21pzXvqpJK+Ce2HdDqH50pVG+toEQsr5K71B018IaxCuvINyiP
rgkznD/v56nIqw0g3nZypNZeKnL5Ec2Gsh1WPAS7wEN6BV73Dx3poqucev651Kx4179S0BqkLAWH
wU5mMeGYX75ZLoJVv8guzCdz+cSODUbST4N4/DZ3Tw9TSBRMMWdYN5M9fM2dx2iBQVTRVr+X1hiG
bo7+QMptv0GTis2A0qgUNOWZS27M1fD+MIbnOrnr8CFTm3QeibC1D/0yNjmIyUoRwZIBLYxhAehC
FqpHo3ZQw9ITpdUkAV98coxCRAFK3zNT5VtbPL+h2R+OhJFy4ugBtBvfmOrYsOh+BZsph2QlfvUT
eMAam9esiFFzATKT0SlcmEpbtNImxitQJ2HR3waBBgHTS+tfCsAvE9iRgsWatfYmvpqTlEMGrt76
eXqCK/zzgx3SBY755U0IejaPkiCwtLG9sIKqKuCibzsBiH9J1tn3aHv0rt9lmeAApaB9F6qf+TSx
5Lxc9aC5+y/l7YdjusrNsflEtWKIdlFvQl5x98UeQanmvRXj+LfJPeqZVwKvTssMZQN5yyAw96aq
4O6f8/WJ/yBNX8/u0+R2y5Xa35g9GrLcimwEQNfayMLuus7Bty7CRa/0xptqV9AGgtbyCO6v0YAD
UeUVyeGWGBPe1AH5osM4G93DCLPg2gm1/VMmwFmqUbprsiKvhF3c/Zhq1LCzcLyAaVXsB8lQIEqp
3n9e790w58XBmj87gnmR4oFQ+Um2LqcuLxUnNgvHq1k12O/Bt7Fer89dgA8vvMe1QE2C2G93rmKB
ucyGBWzs9Ty7sd0QZO+ntplnP1CBjHlCxVT/bFsv8HxmQYl+BQD7POerK2Ezdl3HcEkMdYJOte54
8G6blBvY3aeezjEu4RXbDb6PrJLyjhKDkwTn8byppRMACJ2Q5dyD94KCVUckjsK8QgBtwLzs9b9q
l+Ydg5BLpkyGewPMIAq+0+u71UbP3h+LNxJ93H3ScVtzrsbDXWEwK6hFcLiwBq0v2HzpCgGJAm1V
n5C6HNS4+rjDQWaZxaXD/lPZpUmuOgVF08/BwALMa+1WOzgGZiPym2uaY9/ccGQbsKWI+1KFUa7+
LwOtdmbeATYUT32xgrfDgz3EYEa7+hRjCS8YaQqe1BKJymqVeN+pr6wgAWbdVwUti3uil7mTlbv7
c7S9YDtqpMrQOYM75IMTeQIbt57jFfMjlSffKx/ow6n03wGOasJMcu8ewEanCdj5k3bUtrnwf6v8
LEJb4Vn3OVOtA1UH6d3nFz59zaxqAs4pNHXXT7CUNsqY2VVuUiIVfxw5wyiL9IgfWV41US+iM0sR
gM/Xoef1UdpyRWELTExQQxCrn24UvVI580yjQfB0psVhLPKTJYcA26bbjtcr0rBEBiB1vxS65SpJ
GrXHZSQPlT4To/S96e2e/jfP0AG69nMTa4oxwCtvt9CJi0L19KkfFNBVQZSvrLYXD52JgbkqSX50
f2ECBkeJ3+jczGXTVwqP2rO9fLqBI1OA039B5spj57I0hMTZUCsAs6IcER63F+4pYy7vrP280PKj
8AwREeh24663xA7zu1wqrooxyk9zAvOj+U9CyxPr6R2aWbIEIRoJ4FXhyeUCz4Ly7+LTrg6CzdY8
byPhXE0NhQqhpd6dxxq4bitEIOiYslzOzRAdZ4RgucmX3jE2dTSXgGQwfpBRndr7tYOXRixX9iZq
+5JrZ7mbmtiLkDrjpwxD5hI2awe90H4EsBKKVD648HUmXh7CgweAe8PdhvdFM3Fehfg4LvbWQ3JR
WZuzbqGEHTgcfiqwCzqWlaifOUeyQbDZ37z/AGaT6rZg54/VfIkJnhatFOsnwmHaqYOFHxWKFIbv
MS+MGJtL5CAGSqDI8gvOv2LY2adRk0luuS7Uaozvd4bO8ZEegUFw2D8UiWAdfmAC4P9oKJncP3uW
muekcphYnJyMf2xGQ20F/Q8w/IJfw1Biv5gSweSz26mcsuFxp0QFykfC0W3wDiZfSpBeuwoZJDW5
rR1KdgieKNdKKK01u0Z3Drg1I+cSxqjujWra5g+SV5xT2voECvAidqNCKUgPjsPtPn83lFXmuD39
5/KvFnEEKbH7oMgUi9suPkCvC3I8qzKopUnVCu/8VnyYwejU3BWK9BwSfU1nDrJKPWYF0Z7q/YU6
0BKxUVo+UEJOY67FNvdbFMKKDShl/JjEyn5Zq5ZRcyaHeUioVcPnbgkpGrsYzKeq4DFQdyqsoMoM
0W0jQendIm14Ns/OGwWoUPJavHCyo49CW7Rd7CJHKrDq98H7Ts7D5PoDDWlsH0RsGUAd5xLc9T9x
eBVj/+tJcAU7bfvQXpP6TN9SI2vuR6xD2Vlgp5WzAZBH5K2I3BAXflpU4lB0fjEKACh9hmcyIA8I
H7yszFom57oZ9bQ8UKtWLrg8Ukqd2wmX2abxZ819SrzmOH/W4qxPNZveGi1DI0BChSeU34kx0ZGs
rr/rMovgbcfYnIep3zZDMf+sdkeqsGzlnTEWq+4RwQpwK9hroXYvRkffOxMPr+ptzLolhPxCvqSn
paE8Jv7K8uocBoNwehJA3zlHJlN1DrETmum4it1e0vSZdscSxMn0axhhtDlGpP2XXtgjbZsz4OlI
GnaFILP6W45vTFyR4GuVuWLDm3zieka8y324mE/NOQ0HAnPddfmKHSeGKXuNQw0EMmP2KCA5g+1Z
ozW3DZB6Diqc6okYsgZD0AQ3spoITlzwjHBHuWCtE8lxt/O8TpP+l0jNKqH7y3uMQHdF8dFkvshX
E8YERgHo2oEF/CWr7Cx4vPVB6UY8tHCMSeXlro0oAXTjocmjEM/X9emb61raMzBDAxTGz9/3Fswl
UE7hlQnWKEsPS/EJzM/ZOmZac34nQVn7fA5E7v3G5qxzmlmkgnKw9Jiwmkv3M4jQSk2o15qcsE7P
PgHAWkDXlvqffJNBO7b1PHaZsjE9fe/cdOMkFpAF+HskK9cL6gcKPDc1Eiwy0qh9wJFGLvcmgJB3
rxbwxpOEHbVRmqtZEoBbBuBIBqEN9EU2shzF/cU9k2WUoOLMObWJf2NKTrUgbhIEv9iWcGp4++OQ
BhGnCNf9RVwbuMigEbY4f4+lkkWU4vd99N2lMmxSNrRBc57aPXofiNSx6hgllSxxfMcsETZajjRo
BLp3cw/0BysV/7ZIIYORwN5EUZet7+l9shHr4QzDaHRRLh6Cx8itz50bUGDXxGU+RB343jhLSI8s
5ZhBrGohrIKgXTsuiDH1IfHh4tiYNlfWG7Dc3MyxTXtPjAcKdlxMZs8yVAn6ncHITsVxE9NiMgsd
ljBUcq7tqkbj2pfOipP/iIdQRPxgGWVX5gOWDpey8gTFTuSqm/3bCtg0g5Ol6KLWsUp7gptUz/WZ
xFEfR+OfpzwiBmaMoxbGvF5Am3/Z9dtWFJE9yDDoUsV6e+UatuQU+Vs+P91+TDaUEhhzcd+agNHO
4ksUCXRvvyxwxMdy7RdPZoweQ4pN/RtThQ44gxBvlPbAhIwp6mPVfLGxhP0EbO5o2g9NgR2t6bim
mKmH8KWze33roqhqKr1bo5eixf0UXUNUSIXIy8509w6BQ/BwHPzPyaflGr9h4ByGyv3WeSR6/xo7
fplOpghr3cfBmL/zSq45CPlOIqJFkZkjrUU43mbWtKTIfvwVwxKrQ91LFIoLbwUZuhjFfdZG0y2g
JgrGnGjh4b80GjGqSOvuShUXJtTxRWrWowgRF7dJLLEZk27P6E1JWON352gncPxwYHRXshsI2XQt
JbPz1RT3I91zETLFazuG9AKCaHi7cwzFVsAZOpZ/E8h/mHesx8+qHndsTANk1BBTM0SYSz2YjPgv
06rqp3vHtOkCVlT1psT30AesU1LNVZqWloBa3rvJ0Y3aefMOw1Lv0ri2VM99gAfq8jpnWMWH3YMI
WtPIV3z8vFuaR3noL+o8KlsyCnFyQk+PEAP+l0uCyHQcKjXl8NMBkLW3fiF6tmOYALjd8lyr8SKB
qhMsmSlC7fr3FrLbR9ayuavo34R9VzR/COuLLvTxsNxRlz1mYIv8yQOKJGknwVsvrK5fCoUiA0xV
Ny+Zhv12BeiaRM26D9ddvEztqIFsQAr0y+U3mei0IRgHAY3nD9Gph3sK5QZnbP3RagLaExOiHBy6
jv8iLr+ppSXMSEsaZh3Wh5Ziu/lGv2AauZRce0DZ8bJDr06RbwjPkoELzAKuokNMZFX2W1HO5AX4
Mjdi3zS9qKAoBT/1YBRMG5NzHD6EAbjEfSEiQJhdK+pnLVhnAAOj6xS+dEVWzUvlsYfewqxlGY9L
IZblcCXR3pUz7Tu/hCbCq/Z3y/PHyxm0BJo5tyuilvZeMa7aElF5+xrT56MWoQowMuq38PfR/xy9
TNRZQ9U4B/UmrozhA0H3WugORFk9doOa8fZFH5vTNS8rBOA0+M0XTK6Zb14/qvUdj7gE609ZXq2P
/CiR7DVj5t8PqF2dob/LzqWReYZn57qEWfOO/IywGFeLvl9ofkv9kpWO9zXSw+M0hLwk/nzpj739
1wDr/O7JKNUAhfm32UqKJCHw+XYLjUBrZ4SEzny02nxRt3wFz/zZuH2RTy+ptvjiMTrIbp8kvnuH
pCDyzS7Mctdp00wkL6HDFtQgAJya2eQ2OPK8dzmQFYoHWBFy4dR7ldWDj6t8JpMkDQKzF2xuFKPl
n+kx22PCCQPGu1H63eDTbjv5wiUzLYOgWpYnJ0D9Q0WmS+qo+kxASN931B2Q2FFptaLMexkjznYS
/5aM0F7fmF1H/7Pv1WKB6L6W3ZJ0GlhGhaOF0DG0/MkX//b7b++ny/QG45kW62XwrOoTPyOJtFB6
sq5sPUsKdYBhU1JpJINes2Oq60IRFdRsZUnCk6lnYNAe80MPUdB/q8v7rIK75jwE3g5HV0xetjO0
76nJn7PmjsOBbEpwpAwLQa+MfUouwTajQj8LWkR0aqJ0hi6HUoIqIwJQr9/NqCgRDMr7gIslcy8h
Mzu/1QaWYwSzMH3OGQ404Eeg9aY1IIZDnd0HUHvUKFhyvgkM0JZ0srBVqJJc6Tis52LA8ty3nqtW
SDPyQpAI8j1LEK9gNM04HKovLwkXk2zqlqCjaP2RdemFZ7q/r1o3oYaIcF9gvkpuq1XDbydXiZGe
VUwL+pVY8nXqYrh0PSmX2+jc8b6BWYA/B72orQ/0GvHIXwZnm35K+WxVo/8FFpuT5c3QfOR97E8H
oGFUIXy6NCLCp0h/cx0+uV1RBgCHHbasiPR8tHRIeyvIFlFH/d3kYS/g5ejBelf6eVbs+DEIpPoA
ngHERTIBSYzktQgoN2wr6DyQHAb9Qum+FWquD8MAWinWtYCelDFZu/G9NwBkXRJakyvrYISH6QYx
dTB7c+vJBU0/EtlA7G3H7ZnnUUhCr1eZ72wBuLiXxzdLc8vJHv9jebc31ZguaOXwH7cJQNcwq7fW
9QT/r17CfLFCISUVdFQZONfKhz/bR6x9043kZWjFGo/JW8HIWlRSEoAy/l3amKa8YVWt3j4o7+Bx
4YweykHIatTcT63kwLq0l7KZ1WW9FOXqysJbJALqDmoq5I8022TELb8OTnJ8VDPlVFkF/468YbCX
KanZ94soFr5PYz/v116JrNfs+ei9DoldfAQDISuEZirKTpPLXh7Hm/2+tHJ2Hv/eK11d+pG+adAH
qZGo9JSlMyKU1/DaoVvHclfioJshUo8n0GJItqBuyh6fKc1mGcJrOLg6X8jARLIiPqkW697cLujz
JlFNQrSGTO7Ow/h8HEW70xgFmu5pavAA9bp7KdCyqO/rUmWNmLlFhMYfzzpg5kPd5Nj9rciSZM6U
G1DqhO2D1Y8v8k+tTKMi+sAgNtOaPClH5U/cnHxpESMtuRntpgUg1v7NbsCBaXMS+znBZiwDWo6k
MYC600UN7/ipGx/6WsEaDkoFDtLtyYk5P6YHPCHgBWWwN6KfWdS0MH3mwRoV5YWmcpdwQ1fnDDvo
v9GuijA0XpwxnPST0mmhe0GD6xPAK2z7fyVPphgkKc7ERvnWtJPA9TUD5sJHM8vVxBoFHNEk/Uft
trWAfMugIc6kn4dVZyhcTBGBuAfEWA70C0Zyn3s9P4OMnoQ0lGZKGzylfujhlI11Az1Y2ieVqgIL
jJ8lzTA+WjDYXK2LSehHwf1NRW3KgNE2aFb5J1v8AwnPinHRZvfk2JhUfxYXxRrIrO9vagssbwOw
nHCttQtSWa7BtcjbyMrc3McNliqRrZEjn6nfvYP7cvUKQam3FZG9bQxBWliTt6DFHAk+SXIyDGbb
WYs/WkXft8czgrph4fNgZU5gadOCq5OPlOoY0/LdhxbWRAY2O54qFXdrtG5UUSb2dGNuMpnTL6r1
6QtSUuti8oT+36oHCyp60JcRHHgOmw7DNTRlUWQx47l5KVEUGBzlMRuzMkM0/5nODkd9paclEMbD
W/vEFs+XM6juxfYO91gnIXSAruuJrAH3FNta6jG951g7pryhhDF6gpTT2UwAa1pm5xa29sbTTp03
I/cWiqfT0mJEF4nG07W55YJsfoibl3uGnQIOjqLU6q/XkXGfrEfeUzWvWlaQTaNAEE/ACjO5qqMN
5wdgS+0t0BeDyNDgCB2FMeWQu2lmfVJrvAFwNxJEn7CczuBlCvWS0npFWRTIb/nszCrh/PkRF8Q6
LvS4xuT/kMwRVm5O53BvlyYBd+1vgm2BKoH60/4c6CQF2j3T9CVQM61IuOYG7u3Qdx6cp8d5YnSW
wccO3w98+q6aMEDYIW4SuHp0iBqfO7kohdTtucdHrAYLrpSAzx9zjZ/4fo158X1NcvRjDB0AoYK8
dx3SboBG+krYwk2RWtbqeLq7fVSULaEjknZE3Jxs4pGPU6eQB0WaCF2GdYUco4SgvLVlDNV0dgDB
cKpTSbKlt5VrY1zZ8u3lbHCo88UkU5uOaJOzeS8iBrKQxKjuw4GaQwJ0c8sCn8ZkDHcexlKIfF86
zVNASLklm9EXHqEsg27eBzlURPfhuzajVd4zVuL9lu62JHkzdIVC+LeI2kanCLuVnDi5eVXQHvdh
WgJPzs1cTafEiAfYghNO+Og21XLQRR0dLJ42N7JW/gL0MtINMaZbOTZEf9aw9Ja/tZDzydnN/iAm
KLWYi4bC1wi5OeENvrBEJ7B2e95zt5ucgPNbu/q5MyyDbtvqWfl2f/RRQDZ2hRbQ8QPcVjKGKSbr
u/tj9a0dx/OcU3zjur6hTdyObBf2vxZd9QuJUSdrPTriNmSBNUGsAgQ6NIx2VTHrFYpic1sZ8CTA
0Hm4SU0FjeNRu0qah/Dtl5g4Mh3ZLuuM8WmJde8/oVTZWiN6XDRv5MT1IuRCGwpJAGmi8VGo+/fM
JBc9kLPtQE7beFMqIVv4GlCJ0tSc/OtvZhB9n0VYdXcWNLsREkLghejvmaNRvUM0viny6/coW+SG
QwkcgLt2xmakMSeu8xIyVNN3RkxBh63MXjCzD29Aucb6L3k8bv0bBGRtNQgCrnfffWK7ydiCNzHd
sSZLnySPgPZgd+VeKRr4bZrSkyNPOyaDr0UPAOfa+UtK3AsD2i77uoMWXwQXVxJaOJatWEnI2TxA
8xNG1X4f2z5T+mRZArFAiJVhMr+16Y9ZpArNWbsmY8yEN9/36nx9gR0ANWmayVpaC2QsN3rxlMD/
F7zfI178e+wl/i8WyDBfitN7D2SwIBFYkBOQqKtM29CgZVslvVdfKt3IAkAKEOLoVgdTnw+tBi4N
zgCXB9A6+MwFl2MJCqVOnYUGuPjGsYkD3fRCUpkOJ2LlSFRj41eKL3JwrLXlAxx+j4AdKDWUNnVL
wj0ArVBlsdoDg41MSwZb3DCoiwW6lPaNpZFb0u5THvzJjEZBTM2H2Ew4H8tboySwggqmcxnlgC/U
V9+bljWLSwOjxOtBMGwWRxP3YHRrA1P0EmK9C3sdEezG6wfrNbveCyhdQz5B153ANoZ560GUJc3Z
643Fqyx5iv8Q6tqzU2FmI5845NuX2BQn5MMeGT214W6XMup7ZC+9PYcQdd6XVRraJZVk3cgLdYT7
eUiAvgD0QHKWFo58jUd9ly/9hJ4gJ2K6+K3yuxfF07JI6Iys/Go8AJBbp8WYG1rZ33tw+zkv0dlG
53RPcQvNioxEsyKpPb7Ddp0o8a0dQs50rAijR86ez8F3mZrz6ls8yUIIJgfhupU9hC9nX9Fi/hUO
/LcFqGJvdLUDdkw5oVFiMAZ4uEwPLIFSeMMnZ4yUKWYh0xiOToTo7y0R95hvHs3VunxT5ZbssV2B
uVti4DEPIQLGF75ha4fhWK67oa2nswI6mT/J0YbQ0FvUTHY7BfGS4JtRvozL1wwjMNnZaVNP5kRF
aNRgDwGqn6HMzjLU0cOjJAq7ZMe/oEJ74uHShI2g3JmK25QLl7nHz6Ea4965g6PP/o7RLrZDnm/U
A4looFrSbrVUaek6KrJLxLgH+Adgx4O/R31dTvgLroonpmSmC7tfb1BSCxCXqZJuJsPVIJ6w46Mv
C3gxR8dE9mEQw0MzvXQS+PfclmaECc06T6aL/Fx+OSNGlWlwwAQ7giOh9D4NGZylSUf90wdYekm8
OLqnpRe9WI0Zxgf/hg2OJSkU5IUXr8Yn+dK6nX6FCOipuz3S4R1yoqX4vU42hVR5xWuyK40mvz3X
Xc2h9nBZBgWhRW3QFL7K+teXE9Zk5r9ryCRyDECtFnCW4ZmbI1ut+exGHyQb3BEuul6MdKrbsWgz
ZxD98Gj9Qxk1d8hsavdfH8oioLMRlqcCSQv0KstWKSgGjvY9U6cr67abNeMZlGihFqtCUr6+5+XJ
jui5SnCSdRgOl8UXg3xi4cQogpZnurAR5UmPNOHXahU9BqnZCNVjr1x7rGezzoAkKdg2q8obDDd+
scbSZn769HvBc0iK4jh1uTbpH4009hrhxwidMZwlZ+JNxoieXRN/4zfBkHltfMjsC0TQjbwSzQ7e
KYiPsmBPfxw2rNViQEFtVVftPGAOZfEV9RGfG9dARDtcmaklGZ8W9aCigTqJlBMfBsx0mQU4FT5N
LJ6pH7a6tLmFaolUOyuAHsBlHQqHmzk5smNd5qBDHqqC0XNX+Dpb84tAnCK3qnTPQUayFAtrtmVm
4uaRWPJlR8LJXahD7mVVyaEjgGYfXah5Kz2gwSxujx8awQnZ0DvL+f3Hs0AFdCi/NlsOZ+35AksG
UHRSty3azr9CY6fm0POtDHmeIwnNfKyR4m0RhkdROrUxoJu0hUfowcAw/XqXQJsfagBu3UCe9ahU
l4FTu61YnZxISyL4i5fdZwagnCqQFId4moCMiyke2EliQJKI/y/8JGHIF7soTg7xwZ1dmtmPPol9
C342QUmrTgwgspJ5cIU6YgUWAfABzVpkrJsGc+dGKxXX9Uk6lQK0JTwb3F0UVEQmlvHlooRTmG1l
tbf0asknUj454AtZweb9XJz7GCWJegZ/+e0jbQSaNgScmXyuQcyfzeSLZ1dN/kEjYC2u2BFgE2gE
R9OC6OGc5gLif4uRAbwLhkborcSGZQnQyxHM/Kf/26KAPDW3OL50VvwrjsUCL5wkKDzj8Ko5670I
qCG98ZCTb+JZBDixDR7pzkiVlzidT0iZ23EI84wIyOeOtP/u91DmwmaVoAFR6HVKbxNkwTWOHY7C
vfxGOsXRpixgxcS+PoR8d1shPowcry8KZRLpBB7zuNzMt+dHPg9AA3xA+rMOItP9KfPc0ygkWOTp
GP+SbjAu7Go+s2U7hHzwDxIyR9Qer31z6eDolbqSzMDRTMxRk+RcphZTTSRzuLY3jIYHaXmE8V01
Rx+qfv0AFtZd6Tb4tsIvVMXo60k6x1FNMSKwmBPKtg9TcnVbbkkyj0qMwZ3N3cIPQLxvqBYAErc5
Im83dt4QO2Ahzaci9fh+XdOxqbqqe95JmiTCEA1OReP7vbxbxafUzPBAikh3UcyQ0kG3myekU7JG
0Lkzw5jvi16d1+3yJdjZvLIbaVI+9Tcf6Nb9o5Vc1FG2x/ihcCOpCQEt9K2svgQATGCTu/wUqLht
EXI/rTW/0SC31qeNkz8qEcLYrDa1JrEMUJn9/5xLF9FdViH6zvNlEiOVfo6avT7dHUZYp54/Xwd/
9AslX2m1g+LmeVRDxZKgmlWn1jNg/3gDxwsUJnd/Lm2qEsruoAn5YVT4yaYFyMBJw6GQttXYTOWK
FAHNqLjLpcnoRxn8pcq6zlJ7tte2eASDQ4f25AFJkLZm03rSpeD2ejRKHsn+s1+UuwgZ3PAiCf4O
TXGL4LjHIYz6uGfRLzjcP075kV/nfXgTQy/EomCPOaF+QGoKYs77yuXipTuhw3ru7Ra0BWMFcoH3
Ka22xKtXLMe7BSynhlM3QcmE9CMP2swgAqPmNAHdNSYHlfLlNyIzHfUF7VJQOmwkeo3SJmJf6Qjj
obHm2dZeDd8mLYyH9LsYy0bCpoSScFs7SG83iaraNxYmdMKmmf/4WRR1PpmUlI1cha7MDIgcR3H8
msdaDLWh0RbQI/p1umKXxGMcIh3L0yskQsWl39KWBZYrZTUAkvlz8X6/3Hdvi2SKnIEVvHTOCYLS
UjLsO6kpgeYCRAQMoFKA8jvgr70Y4WHb72UJbAh9klslIiPWDqrJKv5XbNlmG1xBqvDxNicM0LYo
PcdN+6WgbGSjo9ThMwf2ShzCNh3VhO7+341gOo7mwEttitlaxLXwf7a/z2gAZ3U9JiLLUErxuGNP
7Ay5/MbJ8uNxMKkp7Lf7AOQRiBUZLB9+Jyk27BSVLrEOVWdyC+qomg/NlwLkoA+kTMkr0psPPC1K
572niOwikxvzfW+l8MLOGpFfcfgx4loiDdFwYmK7C6neW0pUnqnHyvqHdFbweJws1pl5Vl8ojfGe
H0oROR5HX6WavzCViRfsU96T587QIjhJJi/15OXlKdY1iGeg8L7Md9bLljSVz5W+AS2MGrlCSeY+
7g9DILpZxfP94NplEtpsZ1+kTV3CAfDRP2+4mxFpoO6AQ7VtNpXjAGU9u0wDIcWzXVHvT7p67qlE
mjC7r0lJ3/3KLoNAeRH08dL/4gpHNy6wUmK2c8/KF68kx8Yvbeqzte+AYmeFGkvyvb7fbNA8CGzQ
Jqnmb4Eemb64MXPsbOqtWPAS+ZIcNZ+/95Ik9NN1v6cLx2ZYL14zlmaXPlWdNKIoYm9bK8n14uwg
kLUwoWwXtB/3MjyokdSfoPYQst8sZzgylE5Tl3/FMXwYoik0W0eIp4bAGGNBlGI+MCSGMHZ+d9ud
xIybW+B2Ta2Q6r3I+OQai2SGfFQCuZE8nKD33QBE/xjV/T7u0IaUKzjfz/MKQzK6jhSJfIKuE9YC
J3fvc4ap5bQE/qiR5ExmA1lQzxbWLCHuZVFSExAISf/6PVa9WKgL2YJrz3CIQ8f62/C5A+Ahqj9q
NtJJErTt0LKaynTzFdw9s1k5Lrx/0UL+UaPWJPM5DJqOnLVTzvEZkfeYRlI9S649CrrE4vGxdydR
pgYGYaHscipQw9N+VYggTewc5//rZ9tgeQiQwoQy+54bvxPcCTAVUTIwSzbwsPDXQYgJ/7ZmD35h
xDoYSgakm3ZXLCU1NODL3HC2xgF3cHD9a8qwFBBAnCanHojS6dT2mVLvxMAnqcDl6fc63WxPlVd4
dD37mIzrc1IhLAtRQyY4ZzSM0R70U1YO7mmM8nkUkcYiSdUB3Ty+VuZvhM2HyvTSXx5Klok0GcYR
RFgQrxTK/KSnh029ibQgQP8ztsY8O+8wHZOH0hDBxJpyB5gjTlSnIdw47Pa+5WtJZc9c/w14yit0
DLXgaVZHETcWMn8zEbFBfAA8vs5sjxPBSFEYnzqGOwmus9TOPCNInGV4ryPNzzME/J+KR0CQ6r2R
FV75Zk73r5j2XEC9ox04DVtU7O2TTq3TYddJMTs6iClGxWRUOfxKOxQGplAzsxhE2ncyuwp5CSPA
ayGI5u/pj4eKlhD4bDDMjwF+S5KnvpUpEhiZ8Os4YKJTegExM6VghcAUeTKBq/hLA2UfCJiU6EbT
4erTUAF6RF3kJMJxhFFtxIofIEy5NVgVg1kru9mHOj6wsg7QKWhDB6+YILTTLEu3Vw0JTTlYTRSU
+5wah4d2Ai4q72Uj4mMoVZa2ClRMcGTKNsHT226TNIFOksk5o2Uo3OXFjbmk7jFSXsYRzLE50oXK
L+P4glabq/m8wSRuB5omiGPiT5IUA0m8SGpOZ6eYIqxlyTcbfvzIoxpuyM6eUC3IrmxceTiYo/EF
5PrmhEB84kSh/rKixUAgsFMEfGpQSa0gHFo8CDQQfo1nVAQyEEG6wuxxQd62cXh5Iur+LuQ+F8g8
fr7FwqL5qnqKns2ocj+9cRl4flzCe4mrn+PiM6B6j17H8HsuW3Gu7CQOkxdDubJHTN9fmrvGrx00
x90RteIO0vV9jxLwQc9JS9xf0bYRcnlrGuNSB33Byd2bpPmXvMYT2M63kWsfSCnstXRuiCsHO2+p
2jjEz9A356wimwsxxNg7PRLC7/rdWJFXB4Rzf+QkM4k7gzdEpGunk4MFhyTPMEjjIoxDsTZQss8c
l5VroJtz0buEFeyzdx7FINa2W1mN7YdiRzcpFKJAZtABOueknI0aaZppcF2gOoOV/O4olYSFwFEU
i82EduktK842vXwanpzB3sy6Zl2/K+F1jncPpfHhhz+aSB7MF3qdyR8Wj7ATgK8ajB6VJ1mFIfkR
UxB1tWFzcrJviHErT5SL97XNMXVKtnNongPncgxhHrqh0QZKVaZB3+HWPCnrsQWpvLrN8cUgNl71
TX7y2Ae1KQhYJ5Bmqw4g9d/RiV2sI6iWRkQnAa+alHlKgbdMoMXMhfPlMQfxDgOlqyv0WDSZ4/DN
6SCSTFdi2Z5dGrVPcXVhb1IepUhX5oNLccX8EZcEx8MNsMNZWd8DmHc+aiVgXS6lg2kfncoV+I+y
lwjTJfVZVZP38kZJEXkJ/kxeSXxJw3kDjOyY0UL9Ozgx0KLjtKXe8v7Xx13eh9t4iNGWYNtqCUcB
Hn9TK4cApCxo2uWk7FFUq8S7o5FXZqOpXp6+An2SwwxgY07lSMCmToweYjXBmkrD6aTNQp6o1Qj6
tUZzCCg7yc15nlAfzH0sidQAclnukMwlmyjnfHM67nHMkHw2NChTh3tud6SgXfbMWSObhVCXzH5p
pNcViWvQAfLIGrTb7RJyskm/HLRGu9vIUkTJwmMsLuqUaFhpni8ENHJwSfDdcfDGb5sfkYcNqumA
XA8q0E0qtmmtvPf+M/THqYeOK1HNdTrUqHV+YuIUmEV9/YgcX9Njd3KH6mjdiNs2k3MGyaP5eTbQ
6M1NPgAvbH+PUo1tmIBxfNtxXQStbB/7GGpKS19VJk3MWg3vJsvyMwdbaEJdI1BwUnjauAQR6UsW
GVAcmmEQLZHkSvVOnBf28Spej5PqqrTgS6RNLauxOYcuFo0DXjLtcensaPug/cGOIAXZ5aqbaBIb
JXdNoyVgLJ07hUk9E+PkL8C5y0I7DTPFvkmd+YKaJpIIluCkbbuogMkyqNyxiXSPw8o6nJASzr5w
thftPhrTcJ+BdIwPVcgLccS4hluDl++RCeMJrctyp0JKCDzDyOV2OA9Vls3e9Nqkx8XsV0yshLYI
przb9eNuZpuAVGc6hQGkFzbyQVFTMRboXynlNW9G/PbcDzStaTr2GjMxE9NiA85LDp0HEZMuP7kM
X+90RzYldewEadgezEqmA55mcj/OPXNdX5Xh0W+PUBq3Tmcu3dG+oX77g+nU1DpPUltsKtL5puq6
S0rjN2hlWGbWAsJVpcmmpw9kBkITFUzB4C1Q1y3M80bElRG1pLherszUYuVyWy1vYAFNKpML4vg/
k5zjaEqNaTBc9dqZGKELgJb7Q3dKX/RRg7+g3T7FivP6XIp5iGOib9tnBjymr2qWoQx6cMpfLAvm
C+2ArF3ncfWcBYKtV1jKVW5vZaDvPzrho2vKrtyRQ5zLm2AlxhoVI5bCdWTAGODfO2gSafSPJP1g
cB/e8hbhaWaiITF+prrSDKdlHV5bl+vL4Lx7D6HcaPtWYFm4Nx0ukBH5RSFTKjIq9glWD7AIR6WV
6qXfOs/e1Uf0yoV23phFno4U45lX3aW7p/MYT1Ts2iMU2rlj5oga+FS9WR5hvC3LIljXKckEVo5Z
dNNaW3ZZuKHL6p5X7NnzfU/VC5H1KhTwIkDhqWUcTqW8CGsGltZTlM4j8Ws97+r+e6Bis0g8sEtd
FDUNveUFQRdiEkLdmzZ7oSX7CNONQP8B2SrivT+BdCMZxGbK6PSePS0BRsgk2djLYq6Tt1H0waca
hse9K9OX8V+PgaZ3xfGHLh0+Ewk9E5Q8DqV1guwelwMybGOgCCkNwwCfHZ31731ouDqrxrSwqp68
PDLCZBPEIiG/+04c5OB9+dnwXMp5IcQ3Qr8Dm40Uq92+D29WAnWRFvBNTut/4f212ZXVMtaCAWMf
MdRVmEOfzY0Kg64T8EkdXrPog6+4qDKKTmHuEQKeh9B8MdbxAQpr5uIoWC31q/vAjD0Fj8f0WtCW
Zu8qJXna7I+rJCEA0yY2GdYBdZ7ICQWiEhzrEntLjf2r8VSNVxOSQa6ZfaEb8k4GAmXFMGSkcSJ4
0w1g0zSxllQo/oTX8izvrDrz4d2oBL60oekziKJToeBYn2xXUMQG7mFsWXkoOxjeIVRTUvQLVgu3
gbauoTBExqZntBynsbbQ513/tQnkBNwQhThfo5VCDLFfdSArDuYjlQrmzijly5UWcmj3e7JllG3P
3nMcmSFX5klsZ0mPC2lR98Zu+LmC+ut079oqa6Ej8NaimCixSemAa61Oho0TmBIl/mpld/B36rcu
AKgPiE1ChelEg87qILkc2BeSl43qjpjVvztXR6k/cNPkUhS4ZzsNRvXuQG+epE24xtSPPL9LEnzn
FTAVEdZ5P85Ixau4pjY8ALDIHuXmc+Lh5eObXEWimSekbqcMSaR5MolQGvKxLLhrCur+X2wuQGVd
XUg5++QW+DPVmwDjchdOnO+P9wGKtUQDqlT7+r+dSfLZP0Z19DKV+ZrtmNf4srJSv7vrIP/Hgqcl
7RjypcM7BMRWBEmWww+zmMoDVF5uSgXHhiHfgUkpoE0iYdDYbVC+Vuy8UkO+3wKJ5f18OQSwZfZr
EMVxngc7lrcqcwiBubMtB4mflj/9YWxPkAUVtBm5czGtxerS3nPjM707AQzdsHLlHdEScfZfUxEI
T2su6q+IUE1Pm323QIdqn8Ag7HA+CDFtCp310XhcnZKrgadaeaZvJJHHHtqfIKcqA7VjYpTTQCw6
YoyaEc3neEbV8JMRiu5+9Q9LJexoYVuP3L8P323Bbqx1vqfevgG3AZE8sxF7WyE3Xhgqie0ptKQR
EH5qNfUnYj2E0so6e6/NcTGHBLe7QTZqVC29c6ID+Z9scs0bYfD8LvZ0Ut4XY1g0WFc7Zg1vrww0
6wZxIIwX1RM0+roQayQbXD8DdKcTZ2RJr68QSIf0TlR31q3aIgXVkPMIc96g5zi+wrvjC/6bPTSd
fZVmKqCyZcCzqcaWswM1WuF8PwVeM2SA7+uhpmdM9yBkX0UYKACi5q4iuUf4PtPRXYnXwatcaUdH
/opim+zGr1dSCnJ7/BclaU4FKAr2BGrvPJbmhKiF16SdtsGiiqrt2GOWVRXPBLYwGGGakCUBybit
k1de6h40/woDhgi5PO6BGTJUG9wvKyCi9HM++Nr/kChyRL9C2AFRZotKDSThr9Xd7UkWOgvFVkBx
NZigEtpfPlE+LxocBROYro5Bnz7Y11QOhCDds2g9eHBrXLiMiOURF91xGyKhu3sQ91yE+eL3MijZ
mNKhu0rizXDAerHR+0GiJdVJzZ5NTpgs6Gzb7cxoEhy/Qdi0b+O++DKX+XpyzafStq2J6gsMNKJr
V2BiqapjpHJTswDt3c/Fsnlg6ns4+cMPMDXcpG6A3yjoscld2szLmHYm//fWAhdi++m1PO/tQOkt
1bHNLoYLK56aUhprXyDH1hSb2VtEhbMKYRYaoDnKiIXOKQ73+0mtNnK7r2wqk18fpwt9u9CpK8C8
MP/7nQJQrXbTFXpjwqZyJi1l57yC8snurvZJ0XW6LpK5LOarV1nnvxjwllfOTXiF8LCJ3H0ER+db
k9tq+gEctb1tktqPe1jsLMGgvQtqxnXslFG4ZtISXbkdDzfaTeZGf14GbRnyP6riackxdLR8ZIGb
lKBPOPuMkY0e1eD/dQP28bLX1fLuwrKbElODKcHxTxPrAM+Kx4WmU0FroqHb1W2WAuRqgOveAB1d
NJCUFb8TLCzG2FAQEai4exTc5Sn+Lmmh0nQDCcVd/2ckHmYARigF3bku8PS1udmrnE1fddZibdJe
RPQuCGj1zc5h6/goqf+weamBQNrAjJ3lde7KFcOGIFheD5SyVBBEQDb0tZa0FjZShkqAb/GKMp0d
lmyn4B43xIoVY7BaapnyuPbi85o6UOKIGZYKwHO9AlVnJl6D1iDp5+cUVfXNrfsQRkRRSqWVT0Xj
NtORprsW9YIFWsxCBxvmIcAzM0d8iO7kSN9w+xM18aWu8M43DE0GJNJ+G3Rv+foZokpRe1HeVyGJ
AfLgs3nemrqF16Or6AXWv8rFg8GXz1/CEJXz0cmvZCaxpwawuzzNx4LfN1ytP4Z1Ei01IYqotmU4
H+A9q4upahGeXRM9NmFSqFKCagIVrO13sSLEjFEvdfzh2sDRjGvx8XgpH+VcXPNTKaNrXMgJ2CXM
0l7MbDb123U0vcrBfbKRb/GxAZL6xf/vsKiKKlu/wxRbZtsrWyVzqhbCmkTWG7auoKVKe/yxeDq8
VVTKW2BdQN1xNfh9d2i28dJUTrtLyUyrkybn60GabnsVzh6hQZrXFB/a2Bzc9duMu0PgQwxMBPP7
kw0pxngj16qxcFQRlxLcm6qRrii7PgPCg+EmDO0jo7ulAa2OhFZdANZ9UTpEG9NhODcS3h61q/yw
yoehs1KFlABXiLKXQNko4NEKQu9AQQZGbJ8kbQExSNP5ljsswcBQ/GEAUcme1OtgbMi4hv9GPzXl
TRrpMRi5t7F7e9pxReWk4AfTJsM6+uIIkpPub+Lf9FMcSTovK1xX7pd774tDhiX7C5t5qfAX2Kn/
YZaSVXiziVhHxYo1gw1uiEIjN942l3ug2KVQKR7ZuOcNZMJngdHE7uToo0uSeU0lUlG4qErMUlPA
6tpa5FjrCqAga+xTgCYApGxJ7yHIf0Y8/o6ozjfrANOGPRceYC7bty6ZPo8Kr4EBgsVMJGkFvbOu
0qXYNJNyJm/6v7d+nOKYd1DdDcx4Kp+1YHY8FzDpmIBmsN5whVwmX1DveUb2KlQ+omqHoVz2F9Fq
fksOC9KhqcdhlvRZnEl2udOtYMvCTh2Tjy7GPj92ymp1q/kQjR4HWMXoVsBtAu4qjCxRYLJ7TP8j
j04O5MHDm8YDk523ddqmOcli1moVg3e02wCtMR3IKI5Sbe2wlLGmLDJWKmYcMLrkVMVZHsGUmcNX
9Nfrjy7b7J9Qi0cVVaH+UPN5goc4kPOIKeazFaRolqRb1h+x0kSSuJ0g1m/RIL181QAMhdsXiXAZ
YZRRm1JHc4LQX3czV3kfgqgLR63moVK33R+ngEKNAL2xTAZOePbcf9j8VZL65qGRs5V21H6Ia7r3
XUVJwirsy00c+dtfBmIBOXEC9Jv/7TckS5CID/szGUfEAx380w+ayWAffYapegTLZTkp5EFROve0
+RxBZaJn6Az0995o8TeMGyWol1+qhjFJWv36+F9BJALOrJx3fb2mE0dzgo2HhVEHYPOX0RDsk7jj
PD4jK0r9H5UpHfj1YPUygFRiCNCPtxb7uhj97vJBTt68kvmFQm4fVwyETDbtOciEzE3EXpOou2Zo
b4GhzvUkp4D8l5YoiDH4IFO3p5eISq3z2vIwkMGCZZq177voRrDePUh6x964SZQEmiWcp+CrADFv
kUQQRPuZsZDPaoDwEElfUi/+nFMqXishoJXmEJlHTm8kPuQvkX9edFcdSZN6qR8ThKGkpbTtywHz
HJ+xzwOAmsjsqfXnlxu9f46BQaSsCgu3XI2dlMr0r1RMhWxn0xa6TMslsiMwRspwEbUQi0mTmgm/
YTTL39QDEGYLVsqtZUmX6AefmrriQQnUcw1pyJRSN3kkXaGqnubSXeBVnmJK1ipuB/fxRPNURc1s
SYHiliVCI0OLP9/Bmj24ByWTQDQSaamhpyVcMWREfPItGILkWh0lGzXRYr428ZH40L8wrOsYB4g7
VOy4mUchPJZLCMXtGwpGhF6Np9R6azL51LOdeRLfB6bMQED87qnyMNaBoOIRYf7Vu6Rex3J+lzq/
1QFQsN9+Z70wbuY/A8HU+QqHPtXckpj6Dl6fio6B+yF8OkS0yLPupxKXVEeubZ9LgFRlRIA4mE53
KkSwUxGMRt9nr2BvLxwAvg8vF7HIOaJw3gba0WLelrv4RX+Wqx/x1S2JST9l4RSRDPelBIeNKsoc
RBNJ2N4V5PXhjCBU9Hmlg+HYuQqO2PLLauNrbYBFuZ1bb86JnmSLDYPWusGiWClU3lnrMcxyJD1h
JtGD6uJeIwqqH92weQXkVsN5wwpJpkwrKpZv6yRw4TeRA7kEiJgfp+/QJIKhdy6/ZrmNzc9fR64X
e2aABukH4GnWKsmSmNUC8vWH964FHqpkkMTcf8MvJk2p+9JxtpLnz9rmf4v8CDDr8sKVhLDq90Wz
Q400WCXAJ8cV91fsW6QWMoHodZ6xDcOibmr89JxGrtTprKKO0yyGwwBaNOlSXiQy5bgGEedi+WTg
cPrN9BOC56bXibgXBU7TSZG31fsYVOubPIYZaabEm8XFfNmq8gji1Gf6R3/bngsGD7E0be7isZ4h
PS7NKd3/3XFZ4/72ICW5emf9PnkLGVD8uRSH1yGSWJ1uwUBeGpJCmmByegn8RSse7aQ/PNC7/nPx
E/58Vth721+es18rEW6PV/Y5z0MwNbVxH4b8+CTUfUwp6hypVTN6AANzEWYLGUZYy42g04GU6qe0
4DwTAwNzJd3FnaSP7uU8FpqWkZ1peAXR/Nfu8HsvSoWCrfK4M6PqPzjp7dyjWNdnofnwuhrEZxRJ
R5nfOLP7BKiAMlSKeW8duRwWC0UPPeXCP6qnPzPxVdDGLZPVz7lL7nq8o+N4PIn54BeY3Lx5CCag
0b7Xiw7nT6eVrDv2ZQ8/2bGP/1F5pqKa4nsF38D15KM0IwI/xVFm0i0QVJqq0WMwKM/2yNWB+SMX
C/wQrhnJE63EjogslWQuwLN8g3uFWvzm/AZWW8uOCaL0mu/aUO76ZYliazdCwC/l5IEBhYExN8+h
UyR77ZbSM9vP9Q0Joj5xvzQGfIO2uz5dI3lP82s28rdWkMFBgGAXDAQADT2flOKh7tndfhMNjfh+
oMI+W3Uc14T215u4tWNwvRQkYNvHkjLLxwY1rCx8Cul+SiuvfsNgNKUsLmcaKVLQCPVDYxl5krAT
1MmQub+sn/Bj094IV6o7HUOdd+OajdzCUO8AuDLsLAUa+uZe6J84Wz9INqbGqriO39Pc/qoQRNa+
RiwxlqIRM7Po1gjvXymUsG0xcYE/KpM/2AK6wOA+c70vIp5xOaXfTLMS7ecYnSTv5yUUd01AN1ZS
3FznJCApkdmsF58W/mu5qQnVQK+N6ApCSt0nzTPGhSnvDYxQOhWTpvhxkufcx2HTnT3pvJBdxOkN
2QrkTv5IfOtH9Nq0vVtyMEKDh/eEYO2BCzmjMD8SCNTkbDsPHihpIgvIc0gFtk8ygRDANp6WAIy6
uOQIqeM7NWwG4kjjQqhvJraV686DOD1+5BKnwkw2Jd1qp9IMlZHRq/g7JFaCENsvZ8QqUTUushV5
MRrVj73EDiSFGODKLpBti9Uf4De6bLkNjReLBf+BQDay5MJrLqwAx1W5Ij6gjYrABYvgMsTTUkdb
LVHnaEY3SF4DBvgqoAe9mYi/+QzJaMWFpTdw/i1GtcnCqvpNdEGHuK35y6hYXxInWB6mLBHPB9XF
IIDvAdsjdzQTnD6g4OpHUMU6Fl60a66N1FaKOnLYwcgo0fa3NlUe32OBh4fHbmurP5jTizt4w1bh
MVf8RpT6Hlte1GP21XLuC9L/Fz9GWxtg8zfEQRmMCzTZLzB2Pz1MvjZDZwdmv22R+npI+zG0OIbg
MPJZcWQI8Flh7n1iwTK16XeoMLuFKeQl2oEwYx0/V266Ga2uZFN3oh2MVk7wZoMSeTAe1n6940lQ
vxLbQBFWRi8yj/0rDWxBB0pGfuBaqA1BNK7qXfKSQjfepLZ6aX19fnX4Yd8ZfTW22/AKzBB3UU/k
NrqgdUPiRg9V1rdujp3OTLHbRbvE7tWMIIudjuEKuGze9Yh30nSIF7o/aelhjM9ix1/xV+vbwVVg
8SdTVhwFC4vjf7vYPcigM03OZXq4d6nuzvykAHhWCA9rApzQnRVDYztFQ6epy38MThgWVi/bsf/V
oOEkJDehsnYBoTUWwX35wZRDsfIzu5+cpt/MyeH7zmBLKTw06Kg7T2a+qV0p3JftsXY/Ajkgotp2
WqXWnNe55jqZx3Z3Y4Ip56NaUvitmE3G3ybaZmwUkO17pf6kiy88Ee8uXrDEy40M1cYMi/Q1Wln+
n+p8ROQCS4eUlyCsbdc8DfoUW0IFGKUaUoyUUS95UsziCNUk+ZX3M5a+sWO7dNmkICyPzuXQ4lea
IWXph67+pszglIj4Bukx0F8IwelTGxiDNsNsljcyyp9hcq2ySZhLOzCp8LdPzkCySUo/NHwwKH/8
YVf3Yo2PMfr1+919qRxP2Eice+vstz+qmrE1+S8LRALSleu092HQZQZ/p46lhjgXiwkWRECUnYsT
xw6U4XGqDFootWepWYMSaByQMMhtczXwJbbl9piyHUA5+3XvnI6vNF2PojpYUj4zG5eHouwhMf7z
zGI+P/Cs4LDeoODAvgRyYYpXl7XRXIwW4qYYcE6Xd0HZvk89D24Ll0iEm1hp30MJjpCbB+cA1rT1
yO7DHPKpOIeeSKMP2Am7GARg9KgUb98tVksCxJ/Aw+291/JgZvQTQfRoRVc9NJUKHWO8AKSFL6q9
yfmxgABvW7sSPmZ6flOg1fCpXbjSiG+6Fomspl8VGyXT7Ny8xtZwHSA/2T+flRFlK6J/JynPpQWv
O0ULoIKPjBtjgbNdUUvBYWXUGZjqZ2ZhfSYgtXKf3pX7P1TqYgcrW3kk5Vx/n/jzCmlB2JxIqRIq
yrj0V6S9OwXDrozqtYuU7ZeSjy3zv6v9+uqRfO5nKHI/tEeIBaXza8GeAOlqGAoAPrJTok5Lu5Wm
S1QBddue2w+iqbq7RDPw3+AQ4TXhE41utPHS4i5wheomzeAQN3/TAVMrRd9afAg5kp5hEftMHGKk
Di93jov6riu0xM5NgkdeHD74SLJmdpL+TX6KIxfZ/L8vpJa0+mjasay3saJ4bN+xH4O1eFfMnD5N
EE7+Js9bVitcvYvTGfsaWqZumGBQ3UY23VsmuCiuOzKe0qTcmRcW+7kmUy2TCDNvOaBQzaB9UJPl
UXbJzyfQRK8tmu3ya8+lJs54rJQC2Hr1TiUOQ5AOvs2uLG3GOw8Pn65puB3KkxYnDsuG5zTy5ewf
iD57HCsVHW/IvxYT3u7DmpYQKq81eRfP9Sav5hsUkT+wMeiWezb7wErrMMu9HPrLEC8Ur0FF13aM
MAByabPMioHKg/okAC7lRI3dwO8MTAWcg4Y/Cg1yXx8bjRIiOhIGwx9b2ABjyO4iLMz/c7Kb0eIb
/J3fpplRcbQmY1G7Qm7WWxRVVUNoKLyNgWRJLJBne3ohH7B4F78IPjMDN1oAWv8XbRuKRn7DD42t
hPhnj91GnNWX4yHTiTQiB/oJwqfqZX5FTaLHVflefPoWmZU8bX/d4C3GWECqrUSdkdoB+TMmZn/L
qtu+/E9AfyCnUOMcIM9ePdExub96blCYMFhWq4sgDUOlpic6ECFXVZzq6nlOO0FTkUGrxMxFz/4/
4RYKaid46odTygXYusyQCDzWSOUxEOFMnt+r8UH3N+pVYrIyNGxtTijbB0Fjr0kgc5uu6JzFMURz
ZL1zoiMijZUIGVC9PJ1dWXLQndaEqZGHCNiDTCnRQGuOp6l9fBC6fHfUhTF5KxnuXHAT6CR8TPDF
sW1NYbMKQ+1ddUHQMHNAF3sNlo7Pem6KFXr5dFgdXchmauu1Bwx+/dMwFen5yOPtff18LENx6XN4
xc+X6r7e2LwOcpNaBQHsSHvNEQzWAtHVnfhPVbR878f+S7PFhPJFvz0RV18PJGMaaDzf4D07hqG+
RAE6ivE6b6Bc3QdatPHZvvtF56TyTxivkz3AmIidOCVYtNtKUeax2UkfrsAACzSOLmJCnC0tnM2f
tnCNDjmlq42q3P89rpc1h18ZxqmKpBR+dfYrCac8TqCqqoQT4z4xdNI+FYxxg0cFcuuvAuofAck4
Pe4cTSYcHZQbMBFDaG4SMgvsQfxP4h5E3Y+WtGocWX3DENXEjAKwjVefjG+UQufV5iP6OxfBl38h
lFyMJpwuIITIt7yFKWR9W57FJC3kWxHLqT4PMhUwS78g1KqLjGwjRYeO3z7doZc7ckMiRtJmgae8
ogkBEcKORCxfOYuxm1Z4lVgbbN2vKgZO86vVa17gFBqPUqJ4jpgPQH6m0VPa5YnLe35mPMEI2yPi
w/FNbtS5C3NsgaJaf0fBP94pw///EYkJ7BKClqLqrpRiPkTg2kZ93R8a0RR3u9dAEjSjWskP9IVc
jOvi+hptqrJnTQMP/C5jAUWJ/s/1jH9GlqtnYHAfcopXXwBbpvfrngEh1Dj4apj986QkJ5ZtuS5N
Ja5nzjciZvpcjycz0JZqxIO/6Y/RQkPQolYHDlO9QkFEd3zg1u7eSlO1SBzNQsBGcgdCMJk8U/Dh
5T1WlU9MoezX5vsTFBHVZs8tI9W6Hus9xt0flaZfE5JEw8ksbWhRWhJNkHAzFU0A9lD+mijryeT0
`protect end_protected

