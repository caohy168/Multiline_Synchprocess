

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R+TTV2BAhe9Ek8IveLCAIK+vyB2qa4TorazWyGCbrxCKkVhTBvAD6RqPeP/JqtRuh2zDPzraR9rT
gUyNSWD83A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XM2mYTm+gCT0AhW4S5p7IlzH34WHm/fa2tLSENK5xQp44huwLBqk+dBcYbe4GM+6wqA3pzoUNE9T
SluI3P6DpsOt14ispiaJSciB+VdlU+Q0e63sKyfq++TGO3CTW5OhLIxojUbYrTbdY4WbGkk4yG0Y
qGwauBBx1uBueCA2GC4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M9U+BjMD5E96pT2zTDB1OSiHn8IS+G+aDNa3MIF/jeClLSPAOJwufjuzRcyAtwx0354Pb7AaFOwR
6CcoWPQM1dcUC6avyG/0PRrtZP/KpXS3/9PiWsaFHPYVLfqBMCUDoraXwfpfMxmOy8hD0iI6TtWc
j1xJUXVsbv+kqOeTUloYmwdRx/8cs46FvZfnFpiZXMFMsTsT9zvmCyNxiZefgFKT064BWsCkg2fa
W2IXperFJQzpE9mXVwGSjl6xDUp55esPyEPcDI4xy0T+q2KtBQj2Qn2DJRZ8DKAvjXNQmo/tbweh
l+RGgbFge035kxDZ/t5pFweR/SYowAMdG2yOwA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
absLoVdCG0/WeiZ9M4NtAUjz+XnLze4vahkoVw40DL65GHoB/ikdBh+LyLQ7V3LckxaJp7Ihe1ow
2yXZZfuygvynBc+n/CI1EDwjo64cUTgVLg6gqySahs3D5Xkp8kFBBxARQmdoErJqqhefej6SXrxx
13OxNfq4vRGx7YG4l2M61gUhVtUX9poQdq5dxitmrLXD1kpdnUsj/YIpVBaLv/TBn9G44WiyRNIK
ojx9q2JyYKiWBfcBh+fpJV9PudrBUPMu8kvWsRizFr+r8Ya09D3o9iJUZ6FWOBiFsidvZNgmp1u/
nv56cp+qpaTesLtwmKiZbrhQtq6YXQvzPpDQXQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
t2oJ825g01R4DfbjT3g+VDPmL9PAyVC2t8Ozl94Xb2xucD77bNiPcvutyZFkA0lqWfRMp8Z3kkTE
OOo/FpGS3c1SP04/jMKLZD9E7DL6iVBRfxa3itPHxsSD0RAP4yPHw3yCiIsmB0q25x8+so3h/QOv
DKZh98m5ku9UnG+pY6c=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
koDeaCPE+GNu9rMKu+nnX8UvNKbOa7mKCRwRUXCmZNo0yL7JuxnKQiStr89+6Ws9bOIbY8P6XKLC
WoSokcQl2MIZuh7gUJ+LQSPTB9HIkHPuGGPibAaiYY3e/6TBvv0+QG5gTvuf18Nz0UQyxRzNBFY7
2e0fNw+zoh4XJubbVaqqBBqTNyIM/naqx2G+DBhvJF/RlcpsJUe2eVt+uttis5ukRD1ndenp7rvA
+Ub6MDtoxunfFJsXEQ8QZkuZiT5XfcmJdkquGywSafJqKksYNJZpGleQnak/ePqKq8cYIbfpqOo1
MlqTFX2khe/WU/cqsW+5jXmRAgWueTOvg5hW2A==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wZaMVki09KtetQFaQKbOEpc8bkgxHSc8zyuzh+dwZ44uN2hbx3K7ITnC8dDkn3EMZGwk7C0u4eBt
eru14n5jQ1LfuUg4cKuwRNAgFxc7GaymqPYSRK9OQZHWZ+w6Alh4X9YWb6UVcsv4sCJA8YT9QeZ2
8PJYA3L+OY2t8Dcx3JcdLeVgMWDrP/zfpXyfMdPpwgBSSCqJHFsYdlG06onoQq2DDJ/SpC0W2oHU
JJAOTss7Cf3giWx2XTrorU5k4KbClTaEv4QAsogatkMf+oa9OfJQg5b7OUNbNqSzTV2IvRXtKIBC
N3mFkAtau93JXZzbow8bF+Y708RmUyIR5AX9og==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gidhQdKtgCKZpycO58SKONz/x64JxoYiDvm7CY7FhAgR8N3zqVR49qh/d9ImLGjAjXhz9ISSvhiE
1TpzIsqbVIoSEHhHCsw8fW3eNfjSKG9+5c0qMghoZBwnf9txWcso6wczPV8wSYfFgOnId+/H4w2u
MtSdrp2j2HeGCN7hmduXDeRIcLF+ekxNNZVk0wscD3yxYdFDWscebLgM1N+Cx8uwWvloVVe1fNSl
IBecuxue/tBnCdqw10D1fC8gGorhdNUhO2bTYqZL/+voIIAXkux7Z0BGx6B2uSJYuZ0j2LS23yyk
r0QDrL3YOpbEPBbFhTy9LQz59rkITBRhVeBqVg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lv7TtlI9EkMH+4ifu40NSGcF5VLP+fQr0uBXzvHjgpvggoEPEBlbTyXFtewlIbLNuHO4GjqSxFa3
oGjcKGgjJ4JKEHh9NZ/42sDCCnN1TS1zrfhPhpg3aJ3aGsOq5GxB6oAuNGvsTC7HgKk9lvgZfAiC
9ubfhd8fCUCrbS2jYuGLkpNxtwRxEbxLfMa6l2yusSJt8g6sfH0aGGBJWZjKnUZ1SyA1DmzZW3ox
o1AE17uwesEX5+JGPaqlsN+jLpbHhpv24GF4NS806LjJrXOO9qXbZScc78Z/R2xMBhLYAC0AHR8o
o8hlz9kYq3NSGSCdEMOcxNjVxDMYBrdZ+Lc+ag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296400)
`protect data_block
Pe4u4ug3UQiPMR3O58ns6rfoO2x/DHablFFMC8mWzatiQrMxEAU2cpclVRqWAKky6fCpNiHoYC10
1fz5e97LyQ1Jg8oknAv1+UsUBF/MW/FiFAEuxa079HbqwzioDsFOKmtQoyOL5GfSulQE/uWF9+8b
MTOru+7mh//PAjLVcGVU2liOFpK8IQzXUu90T6eghT2oPfDza2TVBcWELTf8xx52KUgh2bKBhuX7
7dS0YP35B9i3fxGhuJ2QMTWons+jE7uD6sQlQw2wxEUuAZA93i9IumWa35Mvxf7HW2sV0X0TqEFM
+d2mtveWokSszs7yBRj0WZtSwm3LPoLMbXl7Wi5X0XTGgWhFr14oCt/1B5KMdlJMq3GT6OaE+mxu
ga5d7ldKRQTBzZBT47lBAVdd1xezoRtmTXHmzwLXj5te4WHxoOMmUR6nVY+0JaFBJQbFVBylWBAg
LVTt53G7qPgjeCMG3Jp09XbktaP8VPNO4I/lbTRB952heOZRO6j5Yvqbb8S9KEnFQ35MrtRZGAYC
kc8wIDze766bO/2/P+2RhE1i685hbr7TNWuLzHOCwmdBUpKgYXEkURTcfG6IKqYtdZ1GIrYQNauj
Qre6bF6hZyhwPUacPVriw5HvgGhjn7T+LHmocmCx2PKz+QpdfTAFsD8kFLOg+qW6MQe/PJfLCaPP
jIKKHaqEiHVunC+QEBqaHfCz5NvC849oe1XBTiupv38wKxEDnNaJ9YS1EULk2RajukQfFH1FKDDg
dBFbyOcesQWH5b2fK/92JaprUl5OUGP4YauUHWOj2/0pmxEH9nLT0VTuJ4zD1OoVQ15RxYblSuyj
8YtJDN/0QY+wtm2TgBIV0YtnLcQWaLOtFW+D3wmFdx2rh7yJoQkHAUH6NI8qz3RU77CFu534lmY6
YZMONQVE912Ks3XfvHbcD1nmJyANgRPqd4wJU88s/OV3tb0JIq6CXllCa4SgqxYuNck9BLkqKS6C
1ebECXi5z/FOrZDr+L7rC7XJu+NNUSypF3sGJtaEx/lJvrSOhqaRyPXsIzNlViFEawEtvvPu1kSe
1tCX4biDil1f1DUUQ3AnB9fM1O9t8ajG5IVVwazfNZYWb9JWWSUgVmFaXY4CEEutBQSgbHZkncGF
LUqm2LFCNf7aKVUJzevq5ypkgzfT+DVjKbNgvTUgi/G17+bz5A+AFx6LOnF8HPaLRIgbcW7JShRa
uh6W9vT9tE//5sZpZNgPLL+uPycritHIyas55Iab+Kr4uWBqegVJUOWqjPkyv4oQGHNvgMIn4z3k
RvnqiY8epYhpNwXBH3ekPn/v5g+GpbG5SKq4rz/8AzIfFzgEExKLT8WXSCS9FAuNTc9snEuYQ2VO
5TME/yHfLlwBhUtHYLs/kIAfo73QVbF6leC/GYajo0sXkX8iQaoLjL6x1azoNMcRMfNoYHGIOKum
Y09W7gDvfTrwFg1omJKycZhpytFlEymICfQMee9KBi1CdhuHyDE6QhiSNj9tY5I7FCQIN2EG4SM2
UZI+BVo1+1HmgItt1l+yVS+YYKcshUuEn//DICnASpiEl9J4W24E/VXg9s6GbaPPyrx3DeKZvif6
cBy6A8VzxhDoA88aJ/rp/27TRDlA2W8Ojx/fKAu0Quwgz/+uz0PSs8hFIrkk7CkQk7UatftJS0NS
yQMAWXjUh9lhChLgw3raWwxOQmWYT39s5R35SGr6ymBOQyGHsvqkOvvjhV8255B1UpUkErRHAATs
WRi5v7lBks+8Y/AqFPWoUf+CL0fJ6Rt6mYBf80GrV4z8Iej8ADAh3KRaOASvZkW/BBE9H5Xp/SAW
mutQb9WT/S2qEwKWe1buvuHKIY0fg2M6FyWsqdIxU/VjuAJFXG29UrQg2n0LMAu8ks6H69HfQiMg
CP3u/KxR8DLx3CJlxp/9y05HqlOOieFqdnf0+0XpbK1PHo09waHjpDekilbw586jdNWMwJUVjgKJ
7iNWSSi8pc4vySmpQASrkEFL/cVF0TFZQ3dPuRUHsjawCO6JZRLU3V8xxERbGBeGWE4Cdy7fsnhO
6/ZGPkFACp8phmDLxFgkBQ3Y1XubwAgapYKby+ax5giPpkgvV4vsIyc0Sr7iimah7+3slDyawrQZ
60Wc5IO3T7FnXr8l0krlJQkM6hG9Ud9jOB9F7svF+GZhsmqtPSfyuIUSc7gnAH+zv2DkuEtvt4G0
qVIbbvo0cJKRMzxOxHj1/IFg+ORXYcpo3tD2psWdMyWNJtz+XdCsQs49ibCbPEVCqIptszQpDQbV
O7Oel15Y18SLUbiIagHngGuL/RpeFVgInkNVs/l8rTXLhtN1Hjlf1H6/AcGvtAaA1ssMumTkETC7
wPfGx6KSZRWW0o5IGPcOk9zB0chtRMrzajTJ/UOHVDXeuNSaFcfZHYfCC451NwzoJkCdsyptyfkn
Gziq6H/EQrOaK4FPDw4T3IE8M5NxjawjjIW+rqvlqzerYB0riafjjHUa7ObTMowcW2eBrq6K4xeC
+00mM2cqMlaeEN/9KnXP/0R1GmgbRE5mMuUIqsHTsFaJ4HQjydjHEg9sTUAZEetVJCYAna6qWCeQ
2WuHBfEaSWZQE6CPrzBtQwuFKIsFK9MndH6iZUyw+BZi2+o/oloGe1pR7O9CfZUsM7IpsjIO25zy
8qETJ8W3/uRyvPkNj1iLx+8Lm4RbLiQyxNEDw30IpzM+ipJxUiVfV7dPdmQOCJormjsXLSfYj44U
XinAtFS0IPnuPbGMuHY/XivgjhoxGscZNH146QiaV8NtRnxDzpkm7tjWJ4KgRdp+t3fDDOxGMGHJ
KKQNmE1lV9w39YdztCPQD/r0Ee8qQnOZSzgneJzdTTUEoEh5c3GphL+yl7J2ncZXaj1tSQwg+zAV
Qm0H7zR/FIEeh2uC+/qSYhiRnpnQG1RVvUIabCytYRIecC33cN2xOesuqpRk/M4KuhnNsmuomQ3I
yNgsW8BxIqai7fVUJgfYyGzfvgOt51m/kp8xlSvstUwD72952arNBf+f899usovvuPHkVSAO5XPq
OkZzYtoAT9vF8jUQW2LKHAEyVWRpoNPNHvlIN5Le37/8pRqjKFTSAVHgSOpNp5YhrYTJw4CVWBQA
4FIr4fIaKraQ0pmDsNvZOVnsCF6UKkBEq/RszLYnS5Xhiv2IyPGMGK+DnUKtCwtOfjRFv559j+sC
c4t3BxqpiLAjkPO1VRyeQDQDS/XPWaZZWpAq/NnhwkQEYRgmyZOQkr4dhb/kl5DnV5HmDDKPsY6f
L+dRCztbRfNMMxqeuj7slFTofr/gNaa7IBvdpPeqdVIJLIc+Secr0dE1ymrf4/RRVPuwkCLPPLk8
X6ZX//dd/vCioxvepBaegLkr3DpGRcAT1N4HUiQh8Bq3ibv/KFwTqspwO0TbmC4h/OIz8l52vWMA
W65REEy9wiIColTyZUVrZuHTxu1k3n5YOjGMYdiHEETatG3He7851CSyd5wtSvJtzWHz5TN0lfS/
ZNhlZEXY+WJsMxyNkZkK1hcUhN9SBCUinoktSJQ/A3tR4n6W/bz2GFmg5Vj52jyiXvLMbnt2/qne
wGw2A+Syk0Axzfkz8rfq3WyXw/b3aJdDSKkg+xl6mdsWNZ6Q+erPMhHhjClj0JSBJj3ZOS+lGpk1
BdL92DWYk7IoBvClyy7t66JC8DbD2+aRAcDfHbu4kuAMshUed4jBHwd4u/5S61/beBw1eQpz7Qj0
0sE4GHaEXd7LUTHLj3nzuKPL1LL4ehEvM8ej4YcgYKmzdCgwlSSXRtCrFl0Pt7C+b9mtxc5qKex+
b8ApS2Bb8uIgmQWCjEsSWvfKd86Q19jzcrhuI9S6+F8rOdgF6N8kXwvfXNarVpS1L9OgQAJHWnyY
YgqMZNJZB70Ele6VaFPSOCCmFNC5TB8MwEU/oBUV0INU0vSLIYDDG9+1IELbolUidyj2jURR0dX0
QeZEr1DegFINIoRRYVjAy8AKUjj12hnr06T3qankVXps704J/S48BSw3dZH0QnlBAVC5vLe5+dqY
Jq3Q6HmUnkYYnyiEdjzXgzjELeRIhnVt/HdmRxX8GZFxzdJR3PghUyxPj3K22Lx9mujFnbItSu5W
6GXPDG7RkS20gFZXBrqoquvJWpTbQUpEW4P5uTUS01qCqqmn5cbm5TbFC1xIuMjual0Ds643xJCT
vcCgbCR/Z2U9K9S3kfAl8xf8Su+crcfKD+OPaVOQf24C5hDjpeyfeZEq91zojf0LaNBmKdnK6ylq
H0zYT7vm8cax6Y1kSWN9jqRyrJR8zlOrTFAFM+2ArCkU/kILoJp/ta4BZTyUmxSIe85whsRVspbr
FRtULbcbBGR2b4grh+MvEzkj/yQfypxlhVEoWEG6Rj/idKH/En6VIN/LfgDAYNsdrXifWx09qfDQ
WPABeALuVA7cuAVwQrv8isQydjZY/edQbK4cgQVxuOPrN2UGmqcqiGtp3GdTEFJPr7LQC5YnkK4S
kuNsqMkvK37I8zGXa6f4TD9wR8chtkres1sfFiES3mfxcgsgb+xN1yTFkPamB6WR7fBMMoayKkiq
MYvHuDWG7lXc4Ok3G+9TRWp3Dr/DjEyxPHcBOKsvXaaPpMFkwDqzpbrCL8AxtLv+2yNjAEt4JHy6
1m9kC5/IFsS/Kj8a8WIZq2i+yuSnM9jY1biOOhITE1OwxCu9cSPc1XrT78d5Hs3T3bJTjlZDfrvo
2VKmpQ+ITkzpZaJpBbP54lE/tW+wjCwCd8otnFrlz0Rh2wf8+O2HxBKc4ws5FZFh4SjZyWmC3yZ/
XXIlJ5GBDPY6g1r6qleCRr+OJLpHkO5I4WacAP27ykLRZb6dSPFKDbSYT7EEDBHKqcM2qLxG1lNQ
THS+EVVvXCKmBF1cmDkctzAR6HhmQgMEF7I1x3QKV33va/5UmjodDDyYTl27dmrOZabaU1+qXwl2
vSG6wbLH9DvGTmcF/AEdgA8CgWVjd/iMLydTsLKwXgqMt4Qbae4ShMA7LMiLZyeLFoAw8QWVr3Ln
DgfY6c7AC5q17McHrPkTyK4Tww5h9q5j91bbEXZdt7vGmTnO3+ks86cGDcUqCshXb7fVwiRhYQwt
fVD+4kkKx2BTa2CQxp6Tv49LEEiM3IBwyo4Cpd2EzoJmyFCcuukTRJUi1Afsojpm8piBQK7j9S1p
bkYU3zIyg6qFbKiKJr8/Rha9+l7sXY29uNUTH78NwzVfUYfVSD20GqSg25UNIlSBaMii+cBd5giP
qTKrKcW1uh9mlNlNcKSNHBOtiX4GHT2TxQUDQvunrl1PSlqt5wOyDSA0ULp8nDxP5qEREoH5gqrJ
DY7c4T67mzOQ3x1HUFBy0F4txsx37j4IoUeh1pyugaA+C17TvoRQ4sRTt9dInoEI4FmSzMVWxTo0
wptSYpl73i6XIjyr4KZWSFUJaWec/aZw8U1OUtWalqpjhAWQHVYqa2SjEA7TCb1lzY7AH8+LdPGr
XBd8DwYh3iQ3IbxiqAv8GCsVwmS/7BEQXFkqcsZNGVUqGleLvcMv5qyCT+mgcPJeA6i6i+AMEqNN
XsZsmhQkTzUvsLyvGjGoJn4dndg22J3C2HLxVp9HXTZIKH5ChGTRBNMgOOotZeH+fkXxHcVAzBC2
IZbzuG9v76TEbOiHNpr060FcgX3WqS6qj4G3q1VD6RAabZz3XwrHHII/d7l8OwQX7/zkgKFys5Wp
neTmLBpLE5qyjXHhpzWPthhiXWJA3eutkCC145QlO+ZZX7ddKx4vOed1jYWsqsQayTE2OsiFV/dO
wNlgU30RCCDmJ259qHlzAPh0RHx//ipwklbGiVieJUH69h96YBeOTgGljcwBA9x1ngcEnaUQgt1Q
Mdu01jKWaGhMxoPnA0RNjTlBUAoLCx7ezvKdazS8NTak+3edFSOm2B1OkTS2DX49gsBkfSKTS78P
V8HhWQxNqWFGmH4XJKzgVIEZpxxZL64eyxbEFbVNJd3T5CoOUR8eUZavOwMvS8QAMQGdKaAorD7E
Vltn1WhueyQ1ccA+WMKZosmpFBwPySJUlCdjqttZ5gmhdXhWpF2jaVUXd7aXJtoOGPcFi5iaw564
OeuWcspDi++sKMJRFPvOSX3S43LiYXRxDTcfUAhmzRDJqUEuLE6AOa9xWViLgc6HFJxcMGJE/FkI
yHMoijRx0hHE7uFO9PgICAyOt1fPxYBq0QEIO5EwDZPK1ViGIPzVGSp18KKkF+ux2fyfpNBpLFTk
aJuRQB+BMZbwRY9AaP8DmIuHuNRex6KSIDApiDx8H58CtImA/zpt0hFyVMJvctkidu77vUwcg7Ro
VvV9FuvBkwM6fW8IQplDhJ8RDUYwMghsWUIqy2BdQabkjCsrKMem1uSqW2aY26hRPMCafGpfoQ0E
puOyk3wrVSamR6IPjkMXFZqIjFkojspbw9lftd3izWGGash2gPZccoLdkcXNC9NAmM2yW6EEey1I
vnt4DiSLijAQPwGBb+0DkBifbvM/Cb7l/PTto8L/KGqs8FOZjkWPR7CLvqUvA1ur0wxWTw/gFP+U
qKL2nQjBahEG1B7SmzobjT1FhakbCg24tc8hI2dnSMDIhPLa9cn9IPOy4PA44ysC/U6W7SgDohb/
hLuicewBO9xIVFDRNBa1WL9QocXwYmb/jKlggCA1wMQ0l2kr0EDDcpvJUJyoZt9pXcTk3Vu/iH05
t6D2CqkM57ToqPaoGwcE6eJ4N9IUgMeqGXfBq5kFVhMoGKsHgapLhC2Aj98E0x3RBdDSSgMr8Z56
OnRVB2oN+g44sxmcgIR2bWNk8Pkf9DiyonhiF75l0GUqPw2nRTZT+AkXCAP+F0tTSLeHn+C82EWG
OcH79GQw1VWLGg8doDhJzAMeAEbMpcfrTRYMXG4ZwGBB2b9/bi9ktlfbmTwzC9ruGYB2dyVQfDtE
kUCe8k4rWNm0JmGf8TloGApCYZe4odtehD2h+GcRMopKbM7UYrggfbRHE06vhdxwswgbcTb5bczh
eVT8vCnCBzdMwS77oBfzB0W4bz06ezXjA4RouB2sf9UH766BHafNebCQdsFNjfHrakSpbzM5QDvJ
cw+5dNq5JKH3AHxBEd/rO5WqkCXWLTayKDhGbV66CayeOQ4OD98W/LiawNhk4PVuQjASDPKgbBi1
tuKKFwUVoaoiZGYI7pMMfr/kwyqPB7API+pLlW0HqHhbywaeJH5wCsIi3Ep7lVpYzKSFNFmZJY50
AZA/fTnhB3AJfIcbvnpapy7BAEYlQiYlW3yUL/rJLoNwV1l8R1ouocQkGaTDFN3wTe9d1uNA3zgo
3RE9qyPmZomJ7J4Ar7RfnUhTiWdvA1Kl1XYFa4//7CtqUFWIiFGDTtBzvajwk02Yo3G1Xy9jcCV2
57brheLs8b2A4YNXVGk31uIgtHb5LA9JMeCN1pLgfXHVopZQM8a47xOqQc6Ud/yNSqT7528FtHZZ
pOhVeaL4j6Pq1RiTOVOGAf8/egH4LNDw04gyxFz0aMp08iVh97uKfN7VHeuGJtPZ8wacrJJEVKlo
mlvgorTOpBBXBbJooJJPGPbNVEbQGdJp7csx0BBlajEkehIWLzoxCrA93u2ZXYfx9Ly8Uzmqgl/Q
8ze9qeKMwKHxMPx8czSXMdyJshcbQ9aGOdJSXK8914fgrbyTTjRvyIYPChAW7ATtX7BStl4u2G7q
3zYm0qCt2zHLh4MOvvBNcZ1UqWSLgvh64+aEhZEn8cNqs6WFOnOoTL96xF8zenYop+rMPrFSkpzX
rRlrFllHVWiGoC3OmgjPznR/ASUvUnyZBKeeqAvvVvyqVdT1XFSZSTEBIfhPKA9jzJGFMEi+zyb5
FEKSfpKhJJTHXX8Jv5Vcyqr5Yz1KX8u++a9gMspi7kuaWStSTt5C1gl/OJj7awxfPzq0LLZ4qmw4
cNwI74gC6ZPU7dVZ98ykRPh4Ok0sF6tVwC3ChBiNcaa8fNA4FA+5MP608DxSvlUumc9HJl11mxQI
yLele8pn1cFp+TgupKPb8lI8R/3o7OSi9AraLcu1fGjVe+bEL0CedK8Sun6+mktlt6e9Krve89sZ
MsAv3B6IQd/iT8ayXYhNtUVgJZBabsaUakvclKyunqG+rDr3AfmROb4rTHozFbyR0+Q/T4mm+m2J
QxWAh/GiSCA8WcIRsqBO8oKI+ferH6VE8Tc8DX8bxrh+HX7BFjg97e/v3AuzCsUkHFskbvAOGRIk
VZtz51M5pKAGEbykMSfhbl4LNmuT/nk1IyfxydFyJ0zKHxOTmTgp9KdFuPi/8Bk70OeCZ4REZfJV
GpmDqVPShAQtNw7nP94xzwxkA3b3/ZZ9MV0GkoJY8APNHkrYgagWJZU57HElCoaXHbsik1jVwe3n
hqeiXViXW5jmtmeHrZbqclFNC90gk1nCQdI0wcUJ8aDaqbV8L/3wWB17/SUSDqoFrJTkxoTFdN5y
amrUcRfI+SXTmcAX7Yz4BBoNaz/LkqQIii+iiHmjBpyOpOmrIyoLjM2D8MYX5c5zu5ZBHCtMq63d
er+9HHBgauHVZtHUvSmyOVXQnKs1QguYeftq45KC/++HHadCdjilpl9V9XebJR9H6E7PQP5AsBwG
uJyrGy3p59V0F+Xq23Djy/W9j9ubPs0RUnUWtIVzYrqhOy9PqLPmJ8rDxhWLH+IU46yoZ8H2wUeA
WdBVjpvsR73XcouhB5RHymk/JJXZxs0GuT7WOfB8OhlC8/4pFnxilRZNZkl89uapS8J3ZCCbLBBS
PW3JZfew1lruYQWwvqckiIDwEtakx2Nu8Jc3lsdw5Trp6f4bwm6StsEs83TpdNH7o4ixx9bEieXR
vB84UJvTdu5WBEWGrRLlWUlXKPEiesCTDL6OsCJSZYZZhDCIkfC8p5S8FzS+zBsFjk5nrvC+T/U5
5mQT/QdlbphJYf0zyBC1qpCVCnPW5riykwMXKAoHmu4VTHAHaa9bm1gonnvlDpvYl64yDhA/7Wkh
cDvi5knOojTrulbODdyvDm7spkrt2qKYecXM2fdxq0cUZhKBJ/OiTcoBDUKYDp5Px1HpOFNDvmg3
bNS04GHw/ofeDhXNzlfTTfe9SG2+uWsT+uVB+WQzM1IDA8lPG0QQngQ7YpHDyojR7FWsZ8Fx6oMO
HVyW6owL3Zn2DHWIjCE6ix5SFYvIyrI2R1tn2xo6mh9Qp/S1iTwp+yERZFsxtYV6fQYMMNsJM+zt
CyrIRJEi036Zj7iozULlJNY8GUu/ryP6t4TeruutoXEpTrtXB1qgAFTnMhocCSW6pn+BGpvn4/yi
kF3iJEZGytsv7Okp+MyGBRDx+xqXoCinnLaPg1pZ6C+DZa1LKIURmYo9HdA09g428YewuGp4yQeH
kTs0UFgRa/OnK0/qPR/a2qDmPin1TxET8XdasBz2tbL8h9YJb/GKPlLIG1LCqyVx2+v31RxLTNhg
kkkgWkhf2elKP+0mUHC3VQ6IAMrmDsxRvjm0SNQpDxtt9O9df/zVG7yV14UP4i7PTOBlfy4c/tJi
Z6Boynm5WUed84PKZOezebipFJbAhz60/LrQMme2mgUnRsUuh/MfBa+Z2dboKJq1nyRuiwl6fdVE
iJ4yi0OZXIlsGaF0UEbtQOsdTHPjSrFDWPm3PAmybaq+bB5ezmI8Am5i7CpndiO2OS5hy5LAN2FT
ynltZgzPGXeosCGK/4AIVdb/BsnPuoyggdZIV067pESwdkTAAYFuVtJ7KWO9NkNyReGsdxN8VjDX
uuASRMA4P/JNFntABYi1EvAtz6R9PzN/VJf6CGAyh2YzgOLWVo+IopV+RGHwJE5O7ILQZhx0eWcc
+FPsRcwFbM17MLIFcTe4CPI2wjh3/pBCLYTjjEARbxbcrufyFKsO65vAROVeYHbZHbPTmCRQW+ZX
zLOENdeFJq8rMNocl9Bh8tGUH4u3GKM96JD7c8CTkttXIt8BVLL8TyEl87S4YFiGZ0g2zJ2fYxNq
hzu+dSOP01RzSZzT1+dXidvGyx3VO7YC7ejMppWNFPYILlQLGfsQrezCvCwwj7zfH/GHGhLNWUv5
VBpy5YYO/RwCyI74X1NRR8FXwkEl1z/V+OwF9ub+Ti2I9I/h6k9gsJTELi3JB1Luh9ooBCCtDOEA
BSqDiOC5WpovsedBZr49RabDLO8QoVoA5510fukBhWqKLJePCBESFKwbtR3LHeTM02RpmBd26QJu
t5vrIBP+rgDfRUi3HdXIiLEIjzSLpkkH3IYyTAa8ihxS9GlxMhb3YqWfaICnDUoKPcCqXCm/4Yef
xckjJzFxXKBsZLBrxW4fKjJ5QR45kjhLjjdhKAoVNoMyssySBMLAR58ul/dc+G/gpUVGQ7HDmFKG
6TFWutQyMNsbkk35BA+txjRBDP+N3I5R3+9DC6/mcCTL0/8sz5Gv+/pNQpI7xHVPMp+b//aJeosw
rtqjuAhuRQNVmOdFa1RuMS1qpVlcqC5kDSmFj/ObdsEHp985BFeiw8Fq376vfKruQlSQrxtpqGrA
ahLwu1xw0Dd/JAkNUjXWDuqfjiBFZFyybD2go+dLoG8bwLfj0e+70ZAONKJ2uoNCzKQufW4/suNH
OPIBfg4tlKzhzLcjBxxnNow0TQvH3Rsxma+i6OTIBz2Zz4tD2rodKRUqWbJBM2YZuYWwTbdP0+CV
b6Ahh2/uMXAzk1T/mPHqO8eNQv54sANrEflTAUpWIJhEbE4103XkbqtHCSGcGULUG78S6zdEUDGR
tWtRXi2kpaNcDF5g0MZmWmM+VzpHZpzXlVtmeztRTtBC3h+5KpHw5vE2ZnbqtAP9XNaaxtDq9zFc
KyRl77fSE5429qhs6NQl8ybDs5Ziw9RJ28p46NflKLYX6ubZbPyWfsm/rzvpmGkeJ5kcy6f/6GDb
n0J97fmq3wVJh9HIf9t5k/BAYCJU5gF03bTTRztw1nDEOROP8DJM6O8VcG6JyWw+1yNQxdxaGkh7
AE7Bp74qsSMOnVy6duRCZ1Nf4BRsH88sOm2Q49sEWnj5U9VCYudG2rY2dsBXSYQGjEnJn8YRk+U8
FtzTk0s7xI063bvQb+yWuhd8M+Rvcak+397A+/+Vpd2qYF5ltklUTZuKDzZFkkxD19Af7ARgSDRZ
OgWuvHmrW9DE6G1SWlHbKZLXIHwMWhNFl2OjhInDGNNhZtvm1jBftQOS+Xz86jG/Ug7cLMBLBtOe
aweJyhoz/al6MhcVfYv4hOd4gNQ3TDrbaG6dUkJSs8Tc70z5IdpxZk7KqcJ7PoApRMUQH1b9Jusb
kTjeAUMDHN3cYdoijam0sksBdWC98/YHtcuAOIDmb7rAj+p2J5X6WQ+GnEpHUkTy4U5OmvChyzzf
hrJS8lYhh+wPJBLVPUtC6kSprm6m516uHn+ZkAw6LYuiKCr6bd319ZDzFNkbiP9IHYCoZhAGiKLe
yRRvpHVsf4/oj+o0tpCjHTFN3oyVV8s5a9nkfp2/Ze9ARwaKm75DRxY5PVUiR6Li96fw4r73BE9A
yGru51DahFErk6WfkUkBlcufJG0gpyw5PuxNs6YGVslL61y4IBJL5eygJVRmvuh5RO2zoJq38exm
vPAHcP1N8PWSalMZWuOOHYHEQdBrXd9YyYaI6XHt2g8MvWFTyXJTYs0xTkjTZaeFt+yX9Cc/hK+2
8/M9sLGs1W1ZX2s/jkgglv2iSDooAqT4BoFPlvb+r9Z0lptdLgTlZP1PmIExHadJ69gkeqfkhX/M
Qzsin9/JY+j6zRgYpQXO3KcF0X2IsKJfKcwcwbqIHjlW8ZimtGOefgEp1Jyb32GNnk1uKO1CZ3bf
2PfcFJR/6PQ7hQqAv7nR5dUENSb1pB9wD1v0Hma2KvNFgXUDotkfyVFNUPXPMi6EXbsUOwH38U/9
Ny+kN0H5tALxfA8w86PaFArXg/AAP3JRp86VC5drR0/eqf02tDkANhkziAIUGdE1oI4Cg+S3YUL5
huUrPzW7CtmsSluVAqxUMp6jX45HY/3+Iaqzc2xm9WJbFLmGGTJIUcU7j4th8ghghA0dXwGtw24o
pDATqqjmXq8akGt0A54ItkxeMUdjP+B4qujCxnRITJIvzNefZ36VS5ol0FKEpGLf+jM3cpUUdnAb
QMrMzKVP1RkIkkL6InIEIDOnEarPDTyH4Kp+5tNWRMVBTg5/+uMGayDrDG+jMNqdLbMBzR4WYylc
fkhEhPEaQs+yLTRqR5BMvxu7sWVTXmKQ7JeJ5a78KOnSeY9A0wB7EP7SzxrqOBU+bcS/sTrBjkdZ
4gFAPZ1kzemMeTJ6+T0teFz2tWqD5DJA978RqLP+d1XN3sI4KhPEZt8atqEsCy/TSmD32lHu84OQ
9GTlnqn7fhyQhKnSqAZWerhx3bGM3XfR+HLIWNfjynKWtr14miP9JEQT0PpUbqtBwFbxOb0oCdwh
DB39rTeYu0jSuwLlOYPaSVt3C/TRGCjsLLbnONo2COH5GmRGlwn5S9GWfRvb2bUMOyjhJh2p+xPc
LEfxyzb4TZJw62+wrjMUGl+omH/m0ddgUl8JRs//14lg1oQuvoHIxHpckYn0wFxRnZnMaW/9KVjN
/lJJSmkYF+MVXKxF85sq+6NoQrYNFu1rPlz93xftf4s6YdnHRKeGyooG8OKudpNjCEQ+44jThmFY
qJnhT0m+X/TmoDIsi34l7lxE55eK83mi0sC4gYb/uJAukAA2vlVAtOwDHLW4f2CpJkW1GdmrcYH5
Ccu/pkeAf7THxbHZsveBqGmDhNAiNMwTb8+wMPzfAy3nfHZRekvWk7o++TMYBENZZaouCSG+J3pT
fERDqAUDGDLTjTul/S4EoRoNDdLagcwa6Vk/M8MJOW2FeINRomX1znSX5hxfhuaw5VlgEO6WdNrM
06nj7PLC0G2aD1rNTY0IPrKPFFUz4fH7n95G9+lYku2OjsSw7FlVZTHHXPx9RLid2I5RoAC2Wfkr
uXjMKBDq2YhE1GB2+eZIWx219qQun1eCxMyrU/nF61yKOxl9/omPzpZIi7gYnUBl7e6SANeErSOM
4lns130qTYZiGuhUJjiBUfdT+ALQJ3xnjIpL1eQqtRxhpkyXqjGuqbQ/jn6g481KiDGclYLKIKP5
nOVWdqC/WbL7U+hlkabxjwT7Us8YY0Zfn1tkGc/8ad6QETZDTr5jRFQiOfHNckQZpxJNzReiWoeT
wtCW5FIU1wQjC6kB12FqhP+xMxDO+13VGlJreSit6c9qGO0Qpy3CvSAczTA2RJrCRoZfrOkbg8Av
1ZrANT6b2YVU69CjY5QcPDTgHc+yUAO8VoQSKyXND1rDm+Obx5tBYRwjBmmkyqjonY2pMPsOYieQ
4+pBLn8BrN7uAdrg3NnzU6B3AK1FjVxFchU9YyY5ml0lpH/4S4Hv1gSTjvOe+KuvOeyXw5bzMa0h
buVtLdyyMEtFYZ0qkSHUhfXPtezxkVRRxRID0zAjxo6Emg82RCAw3KE8NKyEz/CvVA2DFfKJlncz
6W/mraXk0ABLyDbQJWC1rYOsJy3KvAAMEcGB0CfnxxIRDD23gj120i2cxOVnBX3VOswLsJHL+328
cF+T6XaPv4WhnCOWjaMrWQK7zcIyoHuZ3pA2iMeIa2xki5rrhOriAE6WLEQDGgTZxiJhHYZMQOPp
za6S/7SCUS/LLXpH4EVjPjv1KyWv8r0kjtLRIKOgNR2cKV71vpCrbxLj4bx9oPUcy0ixnS9EiDvy
nRNK068wLhh7Yl7VlzhHq3CLrdTei0YLwEJN9eNc8Wd+8nwpq/EyjT+RP5E8ponuRL+6zl/Bjrbi
ZC5R+XoK3txWocqEMHicEH+SMX7xjjb0EkxD521+h0R0efItNyudQgdDXfj6DYmMlt9hY8Xt+lQI
1EdMZ7h12ZD5dg+EOAcgT8BKthgA37+jSlXt11ZbzLdehz01zrAkQD4NIKQYojsKwG4gtk95uzmn
RiPpHK9oYPcfhH6kQW0Hkmy3tje8y5iWq27A3NtmmVW43MXmjSDnQO17g37gi9IWKIUCwz9iQljt
6r0flq2lD0QjCmu2cT/H2G+7VeW7MjHKWbArNcPf+vbtrr0QoHlmZuPr1SDtMhxaBSfGPWZxf/aM
bRNtYpc9pvZ2Tm1U7ak+Fe4RlXEYzxs/bhL3PJprng6J13VhG6SRQ0e1jF0jJfMuwm1igh5slky0
yKQcoNDoRGflbztpUlY5Ai3VcUYq+r80skJdVNxV5gUnGgmksgD2Te5MapmF57l3S5Y3+adip/9h
NApOJqQeyhLFDXtP8AnA6xLpUXiQxFdzpkivPB67+JsfcYqT4A7xGj06O6ekKtGaiLP+GseyImh/
/HuZKBKBxFDikhUiyrSFrNRdVU+xSFIrxffDfFL1AE2P31O1i48kYjrKQIVfp/NTg2uH8l7rgldt
s1ygqFkxl7QG5MpXn+D9HcJsajDXZ4/JDe7B8UDSHwOx6KeyJ/braZd5dKu75t35c/4ZFFzm1Lzj
uTMKkLV0fPHGRcu2v1QfpCTor9xQVE+E2ivmpbHkPLYC13P3Z/qADqMoYIJz2cnxEMVQy/1whQXI
PgCTTQTkutEDujfXKRuCDNW0X7WQ/iLSe53tZTg7hBn2uL5eUA+4+Z+HL6waA73XU10UYDITVuqr
K0PEMciFQlzeivwVFzV0erL1jaKtPdzpayBzOcSTJpbYTFkwDa2NHQftkF1IRFBfdNsHE3KhFjf4
tqo9G8uKUb/8cdXOeQtKpUFH/hLajgYz1kWfGi/dOuPj+aXuGyg52G9ztcwh/WmRzu+/lbQCBca5
jC2kex1VWC9BYGuLFFI4PQ1/zb5eaqtXcX7FycGyUv30p4UGVMTeD0XHp0gl6rPHnO8THkHPO7aw
pPAHz7vmESPAJHGpYAZWjZK6JL11V0QO1H94KgWl8DbxMcqytpt6A/N4sjhqKt6TzWmTy5gh/B6U
wDWAIJXOwZejeeEpkTQ0Dl1J07ILcodAJSO8DfUD/Zso3VlFYj+b80amJlUWTpfoNgwuW79ezDvp
Yisd4JNJQthh1Rtaf/9hIZqBYyIkubzSiYR8bTnljmy+rxYi6RtC6+o6ZKCF3zr5lxcceppCkXSQ
4rmpxqIK+211GsyEJc8O8yWi//NlGvvMgvwIBcjlitf5uJfH5/wzJ879XBH+R63HsRyc7EFk4vwV
+i1fptgoFyGT4BhJS/v/NJPtc7JGmEI1YtuBYJtPEtuEM2cpzFi5C6pl8zZ36/xLKmA/+iucPQY/
n3mZjx0bP3JynpAJVaSE4Ef784KJKnCfB1hdeW4HxeaV3455Nb5m4a6ridw1Ytj5QdopNE2MQqNQ
8Zx0qqKNerCZtU/7As8FZYUnffO5H5KJb7LrUZzpS0juUHA1NmMhOXxz9dCxMUWEVl75e/9uZk7G
Gi7j8tXTrOU0JAqcFI6hplcm/Tj+D/Yzz0dYVDr9+VCqhGNzXNTZr39q6z6pLla+TkO6VLDkVifZ
O45qQLMKAXNtlcvZFJvN9K22XWbWq38svZl3gkpBnv8P69kPxAO7vuEi7IG5g5vBpK8K/EtzhJGg
u55e4MbEqX+EGZ2AIj/BZPgxPb3mmkykp32tu5EBy9Cg7JKF8yWyhL0VATrVFHaE22RIM07FYrT/
gB/mBHB8IWvFq0HVggIiQzravjDo2vyi845/zvbNsxRnbPYEO3Bo9L0QLCl6eIwZi0RagtAEgjMI
ffa545SW/zV+5hdsZ8PUYanFRQghXeW9rWtxKkZ0xfBvgJEKxFYD4Rv7ldp5qLghy5Yghk1Ynetl
ilL+yHDdZLRRQk5k2iuH/VNyjOjmEMQ+TJYA16z7h9f7GyPxADGZZ73QuwOMEcd0vOC/GUEV1Kb9
U/062bbb+w1gMEVMIqejPVnRnVoGcXyrzWi1UU+aCLuOub2GXmY0JYPMWzmzQ6+nFMnw6DpM1+Ma
A1JvrV1/BoC1PsdpsDVmbcC6uwbK9nxpfM5NsxYKPUMGVy+zv8M1IL9UyHdCPREFQciyTOd2K5L7
uTBsJT7Dp3AkgHOSWDJ0o3Gh+MjATcMJha7b5Be1x9fuKQY0PFFGfWcMVaey61C5ZSzen6XP24BY
KC6cUb7a13pCcFh0RjNv7wgb8nu8WS8A5/v6xJUJySTAzwbWQwaBcVNrmeEQIwLkNz5k//2AvN8S
hmMG42diF2exMYq4+erhhL9su8L0cHoPUiD51rC35tRRglJU7vxNfTn3AsiMv7AgnVQykxJYzZ4C
W0lcsSAGtHYteE9CVnxjhlxerrS3Dpnv1p/Zov3AF8aAuc2BRY87U0L7bM9Q/fQQVLI6DwBZ4wto
1q0o+YCB5PXyi6OJvVE0Pc3jr9nZGBU4pYMjPCxK1vRqv5mmfRlz6Qd/39JkU4D3gemAaed5naNE
31yDe+znq3uynQLFxerAP+vFESCT5In+1QnSo7gOZ5nRQ3A/V2sxwXo3n/8KfqTkT4T11c3Cy5mn
1AM3tepVV+z4b/rjHljEP/HWJwPHulgufuoJOFqeOYOWsS6cgaYvJpa3X/2GJTe9blbUiF0UOwUe
uID39Gj2GCjZBhv4bfLuws7gQVcuzPhb41ECHX1GV8EZvevj6nd+Lf5Sl6fsy+pOP6VcRVmHefdY
1Da9e5QlqlQz1rM6OnPM9KY0t1b1oJNVZ19IbBE6PR55iiF4aRozUZ8oC0aeHZQjL0RAof9y7qfG
ZdmDyqOD3JQ6D7jBJzeUixmEZg0tMrH9FFskNtXWwoha8DaAIriCu2kc0JOqb7vfLmiW0dwM1BoM
WAyATDPItNCVuoj9dXLoFZLyvlhx6m2vPoFi7p3GKHnQYuFfst8a5j0SWIwJ/VQcVT9H6xZ17wqK
euq+fthPdSdEmUDc4ifMZvpWywS17ycvM1/GxJ3RInXmsljJSdIythKmhSFJB8JuDAXdDY3bkmRg
d06obpv/bcEljlb/dRSPWTRN6NAqX/38/V6pBcdOvGBLPSy1m1dve7JwU6Xg2zpzJOIqxhJhYD8t
60KiMiwSH8IwfFqz0sycg3WqPG9F4aP5ld3USKzCqrZDokqvMccB567aUFxJfYagpeqpmIUXjKND
1qQHNlRqOz3UoiYd/ShV30jPxX6Z1kNNGyA6wPIrni/178GkZMNVN1xdkz9WDB/O2GKv04x0niy9
GtT8yP0leTEMu1S3vFRmiFjUCJlhSMbWeU14cA/HUIEGkU7X2aRGdiU1ZoNiPiSEPEGM7EpsLKXX
kSiAGUO6iofIs2GIJS4Va5aEFjtBrnvm37DR33XPZVy60ROIxr2/9ga76/KbTO/hwx3OU5HDn1e1
20GbRbuKIexztn38b/TSU8ZQs/Mx4VNyH2txH6T3vze8ocvii1t3BND6zeP5MnLwZKr1FoJD0yQN
oBnw003M2HrjQ8DKAFK20q7V+TQ83lQZwhwxTl/FNdvu55yAGtxRNdPIzjd9xuZ5AmkXjSfpu9/A
VRPmKlx1uCVj/Zfyl04w1QcLNdyCveWsd3gFQCSKyK2EmJ6JO9oP5bco51d2YAhMAiUMY/KX1tU0
rs/PHyQQHiBDAP0lJ8PHr4j1PGaq9Cx2NtbEcy2eIs4bPcd9OPLc/wPNbyUtbOIOrQLdgEPEsZWk
PRIsfQkGwoNqtOlVyeqAS0qLC8GYPnjDLcnzouipUECzklUwhExHZFY2UpmPzLpA2OPkqa98BORR
vVWN20KjSswO0fWOyC2UKlyw8lekWkt7MdZU/RNdlPunYKLmSuwBgJvg5JW6+Jn7tSswjuh37BjY
7lldEso7F8nT4Tq3MZZ4XSk/kpybnUtpg/hv/2jtOVc6+2g3/q+mGt+jsJfldUuWvusUo6BNmvY8
cuUW9dD3MjQZouPfymQyMjWHBX7ni8683EFx5aEcGVr128YHLZQtzXZqehVAW2nPv3U7VoZsoKNC
2JfYm+s5sfvxA65D8yJkDX2DCpAc8b1mt1clpzuQa15cwh4CBIQfFmUMVJZw+bGlYoNHOW1/R6tE
x6rWr91rDK+iWj9BkFzPVJHJyCwAvnBeBjqnrtgv+EyqIcac6eLa9Jxkac7UlsXYclFR/Nqpxh0E
MHuuIPolZWzp7zYVpsTRJfkLQPsng/Ff4qqna6hs3w1L90v+ARZ8ZjKZbh1VumqIuYaoHe6AxAzC
oubDeFiXYTxHZc7k3Km4v8KJZ/oKpdqqIpqhlWfT6Zc81x1WhDMcxhOHBV+t9PDgOXXGglUAo4t4
aBMQa2pqOWtOvz8CtHbqZDGgPt+K7T6HQN8IiabrbqjPeKhhhk/82YbDxaYiGoHNHAgzHMS9SDPD
Lwk1UDvFjBpNm0yZUF/fVdThwS3IyqLj/NAWJI/xVUNToboUOT3F6U80hU92cHt3BR3ljgvVgYS0
7vlzLFsVVIWufiDcSP+KobVwRXqwI+b4i9DHSETrvlan95K7YHEjNvPQKLguiakkkSBZ8C53b+zu
srxW31jBhs2+XXcggBYcWHhcY+CTXO1Ycw3G015AKX6MQTbEUNytnW5qq5590WWAAP/dpqFmwRnt
rJbmzPx/tL9doqQNVTiNrg6k4ICccmBAvaxHO1PuwFC2fmMwYZqSgeztd8d2ydKjS4mkCpk9Xewl
48TgTM8tppxTVu5DoT5fLtjm22ye83j3iBdakgi1hH2jNaYxmS7lRZCsumX1JY5vN5TDRajx9BJ/
squ8APksGgYUpxv9LeDuasn2f4cYwng0KQ9iEoGGfIHP+ox42+TrUA3Zq6ihfNdGAXSCaJ4NWCz0
rx0fn+6phSK8ZUqIjXuwG2kSS4ukPDklilAAab6Fc7PY1h8iBPOvJixELYnkw/98CQMphblteHsY
/YQvZmNz5zxpO2kQSHFohzIZ4EO4Z4xifZBWnntWPLPkSdm/NVFEB/649y62v7+Ql5Qm7ZTdGXbJ
Q92iqsYQb7WvlVoGIelu4im8QZY36irJ/u/kPYtSiFw8cEE9Tw3B20P6eruwrvJeBNjYigetqp56
fxO08daSpL3ZBP4POGowUOD7qaiF84wI686M11qnGjyIh5nP0bjNrLjHwYChqIoMp4OtKSN1xVRM
l6d3l0I4wedBSeDiNxw8tIIFCHOPpjMqn47nB7MbSnRhZXh9voUIvtvXm1PuSxTQ67cPt+E51sX/
/QkKW9duglcGAlTFirEzRVlb11o45jb3CwVI91eu5CRL/ImSV3b8oG/R88aaGz3k9mdvh270++qN
e3pb3Gnftf72CgSZWxjKWz67pmvoWkUeRB6SVYRIZklCIRgSZjiJkQj6yyIOwMEHAF+BknTUjXmY
LYxZjpoEfoMW3iOLuGUDgKpO9pSZJQENI0pxLgj0RKZ+8wpS9C3WukFT4lbU+Vw9kSXvMvyQ4N/J
lwdoar1mVVQI5q0JOmXsEMRiqtETUVot2wYt8+YYbU7/GU75jMUFvwsX/ELquxJFwlgp9Ho0Ghzk
03jgRGhmkgt0C1yknFXLqFqvNSqf5oxG6QIeWkRK/5TYk3z0+iIXC5pJ5ZO7OQHnRw5yJ9askTDD
iV7YsplvtPFCtFgEpaRVi0xobJx3cJkqSQwD043rT4OwCYQ8iJB1otM/owCcZ8WafdnGsls71zi4
4dWL90OZa81Fe+sLcQnLmbXVrtjn81KyIlYAIySqvG9+4RMZtSiQqtdBI3YjormQbPZjG+C4mHK7
c5Ru3DE28G+afQ1Cw++uSF5qbvyGmeRJOAeNzLAid9cUCC5WBS+h4OZbEqzMlLWk+EqLxsHrriqD
3X7yUw9Z6Zznap/6/8NAvVw61yDZ/NJfUlsdq/NKKNrXVxyxZc54bVTNnvSgjm76UcabsB5YU2K7
XQsEGrNVOZ49EUtZs0Btwf3SFu3N0su8vEOfMqsjmHKPi5L8BnjMw0mXJPG7zGYlX2JAgTf0pq/F
zRe7r6BTgI+VDmLKGU94a2Bey2i9iFJWPRtG1L66s4QiJT0b37qReWvpIi7JmczICFSQbrAUK8SP
GLfKZRbq0YhBXwvJHEin/o18N/9TbWl+zGbEOhf0wflAIMYz0Adnddzqe15lhHEqELaIB7LgZsPi
IGaeLNc5SOm2Y1uUNRT4Pftmzy78S/kfQgr7nPCYiHRJ3nP5G3X8T25nM2OE3F/+3j0vg3s6F+S+
LWhpsP7C++vR65+al4Ok/5fMDB5jjeEHFqWoG5TU/duyaV58t+k5GjWwYiJ8BCPa5NKmeIZCOKjV
k91vPVAu3J804mJQ8uw5FHWBk78fQ0QqJxAi0oRBH8r9N70UujPauPjiTAC5/12WFZPGrkoKY8kj
9wg4hQjF/PzOo4bFQ6+EgehgBPxyNwUaVBQtgbpBGFxMMNGGvoGBs0LQyCJgzsPoohPaLSV+DrGu
EgyJD9EuLKmBMZFbFNbXQLQLFIpt91nHgBP4sgBR057KPx+r2umhVktdgAUUx/qQwCRNErVeD3ZM
Yj+lUNZB1AxOgj9UZ1aGa9Aq+fBCVZQ0gMAyDxsSZsXD58wqAg3moDqCa1Plqf5bz90ZBgkH3jmt
BBleLMUKgcdEdszHvO0xGkum1aJ3aV6fFYP1CopI3ZZ6rhoqmKyACkh6lmFYDOLw6yLSveLbDFlr
bWMbjiXf1q2s6WICPYT4zbDEohPNaktUErud+59ohJwELHk/DN7w9tsNc4i4PoZc+hExvXk9h16V
Ucn0IFqEmWah1K1kWOcbiKoghYBLeGYDC0sxurXNWwHl0oVN4OcMGAGfB2QiY87NJuoLGJlQQrVR
UT3CtEvbNpI7M51dEehmvJAXiFZgy1tupWMgS21RjD3mb33cWyS9xn40DmzuualyPiKHTUe9flvI
zdmOZQk15I0Lj5Gn8Oeesc3KWZGeHX92ryj5l8c34FCUPjl/mug3/y0jv0Eo0Y9EWjajcxUOTtCL
26c6cJsy6y5HYJOSEIOaRRjVwkyvAykuIwjkgoSK3/5ZxW6XfmrOSHFEWUKVQdrLbK0msPepe2mX
1eXEeIQMe4rjZYBrx11jUEEzGTHi3vowJdmxhhDxJ2ZLvFsdMOkABVCNB5Ov0HZ4A3Gvdfm+BKLK
HKcnvUJT5cLVKZ7QJGjQ0Au9PfDC2rpSgyA0D6qdQyYJf+GnzQve2m+68Gk1IUMN/IYhbrYSKN/9
w4WiwHL2ZF4WcDKwNorHKodFZZy78ktUEZWgDza9uQI0gCLSyB7MSC4jnIBBFkgz5skb7cemjlE2
MO4E7QIPAwaZ4/fkpgWU5TstRAZWY5gj02GHFlVkQpuLimAqdq609+nznStSHbTgurNIM7a7e4Dq
KFYt983TDgsWpZ4IDCLoDvhPjSoJidWzQBBk1obH8QYKvRTtQih2lqjr+JIqPBVuovf+GC+6KZn5
l/1hjSR7/G2ny4UJApLK/Gru+m9oPkNYHDihZdBlL//xxTXvmp5R7CbKpTFjdnfwmhmov4axoHy+
jwlC4ZN5R/jvfH/0mJ2MYheQfHfCIbAmbd+K0hlwgu4LMOagEMYWcahysF6fnrXTyIaSTw6bXDgA
lO/+Q/ldVsTwJ7WD0BQ2ITEnbwSduX1iS0UAE0QcfMi1pJY4+dTfEq+W8IOQ7KZSAmFsv65TidxU
stJ7DjGu8hAT71XdD3QZVVkszgye23a/dUEuaMufwfrhJ3pvKHCvjjHOtZv2LMQLHLy/1xf5y+U3
vBly0AiBPa7+oQOhKNwHJHlp7fxtgoQh5wkdL4CBfYp7iOLol+ir1RtVoLI8F6lBD6XhTUt88NAH
dMQsIi4DWJ70HaNLHwlkHBEkoBZ2dlnktQ15GkzzmVmdMZ4djJ0JuMftwbiUBXgNrOGU/gkLXTQz
wxfZa8SaiAT0ICiKY6vxw1HtS1edvJDbUipc6c+IWZ7+huSKM5Xt1spxVMUA2fbEIVfmRI9WtHyf
41dwepulZmbwAafWaPDHsjiVOnKqTgQMC4ezaZ5q/Kn18zxEXXdzEZKhgRJyU/wbj1/DcEe1qTTt
2BJfxx6UtLv5sKkZOprpNvsvJY7I/nWQutILU0Cec1plEK+Kvuxolnb3pqzMdUAo45KgIu/5UUfw
xWyAUKn2DIDqZoN53uiZTugjTofJqiiXyL7Kg+k7etsMkA+99Jz6ji1eWnrMWgs3X3Ngff8h6V+a
nPF6EdgNQhM6gqZ9y1Sg7jYRTDL478rCuWo4L/7/eZydIRbKn6GPORWYz0BrkEvVksaeZ7pIPUY+
mjj3ln3y94dR1EybmhUVXRxacUnhPxJhEILsyOAcmEmGHYN5vchPWSfl2id2LvyxS2HJBqubtl/M
GRs8Zb4Lf/6EUzrM03jrORTqz7q+OkMbipnTP3PPdFWRlNiYXqKi9BU9X3zIoFzbdzSq/eAj5Xtb
0stU20LvpDvyd7praF1a12FVtTQSPeoma3Lu+d8eUralQUtu/5SzKph/DfWTQRw/KRNlJ+yjjVvo
ZAqICYAwGYZRuTRa8nXTJnI0prQhQBS5SY/DbhBP6xRnxprsfjcFV9DgeD4u61EwQqrCeUMOvAhO
7pT5kO5DsaN5nU8AUVRgUjQTfUkgHu2le2gywdRM0OiYvT9RkjGiW5DN0rURusdLiIpufW5gIuil
8DoJWHayRF/lkUT0ZG4pYaeO/82Bib62Thw7VFATU0+BtC80MispIIUwOCCXqk0WLhXxOy+BAwwZ
alTGAF27D2KMf0/g6QekRe10vcw40E7bRFYnZrOPMqnr5VbIxl95va+n9ddMy6DXec3iE0quHgjS
KtYyLXNUC40jpipD4287Dk3x6ZgLJqrrlFB6yP/NxE1naX1G8BOZukvk2wPmwR89Ib8PqzYrJfoA
rBK4wTDJJW7NKV00nQlnK1pLzosJk11XXK5TGnyrA216jyXtUwbLJB3/PpAhxv8pGSdegeLkzzC+
lWiiFEL/tXYa2iqZmtN93MJlIDSXmodyQFEh0cOq+52vgD5QO+wIChFDDe6iZdRDT2dnk9zeV38p
2ESPFm0GF+4C4tICvLJ1s1lu34OniUZ4BoySLaf+3SL7JNQnhDOrYO4xb+cex5l9aNPVGUjom8PX
Xo3axp8g1sK5lOlYb2jbuhr7ntd3k2COTp3HrgtepnbzWFrAJst7jEXZmxfAft/D8cgwf4cwT1UE
gz3R4eWeH/Aeavj0rJCNKiRz0UZZMGG2nDCWT74CflqDJuXscJ2sukq0FN5spfI1pL1XH2QyBWsR
qhwOSSf1X5iiim+8MC6ts8j+If4Q8o7KoHjpt4v1QWkhdFt44nJHnynKLVPU1VMs94m345Yb7b/n
sVxaP+fAanH/7WHzyQaGneUBB/FmdAOCrXjUHdyDtkp9KUjRdFfgtr44M8dUhJZC3GVTXkxpf8Vs
cCtrQ9jw9HwIb282/z2f6yhU5nae0RzytEbLoG/q0mDkKWvVQxH80zmn8p7JJdjjLpJTljgOMoax
kv4FawkgSSvKZ/u6mCPtYLnpmTtyEatm54cOSrZtqCU0JOx2Ox6C63MLXC7fGoNbYBH9HThEvdOJ
vCSZu8EY4gbuP5J/RMIJyF+W1kMNWiMJai04Aq4rCkoNaCfKT+31LEKCiUtgdz0tClpKZRtWNwa3
fBEDM6l/NL/9dhvkJo+SPawz3E4aaRuFeExtoSrL7vwLjBJgIGO7uvVRR/C4YkahYdYv4wUCNImN
M6lsfnUk4UtkshJi64+Lg5oEQ20qG+oW/pDiSpE9w3VijGRJqFpjrw2skD2TTnqfm2Sy2Dmn6slT
ucczQit/gem/HDGjUlWdLeOx+grgJG4cK1pMp3L2AwveQpHiY8L9r4+JBPZDI9IqBHoGuJxsKV9X
KYYrCa1SjjBFt5rl1866F4gxazlNnMOdLhymqFCH7mbn6TUOBnPrcmKIIjMiIG0x0Vsh1FD8nSPl
4BkeUPwBcwKe15wHE2OLjrL5greN1HQpdC8ZdHc/mJtLLxrb+3l40gubuxCHEE+c5m0j3qguX4i9
1DE05Hd9jL04Xjp4MxPViZTH6rXvhIZhBsIFXz5gp9DLH+pOtYh6G8zrfmNc1nSX+jTb+T9GnXwG
nuM92tr51ueUJs9HFF9omatvP7GFWu/07OqH+tI9YoCte26FfjKOVHv1c8HCSl9vzQivEpK35UNm
Pig+azJirHFhjnQtjfX4tdLJgf4ERUff3w2pPyWYHn/n03R8gHeuc5rj5VY1gQBs2fdTFubP99VD
mRlvJ7MosdgUEeKx/bGsjLFLyz4d6WI8Tp5P7w+DBSKUvlrUNGd+HRcDUkzwhudslbX/OfLfaAqC
AAs1mRZhI3VXFl8Nu92RQdz3Cj7o4WFNckvBtQxXKnzkmfHhXyQhbglq3xbhV3ZgfSTrbJpD6cJr
KfeP+g8caJENZLMwi0zEfpi3Z/x171w2su8AEV7h6zY+0S3RpirglDRrOAQ4tP6iM5fCFhDcobr3
DmlikueFfjgFAvC8SedldZGK3+UqHeFf1cte/KV8ZTCu9Coyhq1JNVfqSxZ4QuU8WMYMsA7Ei0Rq
2Y/tTBwteF3/K2nwnRY7pl/aZRM23XRtOaAEkmQA/17g8QAVJR2LOfG8vmNLuqPT0YMnmtJ+UBcl
EoMt7ERa3eEFFXq+H79wU4IED5zKoN7kqNkQFd/Tv8X7jLe2YYs4f+uQpBiIFPfxYNXaUII63En7
zqV153GYNVcFuYN6IJ9MCTgGw9pSn5wA6uORQoqirIuNphhMPScWBdjzQO+f6FbfD0Q1Fbjgr5GA
plPAT9tqkVwJ2T3V1yJKFR/1zgh/MlX5UngOxpg6ol71Ptv/YptUcm6W4geJXNURUci6spulSE9k
0eqyAVizmblvzd+Aqcdr8G+3tACiZ4CPDkYTNjrbQo930nl5rdvwjEvVwBB9xGrMup2ll7v16CC7
aMX+Q4rCcRYClaAHzwYyWIqIIS0Q+M3GIlwzW7Srr2/mUliD94/JuNtKHEs/FEqR8Lce6L+aQCPy
L2wdct2utu0FWQCovHGVpSNtbJdwArbUp8NJcPYcmTfnZYMwP2BycFw4nF+/ZGzqX4/hL/8EnFVw
D61oP5IQwmsXDpi0yIT6PN+U8VH9U5Apm/xHwmgE4OD5GN1RyO4C3Q2xlsH5V0gsg7/dqnE9nf66
b/b0mWGGVgpz1h0l1VgbtIlLveyVfs3FGuVlqDlerkvlJkycdlwMSTYxfCd3zCuCRbYpsS62Ohde
u23Nbsx66lUluUZcd3w28fvXxV1ZotkiRGfq+HONTqu170n5ehLt1/JqpkfyOf0Lqh9/ru5YisXN
qRitHqm1V87IaIDu61pOaicNE8imvimaVda60yZJ5K0xLiqzIRnctbZLGzkLokbFMKD9DYxoE3pN
l9LQk54YkFQg5x3UhQC+hrCC10TrDNhGmppc0qMQ+st5vKfCLoTUo96U+aN027mx77Y/KQDPWuRW
1g2aDx7V0d8XLiPpH+0KAt95BpoYrE7a9EJD9PJHPz/tbez+y6baojnGA7JWIvyaI0CyPM1/FdfM
WFhWsk8qTPl2j2GEahqEGlkiOEk3DYgvrhb3XvaH6j2WdslsZrFuDw2nMltkF99ZywOALmmZtN3o
zCKx1UPhlYQlLdgG5t0KG13pCJkylZYv/mfVWJ6SHtYvEQ7BsLwXGYnj3ACZvo+sScwfiTG8qzWV
N9f3/jEjWKKeoRAiXKTCsHJu9h+hAnF0wDh1JNArfUZ2ml29wsjxvzcm1VUVaGAvXdkRRGXHPQC5
zGyI26YAm2JAFJ9Qrq8wI+2PHhvExs/9C5mRJ5oHaxa7zshacDzUF9CDCBpolxyIe3kKHbrEoL+O
QO0/ybw8bkWjLUU4eiIu70zxHxAGDEbpfwkS7pHyNrD0MxeyfpE3WI2kW3U31gXJ8gw/ca75YcPT
pIlBchvnEGt4axrdxSP0rALX9NerHIAM1FtVfjlrqbyqngWBb8zL5+an2VwewPogrkm8MgbmXbhx
oYpvFoC6fL8ysbcdet5A3+bfFiyX8CwqM+MAy7XpI6IlcflfWRLpd7XkEujSEaaBGwZl2RRLiwx9
Dy6KK2m0w7WQ+UFjALbuw7Fu3dPvstYNtB9t7tVAavEp+xybWbKZPGit5qUD+D3r1bAONuJBQNeB
uN69e39kHZ4p//jHKDbWRtf4liMVv5GNvcUvF0GssKbBP6/+N0byEfydEKKiQLvYDuncGmznrLIN
bE/nmCkOI4EwQkubZ/OAEgPQb6Q4Zhx+1eetnu0XuM0JOcC6TLM/9UT39wo1u/rvY2r0R2djvzw0
Xc/iZ4PXt04Vw7JFGx2yrFR9h33CcZgnVBt6ybQtLmT2xXiA9PdeK8bLmXlJalq2lcSNArjTJdS5
xe1qZJDaE2PbqReWJ6VgUNDJRG1/LgGn5Cu/HOhq+U1o97G8equW98KWn6Gw+p028n6MghZX4GRR
LiWbVtGwJfDLzTADZttbAilVNU1xHhbBIkVoLkp9b+9m+rSK8x7uT61AkBSZloHu3Nz/S2qqvZkM
MmJbOf4zyCCPleB2tpqaMZNvHmr4Mt8msWBSseMYzHiqKlN2D/E8ZbBZXVtr/wy+Pj0f3/NmMaLK
gYANfN3th++2zBvaCyi1r8ByoUCHBJmcLL0KnaEHMQYRelDwhxlwVuZCm5d9mOmsJ606YpQj3uAW
grDshnJ+3/m3jHIvynYt3v9H22hFhFwzLSxiLbROtKKR9XvCc/4J3xy1uj1h0jz2ksBTYn9qRXq9
wXSXtMUxnCLeTE5Fl2OtoNXcETSM5T2mOMXrSj8YqvI8U0bf80GwmtBP2sY/QQ2Ofv9b8NX/zwld
5qbCQ/KF7NpxuICE9PBiTNxNxtrh/cKtFVrV5AvT6bxxN44xwKyVVTFXYyu5TviTdNfid80FHDqL
l+Xlk/AnjU8VZahhi4c4K8JWoW2Y7fUSu0DSIZCwqdR4lB6Mn14ePJkB9Vvtj4JjTBft3qHZ8tm1
OsPM/96At7sAgx1JGHPyAVPJ+yDPuvJtH31JOp4+xSbYB2K104VAa5JHhKhZDGNnWmONI+RIn0yj
Ia82l1J6aOJ6xI/gu2uP4VSqIUCFf75DNgMr2ra523SI5VhKU3LELcFvz02/v/7DKCnbDJC5KEUi
TI+U8yUi1hP2ji/IBMg/SsvUx9JCaDfW5CjxPKzE1xNxGnDGpL2UTa5Qnhe7VA0ORyqAODiAUst1
JzemeAnh/keae8hvblwIK6gEmIT9s0EjxV5/jIekwheeV5HVvZ6MeEyUm5fKcFLVDx6D2hYgf77N
s2EZHihfTRUoJfGrvItveFTlZBg2yvtuBKGh4Cmf2BVgyLG8yHbEqvemqUphPSqgZ9Ko1lnEk51D
e0vMKN6LmCHMzgsEjjU3Qz6HN4CLkcSd1xeZg77N7YLhAqEEYbdn9ooyfBC5ENU3fb9REPTowOtH
3mni+NUtICS0JeFhRYhYhstK/mWGsm12XdzVegJ7qYsIA31wUwsADQx5rbQDHOVevooxz/5ABfc1
gXhvltmFbvXWZY4khQVcvvt4t7vNI97k6Q+Dpnld0nGnx8kLa85KG/Tv2NE45wwoU6QRcGG4QMyx
TbwnFO2vIr7LLYGrjDJDg3kkPLhQcnq9CDbC62S5PgllEJnYqAaS0QJJL9DHa4tvKeqsanpHJEPS
CmRFu7MAOXDbOEN+jecJjuAnCKj+HwmUl+tc16R9ehFZs8F2HPqfNwpC+tTXz1TiAhZbRIcn2xxw
xmotWz/5Pz0Bq/V32BaUKRDkk7oL+kk47RbTFUYvNrRhp5VxrWNY/QH6v0rry2Nnw4naa0dBxjTU
KsFEzTa52EIcerJwpwnEFY3WI8AmZBI4wvK/IM/sISB89aEd7t9xkaFLmf4C1CR269ChPa40DFv0
4E/AAzGDKwPwhAwDDVacUGQN/tMRPK8l0ySReUBnaVFJ2udH1yiilixFHDTCMW5Apj4BUdVt169j
Ug/FmxTd1+aghye7BJtn4KAFP0bJ0DsIbxOLciKwb0Ip8aR6fmIhQXjd8dVmnWZFRmfg19jBTA6E
5YCvsQcFJW98jnFF0u2SuHu3F2Kq2PzniKZtd+zck13Lls9KZMRSkSlbKKHXHXNZiGWygeOkPj7c
wSE6BW1SAqsqzdsbSYekIFQ90JBTf3R2wdwBjOkXJAK5lCAO7pb7ZafKFlw2DqEGY+HMimxhAYhj
wS5duTjCquFxeYftbAmRSHEjvD8gz7+78ti6mmPH6IKMF+V/n0dA9V4F25T9B+UrcBskhbXVv/ku
u7o/vdBRF7WGiF8YQXRasYbKClyanfQwePH6wdx34eLY/64npjLqGeMj/WHtkFlc81tpd7oJaBVb
/nmoE29Qdp1vz4kRujrsj+7yJqiqrqgoPE8a6xKqwuh1buUVRECwwaaxtstnglbvKpKXFFm/VWvc
FvRJtFGe4Ar72dIl72Lvb1rBlXjbfKuGad8f420na2pIHutqLNAs6ncyV03CPRe1BxcrzMnQHtbP
Fa2MH83XFoisq2zD7loMkqahWpItukeq9aTSHMUEcC0dHxMiYNyxJOpX8AW6/TR8l43q87JbpssY
l205wiGMXfBWi3yhU49qj2XD7KZa4TG8NEDn9Lo+5XeOEC1QFq0Y8MeuSQSXSg9ImBGdiiTi60Ah
Iq5sQSNlxBazzPtMHDCSMq7ivR0sOelSWAO6uUySuV6Y8dQEjLOgLpFUOP0qF3fKFsMAXn9ksLQD
RMnYDryNluX+x/4mLFwS6J8WaJzrgEucvJyUAtb/j/uL/1FDm5LTCt26tSdZiVndC6uYb+UUmpg4
4HA3MeSDb1jAl4RfIHWuWcLAt/7a37D7skTRxtw/cLsUkU1DxaDRXqZ3YPvK0TEOuS52BeIAyE8d
qL8sHX5z2bEodqFveP+hqpZssd9KWDT7hEAgK9qOpKuLHU86OTIQVq7UpYdKBQyUoy7NvG91mR+D
/67p9ZAt4/i3d9oj9ftU8CwQw5NyFxkeH5byuwu/DJYlxKdkKVOIUeATZjl6wXrux7RMPW5FqwRc
k6EmPg2NmqZLX/R3F8wSFvU/0CYO8+ZwH0nrTRjxBjdQurwyhNFLnM686Kvac4WEBAPR3pO74mCS
IyYptaVswkKCe8FqOJFbd5hf6Vmx0MlIpbJ5M3pwPpZRIIwspbLcXxh/Hb46jF8g1IV5UmrVyD29
0Ys+t8IDmgg4Qgvq/IrFqGFozEqTfFnqaaIJ3p6k9f+GvV6DfRhZ2HX4KbD6M2S8dwrpEnrq0ul6
gXPB7QAK7UO5vlCAWuOEAJAT7LJLu/GOg8IY0DWQYCPF78i147JZcD6zS4QqHYN/plwGnkDHmKEI
+0SBAitPhgyvsA3p54twrW2KIYz+cRhBoI0c75/JJRuKDOfg7HNGWVTLWICxPogRDMyE8XVeDAQv
dezoFXVyb+WStR9WJk8SZP3JABexWMOD43qV3YXckMcJF8uJD0I+AuS8mMmxxssgSEKmg2nipPaK
/3otvKs6twYYF4Xz2GBBwPcbYPaX/+RarHkh5PnzZXfSpblqS0tQqcRR2txGsHST/dzmn4edDQyn
Y3ZkS4wAHlaEKdafmmzsOc1hSXliQXi7u6tFTVId8+K+nicQVLnKxj5fqsqGIQlEflz0+nZjWs6k
viJA+Nz7MakI8y+17sMYAFz2D2oLiv+8cM9nuo/XISoFWc0O/9zjWsPXA0LRaUMWXEl+XHPkGvdD
HPusbeMjxO6j6YEq9gnivKzxonAphJ4gAfzYRoJ1XwkvMhDmgy+0j9ahA4TObk6RSpJvhHXUKIFR
8whb4L2/YLdmq9Z7i1Dj7SxZZIjvmrIH18nFCVPj+A+0cLcJ6yBzYBFN+HGmQDeMugvwQoNHt12p
RpgRwVSq7iY1uP+7FD/GrEfKEsydbRvJwFuo4fBOVQBfn+4uLIwaie1HgSzGi5wcKtsae7zg0R1/
9NfvPLlHpBTD1rrLeoHlabCnkxvmPw094nS6ERoLy6NCqs34d2OlVccHBPolWoQYk82ER1z0OEEu
JUWzWnup226099TbShArZSZyosKmyHNCCK9rh+LCP2ejtXb73VV140EFCA8rP8SfU05+KJi8af4U
7bFO0iw6Rvobo+mi562hsgp1Krb7rT1V0EzofF25v9UlPj5/4JJbUSBajD/S5XfQcQG2lmLmYAhb
o+Qevf548mws6TrquagvlJDooiaT1o0ALZxtlwzuSFzHG6ftpwpkAYGt6cjPKtRDc2E4xVPnzGOz
49QkBbY+/biKmq5aPKJoVaQYk47/ki7HAVEhSClZrgVWWiRMUKj2yiZRkVt4cDUVBRZ1RyCmhD0R
QdvKWC1HbWsTigMCmeaLqbz5rluIquLA23rHoBf6ftkxojfW0irJeExpAMyc7xUrK3C2zj6QYxSS
vfieZ87S/f2uSt64OeqIrPClHbd7Dv5Xwxh12kRMBGNd7IaSG/Z8k3v5iFVcoTNwRV6/Waq0DTBf
oe0DPahv/5XMIib3aHeEXa/fqN8mQxos4A9irMDZAUuJj80YlZBoWsCOpLXoitGFdFyu0xtMSwI6
Fao8hQfrtNHFyC6TEp+HcqSkLsXrknks/6Lg6fWptl98cGIYI4VIUMPPvOKYMq6FLxaTU85/W/Ks
64nZCtFf6LYiC4ZvWhtDeZiNK/xpN7ErMooPnL+y+qW4S+z1Y3TfxmC8Oiyl9KBFP2INNxrFaVzK
vYmmU1aVmsh+K/PkWmE+vvAQlnwUuKJYeKEdkaqjHgyFDGbCx5tdftR31MEmqNHKta+Yjs5KQeKO
uoDQ+drBV3UEoXUXhiNZp3+tYyO356WjjyRxLX8o7KyIcw8LblGsUsmfObCfnxJyPrmsCExalyUD
sR2ywucv3aF2xazfgvIiXzAOg8NHhKU2ETO2xals4r3uug471NK5iV5g0zUhy5lP9rfvYCOzTMS/
wiPTR0pOv0w41fmgSI1dcVRB9eH52XOXELGSHBH3DnmrRc2iW0nLE3qgQlmlxmpv6GzeKENIHyv7
z5Z4+lD3L0Zk3nZwW6hZg9ojKNTR/9Du82sDfhLpc+vaeIvD7WXYSOBCTrM8hS9LFLBo/vfVDAOl
2OcGsu2MZQqt0OdYU3Tq3r1x7bMZQQpcJUC83PLZ2EKH/6XB0TnNXyiQo79NaEGA13oHXTsO8cln
nmZEq6m/2vEgI5mXYjvESJDySDBsnjpzB9aTiiPMTDWSH+7q7W3NwNv4uzDMp3gCPO78CPPK0Vv9
SVNHd6RoGcm+JPcZ48qmUSRQEpaCUM7m96xNxRsEZdqzslxASlzgoqR5mSdXTfDFxzJCErReSrTR
8VbHX/FE2xxciNYCDZwnqxeP7FkumuY1LnJCcpAW4PrJZncJ8Ph4mB/gEU3JkJR6KPiUDXlymatT
jw7K5MTMTeZN0Ge12nK3Y4uU3OFuLgqIKb32q9nw6XG+cjq+rKccTsu1rIEqPuoEGbIdi79cGWl3
t3mZce3CvqdAm2/TkOeFZV/C+0IlG8q05HYwvWIBc6YeOdJmotHffqV7ZbggVnKCs/gspFKHzHVB
pC0ziNQR0XHrmPqz2+fIiqFWOO6ApapQd3OWEoahG6HTEItm4VGScIgz221czPe+9x6fLHmFvrga
XAC9fXAniz3FC1yKvok+AjnXX9nzoYkyRsSvJF85vFkNmUBMa5PrnhltdMtmjscN7qsRwf9OMe/m
6Uri+vPqv37TUs6783Ygh+zfJT3Km1/c3AL9te9AAd9itxG0X/BDSeSPsCfHp0LNoN3VOteqPPPi
ZEDtNz7FApatIbUBafoO5S9UzIiqxIb8wF3U67Ha8FLHatsSFgHtb4aiGJyapMQU7L75RSgCmxr/
26n0apSaBAaTbsLI8ZQ4hessLadl5/qLbzNEIcHWX9/1LDLjauD6+SoNBAgndRkQ7jZxdFw6zxqz
mdFzQURAXPs/Lzia/R1ABIQ4nze0KrJ6lC9kGXBV1EIxXlLbk7i3UQ4U6r/epnkHeLnSGpjR0orY
/moddyy7mqxxBPO0IGwlRSIXDJsFlgwnSsGCyPzoD45e7zZvoaa1BP2+DtebYeGmWX/8CRllsemQ
pH7d0ubkcLv9BXT5up3XXm2jFdxaRmsk1UxTYz0bLU6I3t9HUSyeHdBAqwwxp57eQ6H9PqnZoKF5
rKm0D1aIjoEyMXSZ22khLihSTAIfBjLGeBFFaVHNUhoBs3hD6XD7ITjQET5MITAc6pxth3GZPl/8
2KLJrWCNflFCeV85JhoWTIVWy4jZyBvZ2QUP05L7Qf/L/R6YyqmTUVQHgO9furuHTxJtAyNXA10F
RTSfQ5wArAmEbWv6Uy/FCSOeYpcf4WNV5Vr9M7UEw1X57Oq4FFwnv864KPOPRtWJNeo/LZtmjiHx
zDtHuWtcal0SECRVrys5g1EooikfMoghmhmSMvpkxMK72XReRT8hZl+Yz3q1uxzITn8LjcBVtI9q
cvhZZfYnLVPHBSszDKn9T6EwLcLBoQsssetyS15l2N5PSuQZS8XmEUalPPeXqbM1vLaUyIBk+wH/
Lkz27blZ+jfpD/bfWIbJkYH42vG730WgF+5sXAKJhB+BQKBxF/z1cnfSlvN93MbKM4U986Mz2P4p
qYwTxVzQEra3RgGpDSzLGADM/Piy1S0TXgqxj7/ZiBAymTrsIfiBI/fTYJR6iYJS1jAwoTSpY428
UFJuh42pSWVsQe9GpJTLX9b/+BVTbQDSbM6EGBUT398NqBUOHO7beQ+W4diweoDbaUymHDT0aaC0
WUmM4aWbhxLwjA1yHj4TuMS9dmO1kOuRrQHKL7w1+Y2sRQklgLlCeI9oUwFRRHQDEIQIz+TMzN2R
IYStWYPyEfly5cVedARwiKqn18/mLbg8VygkseWbEMTy6bwaVOv+flD0yPfm87ADhPpNrshe/ZMI
DB2kmmgiIGviHX1hpKx/nLbeWKQxGfxe0XdthldAmPDIhyPFEnnTM7ZGAdS2J263xBG0SYY+neIL
xehTumMPFyIknKcVg07+QtBr6Yjw3zJc7OToQ0XqLssHCNOpq0QTrgp23Cz0DzZ/7N2wSTmi6KbQ
538DWSO7bJWPKrZ5WR8yNFCyprIi6iZ6MawpGYfaZg3IqHepGlO0aVrNRI3tb/N0NY4hWfcsAUEk
QbG3ttXK69D6gLzOMjT6Sn/KtBn7oAbFgKf77UvyAr0m72SisQFOQOh7zfBQD/cGCagE9HBJ8AmE
CgWUsdpFOrOOBKs3F6lCbBBTERs5nEzGRgBK4Pp+vB+wGC4Bug+JJAevGucqwGoKLhV8rWIbEnB4
PgcXqvGlu9R2/LvPlwftDzHA2uzx5GCozZy++3obGKj3lRFPknHItSTqHa7StRxweWb4YZcQvMxo
JUJTqBEljaeWY2jyUe/axve1ImRlc5YhAvd4yJmbItA9o91JSCjZlaWZfaNmhwty6RfDGI4Vh7xz
rbGZj2TbhAP7hSU2bAIh4vw5BM/wL28dm3LGwJvoiNwaISYfMSNw4tgFC65Nadt3GqnZG+89sMT2
2x+Gz31trfjtwFBz6nTQpPjzgxdHfJK43iVQZZYfMxEvSqnCJIAYd/HptT6qFIMxhW8IsLQnyvoN
GXCnupkSZxXnlZ0RT4bhTvkmcJD7IjOa9c15lMbMrGr0EXTg8nwxFDHzWCwbQmV9yaA/FeF3hsjw
rJs1QSNAB2F+PNShimQI3jucoLoXKr/QI3vae2JwAZJiI+w2lysm+hRqDq5wtsGuA5UhhBrB7X+i
Rp1g7sCe+HswQUHLxO6d+XH4bJdDkn4SsxiPZNc794wwKwmpAVkEjn06uGm3IS8ET3czTRnOu0rP
vRb/MYFop0+xEGEE4sMr/hyIlsqJih70LGo6iZNmhhiBQZfp4zH4sw3txb0aw6/ToAitSasKT/+7
Q093VU2Gnl6+wVbcC20L+3gZMAWWywWxp/+dnlPTDfLSt2LNqcmJd0+doGgfEbO64gzXpthk4fq/
SfT0dD+Ij20B8NSy5eQuwIx7n7NRA/yvaPb8b8znx71p5XHNf0Qfwa6ZIYbLkZvl8UWf1AiT2rUE
GlIeS0Yi/gSw+9ApB9S8KfHaWmHx1uWWkB4C/T2xVjVucNn17e9cuQDXTGYByIlTm54uBKbFPI4y
i0VNZzAoPHCC/PJIW0Lb4J+xsUIveB+kbZqZmL+dTy4t6epHlTKbkkcGizljti6O30nztpqHdf4P
80XRV/tb3cJs1oeruOb3IAfKGugUfzYgnZMlXwrHLEeFPk1ZgsYZh0b0y1ExMm+LKEl1YaeQtpaV
rUROmzZkSabRPEQAtXMCiGcCgNQsjz5o/s7BA3DQgALloY0HAeFruCcI8Qr0cu5bXfW8g5mdiwZl
FMF+PBmZYlpvRuga1dgld6O/b/L7et50XK7p9an8SE/4Zw7k0fwJC3wqUQRc9Im0oF3cNCWYVHf4
6M9M4sr4iq8bzPZxOaDh2DG7OzF8mz/m25YnLET3hiGY3ZCU+xSE2mF8Y3FR8cfXZcJStsVfcukP
cOizi3oz6q+HOz86nlRBEHC6x2cfKHjbPFSaYmdKc169QzycDPoKWr0kqEjkYS2SSLIJqQkc9o+J
TKFaS13/d0s5CkDDULGxlyV0FxiBIFZ/oFwDN+IpVN/ARopQxBvqwbrNjLks773IHIfRzs6WBQWN
ebs/ui77HJV3sP+4674qW+RhvC5gq1Hcp6RTTBlbT2QVmZZFIZ9l0W3z5ZynqnPUvLNdL2kup4Cz
Bc8OYvT/xLJlhjgZ5ZZ+9oPrY9iChto2PaBWj1jS0d1Z9LOhUzqSMXrD366/qOZIkrnbskBZ9xEZ
e+bGt6Zgsa5RVnXw/k5dCTHz4t0GSajlQx1b3zWQcKMnoqyfwsrkAwfhNeHfyLO62aSyX6sVtjTT
x09wDVrUmIvU7qqTmUcoZCRCPIeQfRBSQIKRoUd1qe6Hhle+B+jvf2tdFHjnQDR5nITzetZc0VU5
6GPxwz4uGnLN9uL1piiRzcRM9HxSfNXtpvNfHH7PZC2Q11bQU3EkKaOJPx6dxmdS5aOHPqCkdXCo
25lUba40pOpQz9S2AY22eplcAe5DuWIehUm+itNsdUhUpv4/zBoVZs/qkYD4zJBmQjeL3yR6Z7Z1
nmm/OxdIQ+lIdGvTQlFjVFydPxsKCx5RTidkMREwJVGnf5er98blgWVlftLL+S1rKtw3whccebLF
kbM99v3ofdaTGJCZW8Wf0O97Lr7cDsbag/N6y9AyAsmvx4gUXoBewWjUgTeLJH2n6CtMtrS/jKyK
CI/D8mUbEq//gOUwxxUag57OOFszLHogqTgulskg8z1mH+tZUPyfqmXZGwKzMXDlrHPBSvT09NXU
zCDakct/xOagG68KdiSroaNcqMOG/Jstc4FmAqCwYWJsA66lrTS0Ym/64v5FvciOiKwgsuo6ArB4
snxwEH973FwvrxlEk0kx5g6oazL+ATUsmBh9CaWVPLxX19LpcEnTUBvp2CCQw4itgfbh3QSQ2XLQ
z0cEg1HfH4OUx4IZhRd92XiLPnDrat6kvbvHN1NyvHg0GlI9aui9gr0qrzh982MCHynAyZyLDF3I
G5nutY1E6ENbz69R14Wpby41iUavTV0FWTKhuUtv4kGOl3F2Oi432eyLQ/l0VPn7DcM2HiRoWKO0
aPj6fs9XRqxJWBWnWjGG28XWyHKBLbMpYKe3zb/kex7WQgafd4T1syD04jgC5gVrbIVb5PHQ/dsw
SPvRHzmGCR28dpIFUuq9+aP26zUXswHHK4ngxzY4NgsSlwxFMjRurvxGKMsugayoexkAvLz9j66i
0x2XL28OTyIx/rJxk8h9+EkECczktJ7sHsvsB7DcuUcU1oNvgyYb822olvgEhe0ybpEq496Iq7D7
P1aiCIt44OjTWn3uSEy91WODMtqiDPeNwKa5v4XeMTihyUOEvGRquYYHLlND4uaqSCvdsNwT2rr8
lpMRUKLt05Qe9XV2GGYaXbn8kF3EkO8xLBTBn0ycIOqPk+5BPtsoeTg4VctdLcmok55kKfCnqaRy
7VIUx/fqqKQszQ/CAUeHQnP0vTzF6kGmyTvWFhb/Zh23S6VEmrKCeXWo1kHni7HLZexfRWJKEQJu
1c1qB5D5/s1Ztlc+z488ULRBc+vOZPaaOinQioDMDV5MBRSb1XV2TbhmmhNTCmXHDbSOtO8n2BTV
gETJYJwGWRR6RgsQrAV5fO1B19/WbqTY7Oob9sDhNfECrS3rxC1ayrGklnV3VfbaBOaiJ6p8Zehh
paIWlle24Xv+zQNf9o/Zqft6LLaks2m++RWA0R/NPEJRb5LW/p2OFTD2JmW4f+KkzHyHOfayqi4q
JU/A3eBfxR79mSg8ZfL9kadGonAFBd2CzUR+UfbM9sV9C7uTdIy2JGj9o6k2BrISRmTOF+F3ov5h
gOsPIPmLblwpAryPlFkvQ9h05hHpr6HxBp0lpi11OUFFVXqaC0FKmUxDvU+5MMPEQCKuqNv1U70X
bTmBNIUDPLUixaviiJNqmvg8ajEKbHYDRlRFJLtjCqZE8HYuOqCEbNRumQ3JQvZmXxR/RNo+ytFH
gJe521ORwepAwe8oMjzoiQtHP3Nipzxx1KHG2G+YH/yMEIFXyYBW/hwk004gX0nuy4OvSuUj7lrT
S30h5pMXUFs7e9aSwTrD1AYIdJOvvFP1yEiiwwl5J2Qzvbs8g1Sqv5MMFUWRc+xY02Z/oSSK+eaE
kJm/ssfS2iaIRokoUtnrnPHGrtgNuZl5qNOcQjiU3e3gAUc48/E1+RbwGgG3UsKktDGz92QNWUr7
pBXhBwi/OLmVYximEFYzXcFMgyZx7XstOm2WtKKXzIip+MhVQGDdTilb2srBqBaYbZ9V1CipO5fh
qNIKQLVU8+s0Eqb/zlD2OuOy/8aCnrUroPbxhlQCNAeEAAeGYEM4eE0nGQaUUJ2HdFbCX+JTHJ5R
v3MrJAOWGdYtwOitYZp89HVj232x6uh1cyLVBQo90hhi/vp2JTYv9g5XYlg1ut73l3lYZ5v1N1se
ghNz6Oz1077g355WieBeEIKig/0trklECVD/e/D8SrHxsMizA0ussZFo5W/kvcVIwZAISXCx24lp
zGdmzSysIIz62JoHEL8m+Ik2BDXIXVlb77GEUi+XS6rHfmjTohy1f59/jXkKOV2071CFSwWH7X/F
V1e58HRxRZ8UC5h9JNdY8DzxF25JeEcbyNG+Mvhr9vXpdyAvEpjFa8g8+G7NkQ+gtwi9qre9O7be
9Y/PpAfPwH6TdpQEM99cO85ZNAa8QVo3pvYdlysq8NArVNGUGxFLkprtmDyhX07a3vhyBVkYA3BY
gE1O0Q76i8Pj4/Ox8Pccp1sIuR1xiaiHEB4WrcA8PUOzYXC6HCAgzd6w0BcU8thfHLBK2aGB+FV3
USOQjLraikHLHI4TivhhkeeG3BV3tt2OlzXM9aMwBvlt1sqBbD8oqrXK/YyXa18AKwDU+6vGsIPP
vyFxDbs+w9AiUQVqEGR35tGXYkghLBZD2aDpH9VgW/uNWbQ1J02W/uoNuAR7UVUC83oTMzW8x/Oq
Jc7HHEh5qh/WIgnSNfhcZr7aQfiC1r0KUlYBcwLFxblUQ5oBLN2qSAYsBkewqB3PJsaYkQT8q4cV
DzQA7qJ9CXZloKbZwsD5KOeUnwau23nqqk9/BA1kSvOF8rbJXnxOXBimY6GGitQay6d/lbaGiJGs
1fPuZkHO64ujegQRQM5SiEii0jh3WvIoYNM4cUqbBUasoX9BbvLusfvCXNEP9M+Pdd34AiwXh/m3
Vav/o16nKXsz/Z+mILN0GQCpILLehSw1d+yZqUEx4avdQEMz4jpZccFcBs+TC9DSuTuQADc+GS8d
Jt9WH8sQ3WgFQc4P2lmrmKWf5Y7kVcgP+wxQVVHMceNpCFjaQG6h3i1iZ0Co/0o8FvpRZurqn5qH
cPUcu23Q9evwx1m/5twB5OlXlFGCvZ/Iegd7LZIr48irVUl4PwwU5DkNaG1ikHcPFQkg4mpY1rkK
J10SINeS+UCI/DemE45g3AJMyJi07bAmR9GJ3d84DOVm3/79jiAemu54HzduFApfHQsk+G6SlIMB
X9Fr2TeIkLHOmEq02pZIWH3IW3VINwci2WNC3j+m8w/rJRbI6HvWer3ZTG+ww6q8p+37EIzrkXoL
dJDfxSBepnixJRrRZHSFJdW2/mfx5Q4Fqm71ePcH8UjIjVI4pB4prcbwkDOwOvhRhFbqE8JhIf79
Xstrg6FKUCRL4MOx7saf9HEufLlTc4Uern9xoVu+enxNbkoM1joDZA/I8CkaBsx9wfyRnwy2JyHu
VBGAZ7Ca0zDulEdkd9n/f8Ol398tJu4w+rDWmcweR8nGXfzL8jTKJk73DN0jbBmNKhyOtLP/6Kqi
cHInU4kReA9I4VliT78OIh6YP40TA14kBEnK3M1ljl5nybPSnQ93AHRACSrUZVN9uVPdnBkY8a8A
A+viwxhYF8H7DKJFjKO1r4wNrbSqZZ18dJfgM3po2CvOMlcm1x0ROy/S/gCHwvgDjXrfDpRgTjYL
jSTxiHTR5TrHCsOC+mtPMXeRNhO2nRHGkrNhFuV3sU19TOK0sUUmG+jby9p6D2nWl0mszD94WDTy
IVLX027CERNnMUngqusaQNub45h0UB7pdCLIuFBApKaD3dappc/sK6ZAXx4bohWJMJAV93qfNxiq
4McUMQdfKtP+WC2lSERg4ib5C0lrX9jXzJ3UhvTUa2Yu3gPtFed/c74ojsRSz46UTE4UvSkumpRD
ATi4jg/ypXrqUPSsZxCNdUfs1BAVe0Fmn3fANcqMnWojTfAKmBWnJ53bt/3gLGPiR26gZK6xzhAi
bGhvG0RSbygZg5NS4gH/oDTLKoZlQi2xHO5YPou3HrJ5OZ0Wi/THHU7tSVlT05SPGTlJLzak2DD9
2MCaxTHXt04tDR9FnqMGCPSsNqxQ0YQRPSzW4oJSPAn9TUuFEPx9fttvRenIVRh3Fcy3T3sBWRao
wkTu+smqNlBi5NQk3N6kd1oTF2ei1rFnToYhMTx26tDlVXr/cbOvCer9Vi4ZYWg6/9xRjAwtb4Uh
+UdxDrVsTMSPECMbKHynj7YDJc3v8xk6DN0aBi+1A5BIC60pbKAYpmCwx96m0kU0nigOO5FMRmTp
eA44jEM9GipVBoo22PxcZkIEqW2/15iGP4BPu1yIiPEAPO5psJXVLBgZBPaijwcVuhlKR2sP0pE8
ktxz3oZwjGoMZB8Ul7FRFKVOkLQVVqouMZb5bsivJySSCIEbKnYMK5S4iG9UMoO1sMKSyvRevvRJ
dZ1RJCL9soJRpE6fBEvHS2x8Ymptxv5SuiWwSoutlUXNA2GoZS2OW91BzUgveok+36emR4OnRVYM
ggm0HssVMgfMTWwgGaNMOdNGIckgDBmSIcDfNfyPxeyTHGP77E6BY0v812SSrnafRpeS1+rntmZr
qhgScPso0PyGToLctDSI1sN2xG/InyVgVp/G2kc4Z+6Ra+8hzaKcOorapC/0WeiPO4WvZGkqoNf6
TK/q+oGr8438JAsjaAZalKjmezH+vzmbrsrm7ogr/LMcjh65ihIV/GqxC3OHiKiZpow2CTI/oCNk
4SmX9vf5sft/6RaSjBMD+lmKOqOJmtdV7zar5xrKm1mH83hQYypnVRKlOm4rbuNH4tbo27p3NFbt
4pI+EOapfLAxIq60ExV6fX7xKxEg4ey2ZUTAshtbACeQG5gGX0Oq0kinSJdfai+Sbo7pyymYo8ko
LNWkI+HnYEZqA55v8snnjdoQ74xp6On9hsBe0uARoI9LEi5l6ppZV5Bg2NcoAD+wvjgcTI3rzYzZ
DI/daUlafFZa5sk0Zg3mPIGpPKcOhETM24bTUKkFKR7EkxYCTHl6dTIeWiSgVuPptJr+HYax0vhU
OQ3W3gxjAvoAfFN97Y8tnqkxPjq/giflSkQrm9BpEB7etNPfnCSdd7LqrLbXU95MAIFcZQduh+sX
GbBmF3yBzRBemrKDeN+vgV59ErHi6x9olxGGhoCBV5PrCh4iqpIMWnWfPaoutXZN6PrZceHDGZbk
Gt5afT2P9440iD2JCXdkMSWscInnkWUzA9G9FFRiW6xOpi0XFZZNg299D8bWO/DBPXfwUh7ExnFY
R3Iv41lwbyWf9XJv+6hRmMLwjWoJT+t7KBw2GbZe4W+oZNC+mi2+SofbyCUId0PVho5LtAOcw2Wq
Bhf9hBtX8XYtYKjHlKtvczU/rh7WjYo6foC7k+F6MJ2uNjYs2YJbNMPjw/Z5JLlCSb4TcZ5IPhNr
fptUNFXUUMNVkPQKp2XXtbm1xFDbdDQ3f5ctbY32JinQZCEEhw6ZkJxufHqLbfcquU51Xsk0uAxd
E9cBUL3/x39WLNG+kYMhu7t0zmReyq2YgvFzGLxx1QBiiftRmoQCKq8bvR+jTC+oTRmIwViTbzUx
C4TjS0cy3Yh2ejjQ1Qk4VUTjnLXXMp4c02DExAZvF7UvlE8T1Iy6sVzkdSBq8YCfl8VIOkfjiluQ
dDu11Iipm333MVCYksROetra0B7z80dsK5opxTOoi/u3NLqSvlnOwEhB+vPRF9hrcej5hfNHZ+ax
ZU/O6NnJ1KCx1Xv/Ev9ZvagCWzR8srhRqEy3LNYZnz/p1/9AOchNgh0HB74uhYHVkH7pG9MNfxtY
0tbIwbxtdpt/axZzXqPl4xK8WagI2/AewZl6MNRjPkO2U+kQr6DdAwkpRTT1Vk409qLH1lXuetSn
yOLrGE1dTbaRbE93nS/rZEKRnIxoyjtfnYlsk/7muScNIE430Alzy25Ef16TvwtdM7YhBRwaRM54
bpSnwGipVzRJuWWyKsNKGApquo2mUePRal1SibFRya7J2EnDIMOPenEvwb7NcQpTHLvDk47ysC+6
wMD6IPbQTZl9Ul9KVqL2ymZc/mSXwHHUqclwDx8abQolL30TB0A0yoI+7Zon2olZvm2TUn5nlUaz
Xs/c8WOoacbI2ePlrpvgCE8h9LbCwCC6zs+ac9BXqsdSpW2SqMExL2aoEy5QNZxA5qI1YZuvVK5k
kLZLTpQN8/saNlKSQIDpF73MFb5rJxkf66dI1+aXihD8Nh4ULrzQZMr0pOyAQ+iaFLoeW/bUU7D0
RvslODYGpa20eYyYKqFW1ZN/85/erbgh/9MV8Mkv0aAG/9Bf9hcSZ64IOWsmzFzLYfysn6wbpuyl
tlwG2bRDupENnb/NisxuOdvbfgjBhL/LpMTGbs5uaz/DMI7ieIAWXO916l1JMQv83BrlipPENaYx
UL8HEuVQsN/Wwlbnqd9WxUHTX5Nboo8tc0YFTQASrocNuuKUlysKs80+GPVNZ69T9fAO5GMGvqyj
EeGnl47YzXxKSDZGoPpAP+Y/P2JVPQ/dDop+LCTgR+a7fzDpDQwWCBl0xHcvSG622Qo/49ilUgPM
nP1VLmTmCtliZdfpfku6qDDLKMA0Nf2rSslKMblvq0s1tJWI3WQTBSwwhG10JqOekQsNjJwG2ySX
Lu54vN0T4sSeR4eOHb48GIORxtA2T5X/k5PD0LsHoqcCwBFTN6uVSy3eV8pdpDsrmJoo0PH1tpgs
qQDaWDEVNWF6E9T2z5hTUu+7Krb5G/o7gvBQvQ3XFWhMmaIFW1y6H1mzE31bo9NANpAlfAAkr+we
vYFFTB5KT+JYQ67hREleLRTPK9gZAEG5S011Ubgh0NjQ2kekjQyBG5RnTMdebeJkkI25XvoeybGT
uGfnaKDRsY9xNWvv6th+M6Dm0sMQItG6tw8HSO9LJ8gvEsQAVoo7w4zW8KuoKP8Qv3wQKVGtS5gI
SdRyNbIro+9xA2MseKdlyPeSkanRj2pnXCQHu7JmK7jqn09Gpwkdx6BrFPgdWR0GJuh38hcnXBro
2HF8I/XoIfBCMNQcANoeOk5oV3iKnP9CeOzkiQu3thdTEp11Wj1YmjfvdPs8mTlIarSzbQ1PxfIT
w+vNIhCZpusLWemyCAv0bjcAlQTx+Uer9UZt41YWESwJHuRnLdJ3YeM+R17ib6vejsqwb63Gggbt
3wia4yoSr9v1wvk5QkgJ1qCqz79lsG0AkViLKatdNGYP49gLYXOaStEEQPzd/ma+zufxqcTpaJ+2
nIpfk8TnvFtRrEaPELsRL/HPSsp3ggp4Zw9QiUOifnVUJhNt2y/CV5zkW/E39cLArWSxrX2vUYNa
UdiZ0fq0QGj70Z6qIkQwOu1KAI1HPOXcuaCvU8m0HEg0Rb8wMGp6SEDD277fxx+fWMuiuARcBcZg
ODIAEfinox+di1C2ObxEe5kNypOWROJrYpNPIvbYCfwfKqb6vGReosKKRzxd4MYOrbVjkSjJN4lb
TaELXDUJj4vFBvK3LfMbQvQ3uIwEOVk4/E8bZz68CqEMiiww1r/u1i6x1OMBsaIqucD5zdpG/cLa
f8g+Wuna296845+TJvvtEFg8lhFITlPvWyitu0CUqhBppy4B3UqJ3pCzzsr3gf1ASxDVx0uryRzb
PLUkl3yAC2b1gm8w6643ijRAfaqmUNVeBqFUYfLdctb86VG6WobOiAbUrcTf+SG0qOc66f7GSZjh
9F5bpidrG5HAOB1aer8NGfLZpbELnrfOabOPBfTU/Jb7/K7fDSQQlZoGS2WmvRypdRFyK/ZFYGmF
M5+dVdtf/n8YuvM/fm51UNCitmMhfS6Rm+jgLjJLUrLy047CN9Kk8bsA3GIB1F9v8MNVBT+AFnZW
FP8fIkpEbSmWH8EUbnml1Xv8OMElSClqST9ltATdw5T1lG0lVgGeFUuhbKcAxHZMnSRmAh6fPDnO
PkfXKcUbc4ehGL5pb1p4xlL5081EqIxvq6SquVqRhSADsNVydysIjacBE24wM8ZzqtIFH/D1O4aH
pboUNtB42LU/vMST8sci5HtuYBLIoIzejoao7V5Dh71mZU8KQFtqtMVABKO8wa0xtkcGOoZUcavo
EwH0PyfBGHVzmrK3ka3eGC7VcWd2gtSAi74ZqXBaInbctGaZdL84AyGpIAqx+/lG/EGvt6sjos1o
8yZ/fiY/d+/tH3Ugi6ShLh9iLyoZymFIfInlpA895gTQA/m34UoYyQInDuIZtMOBAmazlHckEv6U
0X4/7s3ngcb2iXW5qPG9jNDmyJQoexKKBYkFJtaa618IIfRR0HBJg3d7ek+tIeerH/DQtVq4+VTi
VxodpMSX0WAbTmFDz3cfD6mfLQvJ6TvnX5uX5j4JZfmOprkNR/pSRhaiM4x3KfrRuFj8iYmqgZEc
jYvj0UBynuvo3ZreRScaCRa3Fu4agNgocI4VE+LKDj1EfOaEdjfrmIeMzJegaHYFw23jNNcGjjC9
tX3j6Hk3zqlGCm69hsfw6MqxvypXkUcurXF9q/fpYJmgkDzTq0ji0m6nFMBfEFPE10XtEfstIhv3
OsrB/tk6zCsWLEkaZ5T0Ra2Xezdfdm4JV0ZsbAwKL4L81+381rQsQ+lBK6RSlzvyHHx5vIPCFnci
geeDZF6E9slWKCPiljCMLGM438hp88GdoUMfoKp3Iaj6IvtiP7gwr8XgJQrsTFNz08joBr6Mfjcc
YMYfLUiyZ7K8Ogg/muAkQXhr+XAR99mqd63eq9PVAeeITffolLV4yt1mvvU7glHplspsShX6uxJr
E+FXbQL5sMINmNCSe0tch38ii2mJsFWY6+L2mPc5qaO8RQNBW3DDZxT/88JZ2/Yu2TpmH4qmS+Sk
0lIk1WJSmudKXM/YgS8OFoP6VZ2pUwYZHb169YtuJuTMlS6tPw3ReDxja/MRyfST6I9zTs3Fku30
EKt7nQ010knv9OnzCYx+kh6CjNmqzjVpRU1ItihP+Vb9naMRYohG3cgeCptvZ9YLFLQZ6LO3LQI6
YUOmq1mabq9P32liHkqek6gp1matBhhF4j2SGWJuOLsq1OMPWPXnwCeoGGEv/c/BxYg8TX7ku4Jg
Et+MXDr71noDDvz53krC+E/JvO/H2AuaLhlqAtEItoIv48yspKc30kY5r1fu7+g19hg6w9X0hv6i
EZBUiPFqoB5C627q6pY12SiTA5CYSTFrB0PhV3+n6/1U4fvGTi6joKXFujsop3vBHiaXyAzf0pT9
QxxrFZvgXo0vovKd0I8vRxrPupqJeB7P2Nze0JusEAaQqxKohHMiUHrUwrhk67wZm6NIm9NZ4d92
Shnj+Ud9xaWT9QlMQVSNbghccpy9npDsOBLgYN38awI3oE85urskKuoZNaMbLbSH0uug4a43e2XQ
4oSJnaewky9mmikoegZbHEyGSL8FNOm8b4yT0HWlaW31si0K3I9m8xdwC/bHLlaQiUMoPp8IFoGJ
GeW//UFdurwZTWFyO7ZEMrRuWNq7pKPUurWrv4uZg74jz6n2DDXv4TmUGi17cyGaXGO+v5IhYPS9
WLASCXYk1bNPgYPKOKDRlAWOltU8pI6NwLigXxKiUmRSYmQvEiMHdRAk0RX+AMi4mgjhK1yUo6gz
3S4TegnJuF1tC0fiNgImB3D+ijnuaddxa8Kl4Cjuqea7nGRmQyk5ibrNd/kbTLWrUOwmzlNqycQ0
s3oG3TWDVE0kZKkyHhb1nWZmydiIhxQaVMfU4yqAqvLPUGc9f/PtGL18UiZ4XqMLaCMDUNaEpu94
mB14gS7YSgXbf0kR8alOTie7qdv+pBbxTivrVoqBykXbp8jdCBRiXOhbcs9ZNsStw2t28q1MffRC
ZqA6nqAHfuM/4QpPwCJ2Uk43vupymJycW2ijvebpEhtbDxg08Q3H896QiVjct9vO2IxbKXGbLWQ7
aXp1AIqsfBkPGLC4AeoNHZ0ZmPaEaRW7GfAwe/dPPtFbWAFTpOjkkoEumAn0y6aozyRFaELEICUb
90emZifn5eDvHiM81bXo9r5oM03xWbdwp5bh9cbAxpiAfCl996IJuHUBEPVQ/2mz/J44BMx+DRL2
2keyMi/THFyRkmUDPBpsgofbCoBOdBeIveFyiMU9iasMB2iRxIQqlD2Uuii9b3w+wXQ/xeg7rkFo
qaYFwEcIj+BZQLFLBk2dMfSD3jLEWjID/FDlXs6vgvep3ek01GYxX09Hg3C6lHk8LZu0KwXMR5N6
Xn2IN+aMDrmXGO37MqSzCcBw9Dpf3Fuqn6mwC6SiS1YsDyr2fAX8Wcv3DvfbMYQrzKMCQgIozNwg
uhWXGXPrNnmnnt52em+A/3vfFlIXQHMIVNKPNFkuP8tE8klPjC6enL3ae1eYJl4GhmzCmsnbjuL1
XS2PxRD+rRSblvK5Id7dsJUmftdw7trul26S8oJLVpCySBI0QdG74sK9STN+YtSCiel+PDt4xqb6
J+OVFjT+mADbJzxwfdEZahcmRpn3sAbmOwv1OJB66mNr5dnUnCqGEunzY0Ug7UKdT+iqLLAKFsnu
onmM+fK+XaAIll6tIOiFFhIi0zhR0GvcEB/8xjH4RxHRFh7tZTyuw/fifmYm7xk7BjQGumWixJ8L
3KCJXMJR2CqGQpUdPR8770i1XMHDLHmifeYAa5FrKYhu9jDF4aaI0KUhqxg9Nv2WUinmXSl82+Rw
C/Hnq2gCgbh6x3HFkCKAbxVVJSVoJoFCmmEryp/m7sY0uhdR8L3xqmZBZUw1fS45ST2qvVtZUJtt
PGHphvt3b2xhPyaLvfHXIsMRMNiX18L8yj4fAalWZOBH17IofCx0sgpLJX/kA5POYppmi8cNU9wa
LklMMyKfQmsVBLmR1FbC2u64+skZ5gWqDFFvQJoo6czyYfBqivLLKrEjkyXmVb1nWXM9QdM4QmYN
Z5kZkto6yB00XCuPBbmD/uuJ6/va63Wx0oGq/LFvNpU8fq/LU4Wl+jCzIXOPjez+S7sxjLBHGC1u
RwraghlTbjVx7JawbAud15AB2K2cDwERePQozg5WcLZ4uVCfDqyqS1vVmkOvndUG+jrXtggOA2Lz
OHIPomuew73oRkkenQOtyPbv4+HKde32XLt1YcNmoOIlWMOmyQXh7K1VjQVNJEvn5KJfUXIwYfp5
MnRQkvWLSb9H5l/LxJQAG5yMhuJoVEbmXtELk0Uf8StKpCHu43cWbVP20usqW1D8aCLkxaq8DBe6
9U4FP7kqmSkX3VA1BMIgklpGDF0DUQPqGZDm6K2QOZOwnZ+09VZ/cfyycYFx9WnW952jRXDMi7r5
bImswFaS3JtbW03Tla4LsMIq4dmwKC56zNrPIYMdOzmBH6XPzfCPhLVtVLCgv6Rpr9oAttA/FvDs
08bJHGTJIyndpOvt/GyCUmrNvwxMK4kyer/2OHu9QfaClJqy5KyTRQQoZhITCKyr9AAmm0u2vQNe
EIVnpAD2QPXdmz7k9Gr1ef4ur59wNM3V4VkzQHo4CPCRXcYxUAWIYaIbrWwz/Xrr0unNBQq8o3wi
9sw9TZJEdHoKQJJ23+0gA0aml6MWAy9xkJPiJ9UzbTRAckE3/ziXiP53ZhbShJTmURqleb+XRiHa
O+JyQKtJWuqPZg1fIk6ia16dq3/lX7rjKYLwoC7FnBaf7sdjYGBvNH2FPunOO/DoOwIwca4sGe8x
qS4JJMDVYrkvXsyiApwbke7ufN7Ch5RyqqwH7MDYJZHmiMLwJhCLfH6luDpMruPXnR65wLf8a94a
P0DbPBYPMKTBBItsqHOmhzF3MRwTUxSJ7IWS3zyG0l/21thBjs8U42StQr4WaZ5wu/LSk1E7CMl3
KaaFBbuh6Zyh3nxTgXp6Usk3j/1rt3ucMVFIUrZOaVds0uT/Ofbqtr/diSzegZuFD7zpm2dhY4XQ
FIR30It2rovHc4KYChTq9s/7OcsHWVfo9++CbvGdCxK2DFZJ62VPNkRDw+EBbIfmbGoiAPIhgJjl
7SevS+un4NxP5xN+LlbZHj8gJVkJJAezKDIVDUh89wZcHldPBK798hsc7Oh0go98UiYgymJedWTW
PUlsRGjWVJeHKAqUrdhhkFwnUrxhys0BVax94+yEpvkVnkxoyKmgiwMGRLJZPckv6Bvyp4XKIGIj
OzkwojvVTWGttSlErVK0J3JTdcyeMAS+btkMEUl1ADm4/GnOxT71iIMdseY70TXvMMYp7juLTq/D
wYgxPzeCQJIFmsCfWPRKrgjvTpOZuGyhDSiW21VRykur3/JIPhhCaIYopumyg4Al7YUix5lFM3+x
npeeMpl6BlM6nUb9Mks9q5DgxAb4BnnlRpMELqy6EfPenyR0xBaU9EU+VDoLOakBIalU6f+pwyHF
4O89oKPLZ0NkC41tIJT6ReWFu3ng+uGRQl9lcx2UwhLiJCgwms5jevLMkDVQu79XdqBdrcY2wC/K
7cZK+eoM7EMBbaI5E5lKqmJHoqJvkTMYOGqTYtfzCaKuMGzLv8zRTuVT/FoFyE0P8EksOKBJ0noO
RlIALwVPaFKsrRZJMYy4ntXcYr723Nj2oCCk1LQbW1YKbmSzJBWt4rgDtaE0AhIvgVfHJXJGOnq+
IrwTUCjX2ZnaGAlKGPjTxVNn3X1aa9Sukm569CdfIujmeVM/25tUSvG5u3Oc3lCP3nCo4kfWhvix
k8wrBXgP/ga1SLaicSK9N5V8MaH/ngrT/jyO0MS/fU6u/669Si/daJj5dljyReDIsdWcHtGN0lYL
Wf74o2lopRKVwBAjFNOFfdIN0E1Je2mt+LQEhiwpIpseaoWnUtT6J2zzmE/XlcBJ8lPtASRkZjdG
41TdJULUwWAW65yRmr7lY5vgKnP/z8yFdqGzu4XBnUe3Zpg5cc2fvAHOwW6OYS6l0w++FUAZjLKe
yZiWuW2nwPQSYv/mqEGx0slhWTOhn/u9/WWpRcEOmyjPeeyYH6iEvazF/f8yJxJ7VYOoah00s9Qp
OCXYQG0Pn9tedj2C/XyqeDWbgf2BhaUMNl+OHJOTjddsgQJn0ArnEdVaXsxQ+oLElPaLczyACVzx
mPyYBfgxwnmbB4rXPm3kQ/4Og9HkcHUtcM7/9xLsR+gG4oSArOMVuMHRIzScrLGOFKa8R07pyAXy
gphvY0PXGIvj1ttudjGa/6NWCk89ZoXhRb15lJoz9WZXJN7sQzjdALgzDLK7sxzEo/utgT0KqcDl
OowHTw0T87KP/JmhdqUkYLRQe31U0ttvPg0GJt+na20Ojr5wH7Sq+iuF1O/5DuJLmEt332kA7kIk
q6KnF5bNjcOrglyzBVTJHgSDhd48NiJKGJIGpnrgYcL0RVCf1X1z2Wy0btweF/v7yD1zf1SrHZng
N8n6doGSgJlrOt3AgMCZHzBqdDFnBY7CqCH37gFgZ+4DFSv4tsjAdzL74gJSAOKDMqrEkbcHpNRw
vGV0TAym/mObBJgCNSbGb8RrF5dYsSVK0DS3hklli05ukHDOt/T2wkK4Uq5GVUH5BP/dAwfKXB99
BmBMu/7t0LBDVE4mdNCuPZnBvV4LDGnbEWHS9VCaFmgCE/lkSeHIvRM1jd7SZFGlw4PuJu7vK1HZ
q40+Akil9AoyBEfu3Qr4Nk37gAdbZYY8IBjT06ycOzjlVqW8zLmsPOGHQW+eLjpzbNKkwoXd74fP
Px35fcGpcBHkTXCib37ivnmbXsL7gImsU4IHGqqQdXRSc+AVtqKc5iXGxhybg7pH5+HelCjZJj/S
UkurZ1M+9g3zDjW6gFaY/zlJdE5THtAiSFJnmgQfk/+JdBvR79zRpERjaPnf0M4ut1BgMU+oypOx
NhYVz8cJeb1N7BqcNEBW9It/9DweWjxvjDxk1+QYPtlWEkZrMR6PmG4Oztz/hNYNraiBnHnbDtHp
4i5UM+42vuVUjZquOU86uZ/8WYz/WZb1+6M3wEM8hK7VDWdIxdY+jln2Ij62HcznNahkg4l483er
XK3ZK5eKWWtUrQEHcm4nRntRvQCR7zKkFmCJzEsXlb8SpcKlNvECkp1nmjU5Kox7i1fB6eMVGfbc
nJc+8PieoNXlMCzR2pUJzYJlR8Gh3NwmqKw0Hqeg7XNR/bIDG5TkwCcvcUsc3x/Z4YGZhTrEme+M
mXqkXstD95by4hcKFwtI/w3/ta3DSUOBFWtmUB9mY4EW7lhHbvW/4YIPl+3sZ6f/1Vf/RKLhfihB
MwfERAM/zH4jR/fwSd5jSsVYizOiOZ6Klfa1lhs6hyv9lMsCGKPEbWJvPZMHBDH9kRbnvlz73Rof
bHy+4S8M+bU78fQmiVDrn1scqxc1qmkw0TtPV9bqnYLBjBIe8JaglxybqkICvfhmRekYby4zpUw6
ZJhVVLi/OJIQ57eeJaPr45wSLoSHveYViDhY36mFKOPXUhkIiVmMpOBLPCQgQg+vRYu/3sBatEG9
UlxPDvpkJEBNsYmRZz/6e5DkWbaV+rinulyskExUxUhUCA+GUxB5PKQnNFhg0G0TMwYswYdTC22P
e8Vt+x92vIRBVmCSrbvzzBhGe1ORTYTMhzJi77/tLtIs8H9hf9R8M2a7FQNgae2/s818GSJdeSCL
c5Y445NQ4m3Od0Mme45fclxlbz/fclIVCZsIT5m5Dg0n5yYRGXbZq9rhXphwh36WCUakpg2ckaBA
OeA7LGFQq0sJdH1yZHotj1j+kSfKzE9vC8oXGuwEdkeaKPzBduXMBa8Oz0dU2J5I6XcS9kapaLQg
98lRwHCjAiqnLME+B9kKUISO6MU+SQRvLE/XYPXIrGZVQE0+MzrbqKYcP0mSUoo8A3ZCjAIS0wsm
dButI2o70ebqxyIz2V5If8ItfF7j2tPnNfux2RNxYiIuWUNXcyZCTm9HOdZh2KxmXag82HCxy4KD
3cOEWKAQv0TW2pHfxDpSrpj6zH0PEQ884MFsajx3Q8BIuB+rHZnFOmspWeNkZbTgwbhpFO+o64lD
EJpRqIy1M2nJck3hKi/DcMJDcAtheV2SJoFZJn3DrhWMOPyX4Xbpln7caV2olkF1iKL47W9dqOfl
YtHpICe8MY15GESg+nJgvcieDHoYJAq6K2jBhQImLskLbmkbP5VubKY7gnC1WL0Kfn8MHkUfS0CJ
ejOpda8BJLb2gvlqgcijDp4429Sp3DKh07LYcVg0nxKaefdoK6zEWW3PLDUA11nELaMDR03NKTne
TZPZbxFsQ7N4mduJ68GgqSiMwSOdzELUlrJrN4PWbIxVExSyOAsmSeiBdxtZriWLavw6iFFt3zL8
WQm3SnxyG6mXsVqbB8JWHqnXtxLl6vaMy/1MpzeXJ9yaOvePydVMorYkcD+1aTcbA5Yc+49qnclK
Iy1d1Hf5ExLlUvdF45MZccJ68MZvRKEdC1+IR2Pwmg5ADuDTTGqXhNcGtXvOL9hOBCJHoptEPvFL
AbP3m9FnXIpRLsZsqUzXQEoH5lGOgU5prTT5z416oL5KSJTIAFJVBrUTgOMnliv86FpkWuaR4Rw7
oECLh97cR1XoASEkdsOMD0bO2hq4lUeCTGE+cTpyuu38C9UUIemnJD0XZF15q/wFl1Md4HdzP0UZ
JImOc6WlLhpDUKIWnMEo3AWAw6gzsakK2Nk9KCicoDtaoqvRQ/iqpzQcBM5jGdpWnyInhbM+Jv7Q
wRYHUzqpY6U9XsrYG5fLTfFVI/j1aGFiftuMLUpzVaDc8ZPjSMawHgA+XaJtXLj9jjJ45q6OonUQ
i6hGiyyQ4gLl8dl209eTCc6ETBJaFJpZQfQi/qV/CezGGR+NYcqVCpUDrwizhUydUa5Af817HG+V
sm/S1Tb9YvZ7WRZfkk4IRbBMnBa2dvD8QkTgO59WUYMFMS6efhpL2/0HIDeiEuRA1MJP/ZWN3gI7
QAJyDKpgMLFzmzelgj22aKAc9O8fw9sm/+0oodX4+zG3e0soF8LjMgJhRccG3+gJmuaVpSAij3zA
oX+ay+WdW1B0iD5QY0XJeJBU791cRS+kIBymxeZMeuv9CEAG7iBeOWSymwAIHBO1x5sNWyvbrkd5
kdQRvqI+kuvEuySEJaLYSrcqsurpstd2t8NZyeQbnTfH6VLrgah2MEAB03DjIvu0OiMFXmk/kpnq
WFbRaqWvCE08/7+/PMw070BXl9mkEd1VpKF6ELOX3qu3wDgN792g0n7QK8YA2ktA6uonGQQVB+J/
iXo8VYKVHXxOpP5IU5pGHV0NzDvOe1OSanz6HqYTmM0XxCidyzlhwyknaUpIPZDzoZq9q5CyScDf
NA331EeQCerNer4jgkpqn9fYrFtTzwP1PLCK1f5+ShJAYmLYK4Ef1s/e1/CuzyL3MUo0Yf1RW2YN
Nz05JuPjU6QVGXbPXKhPt76ok+5S+h0EYlrHtO1AHZsCGEcvHxfl/5iFyopUY06HOhLNwc6Z4ccT
Jo+7ktS/XTfHPBUQ9gEpshiaBcAefrluxKdRN0RLzSkG7PHPHU8dR6NXThMxTt5uS7Q4td+7J4Tx
758I3dKJl3/U/NqYeWZbZseaE3GX4wTaMKiyFkye2IUVfqdA1tSe7Fqtdo11/iu2TaZ23rw1iQND
5OdBZmJTFvxlRUSC1EtR/FxqoUq5br+xJmBtQSAvx+Eg5VzgJjUahc/VmWMxbxR/USVhg22hGedz
yrYm+V8M4JEZR5/DIiARBXUuADKsqKnmeJzeQ0WUNJEYiLfwLPmpZ0i7fD37ZxHM9Wu62OrOcroT
Big9+KEV6/ZjH4e08Z+rOfi9yjrIy3NG/89PBqVFY+gUBR68276Vzvq8+O6TjPYM27An3ikmd7my
/ZY0Cl56vyiuVvchfOwnB3Xs0DqQrx1Wt89B/Xj7RDAZvUliuBE/Y/2ddmE9/HotXGUPg0RP1hY8
G+PKGiFKD7S7TY1T96cW133O7GBuWvkJbkLFpFLlvNzSx3tBRdZQN3mCQXg/3wsl4taTKyefxDpm
oR0GXA4i1lVKIOSaP8pYJbbdu+koyDbqp52nlWUSD94yNf7Ytn6RN1GvzR8fHf0sc1e+TQyfhf47
rfvyHZGIB6rCrdZc8GLwlmOl2PG3JOKQVafLb0fBkqZ0iQcISigI/OvrUrhvGooMjSKSq7DCvn0H
WCSy/PR3+c9hp4MZIwK5pAk4S0N6qdxOnhvDcmy94a1NkAGpAKf+ZGKRuTcgXMXa4jEPbPiN8h5A
MDdZg0+q8mWzVM4g3uVVwoXU0rMBXWdY6RTW9dCqhHj82P+NL7p6zcmWsTSNSkZARCiEtOixmCRR
0OPNjtzDnqfVqx42hiOsDuSX+cSWKCySzbx4tZEfsBsB9PgBQMLF4IbNgRwzh0l4WXZ2PG0OD+T6
hv9lN1nbtj1raCg2OisUJCBYgsoDL1+kJDmFkvVVVPDJRzH7/HtjloI2v1gkPoO+oC4rEYEhHeQM
r9pBLH3RJxDgwfR6ylBT7mRoHDVfA3K1lWWgCrMMCWfovK86brbLFiTz8iwD/mNb7WYb+nQjRjEn
XyzfJ3W+DcY5e7rLGdSFyK1ps5jvmFJ82WHDAioHv9MKF6Q7YLKTcE/+BdJkY5T6u50yHRWA/oyS
EoJ3ZBREOXLoN9QAtv1UVeV4eA7gCxxsH71iQ9FtEgHPRUiQtK6+sXznuALmCrJq4S0IqwJ6kto+
NEJGCN5bMJz7ppnOSXWrrveBiCvWn2qt+Hw73gB7Zw15FViTNES5x15ymx1lgkR2w24bY4ja9uLN
B5bj/fdZ8WA5RI25X3WRk0AC+YAFjb0VW3NdK26BErXIpu4ENhsA+XCcVvZarvhBSV/Mesmh9R4x
mB25+iFJk6ZD4Egemv6F1/Ed639NWEx5SVvma7lPAUeyz3DlAlALO9PRl1M6ixCxSTHkGBdrVGrL
HAiQGbXI2DM+L0ET9DutfpMWQW9s2wireCwRs+9eGvOTcKi0dmV8gbu7i2gVIXTc0Vep1fB/XQJV
MEB5FKX6SSbHs4HanrtlEuJ4EC41VKYvo9u5yOGjF9UDMEuW+567b8+21bgq4wFXlzWWA3/RPnNn
SnPcBgr1vOaApKp78mRQ6rBsizRXYsI505lAi45G7mGIzUBxFDDaGq8Ukx40UDofZHQOxqP4HZXz
R3vmdtU9xgKtxf/s9o8b2b5bALUEq6dSDA6XPk1toek7ytXc6h33kFDlJl/fdmmRIWAdgx+dS8Pb
0Ke/nz+pbwy/DqVF5dDY+0XET5iCXO8yLxgUhvX089fzCHTPlITS+UaQe+DgM+pnELJtzuPJvmZe
DZlEomt8wEvl5pjR0DufkUbCCurFLo5jQdk7QXN5+dzXALI3N4cQ09R6SB6iKYm0GH+jtXKLJHul
HmLJv69lTaV+JRGrrOe+SNFPoTkPYlotLDd3/QRurcBaqTxrqK/MYoFOGNd7e3MVSdGg0zMfI0Hm
YXyj0lUDv3H1okTGlR1eTtIgmbcUf5hcsUGAaP6r3DPpJJTDS5IQwgY0fO9t6Uki0iGRB3qPcAQq
TNN/3JPPXzVkTuyzLAiRqSrAEMmoAN2LR9k6zKpGsr+sQPFJ2ELtiYPO3H27pVuePESt4xS5HzoN
se1zkyLeCyBzcuPuzrkh8QjS7QByZtzKy4zQhUxbnaaVSIexQlKN0px3krvL7IJlgCDAmEWK1B1u
a9J/7DJYQLX86jqm5jkbeB8X2+XCAne6Hc3q0qGUqMTvpBWbwHCD65sMyuRaf9ZFuRUmM/HuRege
E+JN88dmPfxUzVHjVXbCf1UqwqWhrXvuKrnCdHnoTR0RRQFKoKMwi4E8FdHBQ6Bln6BJuYEj7zN3
sN8tRLbt0JJQtKQ7zqX35RkocYg2wlhW1utlAZrIVs0hhJgiwmdBJARoYTcvYmSL4ZPzCP6/xnXd
rX549mFPTCfUHNIQSNyokNpsiZ3ajD9XTxuCPpe+UqnwaIdHTkKqm9J3APXY4z4uNZbTzg8Fm59h
RlShoYTiMqYdLfMUDw+q037glOx5WrEKo2J0oLJlR0t0OT8eOrfIEexkS9lUx5uhFZfCH+bx6lrC
/KC5hG79KmCtfR+/nouWm82Et097tsyMxEdhJfrxmx218mpuCOLp5gWWPiyktrtLAtUyspNV7k20
BBShUDnoWbVbJehbx/UAsj4gN14jV7Uyo6/oxLu+UVoPVmpqTvSaKnKY0MoQZyxV1pMY0fAsNuIL
T6Bo9uC2Fpzpw2RK6MR4WnaXUnScXAGRUfZ1TZoGOuCLcbFuMCsj6eY3S7prEE3tM9zXIdt28Gfw
UVmyJEzWcPXfiqvBjsc86b4tOzN+OybmFNUUy9OFpIVJOind+AFTPQWX5NF4dCeYQUvy21oS6qwn
AgOgy9AfDZ+yv24MPVFLlH6pUssaK2ok0+4Ttce+mJN9nInF7Remhd8jsLwOhh4h7FANQtSDQ7GV
6SA1lttjEOh9L+tboZNvGi54LgB2dF9afsVt7XqvIfGJgmYDpf4NJ30bSh18e5TbIKSxjpTaeVXL
7TJMZeI4lFeDKfXbU3g3z62qHZ8u+1+CKy3Yay41hSnCA5pBE2spIkpJwRRBfZJw/t3Xw2RnKY2C
pKkAHuJ7mqv9ws380brfusxj153F4OSJA+gpxAfWanucFG+dTKYI+dospNwhoNAiVaABBWSgMVsj
glbdV2fw46iRi+Rn622gGDT4bWojQoKameExjTaTh0A1gnxZkq9uGIpTFSfvCRGhOB0MqIkMe+rm
VxPlo71VNDX6vXKgziPTlU/TSk3p/4r9AZvTGT3rfFqGrJh3Odb6VKI6h8dPJeCRcJA5X+jl7uKj
f6sTGko9zrd+PcDLu6GIo/YL0C6h4jbgUkbX45luqBGtlLImB+emtM6qO7hY1ZRPM+Sl/i4hxpRI
LvFFvsZ93cMvMzHtqtJKs38UuIlR/qgU2dTsrsIb3B/2lnIoMZiUvqo2l/FeIs1ygndBrvdwrfKL
SYFr3T1+nKE6fkVS5WCeu/Y+CuT2FeoCr2nYU7cREDa3H8VpXgJaK6+Fiz/i6HJ1PoFC0eELQupk
cCeWezLPW7B2Mu0BztCEWzY2kONaqZYGe36EF6q4iUrKwmXB51KPYajTZDqsFSUGmG0/Ofmi4YYD
buo9ZJTD83JajkrfpU7AjeqeT1w0jfKL1+N5aCpZzjNZqNjTIbQuop4ucocF7FqmNDOOVy5incNl
nlXAyd9HN0U2yzWMoTIDt2GkhVPT0gWPWJnwc3Nea/mWTpS/ASgSOSqV4S5YvmCDLsaYWFexEvBe
1Tw7Ta5vGpUzH5wmIazvBxtkflDfQL9HgfkYjo337sXY7mtEGdxvhawOr3jtt5HERupQ8Bs6YTJ+
ksydkR7ggvDzdhD+Ep8B3YCpwEqyxGmMZzVujRzfOiZdtl+lsTqDO0FnpZc/Y8UsE0mF5W7hsPPV
6XSb2+JLV1o4k2Fcu1tPU5TpTYSwsHEVK4zKlshEFr7p5D3h3C76KzhH1X0VD2tWVGaTBCR7v3CA
gRnrD0LntoTZRZJJm6dBnt6t8QcZrJ6ELsiy+lqpaoF1Mh/x9nhSKFuaClj9mufBoByiGEBq3djW
7ihw3dqTaTgGMhPtl+RK32I88aVaXUyYxvS4LyPWdmBSBk0EUAzn8K4Ug4iMdcB+hdvRBDny/B7C
dlnC6TgBzOKg0ckfpPmiiuTRflM6uFzslP7Xx+UT5e4WdymeCNE7RGjjXcXRtEBKfrLiAso/wxwo
XXAqy7cqIwuMpGV9EcnCqAB+Z/T+Q5AXBKgGIrCa48ZuIaJx2PI8nqmQ7VLn5yHyCE6/YTJpeZmS
i77uFJl9R7nni+wwRluIqq4wxnO0Xgd/DloIbjYjvtv/2y1Id69CbU8r6YCV5XvzWxsS/UjuJyOB
gcjccsq3+MgABW49qVuSAiXaCCqETG27E5Hj2EriP1jYEeZqNwOOlw4iICVfasqFj4+cBAsq+QD9
AUp2HzxZp6tWmeveDOg9NQG4X0aTip8EPbA5WJfEdny/zHKcZpO+hR7FyE/4w6belYoc324BTQSe
8KGyLNGtRCtcseS2vZxcRKj2M3GHWNrqIp1FX4qt566EbQCUcW1i8PitfzlqRKMT77c90v9ha7NV
y0nCbs3+pgdT2yz2iwjZTc1yjO3iYUPt4fr581ynTSI1BTpoZdDHWsW5ONoaP6LXyRDx1xF0hS2O
uEJB1ZV7R/HZ175v8p6kESiXOupi8iRLumahsJXlzTIS6HF6bsdI9OSluEEdOaLXQH7mw9p/mSVy
57gYegNNMVtNv3eNb4dK3VQfUwWLZbcRI5c6qZ6SLj73TaZcO5+0F+X+oay869JZJR6ljX4Cf5q8
fwowDfn17ayiCH/yTjdHA/CaWtQ7XctU2ZoRCqhqT/FUyQin8n8Bj1VrXpFHonoc37wFNoTnWzMy
+SfHH9fDzApULQ9aqPDHkokviMO+eGsehWte6pkOjPqdwN5aXqFJH3dhyChEp1t5jnvvCw+LDaxb
AKpIL0GFQUloD1ZTEaQuQa4CABaLSa+BIyzpvIFZcfjfGk+ppwWqO2uFiifjkjYX5C/F6oKEL80e
O31/EXJJdU3PkxlJVcIpNZWDtMtGMhfNNLWXjVtPkP0NCj3r3zkXhGCWS6KskJuD/IzQRyruXHXY
Vz5E2n5Mvag1CV0UNDa5XvuWtx+dvJkwGLH0D1m43Nl/4P9s0FiZGJiCHHZIXgbiSuvVglgZXmab
p9nq5n1zFfRiwJ01zKfhSoHETM5q0CqM1ljwWQEite6SzyockNlgelcmcDRaFgN3rnMwqkg9KsVp
L7BWuisEKuuDqMVTajkGwGH6n8fyqlNiYpZtU3K7zFDpqdQ//3E9xH2Ugd5VTkSJjU/hRjaUuw4S
9U3eER4EjP1NGZ7iD1+OBc+H6IUfyvjhpgT19I2Gp+t+V2QCs96otrnEgcL2tQEM0k+nTYyIuh/K
jiJ16kqm5UntBNey88BHAZuznIe5Ke4Spv2YVlIBhAcJz4nXff70j3pORb3It2n9xbkjwOh5G2+4
fKmZGCN12WrxEYCUeZZaeMgpC36nSZFDrity0qMpgEU75gNAOs5J4Qk3Z/qoey1EwzhEukiPsoi2
znmRA+tbabrE4S1+7cPu2WUCcW6XUX4Ifah8PY3+1VlZxm6/AVGafh+fCKfOxiW1sDg9SVENZXj9
W5jqUDNRr86dKvpUIfMvYUidyV+gvAhxaqhAk2ATq256LpIuRTOpLYjtxzQs6aJwvuv0DsH2wL/L
ptFDFjhy28ySHtxHOgfdZEANh+EhVe8iKgEZdtlOr6mHL/G8HPX+YNwEXuiKfALhj9W3nEvc77wX
2dOsYl8LSneSpln8WbxdN2Lxw638PWp79PedwvOTf5PJ+sfpDhu+rO4Eh4PKBl933KAy8bRClnII
WLjrrSU+T48beb+EGhofA/2VniiJHKB1fO3hnd1fifK2Pg3qOmYgYDAX18R51S2575gokJJQVFa6
oh0hwrXfb//YOlW5uNli40PrGKz8QEWzYpXIgCARZzPThNkvpTxcmBdbhLT1Bj1kOvHyEFxw+tBV
FV0Vh/WNhwE2ahtfB0YfUI3vyCKFayls+ja7CLkJvALlRtj7MvP1j6ego2yvFzRsK1k/pj5skA/N
BxCSZwWC+XgDb2wQMmqheNF01ya0tuINMC3GlneKsbotH4Nvtus8QYVPxUqBffvQc1H+6CI8qEqK
Pknt52TpYCbPC2h6FTo1rbBti8HMhjfgS14GOT02xL2asyZLpcjRJbSPv92iOE911XCAD53MWoNu
1C49Ah8X0mU1ayF/k54fwRTyNCJD0ij+RyPeZpPGMutj42NnNQ1wKtXbrH7Da7A61kMQHuLgQwgb
XS0CkA7/JyynXl9LPZgGyIUd75RmKldCyOJsSrz8IWNlBh5xdc7Bgq5Yeb38qoK2pImKqBs94U5c
V9kBqjMwJ3GnhO0q38kUmicZt8Z0Pbyt9Tl8/CFJtDdJITuY5IHP0n7AqmzBscluGbmo/A0v/pLP
PpC6oIhuc8h6yjV4EJGhnjWj02/aQ8w9Oe29lXYF8eBotBRz+jnfrrAnWcP8uhACvgJQQ1OIbEdi
g6EiHiIhnoPXaZLD/9dQrnF4OO26OrA3uTyYIzSSj+QNTwo1hrDvIZU45ISMpis3IyxpA6px8GJR
RoqSD+FAR3mCooKXM2FHG7iHgORCzkJRkoOu0CiFgyab7bz8VLyfRnGYd3XfPA4z5T2bvNNiKMzG
laY6tF3CTBJsp/DCVvG9aGB3ViB4FPoALcC943QzW2dt4bC/dcaaJCtW82ZMRLYNdnpLIBFq6iGR
yAqck++xOsRyh4+c6LHI2mA+vBATaLf2DEgmlVL6HP0OrlF79SvZC+iJth70ok68Ka4qABmecLz4
dYkIU2ObQsQVz1VNV44YEDk3hJDVN+b1cq+CIiYXoTgQxREPf42aBj+xXf/aGtEB5U5uFh5eYI1j
vPSExcTeHBPOD0uc3kf1/nfWOog4bpKtnNghfahxeSSKPxW0FC9zOQElgVfZuvmQXaprVl7PEw+2
vd7eVlLYV5k5NxJJvaln2YrGdENgFjYeFHu6DRNVCC4lYP6xUwlH1Rw0ig4v5HMQ9nEEs5s5mzXU
bDFKjXZadid5CJosthdhYgEGifWwpdgNAXaGzkm7qzEGet3IHyifaTTcQ3zrkeJ6BzXqkFf2bFmD
7yXBiROM3fQyshiIo0mkgHObAIOz7NEQVTNkwCRRxuc3U1Yt9RTfDyHJOS8LYBr536KSFxFhrDbD
EXCPPWP/jqQwjjtJE4JTH8ocg/RHaaJHw6fC6zMKUVJHENiwhKaiZzp8WPLEu/ujevRCna6c9jYw
MAUNYA+JBhYQs0EJR2sQGSJCKw7NBCMCmpmkAZnuVEp7EFvO/or2RoLuoYGGbQGehajko3GgkHKV
xhW49/X06fFhaYH8IhwixgQNLKVd3ZzYOk4Lh8ESIoMBo241wemevMyBvhMtuWB0ir5JAAiBC9n1
ySsZw4nqu+BeVlHXmGf5lpm+/KcVEE5/5MPizBQnQwJ8ZRUKWA+0YHKFOkcwydj+YuomY2us04BF
8lBwh9JcglbZivbecJQ3oErPI2pniCzQOP725Z71yIz8WcffsnHeuTTz7c7BveN+WAp+9r4YENCm
o78riu84poaaA6yLG16+GGFoTQg1ohytk3uNtvsCACPpG1Ss9xc4auBzhSbiAmZ61E/1PD3MOEhP
LJJ7hQyobMkEOF4B5ouo6p8hhiKbzzivBbABy1XT+DQztwLOw0l3tUvXe6TBxbGjeli8VsR+PBb7
fifQpLL0WF5lZs/cJ+sMnv6ztWp6W4zIM7ZuNQ7R+HJ1CzdHVyMj9A2XJL0CgeXvedXvmSy1fzlt
xn4s/ta+a3yGm5Q6EgWYqerpr4U1XBdhBb/zDTPjEI7dxpoE4Y1C2RMxiker0tSdm8gzK5/kv6dP
Z9GjetVW+4NBhLzQx39FknXUR4UJEJrUH8sKx4/+Th0YSBaxXyd74r3o34jXUOPLg3Xyvp5k75CO
fhi5WKyfFA9JaVgu+uzniuND66Ue66J6vAW4b1DeonZG+e/YrNLuaFNjT6iuo2imfFghuEPXSCNW
gIdVrR2rLV6EnRuKolCnInhifAkyiLqGQPNLMOARE+wwe+pT/0sp0TbtT+y/Xorc5SDA3GjLBebZ
KRK3a54lCGk+cqYodFUbrbO3Ou9jLLHugWksUE1X/L28RnJEkRvnAZ34OZisKVlWW4rpVOsxDCVq
AdzAQtmSVJzKtbt9mN7HdK5meJ2oFFByRwHxgXEt7Jd2lR4m3o0O47DpJkJYpNsDCaK30e6xrFt8
Zkmh9CNPYngfkhOghGA5yM1x6hlSZQHuDXkRCgBMp1pjFMvWn6JQb5oY5QFSHHJAGOL/MGNYY8Jo
ETJOxWGB/SHcw/F9taZg6+p+ZXBsuEld9EJDZEduT9ZJC2puaiX0rf82EawNILO9JqMcxuIfzS4i
KTZEPWzhGZfTam3dT59IKc2AlbRrj39QF3oSgrrZVI9KCAAe+p2YQInoJlor8yAtSc8oZHvD0rHu
ozMOhPTfj9/dlvLyZi24t/Ny2LeFApJiUceUF58JU9UkgVkxOMD1Ton2hXT9WXJcXQ2gD49oS/GX
U8F4XCAdDD2zBIjpnnxa2V+5p9jK8FsIH85bKgQjkIzxlcgUePmNoD8PDyi8zsdv6RYGhqSv6mgt
2rJFK9G8ey3yFFidUZxGN+JNl0U8hRnwoHWwMwvIGDEXw7+3NSH9u793sBjOvYJrQ+tTtOqv9Kdc
CcjggogUmTlY9t1fNK+Lkk1x2i4mM25gq+rZVzpO9lGkd/XR7YI27jr5KgZ/pwlrnMaJ0+BaNaKD
ceArs/bH6oWmBEDUzxF836gLGtqg13ia5B0DY69oTo5VVzzNoSP5TE4cJ6BpOQecF3rROxIo/sRu
+DhvxowigUKUFz2F2heRuuek80sDbOV33Ps4CLqLnTJ1WTW5tkSDYGQeNNzdqLO1LkpEslF0WCQq
jUQ6W7yZIwE46x5ogcSyZWtID3bpJG6z55OvucK0/Q9xNLmW8HPIGTv5WA1BWDkkVFdjNKf++Gpu
GK3NxectvzB+r0UrIr84QwnXbM6o1gGosZsoVQ1R5YG1Cr2HG65g8gZ0LiHlXxCZkjpbV9NeU5KI
V4b1/PcsUOY6WmW8r/dtRRF6pDiMFF6FPzHQ5kvJZcaexZJdnIF9pN+lAU2BHLafid/E+4YpjNvo
xcP9ByccBbFK0hTnCOX4LkzE4J8UPVP7N8UNTctSUx1sHUvZ4HJrCl8VLdROyy5svv0CzacbxxX+
7SmAxpt3Hf+ckQRAmySI95B3R2qgkX40fujxCgjB25D1blAmVadToFeSb5NFX/NL9/H5CGkyUHKd
P628U38baj1yQSEoBOqjqpmkfKtYH3SrOIw8HVdVjglaaZZSuGTuYt5BB3mmtaEyF2I/uqVwgoWh
71naUE7lkNN6UXhu3YzUREAAMBIlqZZwc/9uZg9NUNqjqdKYElLpLiiqL5ogS2rSe+Osos9DUhzU
L+KZiCT+J2v0q8ZO6LIuQRGvK0TNEpq487UmKQ3Gynfy2PVTYXLPRtlA0X+cG0wYaH4CEtEyHbXw
iLADYJ2nZQqnTu9DwzhM5TwfVG8qxATbAgHQDzUlUARguFhu4iNYYQaHKdmThKbHDO0ELTwOeqdZ
peHs8MVmqdb1UVI+597XLKQGLrYlBpwudVmE7iIsV2qMlmPLAXZEsSGVsug4w/Hdktj+3zVHRaAP
lIYUVLILLF538Oq0dQEVrWYLHtPZACtoGGEm+DjXacJrEanp0QZNPul6Mh2pmFEuKbXBst4TJguw
3KPO44ay6AegVZOtYuNlXEfj66NhnOoO9xiZK0SqmEBXebtrHyAd2KxBc4onW4IVd9Uo6p/IP5Qo
FH/+dvzUdoDQ+WxvL+0jXcV1pegvUlAbHkIawZOBQJJTUHfqLb8bgeuU5aEppSlDwIZmebYZG51A
QBfYW+GPZ5/qYfnURT8+/2IKLf4L4v/fgaQJCyv0h97nSt+6QspNgki2Dw2PwR7g8aSuZ9wMJxNz
nCWgoLtedGSTRFAfFxGcmWGucZhiX0yaIGlOSVhHeQF88V56oqziZEJ57SRXPjKCTUgP5f2AD1VL
DHlfFLlNldMFT5irapJoUvY4V98qHnTnBAtbEWEU5Cqxs8iRalAH+kJsRN9dtS6yvTJQuezU6Q2/
aQJhATNOBqfHeaORW8kCjDdNWDy+TZvaXMxDTeTLLEi7XHlyU0+lAiBDvRouK92HFVntGGGCNL01
fi5KPtzVDVkfyXxQ8qD7z3ylwXZoqgfW66i5DZ0IVER0JPcolRXDpwpgskN5+TvgFNzmIzY0uZBS
jMhGwoU0V952UPvFre2yjA1C5q7u5GCGlaiMzXuuSoSzNC3iX1AjP+FtKyTsRDnwNVDKCeJH1Oa7
TZtOe7ab5cmODRlUnLu7yi7ELwH6LiXtkl0zRKuYxmKy35ts/e1Lckj25Imr0dBTBgopzquRWMyO
Umg+ajjFlpaX1TkShP7KdasgSVmCNGIlUfzfwR3Zt+xrkrDC/CafAnt4F/tZFYDyWoEGW8wPJCr7
xS4X3CMbRl88l/Mepn67rlESiAyJ53RLTsSTtdbBPH+SixfZjhtk48TbQBo6oGTu4sT6qRuDvVOD
dy4V7IopYt+uKTJ7fXPKXTJFTHCJz2IpYgB0FC1qCj0lz8GuOBj8yY2cTgRpSkMwjS6bwMPr3o0t
+6KBOum4BAeNKumYoqdhKK0UxZTAhY547zckT3enZqHLJf2bhm876ilO+iMuZqa6zH406z7IOeTn
zGKOOBDPE/iCqyhdd1tKQPfCcnz2awrEqJlU8QriVgN7uluoSNswE4VsgitBXFsGtIhUYtH0DCFe
V+cmxHmH5VaCwxYuGgdG5P2Dv3b4n0KMYTTm5jL9O0mitqSFyYcyyndbqPOfmWYdtbFhChQoXX6U
tPq8IlYkM7Z6wKAhQRGRxYG7oSiEifUehNB7ZpAlSsWJHSZnSzd4JuQWnK/CPyio50RPnVP7GL5w
oG9al/eJMeAkaoM5WpmH3TB261drsI1YzXfRE3GJtJhH4pWrVLQwiZMKJFmYF7o+ybQuA9FV1Bbp
rGxEnX3uflr41j07GkpX5TQhNjnr9JUGISISUOlnuYjZNKxv0biOEuO4nyTXDOI4oKlUkPdu81Ud
2R8WQA8OQK4Loaz7dYpbG+23GUUiVF3e4vy58qYXmG/vzS3FCRsMxR05QZ28La5PZpiEwikHf+rQ
P8EXGMnL+bD0Eow++hjZ9VdF0q/dMfuuXhObrxGT6lYZ5fmY1a5w+EklqAOHBZAaKvhkE86aTUJP
9V9A6phgkvUH2mdeaF5TRFbdJhJUfre+en+SaebmwjVAF00JRL/i/CjS+AOQQaZnva7I7NSs4Cte
sYnb4jbpWUuUgRRVVI3B2kPssjTT6xkYp2+4q/I5RBc+lvdHeNDQvSGISV4MK51elJxekA5f/Dpf
eP49PNpzRLygLLTxpaV27bldFZvj4JY+OBKF+kDYwcniIU/Az5gECGI2t5aBhIipG3peReCVl1y2
yWeWzW0xgA3NUemmEvebDERAwR42Xwwe2g3YPguTbzXxjcMZKqASFteatAsAwRYj9mRwg43vh2DM
FMUaI/NS5SgcOwZHTDvGOtyylDEsQx9q4YZDL4durdH/kWn6V/OpTuy0XfxiNbOBcKpjMvQfJ29B
Sob2Js/djFdui81Ao6nmpjTiC3sLkLxUmlrI3EX+lRk8ezdPRGJy9+/6eTkrIzBSdQgpY3auZjK9
2XnDMj/6tuUmGpYvWUyfaMTWGGSCrh4pploHj0xJu3htidb5kSIV6+Z93gbd+Mp5e3VcV7eeMvZO
2hlZCKPmH2owx3f9e+IXNKMeAD9F18F8sE2rwoewGXdlkhLTlc+DKLTbEZfKb2/1vzQ2ApSvYX6s
+r4LMIvRGG6455DYwd42r54q1lvsydCUlGkGw9BZAuSkZlsu/7hbgAIsW04rLxVsSBG9m2t5Ydtr
AAlIfyQfR7ocw1iPLc5hrMolmzgxqR5owvdTMs3dNURdfXFDue6uhgakoL+oM+RGkhxaskg8GZVq
dHWFy58ivdFk8TIr5jyhesxfSrURU5hYBFmMZF+8/cs9eQWgqkJR7qhhSasGAvZO+v00zKdHi6G7
IyiSX4dL8CmmlJW+9YbjEcadwzhqjjh5cRneF26dL8TL5ENqjF+6JbLAIVKorlNFEp7QoC9DIguL
i7yLIc+AM5J0A9mRGlzWv7X7LyG0ZPC81kBWXg8Lj28HFEnB+KO+83VYUTVqEBAuZq0HVvEG0Fdf
vO38ziUUVtzuX4cYZtetF8LGUlMT64+6vj85xKGkaE5KMWCBmBzH4dh6Ry7QD4GG9mcjVGpeCS7k
2B86hhw0+uqgNNQQ3KVRDmbfKuKUH0Pq75GrYUihTxlIwLUQv/tNEV7ThgthJMyKcxJN3PDIPhtI
XivrQsK/RMVHYMG86N9CZX9us+rqYq3fXasSzfJYRFI+upTcuGPumBi2UEoT7f71zD5WT1rEhjcg
JliBYfOq18HCzGNPQQbsyz4a1sEpyWNxt+nQSZNVzUcJGcaE7a2sYa+MCA4+jiznJFMj1Q9vnlmC
0hGKBotzvlbV9VnSYeWfZZrqgP+bY1DU84ArG6s5FC4Qo+8Q9L53AsLtkuyOvtBE4izUYwyg5uny
Q2u5Q5OQo8IzgfnOM/7rvXXZQnZ9GNIfBf2GZARTIZ03Ry6lH/unuzILO5VIb3qux8iCqs1atsIe
Vmo1GW5+bxCB6tkQ1uGJbfzPyN4zLPiW/BgFkkolopMAV/z7xxKA/8ebgBs3VNQS0xGV8XsVxUUF
PXahdUSS3p2PXrbv7ljw7BNVQ9BOv1MtuMqzL0tXl2wfLv2s5ZFMpR00Qhq7fmmg/e2udDP5yxJx
aRe2BJDvUWJaq5iznj4GRX+Nhs8XdOsvSPCcgbMF/v5Ui+PePKfkFQndW1ij7gq0QW2zZZaWa9Yj
zaPtNhXjbUjD0YnGtvIfi51cy2QkC5tsgQA5An35VOQW92QVYsUC3LTjvRLVgBOOhIsIyAwojCDA
ifiB/7u55OKsQeb0xagxdMj1VGjuFYK7LAhmuDMFfLOHHSfu4iqICyv6NEtvZFNr1b7/9H7nRkWe
Yk/THPp04FqXN6v+0t4ZC/wylqnOBBjU1Bn4ruOVxgAUagTTMRSJ4K5n52KDfuWq95HC1wPx7o6i
ppe3mIGkEsHONh3/OHwaMNEUHqnbu0xcDESplL7CAP6FEQqphchVM7CCBKjRRMoDZnQsaJXi+/Vb
Eazv8IKZAQYWnGVegpq39Re6AebifccQsOYOMk9Zn/VIsAcWC9l09iwkLwDTwIRfkOYic77rM7kz
Bgq7tvAE2ciw/1xkCmkRcZGW0fhlLjC+RF50o7SwniXV1ReiHtY9StJPbyjqloNEQWErF1pHZA8/
hWX8tRK4FPlWGwrnT+nfKsZ5AWR29L89gBM866wx9KuQSAA3Dx6i4kTDlRr+yfFt20dL0BuC6F6H
3sEwPy3If7fjtgE7jW7riUuAG4VfocOS+4uKp9yDySP8te+K+mOnfgmD9oCCucv3MgkxnUawHm3e
9JoKVv9gKzZEuHlCf0fkl/bwgz/vvLhG31nDY3Lx3tUZpXA4r3UndIJC8IRbO2+vHIeRji3c/wcH
L/dZkgIl6s2mi+ztUzOAUnE8hGlDvVgiTVdxM2K6fSG54u3jGbE9QBhCbHaEY6EjHMP51+mvb7nS
SUxQJtgXH3sW0sx/6mK51OfJ+YutJIDM+4BQcjN655NnYydeJOk9SbJ3MpaYE/xJL7wto/PA3sol
GD+UYuGuXdD5a/AQd4tLWq0YSHCXAhP1a4zFzIrRFN0maKu3MkopnZqOgHY3y3fUPZifZNAsZO1E
+Kp5KiDlUDwmPZXw5MWZTVhBbnIWTUAmX0IE61z/ZaaDnCjMuuLZFKJOq0W8UJtcbjQ15b4IM2q8
XOzJpTRdAero5jzI0JhUoi/c8OQIsZx5OZgbCvDW8k3BYnQbvVzSoW6k6yOjl5Y8LKapsuHElWO4
qHMPNQtOqbfGEq6VMbYFI76gsOJZc/uLW/TU9BHoEospN588/Vblk4kd5JV51ahP0HBiL+Z20piX
Ujmreedfpl6x7WDgsAi5F1yi2qtp+r4QdH23jOtcWySdodCMmAuCbcyidrkQSHYOSFKx25oYB3eS
tcDCQqbDdWf7p4om7GFhY7Tj2c4lh7Pa+Vk1JTBygOEd4WlFDRNa9NrHy9MPepggFCCbvcqPVcou
i63MUQ69/PI2KaIjuHhIDDeSowWq/ekRrBQAMD9N7oTCbaE65pgg/Unpnz0ZbxJ/+4cXjqJMVpV6
vgIQOaH8tg09aSPSVJgSQ8Vlo8fOhfzxj3mH6UE3rRXV26o5e6f85T6ELP2/K16AiMHbw/E1q/Qq
Qe/K/mbgZxZ0gfXdr/40dtQtmcjUvGwpZ5GMmHlsoC74wA2RN6YJBe8kB1JtqFgcvcn2AEAlpxhK
x3NR7ns/L8Wg7CmfQmRISOBetHImg1YlFk/2otIF+fAgPga44KqMS/LeeO0SJ/w05KF0wtKITOkW
u0ZtR6j13zoQKcSme3LYfJhsmQNF2u+1qf5WwW8m6DPFI8u2BGgpz3ikGsO3Co/D3oiaWmjU80GZ
/x3prSrai0lpnKWEs/RnaHgxSSRFW0q3DY0Z9IwI9+1WwT+tpD+6WW1QZlOkF18kk0ShiTVpx8LN
DDtt0mwiqqPGAFxZgtwuK+Twjj6Z7+pidU4LG5AGGgXkN0fsS+ZfcUr25cbup53l7Wihh7xsSieV
kzGFeYUk5yxuM7y0PFMExBmKRbGBh8KLhKtlNXi0EtiB6kPzMtNL/s5sICW4pMUVTXUMVa0qzqml
6JJHVkue9me0LjCF+KIqAbY1PaExXni8dGTyaPn3acSIKmYoPExQ7lEhv0HeLCymFrGkAlmc7Ya5
WqK2k91a3uWY+qfFJPuVqH8WhPFoo9Tw/Gqqkqzz8GlsfO8fjo8+TgCExeYVXWZunwGrKBYJ2wAv
pm9mfOwTBpZKWOnbb6yf8OQKNwzctOP3SwI1twj71vxTvYEcmuC9nyLvlcwyxpOUHRQGZ8BTgsfs
dfCLp6ijqWpiS2nFqkSngBj2OijdB+oMul09Yntydb63/rffDWjCq0h4ZVBEp0j5r7Vv8H40i6Eg
bbdQpveRhUJ65KcTX3nIEk2JxRI10Zytyji0RPb/0ncQIINRZOsseCWDuSuZoEvnI27sVJNM0gYE
hPaaGQFKPm+2h0ChntmPvy0bHv4qlKweRVWfm6k6q2bbXN4BpDvLvttEB2G4V7WDOnEVDmLGgshH
9zqsvVH0K4VEdBPWrA1jcr9vjRc70uPKLIaEjm0SOB7g8dwCl2vUf4Mfpwg6v5nc9qJlfAxWMDq4
9bBJt7lKSnbqZJiY2QWTR1IKu1jWyEA5EC03+MMch8V6hj94Hjb7pK9YMAyerqzK2iEGYXnKdKQ7
hYLlard1TTa2X5tRfD5ajFaYdVbIeAZoAPhL4muFDEkLadkUIla8bpg2ca/3JrJWfC3g4O3zb7pZ
HgQffkIaQH90ByYq+Jd8BDDgZtQ62LlgoOr6yMIx/o10gpdw7w38cFcDA73XmSTJAcJ2nzZPYRAR
3Skdg6QCoE499n/URui+TjygR8vzXjfXprE4k2lvpZdWbDVR5Dt1xCZZzFKHpTq4Xkj0rTqHnBpy
fi32wgOBDzpxFii3Bz1BuYDQgdhNTCeF2o+XkmZIiD7GgyjZsRmF0Z5Q0x/L03LnrALxcRA7vou+
MAbDI4rg19EBK7pcelEpuD5BnUc2vqJuGuSitVVaBMCIbS/MvEcYU0MuFZfaRCCM9wipv00ZQ5Yg
PgAvn4KL39+rky6ufmjpV5SMxstaMIau3uX0ybEJ605G+S5XqatWnbfq1kRv18ElJaaeozhfw+Lc
wDnrkv4gu13qGSb/bZXG8FE5J9t+OmWZkx+VumJ2Yjj6uOzSEs0YRWaqIOvKq2+Iu6BnjwodxkCV
h7xH5qe47oQcCo+apLJW/vKyREr9jaS0f/UJO+e51aXiiHyFLzZBfF2pkUDaTcGtbTNLp8xsedTG
/NAUrfq8Hzv6LBMIzhdOQzJuj2qu9dPHLsmVZ3bFFqImUV9x1PsBqhjNqL/lX/eNVhxFd7w67j4x
38XLDY8Dqh1cfzFHiaEtC+Dx2KoYrC6+WAOLsh+2TOkI8m2kM8KUwwtN5tS1q6/VPbR2KlEpJJsy
4JMD8MZJdDx0v4q/sxSPpePUq93pkqh7fbYnJd+P/txhDvc0ipU1UIg8/WqzfndEu9aubYKKNId7
PcID+MvSfs8FH642N5okvPd9rs3xSb6b9ayQ1YmAc64nDmi1WGb+K1pT0+zr6VJyTa872syOUNIw
cEl4mFYSOw8dOlqL7cqhBhJ3Uz+5SN+gKhyaCL42VoXc+REgn73oMFTkq9i5/XSai/TBVUrKU78M
N4UbKqecdUjrYzXpJFcskl03UB0dPnuZZ5QAUq6csdkg00HB86vvbfwo4dJ7igQ/0SRErMm9EdCm
D8VdIXgQQIMTbQztxsRrVuIM9yWrFN5MkbpATE+SO6HQyF/gmhu8wuupx+Lv6aUErwytpWDHET3k
HX7QRNRF5NIq4VgwALetb9MWtJ0mL0Q7lztdnT1s+92LyTo8olt4jm0F+QtptcEF6OsgNzK+PKmH
0AZzndqnz+yekHsHdwU3KFdjoPV+7vj4MDZ0vBdDdfThWX+h77eK2S2os9VHSAvB3fweHRpBSR7o
ndk7a5kqT8Yd+qxUzU1c4YcY3fLG5+JynMQpuIcRTtJLU5SxN/JWXm+EX4fh9c7grTXRDwaeFgf2
BfxJswq8mHYfzzhvDOg4nLHokX53B7dMQDMfPLw4MX+6RVorZ5UyzRSJ4fLKvePwxSG6yWodS+yf
oqBL6u0JB+o0mkZAgNZozL+lolVSJOGc9wH44OMGqwnQ7yI75G423J20vQ9ksDtsf/I+Yv6phTsq
FLWvisDE/WeLyuXGn5N90M0kzXAFGAYfv72NccC/vES7oNjEwuGBV/1GkkiquvmliN2w0JOec7qR
4OleNGlbKOObxzZbcWYTb7J6VnG5+iGRodzCu6sUq7N+rjfHRFHkqiiLMmGo+0bev16HeTqS2Mih
PYs8FLP6GztVBhcqxlkY7dndsc0rwkAEEyUa184k8W5gUdKbmxnKIa10gd4yQ1m/7UfdmOJexJYp
pUUa0hNBs9HV9wh2Dak7QqIScOveg7vBJITHF+eVFSYfPOeDLn7GLFLKhVJYu08lrO+5Unbyqwg5
G7dKoJyfp9ipI9/d8MORyzVaA7+HtWf2FxiNakim1tLhVq/Q0BKfECdPUdAZ6QGRm8is5AGMvLvD
Y4AhlBS5UjmrTi3S2sTcsN33rCYcatmtpn9NljW/+qKg42UeNimToP3jtPaK0IgqYpnkRUSnhfCl
RG0eZE8BmY7I/55KAVyqBqoiC02wMY5pieMJ4Ey5t8enquoGC8HeaJpJOviwVRBfTHUBHYK0gyOq
qfgoe8Elr5xQlKzeQd6QReTlNssDN1EgScvFPo13pKNlOLv2h+hWIU9ClfDBKIMSo7aBpVckt+5/
PQQUOR9h8XdzjtwM4NK8GzX7TOMd7kDuBaa8KhoZBP+57kVfG56X121fCJhKFx3AKBD0trcD3N+4
M36Z7NRi5WR6hJ+benLHFRNGeE7Z0F77Kj2iBfip/oxmNoeGJszoht0P8ZetelcqetVUAVoAhgvj
RlU6svS7EGm2WOy6djQZQ2fPZW3n95/q8YUjFLJj8cnbi5lnrUejL6Lcj4MeARecmPLxqFxa62mC
ChpLRrv6ZWJm3DL8JAGKTh00CZ9Qph7uBfbEAq63zXst15Ds3Q+1Qn6dt59y90EscY/DCVLEZpjB
0g2MLm/cypxcuYyOl9jjHZPRhNtr4sHQ5SJV6KlD1kR329WIQ+nmNScLkPBW+kJ4eAOpDJBKI11B
88ByUJ42JkBYBWUV+wYXUqJhGbkceATf9nLKfnPdsTmHon8OjQfcSgizcLKVhbfmL7Qz9bbnZaod
6HHk1RSzL7A7RbUiG8WYZWBR1Afjve7pAxhkSQ38M1R6n2laCvvsIGvw6y+dLr+uhEFub62QN7V6
H6NMjkC6VnCCfkaaik+N4EQTSH76oZJtlgCdhRXkBfx3Qpz/AEIC5pVCsF/o0YEKZpPCMrMrEUQJ
i9CYJ2U4dYVvi/Ds+QDNeuTijuthRHzCbkyjRwDx1PE/FmxUyoqTGhzfFyMA2xHOPGydTlnl20mR
DB09WdMgaXOMNzuMLCIcfAZg+4IaI7MR56PFqKMmPlGzZQMXXlO5nq8Wz3cej8yB60c+b4QNFI1L
SaRwyhu2kcu3b8Y0+QUj1/y6D8qeYX50vZmVRynF7zKGcmsCnXZA9N+eBmDoIcdimIwb9KfOmHbk
P0aux1ZMcNRwwhigGZTd1Uh2TTsowLQcQfxTqhgEW5b8hhx2qBhpWaET2GV0AHzKgGS6UBgZ6v1G
EQdMNvQbK2BzsiStoYXIA5IeH17CzGS7lStP99D4y5MD9fv38ea/CRaJXOQ+vfvel/S1Hy9N8Id8
fmHkZ8R4flauMa7vlfrSVUP1qilPKvgBX6AD96reguMAYuT8kLEFE3UTwXCXu/8MRlk251iFLs+w
TEeZgmma8J29xYTVwohzkUzZBpoDl1lFVR0xB0LNg69Q0qIoJgd88YsTglxYUo98Oow4TfnYaGMu
7vXtsi54pxwwfvN347ld55BA6FdVNSMp1g3XYC2feh2bV3B3xxlS292r1dbQjyGk5HwohNOkoTqH
Wz2ieDtXtUJ22wHEzelGh6+1yTyblAYifpE1wG8BOThpxmnoLveYwUoDwPhA6UOvbCUo4Wb8nKD6
5s93uJ1dBoLWP4uFcOH6EYOhOohbC2aUTtUr3TmbHMq9K41J1Mad+BfQmdk/90NBeE4v0n/D4h2f
iya/IbF1Rn27WzL1zLjoy9MbYMBfhIdRCHTs5rG4cDcidv+6dPumdr6vKnMo8tnA3RltFSZDK+c/
GXcQ4F5OAIpYUoYE8gWlagboV+3NGS1wM2OoQ1Di7WMzdUaIghTsQZrpweJR8vD7IXcMtvkgIMxn
J/NMy2jufk7P6d6bxGnmxlX213oe3GIefHmhRFpZBQMDcPU9tz/m2qNjsc1cyaocMbZfbBP6sXGM
u5h/89No7gWll2WkLla0MoUFCYuf28fLGv5TSzhaWMGD2kmsZ0Ee2vxq/KcwbafuRe44KascnWdK
0enfGS/rR7pXgrTydDjltHbRErdZktsbM5g1N7a4A6PrBnDwJ8uKDgifa5qTeIPKjFSM9i1c8YAF
K+btUimas12HTQ1IOg9OJrqe4V6Pq+p3kc97ScEx6gtQjtveCOsPyKSRQDomEDNSpGxNnJbZm3zX
nJcPScsIKG5FCft9MDlhJCHVmpNK+lq4q9fGINgSU60R9EB14ss6e7t8tu5CU2hf7tM7+0dY987t
Na7rrWcGNw9xATpXZkv+vT3pWCO4p9kyLf5+kvpMRuNrJ672XMU/YSel53meOW3eTDYTZwFkJrML
0ry3Qnu6xXDmJniu1b+E6ddbY4KIUtKIgvBtj+EwXsdLygat0ivxHWvTIS1dl2BXAWj0eLdCZFVA
HHewyMe8EcO3rf0/6bYgE6mWWhxy9gRfNgeEYaNuOBrVUq+F8LL1b4gWQ37SFGhqFaMTlXMzz8Q+
/3Lzs9hdTmEsG32FylFJFOsELuE2C6FIw9Gg0+EOi7it5/tTuR0YXc9xnoHKPJohxprzoZBGJJWi
9gM7zOuG6K2A5Fb5lA7rwjINglHVeWrpXaO4SoZffrDK1ItpijvTa79vuZPDRVPX3UX2qAIle40y
HE0XUE4t8PFmN+K5Ug1tfvGHVTDW8wjuwCm9MdW474N4oEykulWviRse4Rrr5PbckuXH4yNQfpaF
V+NuzphQAJml17R4pbfxsG5mc3+QesgShTPi0WzDR96Kne4MR4wdVkVCUmDxnhBVqBqINKQ5FRMF
XZk0eKsww84nz139TTsEv917h6c/jlGPUuzJimmYTzTqJ0kszNCjxu3rOGZP/74FWgeAgUERuY8y
gxvwR9Ul6GA8Y3iOhOaWv8XEDa6YF1VZRAlSK/ux2pUx95JozL7GYNH6uoh8Fr3UdsEEpSN2+Sa8
J7m34h8xU5+YlO9w1tGjYA6TD/IbAGB7uAHiv5924rGe/j5rxskAT8GFDzCeAnum+pfScKW1Ylda
aTaXRK+B5mcjFl0hDTbWYpSCn37I2fB1B0exhrWsNkVLRnM2Kz6qiFK7WXx0tvGZpI5+5s+AMTUS
8ZeeS7X9xQy7XJyGuO+OZ41Nf0XYbeHsg7Tn6omKRxZWa99M1NEy8KsBf63zTWd6+844YWPCjexw
aoskqpRHF6cqB2Suw7yeYqBHxC51CrFsCx3WmNZ2FhXcjK+LEiWxzpbGb0m1Gwkt4YWDK5P873Uj
BOlhowwg8vO/jcHoPOGU14Qe9cMgckFTlVYmnB5T+bQnMZGsUH8gXf8M9X+craLmoWhPFVHQkiOS
3RS2To15E/VrjhLxKEqo2fhGfFXsS9ILpXQxFU7Xe45q+x7IdZgH6C2h+ILjRlnrlSrzKnXjPlB+
Ryne6LIfeJ5mPR7EWo6Q4ddwpPfwNbDAJ7Bi83uOdR1/6nyvkdIM3p6R+asct8nfkZ16Djo5vU+E
CiQDxZMupzEtjf+czelAvSrNGIXYoySZ9JmKTnVRyLT8zBu2xhIIVLCAXUQgsXPGHEx7U9TeEMI6
J4dXK0YCYbpux1OS2r3R9lIiuMaG53QJhWQYdVfoPER1Pj1Vt+1V5P4Q+Z7tUSAU3URp/ITIpwt7
CUr4ZUyPmUrNpsw1N2nDE9puE1LFARMWDpFVej77yziKr112+2MPJvyohGEIaxzoi09m0dZGx9Lo
Zoo6NxenUWTUZMUAl+Ib8icGDo7615NpQ3i1xXxVwewvT4hNQNmh8w6PzG3T1xtpaNxXXFRRZRkA
Yz8Nwa8QtLxIBoeG6w5qq7w3+cOQEenLXrZy9E1kvFybH+NQCyo2QBGCzoKbCUCqmiSCNxZ5dIkt
bCTK2aIex6PBLCOEXU4196cY5vWEqr+7+XhK/sXBPbVuZBYg5xAzH14iZFvmzfGDL7ZkUkb1cxzn
+ImjNM+vseCgzahN4drsNhNsidVvB6yxIHWRhM5FbkxjgqDLa9ceNRxq5jTbaKiPNSZquM6HuOLC
DLc2gXQw8TxczoWOAwl5+DEooOZxxU7UfHlgUfGcPgrrTfomfuk+1MZyMJNslWTJz4KynbjM0yw7
4YJhg8UjYIlZUQAgvMNvJpo5CU541zQS/v6Bn8PNa/BK2y0TRMdZpw62g0IszITWHJ6EWP5SmPrB
DFi/cdywhpEFQ3ymRxoPyc3HUD2D2zwed6Fy/IG/MaLYeK5y8G7DiB8PmHYJMwTLPnL8pU+dMIS9
4IAI7HCq4bnWB19Fco0ay4xKf/Ow/MN+YlKuwowBtyhuGOwFyT3BdQplXWpAinHTDgQDlJksISIs
OiVMKlNzLRejJPeGm56rdwj6T7ZMC6E7sW8Pui/kBUTSfvCgEhrTDdL1eAJhS0wSXTwxLvuPJxk/
S8n+bg+aDZFjNf2Eo5iKqqtzBW5wMja+BShs2TmD1LhWkHVG3qcjouTlUPp1AAjL/sjzeN8XeKLu
Kif13yn1R+F25qmazhjN/oUx9ObzySsM2aw82BTyGD6IhkQVQXwh5Ocucrk8s4V0FE95qkMvH3mx
YDUddXb8F0OTs8Ogz1p0y2YfFC77sEtxdb+bylL5c1HVm213o9tQjsPpAaOoFJghj5MgnjWSxxCD
xMoWEl95bSnl3R9WV6NNumNe8UvayW4w1EFkGNNUOCaZ6AhRIn1DLFKyc6P+EzzUz11c5HOizwxE
odvuw2mZWGgpWezWMjZ8Bl2DMt8Fg48n6YRYwujb/uw2+s23n0alYOLOiJuBFfdQGGUfAZvwSjVe
GJQcYy7OumhWYu1snfrNPbHVsPkjiepif6BjLM4KONJnITdxyj7363q+v0Z+SFDZ+Ggve1uVLUrt
p6pxiq0O6lDjtlGoXLJDn3cV02+lv4hnZA79NFHKdWkvem5Y/RGXHm+VehJktYDXeR2sPF1pn9+y
MUcJIDXlH8lHFRJENB4voK728CRkQveBv70u+yC2GSg6RZQAdtfc2uiHbXrFT2ZFO6U6k/wEUvnl
5bw6x087Xxzivek1AiDgL+4w6KtTxlMWwefD/23sSZ8mMXY9aP5pR53DPq87FjWAf7Qxdrxnw6FA
nCy1FUtqiVEMLY+X5tssjrKq6tLrG50HVeEOLf1KEGSgD2TiKFwcvCi9gMP2f5woVizHKE8g60ty
Wl4cAICfpFvgLXQ+LFOPhpYzMvu8LMCwCiWrzDH1QpFiCLS0X9AoStVA2jLQOX4iG4qGUwHQan56
mlxGXAFEd+W+C6Ms2gTkFpryD5o2IzW8IC8LWIByCl/iKB0ksFhBqZK6jUqm4i5HuA/cSSJfOmt+
HkXunnh8eCbmDRCkpLCPEu+9/1UPPPG6bx0qSgIWJQsyh5mLvOlU7vKIWHNfXTSWDnU4ZuMF7FV+
X6BRFI7ufmNjga4WG7eHOimYX8cv/W3wonh5Y7971SRA7gMPtP06mdJJG+N/2jc91XD80gV2q/C4
LRTS1h4Xm8ZtUNsEl8waCZdIG3aRZCYgY2euyyMnbwJ2aagDz/YYmAXX5D6NTpCZ85PeNpYd0UR4
BVVGSpGt9olayBpa+CTSHf7j0ADwgVPoEVoEvZNMfq6KvnE3YRvEZYXeqwYVbO1Jes7sN5nq7S5c
C+CLBs1+eTAtFRa3V57sVtc3iz/sJgkzJMbJmr+VKJIXiDYoBW0Vk3l5NBAwnJkP9emn1OISpc49
DZy1Xyhty2p8pL7oj8Qy5MR2fx7dxqH+v4rrt1kxvwdJ/jsONHHkxVypxYNNX57MfwXNZGvu/c/x
zQEnsra4B+pjfGW80auEsBXZQMdoSFT9wyZ/g+v4YHCLrEHsLymSw7ve9ayWHOD1DJ9nNKv7f5z7
bsRFl4yeAKh8IYcfw+K4VPkJorTPhL8MUZ5peLmJ9YonvwutVUaQwijem2NzWKaWfxyUbayIqqvt
sqdcq6BckKoFxWB8kZ7x3Ocfy0lznDV3AgNEcYkru4cCEGjF7WI7XkpEkFKoHK0u+9UBhx2Qu+Mv
sE4GIlaEnvyuBqIINlIkkfaLE8Ol3QSQeBs8EoP3+lO8bCxmAJSokPIVm2r3Y6mfD1jhMKsGKlAi
O7hK7AnpWHBSVqlSGUVShj03BkOn9S1DYRsxiavEdV9DxJ064Lu1OfgTlGFOVg6GnkNcTJrYrPkW
rYLrEIXdTGcjfFkYTW8DQw0nAvr+DlpSMFgjCeK6uZsPIlUYUvCQJhIIdw6t+39GN4s+yNt167M9
Pj94OWVteWCuP45m3QZZhDyCiJx7OggZqCWfpoYg7q0/gqSaZ0wr/+NVl30BxidycER4AaRU9iKE
dah8teiiYRQ/kYEfMrMILLBP+CmVcmRKDsfjRq5wuK1iu9pUzk5FL0cFglFUnYOYgDX98L2AOQ8V
1J/vPMO+GGq9xwNR+9+z/NWwDGL25qLt6NToeg5+6dXDdoV6Ow+l8zzUt3V6ZNvRqlMu2PVkQj4B
mOVjz3WlCAPI2v2AVVydwj3G2oRA2IsXl8q2RNV2vXLpRb9E5f+8Yvvgm8/L8ygdAHDFYG/LU2rU
/yOd3folnBRmD86kDWuvxCDbdyuB+3s8VyGlyhWU6s4C3IOYB9LgCIaP0YQGuiRedfKX6iGTOfnQ
ePCMN4ZvePSMYEK/CjscOjjrkIDsxJYXQZi35Lqh6zvD3fKr5bZb9ZdkJj8ke4TjHeWXATvNYGgA
UVWbS15Jh3cnFaXHwbC38EBrhB+VTUTvtwIQ/8BnvYS+l/f6T0hbOrw6NnbzJwHl/dGQtl8tD0Rf
my5pF9/I3ooqPfFMMLK0q8Cs0+rq+ts0OBjtKeWQZlOnFUGJjIE76/cn4ja8H16V98PapzFqfrIU
YNwDnh+ks0HoB3hjmC/gbKEa3bGcznjHCLnWAbPEiFuD4W0obloP9UywMMZyVX6Sp3HouOYUDzP2
TYJaw/zgLoJ0kuFqstE93SfXVAz6TGED6O3Qfp3UXNcGh1avtHQkyoKSdAAdhG26QXnpoZIdgeif
JjkkBxUAYiRmt15A1mCo1QoM6vm+dojwmYn05zb5M2NrA+nAuvj8Z2OYs8Xyp0OudAzQHZVLWliS
OuOLqlJZ8kwrucwFuYxMeC4VtyBhK1pMUlazPt1XsPP7g1twFjIgnTZp/PZlikkrCJUHgbcuQTrS
GHY5qEoTD4R5HHo+G4ycOc6CkN7Yp6EEkFgYUr59pcytMOjF8lmk6oVFWPY17aHILjCbll9WiRSw
3cjQnPps/oxEi/Nxq1j+UWhAdKnNKOI+EKDZQGk1vVKMreH1DZl9XXnu8YexaddeMlHagz62TZkT
Yb3g+YU3CuML6hzVT3ROpIpij9a3dCwx1ojbZwpBoWUdiz0+C/eauda0545tUz0Q6jf4dgVAvtqX
sP3MnppbaEbi4YwTovmiKYqOqICOA4zp2596qMCg0z2JRSKdPzxAdK0ShaTYDKEoduOzKqlS2n4d
JIcYu8XG3K2KlCsIsDv4uQdCREqUFZ/CCbGQsH3jHuv19CTJmfeubABuI7fCICs898jDi9WNdW82
oli4eFleyrTCX1Dtx0Gti1TkOmvSqS+GdjA4Mv2AAkfc4gvBdAIr8z9iW3wVMjOKpz8Vuq8c04xG
mvxjES7Enw+nuPsBwepe0SxuenPXMpCCdfU+X/3y8VcPR4KF68lSJzWsQEDlqH3V305VOBQHlL8L
M87dJa6O4xpc3BE4HRLY0AncQ+rcl/iZLX4kM7UcN1vtpRGqtnaXixnOE3qg7MXH9GvVekAKJMoE
XkDmuIj/KGgMESdoAilzNBky8o+JMWnzNxkmei8m4zCkBsBiVS3zD3vl/XgbAjk5KiM8T1ANADSD
2Rfgg6/yNDf/IOZkb2u/ALGms45kjIzhojJXRD3I5hH3No8aCaLvlJto3coL+Pb7yBzbR9XAAh5b
+cqN/WvCebMHdtt7B+1mjRksicN6pb3OnNQsdSH6BDDXRjpWU5wsmIJx0Mfcnvq+By1EHDERq0dN
KUM7IaTlJyuTdl0GrlqyQKuicwm7LJahbwMos3EFi9ZuMVg1b43hE9sKaZfvaNKlaIsWddg9mTNV
q1Pn6gfwiXAEL7KcT/DqgMduhNArsFXQ6WEKZC2zSRWzwYj0y/+ZUlf4oeA6sZCgBwFkH7/sTIVv
MfUtMBHUt+xG98f3I6bo+O4G2J1wMK5lPaMeOXeLNRRGs5lTtQdYQyqOU0cPqznU1YFFxVdIrZUN
2OphnH1sEkqq6J/nmBSDf++TRlm7ZqhOO9v5JIbXXVBVwatuj6gK5CzFwFlK+Ihbx68LKR3/v9S3
6FtN54cdAPsrhDrbba8FP2SBKDd+XzsO/79pxugkwRU0xavnERwp4639ZjaptNN6rOIwcL528+Hb
494Ev/t9Ui8Lj8uPGKSW7hYSn8NLCwkRHBUlC5iz93XivQoOKQemGNIIuUcbYt54pXGOIBvHIMSj
szQwMAWPEiNBAtTYTY7QuVw6t7ek2ePr41QCUfnpIPq+kLpG4kB1VmdVDKNZdwODb5uUswqA3avD
wtgHi51uexU67JaH0Do2Ika4NGAl7YCbcYRUgTC+G/BC0I9nX8g0uW8DxLA1SQjWKBJWw+7CHV5Y
/bMYUdYtKhax+xhKTVUPOa4gm3hrfkkOaKHoaFPxj2IYzWltcWk6lt8Euq7g1uGh+hCTAjyU/NZb
2vs8lbrxK1VxMZktWmlxFoYm3iHESAJ413lSHr6/ERbz0Ud6lma6AGDBuLVdyq3adDLXPfdLUegL
MvVPEdiDda8GwYM848a95sBr/8DigV9Cm2erhGxxiy7/boIVSCqtvUEv5Q3jE2w5LrP87yvoxnI8
cZeu7fpL9DhKSwj5tK/3PQHa+QGMRRhT3o0jflrtLer2xHamFyNhawavkb97iHuU+TiNtGA4Wfl5
GHsWRw30/vqiXpIPbzgScspZpqwX0CZElv5ciJoFMRexawM52Huw98akdLEh7PpVO6VQYKOu90V6
ucytMXcbAAUEhT4ApuQRkXZEm9inQBShHztX2bdug9hiLD4L/yfQcSAni9fRbtwcwPMhGn1xQtju
gram9X2IOT3KVtJTvijlHB2Q/qD1VWFy5zHnPq7UolLAo2QWDXZos/8lZ+16Im08QG8VqgeEfupp
e5PD1N21iTiMt/cw/HyVAxRJr7mKMTgrC/drOaKpDpROe2vBpzW8HSmnRDD7JTlbqTsESJS0mJD2
hHN/FD5v7zTgnlIClQZBgu3ebBYTjOIBdOjEnvUQwykXyglPfUiRDasKThTo4KZcw4AfBGTQuUS3
zXBw4g0VK56KnYyzODJCGz+kqAjqa2+HbO3QHt/KiG3NzjfDbtl8QC03MtxfWj2pbp7DjQzmspg0
7pNUQCfeReMc+Gt+D001RSO/Ed3MHMDNSwqBor1JNNoOqg+dnFmC5Zz2MbxPSWUnPYfibm+yDoCi
0lqFBHR09jyXSpskGG4OYLMTphEwREYzbrZfWfSjCCK9bIXlkVGlsxPGs7V36xjwLpNR2IqW3tU9
anibJv/78ho8Zi4GaUQsv61s6KRf451Jmr7156H1opSbOW3KlZDEsrpncdjOUlXToVYHnJIp2Ny6
Abrx+b+tho3ONxXeVRYewoxszZBr+ZNyJS8n6LTvLK/kwKTeDvovNJk6dwVp/DFzBN07spR6zxYZ
eP+69QO8A92irD2vKAlu6F0+zF1hFElFzRnxIOg9bMgsjD9wY7vKHjbCuJRy6rquaTiAw2HcKIFQ
lZCuDuqmsm80tYgSCMvp9ul482Zs1AueqWH7IRcFfzX2m1Mpi00y8Hzg8XDgUdguiqVxLwPEdcZP
XodXiqLiT4wsnbcwOUs0ubviRnUQWMHG6o6qXQzemNs/SrrU41JOZYRMsboLvLosVKv7xRoKCldA
bOfxuCKe1YdHj2Dm5aBIQ2/0ea7hNAXoWU1q8zfP8UQfGIlqH7CmrFXWvwOl1pivdisIASAq3mZO
1QajzzXwiJDDnBA1He93EIy8n3Iw9cXyY97wV6eoObZKY3gK3qDDoBhqqfew9XxOcZsxMEGBFGzs
0Gr4KHV71L/FiBkpk0mwJ5PTFR8uYYIRL71Ix5qbsAe+R1LjGjAiEZP4lzCw4GvB2k+sFKUsr0Qw
U4SN2I9K49NbAKAYDEmTgoiBZw4sNzSYUEuySI17hn3d27Wk0SGfNm/a/1IN5UgynmKvNwlsbJ/z
mJTYtcdEDo+8KjnkBGZF6Gu71DfeAow3VBA81qsvVKpsdD/K5TnbsYQBNLjEOUV+JfDxyaI2E8sC
lOBLK3pC0HCi/WjkO7nDIopIMiX3XKyNU4VBWb91f51fCEvhZWDJXLQvsJz1g/7bq+dXDl9Ew//G
75HLzgIJIPq0zHrEqMk+4kH9OGsljVyUZt7tcwRIb5kIICXQqtpTplWqhMsFJTGv6SXvxhrtSbX1
p1cpxMHVQFvconeonMaLCS6LtMP3Bi19dWsJc9h3z7vi5SfPk49Wqn9XCEamV5mvNA7oeUK7XLL4
bfCNxD1VFEjVqQLDx6k9+qlv8cgOMQnDOX6BnA5TOHBYnaW8pVhRWqjz1Wecc/sX4C65OIRcuo+l
9egmYEHcra4gKBdzL6IiNvMq46/yuRkhHa/y5v6kDxPYDJ9g+dJUpZI/HfL2rpjg/ml6a70p4ANT
O3bgy0W8ulLGAOrVVY892kaXrjh2+brA6+aGG1gBxkPeYiMsiR8bF5Qe1n/NdWM+3tKgv2TaoD4i
nxZ1tqeyJxVCMapJWPp1DTg9AKb0bHigcmoiAv/JCDFCHHlBfecYvLNod7gNZVnVobCAvSlcFB9/
8wjzUiafrNjXUmOJ2y/AhCYVimGSM8CezQ01ccmItRyylvig84/hUgpKduqQBWZ2VmCtoWjRTrY3
FOnLt4s2ORVO7hXX5tyt0Zn2r2VsgRjGRPjyoAvlCiU3b6+Il82IqL+5y8dDk8eMrPLn6NBPWMBg
giJ+/HZk7g+gRvIpYFr/lMGTuqj8f4PGUEBBdoUputTrDspTsDAf612WIB27qZKzqmv2RTeeTwtj
FgpnF4v4kmZWxBInLYYZnSIOBFpA16jKYjH7zOXkMeKFC5vKtjiEtapNkEXxQeRKVzGHItJk32+s
yHfDQXLfNJn+NpqFIKhbv8H4nJM6Nd10zRjwX18cDstm93h4tX3G+ZIc2vKKkilUStT0yO/iPO7e
jGjHcVg8m+Ll3mYfhJMiqm75CxzDR+xXlQ/v16kxKllFigYOEdOb2Map3pKI7f1SlhFQ1xc1vo0B
jv0wAhyziAGrMMIug64eou/qnb6R8Km7TIar7Xj5vDHb0cZQ4tTM0mtkYPX0tbpsUKjCpN/LIWJg
hJyxU0iZPNqTM3Mtwubbm7aenM60h7xW60zoryNCqqVGI1vGeG/zfH/FYbuTEZikR5VNn5Jy6C66
uYUl1EmnKnyZRqR8QRlE4cCVZHNoCm2NX0g3HDzPzMjhqMDv+4rtERfHSiQgzuoMQhk+tirtbgJ0
jiprHSmsstOBi9JjRZYXRDWLq8zFY7hHt3Dxai/LhXaduKzX0LI7W/K26drk/dk8twRfH+Xb+rnh
af4duh8wS59FO6i4VKTP5a2Eh6GukCkjM9t4sGrR++nm+l65SRjPxVmc88P7WOciYAsNqwZdDRck
2T/W51HBHBwIMak+QvhTl47GWmLz7TGx4M5Jk38wX+70HT64BkJVup8zJtJMHEdDIAlmHHTCthU/
Yv+BwMB0Ses7C7OUhOhX148kNQ5QrBBt0jzRjr7uIN8J5HLgEuvI4T1bZdKsHZMTWVUuZehmqdhU
XH3fWw0C4lsAZwN4C9PC+lO0kYqfPReeLsub2iXor6CaNwKyrBLT964dUu8ebeH2lcewJaUr6tEI
NxUaE8b94psx/m4HGJfNB0InRqnCkwENCypYNxMSI/nxEb7bTxCRn0pNdYr5OyEWYMaw2yM0mGEY
MINT+9PSWBhzNO1X2WEyQvgKK9R0XtZ4yPtYsLSd6bBnaQMrmixaDIydTWsWU4qPQylUfZu07/MD
o8coslERBjvBIOh+8C00VnXGVQqGUfglb2xD1XUAtFv9LuHAzNgrC0OxHQduyS1VfLIGIuZll8OL
jLRsnmzY/LZwZanG/WdK64jgnu0ohwnOQckzuuhS6cd0XfMUqNrUJ2rToSEG7/THXDiJSM2Nbh8j
aWFMOg9QXauk0b+gVcBUPMOwNm32A27j+/AJuI9qgyxZu16TPdlDt9OHwYtq2l4275558Nw2o4Wq
hvZUGrKTGclSvoBlOQGJiM2HGGAmIEMSlPkKsh5J+KiNurDDLfD11kZqWKrS8+Us4TSf4gxVAvfi
juU6DE1aqjQv/qTSoN9f5mGsOsZa75JVF0dsHh//OrRquBnZ4XIzaF6HLs9D30pKAQUuBu/pea/i
QHKJA05xjVektOIufOnNuxT5R24pAmL777OZj0MqwpGwmYu+VZQugpVEbLaEqFc8VIRr7LDtiR04
26EO4lFvrEnX2tw8yidlgvqWphn271HfOBVgxKV7elhoESg5RPEA1+ON2a9wOP+6wllIfggogotj
0Qf6BVZjLTUQSKbKXs97fQ7tMILWVtLW2f0Z/FcsOtJtwtsbYMZpShsWUZ6EqjbC85gKWpsZ3XzD
V6gZs5gDeTkpXYU4kb5sOSyH0xxNhLm/P3JjOUFXzJV/+eV0d9gjP5ReFiFoVeirnvR2g1h5MzZn
G7zSfVTu3of2bUksEKHLtHH4UwKxoz/092hyLmVQ/WISsWlSaPKlHHVgunpqZ04Z5krdpd0CM8Mf
iWEdvem/TyegJfkxHlTuurmc6s2Mu9Nqc6Ik2yWBbfguEbnpxhGtiTtMgomDTdYVuds6OGzyKxhp
G1H6VlM1exgku89hzkJUgub1wIGOXd2XYfnCB7tuZC975/NDs+rucTStcKcPAbbRjTt5dbOmJb9F
j6ACDmdz2ghGMQxLeydlvkORDVshNKfAe5rJ3870Z92A214BL5PGiSeeJx0nxyutNiZLP+xGnFxQ
9EaWsVlfkhEKpO2FqRcLWjSFnDn7zUvQ7U/rBqOJzsesatTwH6AZQEIML2ZPM0tgvX1xcoACMolt
hLZhZZTuTQmYS04xtRKqfWcx4Pe0hVRXmjYrz5twvRtulU3s1XZCc4p+P9GcHeqOAozwolhEe51F
PliP6UW7SYsYT4nVp+2R+ElTYJuGN5iQ8+pPKkdMiSX2n3qyynHBycBt+h24P1Uk88IxjI8Rwc+n
/ywD3v+t2eU9A0Tv8/r7eulOWlwtsV7awEkkRijYiDQAXj5fojS12mNMaq7Rd0UKpFKYn/2O8Y42
he2bvM500dvry50e5yIePTs/F6gD3VFMHoCYFFcNiC5Zi+soGFrDLdtQ0N59KYWflQ9R0k08SNrd
ERolPAyQudJ+Qn1/ScGrHTnKM9IdRoWH2qFiiHkPS7itza6HGqnb7Puqnrlxoq4MYCpYbm5IZbxO
4EGZ2qOyjcRmKOf3qxidh2E3i/UR7bNx8kkHlYJd1rRGkCN1f8LpD8y+tjUPeuevFwF5Sl7yAUL6
YJQKVxulO2+1ZMK7dkPuomDzoFK2IA3BnH/Ug2yKJsEDLSiNDHJgX+ygNOcXqxdhozYTPrQ81FQB
UlM7vDSyeOBW50CNwHgCwrwKxyOR3Pr6Mzm/B8KBlQsXEnDlGXLzSjLqM19KVpAZp6OrlijBrkF7
4rcbUAXUb/x8yvaPQ2VzjUUqjjNzDMODcKjwGmjuD78cbwtE2U7OXaMxwdUZmxApMuH1njjzlbQ2
m6DJjiEYiCcHkO8FanRRAlV6p3AS/bnjI7NWg/Qb7zuh7gPtGyCThKnnLkyHrhDSDKr1cver6Tg6
ZYV6k4Y4B7agI4HCg0fBMBmN+0BqV4gMuzUyln8eWBUI8GwpBx1VRyZm3YQf5KC7qIUp9QzzwErJ
UZIf/QU142qAKpQN6qpMbl/S3tMueT4MdJbLsbM1x0WqUy8KLAX3T/o9RMMT0cWSeW86qNiYmpKJ
t69/nBiCZnAhLkOoVQOQadIJw7NIGHYucxi3TN/KiJMFEnd6P/rrdTwQ4xI1sa0OGHS4FQ51zOZu
6ROR8LIwD5oRo0Egjwvbl/RJAB6bJcBBX360OMGrZPhoSKNGLmYM7IBn+wslxCe1CNsAYhfB9HCs
gIHJHuU6imZb089xBAt6mJbx7n9yMBlnfycTvINZFXbBrgR2OyP9m7iI0gGN0keW43lY57EjhJLO
Wi2WMaOBPyU57Qwk2ni5SHYlMHQZwWuEKwoOlL6EOWPvaMIG08AQrB2sjF9n5WIprsBjWHjCA08l
Zm28ehLiN7haGhwlurTkNIJXXDJ2Hwu+/FvPq5hEZkGGMSnClncNSZrmYHCWww4qr7Qcda3T7trm
LrlxjdjP6w0B/n2OWdnNny99NcQ/uR+IwCuiEzgwaVVHTalle9Zk+HaKDYfojoCSJBTYUc03bBRE
0YHLHP3WrpJZdJcgJdsJM4aRdqAI+SQGbFmUinGepMVwEvNwy9xnQ3hDDxqg7R9PK5R8HUP+fnL8
bQtVCFzQjpcBS71qhSmEdXnaMkWJhK9ROdOvoasNUDD4K6uC8opMlJOmWRsMveE9f+AwPOnVHaHv
P6uY4Et2A55dNCVIqfG+YXskyUSwWkOajArtoAeokuUY8Upt6ZSBDB4RSse0rmjL48JFiyH4rN+z
/X/GS0YBviG6ei4FGgaepsWD+eY48S9dNC1rhh97rWX/Vm28gF96OwRwDsT9+x88DjwUkIzP73nb
2BZMyZbZbGIlZxxCSYsQ925pdqCnzfnTRabQEYpTaQ4wXmneSLnxAdbI0IgM7lNSqpqiWyuIJ3J5
UALuAmFFw09UjAvhz2Cv9SMxmzT5wGwrbhveBuAv+b3Jo9xmjT/9wZ7rkfEvyN3WJst9qlVhWdV9
xC0rnkY8wx3UUAxz6VPt2RXAneSN7T20Xk1xloM4e/hOgaWRf4sSY/GkhQPbXAiWH4xj+hlUef67
ww0ClwpHpC+ROLLfksCc4JTG2l5UzPPEga8EE5rPwiMn7fOuus6A7zur5KlFxaKdcF3WRnyB9YLf
qTPoFMiNQ8eJWuE2ryu6UUCIs4NsTaFp0dAMDlKpcogdh3JqcYtGIxsYp3bX1+S5yk1+M9zYr5Yl
PYYj7br0zS04ltrl9zT3Q/nnn3kCzUOH1IeXZcOHLDSH+9ADak4y/KhqIZEEot1ja+PzvlLoFGWa
Xeszj3cjyKbW7urgI18mTaxW/2ELNhoDqv4Y0vrtq5cGAxGu0f82VyTfqTjcHooik+RPdH1ZXxIU
cKLVV/LGDw9vnp3Uqo9NsIEqHnIJ89oMpkw8YRW3PAQf5WvzmrgydBFyhIDlIWxcsU6ZqNob0qs6
z5o6Z7tgqgNe8dse+FG4y2mZjav/wmQwsaEYcNmJg5mnJV6aTbsW2qpD0FxMjmEhyTuLl5/CjHeS
qpXcgKkZr0aKsQsS58d1ZeegajRERv9l0YZMTwbdvZ5sQMBJwkWDe2mXm3ePeAXFaLqGo3SnF3S2
7cdNXpLd5DkZYXSv4AlDWezsn6CVdZiGnT+uFmQ9OVpSmCiFxk6bgODlhzp6IwsZsh/1mWppDUVp
CjPFWLW9tSLyxyAV3CdEJQPGdU2mkSgj6xXU37COncPacCdaQShiy9wAEl/Bz+0HQQKaMC2+NuiJ
icU1fnrJPA5HV6Z4mB5SnnG8xE0vP6Z0FQ7JIMC1jgq7ZK6FMW/s0PrkZN2Syj1r+c6q7sRnXjt0
hPaOaviCTAWD6s5S/oEqmCbvjdejVjbtEBM/mZ1tWJZBccTBs3XAuTHW/fuN9uwlKcTd5zki4H3Z
baD5kVILsvVX7QZwKZaDxYc+WMiuDMXkQ77wXC4x7x5WnI7wH1OFwevS2BDOrAV/8GfIo9fZpu6Q
/VlPM1wESWqz4AcApturFvlQJ6lFy4bj4h4n7trvnnx4vkqQGwuACShuCX/lzkiNBtUNZSRj2Cxd
rZoEFEX/xk7uPKJWGflyQkf9tF1P5hsaFGIlTplOvtfsnOhyTJL/St8es8ebKXXsHpx3LHE8oE1F
4FJkuqwfowWQ7vnOrHdGA8n5gQwMdz1sgB3DR5dmjQCcTyTR4kPVHI1tIC5Juw7GL2sfL1m/YOCc
lfiWOhP0MOPYyW1r0huPiLAtMI6k9zZxQPspvmey3+8pE0jpwEz3dADRjVqZo9FN6b0cWLogow8m
VJgPNCrwf0Be4tLMJmYYoV+Bdg2dsOAwnjEl9JY+RRmXacb1pWjC/cVMqCUEJ+9MMovZtmQoukYr
a/x3WdbJzhLLEFrufOo9b63Kc11t15G1X5fEMi4ki1a9kfzU9napsye2r5KeUpQ0TfvYOujAwwjF
VULXH+37iqLeKATExA3tufcQ3UrGuZMr5aXINL8rXtXX6ZsnwCT8GKcY0C7AYR5tpH3HeicWPOnP
pv6i7xC3HuvCq/iI8wJ/1OQwkXZA0z/4xHCmt7W6xi0sHYCqfUUmhVoorsEwx5ckjn1FwxrXbyyq
r2ykEf+fGmhtdcfRnVpyVz5bpo8R4fTXbHcksR8d+0JXf5MDfqjC11R105uYxx+8k31Nl91cxLf2
UlG9US05scszN2zcN/djeAhWjJbuXIKJH8FgVOfaRBVXMtzDglqZbg99U/A/dnClN5nOozbu+v4b
YDoWyLLQOmzdxKKsYuX37AEQ4v0jE7R6iBWFnEZLFoKnRLle/cyUC1PN/kVPI8FQxMrgSMdHfxOn
R6Jp/nLJ3XlbZrAaZ/LzEcGY4bnXAUCJeTT23NKhcQ20+2pZelIrzg4YNx+mTQoai3EOMW+yXcUJ
iK49Xdy81p2r+jUh61ibk5+yClCl1IMGQrpF/ITrsDxjD0XKn5v48AvjCysKoZISugQBKWmFWp3O
724F8wIpgtu3fO67skQdb9dmCSaKH5B5Y6UReSVz4akWV+5ohVXn93DltCLBG8NRRADp+A6rRtX7
0osihIhtIorDdDUsW8yglbGAgtmbJNBxRMOBte1pgeUPCqZtgiw2os7tG58ECheYM1E/PXE6IAMe
Xs3KRqDFVlEgew24UrLIDETDXpgL7GBYjP9DZVJ94eAXlL3FYMbmcw4iQj3UzHDndDHVHK0JeZFo
C+QdQCIoiilHc+8qajVBteBNOI5FJ4vGaJAxVuIYl6dCRGtFXF4crQ5b08WNcYCypo/yjBlFRREt
n6CXrjZam/h/zdKZsgd7UXJupT7bk0bWa37a0UwVmLaqR8OVphm3uEm6THrWr14/ZFb6HeeJzXkT
qSd+4wtk7qk+KiK46PJm9fXcjGas0vJ4mK6DofZgKfrsiukG3kzdqz90Pje2fC3iUNhEBoU5Nn7S
U3xTKLjbsrrX6mjMlfzzR2Xodq4hIvcG6+qMCP126WzFKUOzBNady2mCbRFz7Ze+jmO23isL3e01
D63+2hc8Q+X17dKbltzLSDZ0L65SxVr6XJzhPiqJxWq57EcZKgA838TS9ux59J262ifG3Ocrzc1Q
E+UqGsx8/7xD+r2dv3K+kjpIpegPPzNDTcZAk0h/7liuNXUuo4boNmzRs/T8T6mhM5f5F28rmhcA
Ud2xAApm50hAsTWFIAPk6NZ6I+Yj5ukOhpdiYZyyV+1EAch8qczgxrSq92nW2fTKrUMy9oEERATg
W69Kfxmare4mxj/OfGi5FjPJ3GAPSvz8zwnaGjVW+oLxopUvv6BwhhL44OdPoK4kxNxcrCXA3QWF
E+wI6MjHoye2PAzEysUdUXkfg9xxoMVbZ8sjvKDl/bXr5CuXpUTSYFo1pHpMj8+SnUS1QSqbmPeC
nNhiBopcN+DFcVhRSNXm865oFurQMPsePwdvobJ/khElQvQtbrz2jaRQ2VjLREBpadDThTsHbMg+
Mw00aXIGR8Z7I6shjbKj4wt+zj6vOH+bnd2sAKjs8UGUJrOGRF/GOBm41iPy4zH/a6Qzulcja4Us
ScM+R2ra0eFS2QLDzjifxD8u5MbNJs6dCzfQfUdzqs0fpBc/7VYL4teju961gJkhm8mE5BvVzo7N
mZDrNQxZPHPcF9PtzOIks2/vbugSMu8zZoVNjzti4Yd3Cpm2G1PjP8/NKLVsaIzSXUMBUExNrCIF
eOXfLVoFG04oEGlPZn3WFHypw6GuNfErwypuDDepO4k69+5zEQAn/6u2LrqmgNrK6Ulo/GSXsV8H
+us09dC1NV9kfOopk9spsq53zeN9n125PVwJp3+HhdVliID1CmbRKzQEywVxqPoYMP4jLEDrqSLC
FqcVCY/YFiydTGksghUgD8jhiJrcTURdnkf+q0EewQjgfw+Y5/DxiW01agQcXn5Gk5DG1B7wsDgY
7gnxp8lzbyEvhPzLxEs71sIyrwRdkv7vXEhBJ/0S4V7aA3XRfZcFZ5sDqGzEVg6VVE2D21/eCOAv
BBDNw1pNVrIKcX8eRjJ73ZV0jXqRHHoAZtkkxgNpBeCKtJao6Bck7Sk7tWaMBMaG2g9T27y0nrht
reENCfyTcy7bh1n9I91RD/2eqztyyXrjxyqjcQ4/VKgjrSZsIFN/fPQS3ZlR2p3Pbaxu8235Vwp6
f3ypw+BRix7i+hfauAx3FRSebMz14sj88pJQg8b9HxklXT5R8SumJWTdRbag7zWLRWBYgahOo+Ct
ClRcy02hQ8v8HHNEgysybsa25CacQPglMN+l1xedACdlxRZMvVrTS0RXgDUuCyVFrzOKzKiOisvb
jJ61qZoDUG1NT6wRc3osij9sGdhQP09w//CF2jcWVsvuJh7BwprVbYvHQIofccLcjZDKG1WOpSCX
mF4WbR8eL0Q00aY+nTIg8dAjH6yZCnbv6ThJNsfZ4IxCuqvroxyT0N5qM3t3V6GsumnAy8tilttB
JV+QdpRPupjikS6jXELrmMC3OOFcmp65A/9UgrYPCKErnpcKPQiRV1CIVWLneC/CChB8qwe+yvqu
jTzxlzwAXn8eix+gPeqRSuJONL6RFOjKYWuknphnAjSG8LeBlqnc+O2YLJgHJbToHk4hxNOBZpMQ
/YzPX2O5I5Iku6JLra4TknTH5sASeBNNYPR83Kvf00w1aMItexTu+hPpx3S8aaMWi2jkQgseu291
tfoPiWQ86fLFZ6X5NvwiwEUivAxrHWeMBkieN0Qj5Jvg4dX8jmEBKKeidheUGOCRJ06+9ZS1BLko
rOf1sJ2PfEkVqai9rOBepZkAlfEa9hqWdrmW+ZthEMFTzbctdTq0J/5D7rbGZoEr/LY3JcC9rXia
XSEHpW1JxBPC+i5yNOr3baddZts4fCIn7O1eIa70OeYYIpdAbTptlE5okc2kyS55NAv93ImcbD+1
XTkJFDTz9x+JwlHe7LFrRQdJ24RFbKYy2R4hjUwtuFLvNxGTLQetVvISlUtbPx86vT3237oQaeHs
q7G7dkzdHXlkWVMOGMhv3PPqxfwerXeS296zUxrfNNhKsLBx6/9bam4h9eJAngsJY8u/yoTIyCh+
0Ef24NbnIJNC2wOI80jiufSQUUVqXwNziyRnLrwbZyBxWPR1VpnkX8xPqiJR+3eGPzWwV5V/fmFn
voXuvZ1zbHhAEmYU0XQj6GIf3veTt66sPGnDqJ6+VkMoDK0K6kbMzwcceJUutsquzNQvlI9cJiTk
5Uzj842eraf7NERJfBQhO+JuyeCMwym/FQ1W6CSoeDhfga+JUdJvvVsJRXLI96OfCibfwMnyQhct
LtgbG0LKvLVg9l0f1C42nNPjlMrmVFS7vtz+vft6Kb2AyDFjb6lO7/YilaWDcyBNlvfAMUZKQcWk
2DH02kM6sWV9g5v7dP0a3lDXr+GUqtVrqdvsYw5cUTpwcaboTOQ6O8+fdci2Yd4eHTwEWk2Fg70q
REa0Myas74KBH9x7r7Nnk6jsBGap1cv4zhYMKXbmeJgImpKY3cK44ua3BLwoBGuWi4qDGA6dF87g
MYqOcbjMXTf5g+3NtgBEsUNetdqRW4lj4vZHAlCXGdnSCUOJ7Hym/cxTFvuFyCFDbGblfS7VYR9Q
8yXU1jtdcvWaRqLITqS6qvOc+qBqYhKQAQuwXZV6YwKGoFESRq2HU87nfp73doKhlilmP24x06pu
Ek4i/C0ndS/lcQydVvEmp5HMrrB13ehIPuEC29yQbop7CfKbXuLsQqRu9Xxtae2onp6vkmPmRbDU
2DWyQKfWdP9t1cU4SoN9y5A6NXvqTvpyXGFMMUVRxJS4DseO6xTbntUcXHbWabN4ynKTbGQhp4z4
5qNQHRoxGjOWXeOoLve2tVvtMuFpdISuTiRwvpi8EFuyS8mbgZ5V+Zcmr3q7M/upJ5q1eo9IvQr5
6KiIhs73gCjZa6ck/1ouOX6H9ZgWoTdjUaCy1GiJ/q46OTYJ6AFu1JBN4Max3FMQmQIcHtjYsFAE
vNySonY+rnROaZdZaBCZZgtjCAbWr8YVUq+6+xW2QhJnBJg1vyKDAlPWyJUVdcUSDwQZjbFCqU3Y
BAKYTAZ049TF/B4xbM0E2NuBvjV4cDzvrmCuFUqYGNDLvT0A88b4QMvHn2459vycc2os0OsRLKkX
jaeyhyTaaCq743gk0vgCgByz9skP+NouwF/ZtnTjubGubwI/KxbNSYA/b3u/uBpVE+I5Zo2A68JK
rDr1RB1XKDLBwHmFpG802f+nP1wbPvkI7PXl69xkQr+zEYhbsOTlws1nhT5eC2OikX9cd0AVHEjM
cSJikqs9eE8ld0NYTbNsPHcsICFosOFQqQKtzvP61JueD7udqlO+M2yyZ5/zrkYQHy72VMHVVjKw
/N2uoFa/+uhU0TFFnCHZ/DLPLwsX/IOQRE7becAdW1RykOffxC7tf4ZHP6q7SYiPmgKiUb2L02FE
OsIn+zGHBnnGgtFzmJu+vhG+EpenTKZlj0G2HQmb3G99GDvHvM35VhR+oQhXO7dsJA+N26Wo5gK8
nJ4q4u63tnjK6dlzMhzClcBnUTtWyK6Kh0ygmSAWIDDusZmwawbwPL+2vKw22jm/7Pzsyfe8DEIE
dU/OOZQ9DhD8WzCc9+Yi9H2NlxI8PURvCJQtT7gIT6qtoxiFMzHBASgV6ZxxeoeoXxvajmXDnR45
5I0Ac1h1e4yt/Dk7T8+oYY3H+/mTytWh28zAq8mF88+4ucM6IdRwULy9tzkrtf8SRCVOl4HACrE8
zwQ39Ed0eVXKxthAmhK2G1oEIUu9Lp7XP2F2dunfor5O5lnqDTa7fXpoBa1cOKwzaMrI2yOX1+dO
vFH093R5AtDW8BzIaiVIZBKYimB2dB2rVFD/niGm3Gl/c5j9ys0atYDRa0PAPyL9LTsIz6nTEDyP
ngjzI9Yot4fjCtiNwrq6FxWzBZGDBlmWy1oTzZ32Nvj7v+JZbucQGPKn2ql+FXr4jNVHwZfbivTs
9Ie0CSBAbZc5bMWdPSgDNV2zMQv8uCSrYQhlBXBqv4d6dPvou+PX0Fh7gPZwu01B2cAD8MI/z8cW
9L2fPbtoQKUoRCCpMSLuvGJG9tbYUdmPFU8ZI5pFtt0qDOxV/QAB28jB28oT8U7Jbcogy/ABLxjO
x3ON9Syo8ygnW1eIkn0fiew89RLy4ik61TSYi8z47T//K+wVyTvz4bikfKz9EBF6OnZw7gFK0vcb
ChULIV6Z9Nc5IP7aTgvqnZi7u9hkNJce9rGI0GYZ+s5w/ty9p81njufsGo6SiNm0WGAlxGaKU0gh
T0XBybIhHAubu5ThrsjWaNvDjqvFLcs6KgKf7KqYyuE/eNNpH0Pj1oxFYEoUzzHWIO7bCMHZ12Kk
DLhKOGoKDHLqkL34xCiOTBksYZAV3IpjNvx8WmsTmvXCC0MFT4EzS8+w3nyaZaDVw1Vfh6Hv2t3Y
m/WLq7B/t05hDjI5i4jU38R9beKAf4hAGDV4u65egh77cqD/7J5KqxT4V3CbJldITUDFk+uHZKAs
FzBheVgQEBCvg8rquN6f8pznFUFduieAt/ckmVcj24psXceQzzDzCDLNxV6+Eco22K/hbZlUa993
VJfrb8z3MeiRaKOpeawnoNFM6kU6XgzHSHBkdNzi+WgeZXQAg7i5YHtm7/7yb8of8apOtLDLnln9
UB/5OGwAxShi2IfulVKt+33Zk8VavDU1IEq8cPK8x0kFsfojiX1hb2QbRgj51nXo1CNWfqaGg6C3
FRG8EBnEuvCTst9BXa2JXZ3RjrB2bygOwdErOOW4REzor8mItHaM6nq2spV3udGvzmah9Yf8/7gn
b/AdELHnTpXtD9bgZNHBlOe/sFqjt97G3+dZutEswjBTglHCa/RuoFSSdfRtfcXHDSYQJOAtPSh7
17sHE5Ma6t+5m0/xa7y8BdPwfkYFx1wVUd7eI4eRJjsJrD2ggp3wid9DRjwPSqSSNIhXs50Iz7CU
8zQAJrUyG4oBuz13LxEOY22KTwGj+3H9g7UKYgvHqmTdRUUB9SRhCr/H8Qt9F6L3mVeKjIgT3gAr
IGx9sK75vN7kAtKfH2Wgdc29hXxeQAxbD9iRz9+E1NvQR0t58ASLiA3Bd7tBXWTdYUxSx91g5U3b
TYygBJM0h463gdLEvv9hpaEc39Dxp736VgHFlBW9hDh36r0DsaXkHGATDAG986HpkqHP0wz4y1Zi
Sk3mVeHcDgc5PHP2+WaJQt4Lp8nWN1vhuOUxZLsRnpNn46EpYdu022VTX6yAeV4C9MqO/0MxU19W
YR+ResDHP0RuuHDmjH/GFguFj31jmAHNV6nEq5AyukDl49oPkY0WiGp8I1ymJdbJIy9ZaXm+XdMC
nwRCcdwIeJLLEWM8zZtoh5NzHELYNen20xkJ6/OUz86UvysAHdlL43tOdXatgoEMXVYVj1AKq4Cd
SbHyi0HsIF9l5unxmgqVn8GlgDSr/XJ2rbeubpT5lhKaYfB3nnerNHvw7R73tdEnbtKbLHGIf5UL
3Q11y5kPTnz3CLw6VlwuDMIKGacjw73yG1Iqi6FqFl1ASSZHryHVpGFnZLwoIDSSCPipRuCOVv7c
+9r8LeIOU/+usJpMomnnUiHf/YVklVGg0qujQIYgCEhQFWnH+GSifaluH+1B4X+gSGKQ83xh4gmT
gBP9RLIOV6L5QBNSgtDhGvFqWO3iPG4zZvFqCjxSBafKHGK04M62o1b2KeeAVaLa1BXk4/DgM9vP
s/LrL95xU2mQS8kZ1abs3Ogi77VXhyA0vYp1u12O6C5c/somyR1bYPL+7ySac4c07o2/w1hxu3op
McxG6f/tMtHPgFmdVloYKQcE8HpWsVzlxJhW3QgQH5j/gFpQ15OsuUXkECLw1Nhv4t2S0ser2SC1
MimAWrX/xOgGGHplduJeRUki0xTQuz64AurL613MvldDcUHxu3zyGro1/fmcKjs5nH8cbe74ZA7z
xchd1uGsihEp1RR0COMbxGnmlcCxff6N6ZOPG/b7NmgmDDm48meSms74PlKvmsEycUKFXcQUbHME
N5tY52jAPuXkGW+hbM/+tAf4hKYNTldihORi9uvycnNxe08mmI7xNh3GrwJCuqklAY6V+aAYgj1R
H7PK9mwXX7kLkjAQHGaeKBy7Rbf4jCmExISnwvjhjIV31Rf/SjDbUSA/xzakKl2lylGaHMtaCVnu
sYVdQ+9nptvGcwS90MJzFPZ/p3lnZQqhvMzG1Y4pkXm2ZYxWhCxo0OxSkmFf3yrE25Y5Hno8C8Xm
/xlP1iA/2DHPeWVqXiR0mMX0yKaxwwA9xS9SNwvJBL7J1ETNWqf833GXQvMR+MhHZjwMa3oehrq2
tnkXtTfJgow4lV0Ibk0N4D0QqvwZ2OdH+53B0h2cCb4ubnJ6CWwDP5lzhWlMHmzvQ4NQ7fwCVqOG
NTrcY5M7ynvs0UgrgR2c4UZtQUc96gNsNFH+x1U1SxJVIWHLfCabQCorhtNJEENAQ2RvlAux5rGO
T7btEGG94U6JCVRc5Vc4LxQVVDLr1Quwr/yGPGVwlmMDjs/fTEg94PSSRUQOnpBYZPRXgbElv6Zm
drZbIAoPpW5abFAix1gEvfLnE/6fEYABMptvWnNJpTWK+hrKxNdkT8UzkUvcgSVpcuz4ebtuuxs+
dNEaBnJS2hB/uwZof6FhaoPSiXpDrFXsp66yaWL8uiavk3B8SqfEJ/aP3fXhxl7Z9dxJgx+XJRSZ
8+e0Xr9KqKZnTpAUfszVnPoRpjbjtBwBWJSQTy2QXaPmvjdzYNDfV9DsyAvG9WJo+temQdjHdfcp
sAzPdxQrrwcjDzn7ailZCW4pvCZu5vjKfP/elF09bpfmpEbxSLRfthljp5iRlsAq0G77pBQKFrU9
tBAaVhrpU+dV7FxOWX+Slfd/iDch8nO54hwzBi57xeUTcvZUo+9LytUEszCNtE5ZzLPwlLipev2v
N56FpuNPGZSxFOX2r5FGXihmmfZZvm6a2MTLVMI63Qe6d/VwuO18yWAcu8aEHML2cO+9t6BG89KD
a2Och0mHEMxUHWX1WCnk7j6FXYyci7Zqg0AKcC/tjSdSeFqHpJi1cDvpKSE0OTEAz09uF1zIgAgw
M0zt7qzQF3m6GpC4qIMPGP+sO1U9eh0npFVWA7gtIIjGROgabp+78ejVJYvGCVq8uYnD7bhCraJ3
IU+NMClrotVHOxAc7ztDEiPD4dZ/dhFojJZbbtaF/IxmEky/Ozn1iwW7W5w2MOpwJN2yeOycGJii
yCII6nJsV1I0MPeVu7fLrIDqU4f6e7KFApM7FUW5EuiI7PEY98nZ5lsNUAca8bDscZFZhRfTWO1d
Ek91l7FqJD+VhIKUW/+F11JBLZ9ZAVREQetv7pUgxAuCngUznzD/23f8pEkvGeOX7o4qTl7cgybX
5Wy/xUwtbKttRwR4GSxGkunJgXP6sQ8i8MtN8BtmE08Ti5YuYjyhydNFKrT4Xmb4Xw5B07Gi7czv
unYb8TrGRSnxDZdyGmoGv+Hdd07c//1140Ob3s8eMyea0wzv50e+ucXipqYpeY1IoDi/71lJvkXx
jJPd+77/XI45Nm/kl4tkVFQSsVDWQBHnhhv73C442fHmNUixHV8dgVJ8RFAE0ujJYZdP/qzQR8Ay
iqDrhzZGByBkpjkl5wfSJGRKxkicC7cWUT5GQ4ko3xQcU2d2C2V169HIl5Nmq+0HjqFAmSGc2mgr
qGQQuuMd821HJF84uM1mOUQrQJR2RsnHaRGUb1QSl5V+uXicAj9NIHaElo6qmRwrU5rOqUlujosJ
XTyp+Os/t3G/WxWIrqmkZkqThSIoi0runI6K/zXwZDqV+1+bmJS/6Y12etNWtz36XY55UZDV4xb5
oyFUEcrKeTiejQpclk3ANPa1zuxauAFXTX+musjewnn8PwaHJfSVaM+smhA4oSZ/U4h6yoo9u5XQ
gpFgtS6s8rl69MOZS7NCAlI7ex5HadMpGkK6KVmlbO+zQPFuYa2ZHcGmuF37/Z8sBqczrgGOQhnI
1Z+4txH4VQGBpfxmwHFkuTQdEC8aVgyxSEsqEcYAlbtw7oQI/uv21Cjw0Qc9x+W74WMpSBJwQ99l
ntJkolT4fogYTO9i6OjztyDDGlVQPHksVpSlkqAihbRmHIwjA5zOGqotNxi87dIP280FbCpXsjWP
eb+ivAOlpzPBo4tuiTPS32PAP03rIbU2uYqPpe+kPSlTj35qtXhQOgMEKOLmgGCZCyasBIVN8LlI
7ArS1kg5J3DSTHN2uoHAojbaIojF8beiaMZ7YH7EQjKPnGB3LsBTD6ATEGgL45es3ZBxtGMqzAly
yHIsTHf7kMFW6IrsZ//K/eScrAARY9mn51Se3ajgt7aOOYHbs57sTSKwXznJrGe56QbWh2276doQ
esRdfTQbQl6EbTrVWYFiOuSpIQ7JArF502PVOYzQZvx9zHJWWxkf3vF1slJTACCZWmcmzwDFOUbo
2Z0RuG3gXR0I6MreEyYNZw/aQpHx38uDPed9/rBMH1QmvJHm/PFbGh9DWP+RLAdIVPJpmmVJ7hzX
urssqHfrDj9+d3bEMwNe+5C3S1wpv0rWN8DXwagjQuGHFfspuouDu4z7/MFQG5lP3bwRynlNGq5w
fwrYY92Mu06a2qSYPcj92kt+9SRIf62MwmdimrLda95rrEHx0e2EjwSVzzSp548Rrxn0JhsJQsbX
VIKYUgwpkuK/zsB0t1KvtxiHhCN0dSiGI4dKK9Fdfnd1lcddKaU06/Vq87cYoX+4N67DegUCebYF
RuZhgT4j7IKAXRkV7Lrw+0pzubSot+Eb9welxR4ZRhInvctxgrbrzLmxK9K9csAL9Rm+iF+7Gv45
e1aaUKOTAIx0U88m6OBszKgcvaZ6ZRFL5Yq5LPPFYmyF6aG2JhAnP/fIM6yg1PmAQFb96HU6GhLA
lNI7cGgyhUfZhWazb+q7A9SkNVp5Pge28a43p52nr1GbgweqegyhSgmpCwiW0zMAK3XEe6ke5WVr
+N4jQ5Bx04zrQzSX62otV0t+CCdkwML2Av07ZfLGh027yDa19X3bl2yCQKtfhWrJqlC4Ui9F+RBi
qNqfywZPlVthCJzikr1VKKWbmFD1pM4YeEllmRONW1Pu5c/imPvD+pKsP6JiQl6LoaMOg5jK2i/S
JNeLfGoKaaobBClBiItJmYpShv3Yg8imGfcYgDCYwyiLVu7EXlrHVRjXJLYymUqqsshctHRrUgn1
WHAGPesxZ2+xBAYRPFBO15WuH1UnyrDRgE5by2+faZmRGLJNGChbAzwiq/L40dOjfqEJIgUaLAdZ
i6TzQTO+vCElFfQzBeEL34joBaVN96UGZ4M1H5JRyea5lSSnDorvR7a4KFBOYK4VEszNbd92P2//
XdYtxNFsfdJKJA09dBxYG+t4XReQEp8MzNwr1737ZiSfgCpNwKPdAnn099nOnFkJN/5O+ZI7ErBP
OlcU6Flho0Rxhm28NLSfSTGchDqNmHw5k0PCg7ZtbrsF1G+ejmEdR+yeXP4GwsAoY6belbRlnFaF
7mC7OW2NOLIzc+vNU3vyNBpG8bmr0uEqG7pE7/P4BVHM4IqC5IKnUEJYZ0ejCNI+eKbUGSe9kdOF
LX5Nv/GvAQktv5kw0c4qjbNlOMiNqgVuBLsCLtpIV2zW7JFAv5ahRiBLzQ8I0GZqQJBfqFiJUetF
Uj9oIMce7T1LL3M0+j+hlJQE84PE4UqWzKDhjIYPrfQOtod5Bhh5XAw13uaym1ZmZiKkxBQVLd4u
xOPuXJPk6YKbYEzgxF14a4Nb0yF9RbNQFvTaWhf6iP8aWGbKmv1sr+5RR9LYHrK1SfRkoTtn+NkY
oQoC5CEfwsEUxh/tONrNSyus9Tyj/5ACp1U/Re9dLF5D2hvR9rzdyZlwXEoQ+vfKIvFueZtsYtzs
VXS0nYavXMEAPe/fOTBIeZ8489yHff4uFUQPzkFikyBq/04Os/9OrQV49KsTYiAXMfcri6Q1Uosi
m0HAOEPvF1eIEDkODwnt/oFAFHwG8BzzXN+BNFzvASfsgLDk29AnoC8bFuCBAsw9Sd+yF9ggdIF0
79rC+XWv5ZigposRXW2SpHJjmT9Rj6JC4KuroZ12hO4czUhVRn4Sui58a/Fz+XSCO8bTAG0sMpa4
V3WmEWvHmgKppTnzTT6C7umNy7IQOMi7eAEZ82ZKX7U/eqK/XuE7vpM7mHUL0krVlACRHTIjaatz
zCyVPhTv3jvij+VjXQGG0mLGaP3amFCPZTjX/ZnT0X1RPqAlGjvkw+w5fsdDMP1NShNdOjlmZQXg
hxn8bcLSBrVhvociPsxvLHFRKkhK5mu3mhWjG3ostZUvFvfapqOB6s3lsLU2kuio8Ll2eTHFGK9o
nxVvh4ezBW/EpuzH/fDpxK2U/WNTqjgNrUOF9Xfm/N1jevLWMri8HLPoG7cQf6epy65t2MGa9hLU
a4ai1szl9bsFCjOxVOhKUlZvge/m6eJFUyCme8RISgAtEe0sWdKXnZce7hdTq48DgOEpeVeKhPHi
Po5Qij2BMTOLSE1dGAEzqR2jZi7A+qX3R/owoN+QK7PwInP4UTu3GVebW8LPKlqQJeDBwDxkayrR
4sNDrPJ1/WP/BIUUNB6PmR1QHEQMn8qZTxZxKL+QeBYaAWUatZ6c15chfGUmQ26ULjOQmu/p/3nT
0IBk2jCgL32UE4TsYqcmFUTTDUewtLswcW40Xz7VcAKpt2KiasmBd28W7YxzRyQn4mubU+fFlx8b
FnvHhb+tyLEaOzZdeBZh73iiSUiEOQN73K0WvSGLAKLJGPZVgm6rCRWVnyaHZULQdt74ivhjBuxO
5ospi6RPru0Ayf2hBYUqCxdD2jeiYwNOSdL7uBWcKEHUGaRIPguI0+0cwPXXNLaXvGkAV6VFzb1l
2LSDCzJCgvfkrdH4cnaJAVfzOqbb+OsW4PUWRgJsXePWzg1eqO8BunJ5HYD/QGzK0qh80tgJ4Ekl
j+1WxohDD80uepP+Jd/57AQ6oQJSa0z+JszQCcHxUPFWaIAS/jID7jY2ObDp+gscBwzTErfIQ+5Z
/lg5QBJ3vOVnXWWpz/T4MvHiU6EFl39zVplL/Y/A7ZNf5lXfn7WaakKJat4W6CsSzfwQLJci8vl2
WVVDzCgVajR5zJW1uPk254OF81JpbSV0eqlMXjF+rQvWps4EEQeW8UpntArHyDHOrXKYhM1t6tN7
7g3/LpAv1s9xsxnDBpP64KesymI3n7dBUeW5khnAg8aZTZuBA14fM+5pUIzwxIMzXKlyrB9RNr0d
+BD1PdivJwetW65+r6bO/t9ruuUF8rLYPEIIodkrX3le1iaiDH3bLmHikD+9qnycul1sWevplzzu
ixsd+JDR034L3AiGtzL9cCFQZ8uzIwrpvqsX/PokW84+F7tPcWBAKLkZ3n2ix+PsI90jHNwP0hOX
feC0w9HZtO/1J+OEbFExoGQQotfm4qOY62kNAsmYEjb229XZ3NikKRnB9BXMSWi2Y1amR3l/g3Lj
IRw+8JVPQzMSTF+lupGDFiTwrGQ8POTANbRytzv2WOdl51nQde2YT1Gsy1SYvt7TC0+ikRZ7DaEU
14bnTO2831OIFQ7Igea9p+3klqmBPjZ9ARJqBO04MVdT62mPU6aHo7sOamRo3SjF28/hKdHjWegR
PuRwnQi/3858yGjSektdsgpKxBcCcYGO2bOggk4hfTn2mrd1JcIIVN8AkJcKyhk4LasgkDU4IZQX
IqLeIf3jzVvQNWHLpsoIrM1F0D+9GTjL09brrxt4FkVTcJWcQ1amfngZ9ZdplSPfVm2ZAv57ZC4z
TYvm6w0l1q/0M+GOmLfoyQ9YfXCqHfYEQoiG9JG52gT4NEMuFIHv580l3RwIJ8trtT19Un01GgGC
DISFgQxvwj3B82Qg0umqL8+RdOzRdl/2FljIg5kjC1+YZ24lXzzzFyOZtR14dfIsftPZIJXUFDt6
6rsnhyw7GKDMlio/wtleJgB9KAFtGzq0lcXJ4UewZlQSc2dn7E1yYdOIX+2nWiae2u4rLvz1ODFK
YKhnk4NYo2PXAaVhYlP9ug8aFpM9qtC9/BpFuGLil2j8T/9Z21z4lOLW7a4Asr0isj5lfRYaVIiq
NahgAQTsy24JQ2SNsR8yNd2WICs/KZpyAOMjq8I0Nvbw/9oQLXmXPExfHhIyyUVIIebN6hUazTkv
Brt4429b9K7OKy3fqOu4YfFDWWVtz/wPE4W/ZHtnP5Cd+o8vMpgP96aqkCi41x50eBGZXiOdtf7T
aBKp3/ugQdsrt9SK9I7BIVRhHO33QBM/oGq5O2ShnlFNiMUhUbdBLPDTBBzDvcX1oNRKmdeuAlFq
w//bBdnNG7LyOvEX68WHGtpA02Xkr6/EHaP1ploaLqkOo3ZcojDm5k6vErTIKOHK1eUJCzSlQNlR
a0v/Me8kk8FP8gO6pAh0nnFOPY0uRqygjco0ceLjXARYB6vB4rCH4htc47iV5BBR82UQk9QvyYY3
xxauxfsJs1CMfSOqKV2f903XhsCpdGakU9MbkjaV8XX6tHT6ji5s/3jkpb+xJX00choy/N9GWVMG
+ccmfes9WpheVHgnG8TBIolZcqOxaPPKz6E+Pxh+djMhWLlft0tvAXAr0hxWronDHysiVtzdsKoQ
N67GKwc8KGHT/xAWqQJr5x+ChK0BVbmwc+zAMYSxEONQTnxqMCs0Jh9T5F3GbzBmvbzg78QsRIKZ
tEsjYU4BnTzBFoGl5pjvkWXW96Cz9L9sx5KRaiYVUr2Oq93RatfY0XGk+w+i5J17GPnGuUuf+TZb
s+fzKcsg2cZD4tH6qUZeA/ZEfkroLjUN/+Vz/6PX4EiW9GBakYTbesxyqxP8gGq51c3ZbXknkC4s
uRBDj4sD66cwZ8TaovfeDD2gJ5lEVkNoacgFaAykPFDTw+7obvemJe4ZoEqEDPJPWTL03+ztm/Q9
9mRSVUNhBKtHaSm7X3h7k73JZVm6yoYiWUGARURXVnaMO+gLcAu8klspUuoXF9tbZnzwD/cgAaa+
A2HkcVlc6TpmDjfg/YEcT+LM5tFFjx39PtlkB5ZHh3ll1/1t624/sMwnujUF0Xortu9wQpxv56uX
4bcljaUI//LksJ8cx34ifw+6wHbDi7rbe1fq67HgCRxp/+gqgzGltJa+shyKq1s5ZcsvRlFkh3nR
N6Qt62Quy+ZNBsEKraEI3aX/rf9O1nqN2hfDVcW1qovyKak2Uxa+qHIT7kOtK+8k4X8wQx3qhsHP
z/J7LK29gMa0WsO5mIShd1TlV+rGPamHZg7m1aIzd3c3qc0AIDSci7W5HCxFRTEf/mJ3SyGgrJwy
xGSAlRHj6XPlsplD/orHOBclrr6yy4sv/DccP5cXzeUrtBoYBvtgmLLk67Wd7Sxlf+7Cm3UO4Qmw
hJDqBA++StN3GyPcwVD4wPR2mm3DV6V/pAJ1va8MttcXToweMDvL2F5wFj3N6a0cMm6ui9Za4V+t
cgeEWdlJaJq9sLw0adCzkFPiv+WuarZKqWq/4tUc0bRjVTiyT/oSL3wFs8JBbf6hDm/bXMrmCZuM
9gLvvwxMzHJ1/WaGiViohnpm+hvGn4RREDIXmuxPj5q3i8UjT1sv4ApludXnR7q/itWq/yUYKBBF
Q7dwPtDi/3tNr5bCYBlof4eJyOWjC2//NuxTKU8bjMx5b+eqIkaTiuFl6ZEW/mRPxTbTQ5S+A3UT
f/8gB2R+eP3G60Gr+yESIUHibOPu0MXBgApRq9DDgrF473ytFxF2M1Lu+FwmgLj7iVPbbL7Q/Awr
Tfkiy5Mak4PW+nlEjk9rlaANqhSJ6K87/j3v4Ap2nFluraCrhNV5v3+Krtfn+2ducVHf9jWbpX5C
8fULUbtb3sKTM1XWOrFRxRJVDxZwBBdTGsYAF+bUdJPY+AZ/mqmcBzF5i5aIHstX1TYDFDbUCZxs
en3DI9sKF17jU1T0v0p7SLAf9Zh0s/rCSEl7tgy/WBhMPcv4u2fjWea6xT5JETfghx19tJc7C/AW
bF6DVwQq2SDvI9C061ylCUGIJHpqD6O3IeEy8BBC+N/3q7JadmsjmNqq7Qm5ZUw2Wqp2c1uD4DsX
QgbW8FrWU3aVjBSIpTiW5DyPyNUsbpADbz+LvIv8V9lhqCFiEd+W+RyLP38CyBDNLtETTTrJMZiu
wcpalMmrZIcfT8Wfdy0zjFyAeeRW6XLHUIUJgtqHULIN4NXOGIAo+rSIoyqYCN+tw3VevRdvrtMf
7G8uDN4WI/pN6cSvrafIvMWVF8ofsR78bfXLoarnHeaNQTdIFEW9urGFqSU4F5rsaLyaFIxyjrGX
3dwnOwQiUEpYO74A3avqB7ISuRuZrPfprMI8e+6czyfddHSbV3OoRIJI58YhAnG3NECIce82P/9h
0Qm4KkoQeLrJRxqQ2EW1FSdL4cx+WxrtjduyosrlJCK+8qukVkOTqToDoVbRrNizCIjQ90DOG2FW
qyM1O04iZXO+bbJSztt7IllqmDOu9SqTe+VB5f1qUAijJiFQkXG2WJrbu9hSgsHXJaOFOSYHCTV8
oHNIdtRJJk+jB4VnyC92u5J/n8+p4kTJchTTwPuAXzQzJ1XeTp5r0EZEdSTGIVrDtC5AryzS62KF
XHcQhgXge4OzIoDEDMKi1EU0xdqC/L0Yza9jn1/eth7lMyidYecBZrts/DlJ5JZV1xx4D3+aqA6q
pUgMIjIRuBqJ2U4Ww9Y97+yINTkmd3TKCNRYl6mvEANmf0S3C+FlK1ptL3oitoXZaVF8GZwNlZjd
4tn6LDbc2svPv0oTr0acz9uoz+sKRhNLU7Vsa3WkFEfq1LN7Iiab1zgYXHe6iSvxpBJPdDWjug+F
+aMVWgmYrFC6gWjsDwiSWxyBwXqnns9ImMyO1lVSis+JJ+NJRMbCOPLBYRUNQIaRN9PRCIkkjFSo
VqJizP5tHDJlfRMFyioA1lAg4okvfYNfA2ph/ybQBj73aHs384/yLjbkTjZzfVtB6I57DmxUVSsX
NHptZO7LtHJacfM0DuuFtlcfrBI1na8yyYWeaxVBhH6g4+Fv9V+RBLIoGGFOAUN/jWkBn/uepk9h
ScpaMoUex/C6VNBCWdmTI0R0v7f+RYH3uTe3yjcuBcsoZqpRt1U+ExsXFlQgabKMQUWE0SeFqCVR
j7rILBtki60XmiWXZOQEe7OsCGlK61Jib29R2fIqbEiq1x8Mg5BsevKHioHZomH4t5wTrQoAPcSc
l2NVyD4Hlemygkkl0iHGoPhkda+Xbt0+t0q4QC5J7hO7HUvA1CV8EQ+fMcYNmPNnZOXEJVYjHPRR
VV+bKcMHpbHZeHnxTJdF7S9JbGIGdRxxzb6cd6NF6aerGnKBDcmvFvG+i7lK5CusHyKZZUaeepPC
Dnqtq8En1tHCXQrpJ8meHih9p8jiSdsyKfyRJomcSLY/l+oGyE8/9nrKlRLTNo4vlj8PWGRtPNQW
KYH8q3bKYy6LzDmjduW8z85DylF4kyBwVcuALqgu9CVckGUstpkJ1w65aYYeyjPNVlSHwOiKEgK2
K2Q2AnC3cwMSUluJxQcUcfA+GwSd7BNxaW+urkyXVrll+IHVAaFw8ufVQhyXDGH1FBcBC0YKQ2DM
von4JwXgs2VsX3H2WqgE/YuwIDmP9Z29jCcXnAvGeRI04MBRJFaqLDJyHFiGfaWoa9G4rf9I5W0Q
FeNQLxuwWqtPhK609soJhh9iEa5GfiHsUCaPoLWPh/aM2ZBdr8aL4ZqX2r+o7gd6iDPL4s/srxap
Rv2e9jVBt/HCqrj2zq473l/G+fOURbHCbH8yg6bej/KWXeLd2B9BIwMRul32Yp/gN/u/LPVjsb/M
FIKS3TND0b+RtxN54xrnntfoWU1K9gEf8zWLUuntBScwfAXrGdF9DaeKx+chEilAxMAdOoTNLxq5
aHm7mnYsI+E0daIzyXPBHlsI7iY6yxQNrauSB/Ihs1MvD4T3CxbNDKY28U1YZ2/of91GvCCCAcIe
PiUghrHmUyPc38o3hImCfA0v3x4MnFTTTEAu5fn2cePFhw1LXHLugi3CWXiFR/AoWREOHs0P5FL3
T3fLf/E9xtNkWGuM9yzamv+HUl8Qjc8SrSBLAUUV2L6taF6Acyzj+pwhnLE/N4r7wlnV9vKM2iUq
a0S0VV2PRgycvyEbiaGb/ZkERZTPLbBCqgdDbdQHfHg64uqL037jymc5DsO3U1eVc/4uDD/fM3FP
uAR/9lTjN/nUP4/TiW30t23ikvUNyNZIiRWJfdQtXJzcTSGRZGbIBTzvnWTmFS1hu9UccwicJ00N
sspS/i0P2bPAmQzYQqlVMsMTV3NdjcDonSaW9/imYIL0beK4IvIolTZArorl+uJMMJjawcRTJuxp
0zJaGRfPEbev4tBs55wOhGf0bq9bCA4ICWVFeJuBihD8W1tqtY1DvgbUH5kduTI0tGp3dwRIeMbx
15w5mTrGhhJez5Xvfk/5p1I+UrmRjNOpMWuoaCqIxF3DUO2kfouFvmGACIosdOCfYORZz9AHlwi9
+w9N/c/JGMdihAGu4fLg8wo90aOwk76VcqAoWCVvuYIt8dSu/LxQAgo0nu6zZZJxk5FuSE9qKqNb
1J8GGbd5AywlQj/brpzM6SJyyKoH3VGUGyovuNBctwkS2kWQOBQ5QczVvgFWVLlZxFAQN0R2cYgS
wujzsCXvamlnOpdWoPevRJyWMnFp/Ts4ptRc7iuOv76/cXTPKD+8NRl4q1SIcBk5PJapO1mL/vIQ
13da/96K3fjF4Oiq7VJjckC6iDLJevgUc1zs3RTQCLec4R5Vr/ukW+Z5oicTT/fPmCF+jfm0H/7/
Lis6NZsCjv9OWBKoMhOmKwYshy9Fi7Qp+PClsP+wJWohoUrv5HHs8AhtCoAdd0DDdKrByugs9bVN
GbLdIDIrd+jvTzfwomH4TYA3XuGM2+sz3X0XEvFCe9tLcdfHQiC+y6E4OwwK+N6np5QkPzutdPgh
ymw0nEuQh5zZ8YPuRbWBx2vofvtkqy1+ThObbTRxUlfwMsPCR9ydp2tkvSAhDYq6KPLkxNKEWZfH
QlTBBVx25ZJnts4L63NJNilZT4okFL0chkY4FH1nTfneQCbrUURz09KTYNe5SliLUcRzB5gmuliF
BTJSYM0xuQMEBmkyKZbuVVOyqZmNZr1zD33VDIqDO8jPfmLlXSN/MlKDKxrmTqe7vNeNODs/766V
/NYzz7F2f4Ab8EogDYKwYwukbNs+fU6N7pg4uuhrE9BXgAn9bYr9j3HmPGuw7D/EZkYT/HBd8MbR
tsl2jWHKhZqiZxOf4TGI3itC9zazr9pHwRo6eApBueNJfvLpEZR0BcdGbyvXq/kn9r47EfPBSuBU
VkKBfuPLSF76y+FlEnmFI5ZMPCu5Ppd2AcCdnbVTFHB2dO+pPQwEWAg6tRoY+QEG2x6CKVWGhD/x
rP+RpwrR/9QDJPXCncNCgOpH2u8hTt8k8vUypcVmXBEXYZ3JgUln9g/H9wNJmjVfRSgNtO+fp97r
H97m/EMMKYrT8WgX0RdOxk/yhVuSIkXhv6PSdk7oDLjTl0ryPTYGLpEK0Ybk+XoQQ1kwb/mSOvXS
uNZBr1FC6b8QffuLnn+jV9ZIzjW8Xqen2eSLZboYtUyxEW2vDtVPlqMgWLojbFjg62UENdf4iEd0
FabSfEgKHGy3b8bhfrRS1XvLd2aD6Mo8yBzOgxISqYf2LItMsNMfZiSy99ESrjSb9GIA40vEvwqm
SchHQt5ibJNOKctpJXBlmEeFY5Q2Xfd4pGM32NBSSK/ePvrGPdpN0ygjLDLETHQCqWEV51Eu5EMJ
CO3waHN8kAVOEx847XJPIzR8tTpY/IqY1/Swia7RC37a/+8XIvESKNVqqT0kRdSEq09CKfOFjDze
oR5+uWI7U6zZuVyXgKEBmaxqdJ1XNogn0I7iyS7hMqkpyN0gOES29j4apMWbusVGDaq68rL5S4yl
BW1rKm6WDEhCEOREejLXmKtx42f5SW5now+fEXDiJcmxW49B+JTbZgiIZuDe8C/p8eEPA8z+/C7Q
vMgeI2Qm18BHKHbji0nQ3F8tuwKw2HwH0WOkPSN81j1MvdkEkiS4hvrBQY1lHUIxwmWdhMWzqZCy
/7W1hR1RyoAfKcL0fPJ8SbP6Gzuonn8PDhiUuP2rRFJmKgDhmeus6n20YCpxvjCf2xuXGpcoPzae
Mk++/RItqfdHjTy48ndcYNdUUCG6r5lXq7lW3LxGYAchUqFvmfuAO9hdNlD4iKhqqJMf0eUoWjVF
eEZdiZHGf/cYw0B7otTvnHPTiPv/98Fp3Uypv2TItEr2GEwXf1ns6C6XZzxKze+Y+cPEomQk637Q
WghdExuXMlJrNdXOWT5aBfOInW3KK6PJapdEKYdIIlR/wLGdwHs14UkOzJ8pD6DZiF+JL42gjx0F
/s8E0QWze19kLglGvhkeN6jbCPcTx4ugXPj0KU7DgNop5/J3/Hgg2mM78Q03XuOpAyaJLVoyzhC4
wQPh7wfdHaP60on+Ol2JmXVkCPGozzcSa74VvIx1tTm3pZIEmT0Mnwpx1KRZzSxpzfoctzm9R5Pf
NMpPSrrFvY/2FXiZy4xLbBJPJGWtcMhT7mhI/saprog4xdP6FkUpeFQbEf330ugL28R8raH34Hr9
aQ2CsW2X3nIavG9PuOyIrohGQE5I9fVFby2Vw1FkyWGJfzWanqgc6FtW3aICr3BH8xZvhbY8qxqm
sXfvprEefNjcak5d4XO8dirRcWs2Xzh2fM6L3e1ItehSmUTuBjUYCVQBQPU9LhYEZNkWqD0MfMXs
KFJ0peKt6jlwGwuHqb2hxagx6vRfVObY5n4NsEFnxQG450+fPzajAR6D6FU3GWbfGqv1TmCP5PIh
B90Zj5vhlTmWVy8fi8yUsy3GQRTuaydscUz/FJ6KZhbiXLTcsdVJAJGviMrSAGBvY9Y++TMOCg+v
zGTPlIqJKaf5NRI5HdZ1WIHnOI1O/0UjfuiX2DFHamb4WEkEGY4XhEsU2pWoDA7ikQFNA+ce92Bp
l8N6wyi1PicY2nHqj/rhsYoCtBs3GxHlRnMl73vMbemtrEMsD+SkhU9fuFWyDxTWTJNINAG3joeF
f/ffgpQOWtbO9HUlYeRmEp9k01C02JMxfQ8mZMgBYFEK9N9hGbi/XpqWsH9bcBzvtiZis4Bwsul3
Eu+9S/G/gw3i6WG6KQ3QFt9jwcOqU4EO4LGPbJGt7z+Mni69OD5KkMugcd5N3uNKp7QJZHd2k0pC
NwrDN1TVc1g+nLbJZfgdcIgIWZCXcj7/3mRnFFqdUpfMV9Vvv5XRxTZ0PURkB/vyeRclCjWe9Ffh
nn39q5KoinC4q8Ujy0UB0n6CHpU8zMLDjngnfDdyCBhhN1QGIn0MFpAcuBDOw6lSM3wPvDLun3/T
IplnEYAGr5W5tONpJ9VC/zt45kjMZQsb8ffU84B0nBq6z+/C1CIKYRJSDIYj8ejDoUEg6R6v11+y
eL3XxiJi6MIz320Es/gc9aEQqHfc8aUK3p4koUAYmfVmaMAWM93EAMq106UmDfKKg8tvK9fe5otD
wG3keIWGeB1hgzsoBXVhQ5LJb/lIgsORm+VYVQ/cBYo8HYIAjL/eUD8QPX2BrbI+nfxx0bg8j0N5
M1KiIfD4Al2Il4JIPZpC/0Bhqri+FvPRxKH09ajjswyqYYDm9lvubezAVb1oZWcFwQsafAAdoMmI
1+YpEPE5yxZuPHv1awANqZWxbcFUznLuZhG/DNXPLEozUeUPhICx/imjkv7+mOmU85KctqhZQd7G
yFBMEOjkz0dK9yN2xHrxWSgthXTT9WROqK7Fh9eoPONX8wPjo9L0LeW+V14wqB1BjX+WZrRJXUOM
pDe29xlHDOZstRJovWfoU9x71WSSc6Fy5ck2ASljNMSCjM5+37podufN1J6hvz8PJ5E2egfHwIwy
e0y/gxVsrHzjJf7QhEU4VnN7WGLjEmVpHEjGwWmvZRC9xW4t4K0PD0HkzSX5YY3961+oHQNt0qiS
c5ACf4weFWrtTBxBYqhTaTy4whhtDSnIaYww5zMHVvE5LgRLuikioFguM21StcaMfCsS/RRNwWEk
VAK9RisyNyyYNFmj73mii3PhYFI1Hj1Cqg6WavaISY95QKqpukTpGL2R7YOcxy+/g4eVRXZoj0fc
S3akQOdtZNu8B7WRgZ/tGeLfkkR2fHmz2BYphpzj8rpgIzxkyx/PUdT6WJduyrCMTXRCT47fYBRf
QbaLJ7t15GNB3GGBWJpiH+pjE9etLuuJxqaaLJMCzlffAwd2Uy9xQ9OXqCkGOeKC3TIaWoqdjFVm
EmsGP6DYhVEx3IbTNfTE7wpmU8+zW4qo15R7NmaCbAhaZcCrB5vsrJpxShvBPSZTOsFFny/iHxTw
x2gaYBeVjW+7jvsBx5yvb8krq/dnfTnBUQsTxvYAzVD2Cjo8o4T9MgJCi9B7XuLzBpma1DlqCrQb
SbKzPK1nF0UIKFfl3mZY2hUr/YWYTVj2NmGcT5MzhMNiQHesiRPeAOsNUWbnP1GQk2K++D2fS0F2
iyekDIRahj73MXV5Y7G2BWhp/W52gOmNn1SZGofyB3GzB+oO/ts5livFG5wA35ATn/q+uvi8Ph9v
9qLi+SKyrrddDKd0dgyBL8LGI9lAYxd08ttZjAC5YnZGlurrEDqGiMf6KkNwbxwxSJjv6dRlKGX6
U37uNeqKt3y3BZgES9xjDhLaufKftk/jH2LzZ6nlxDVg+2+V8ToO20U7etrROhILt7V3uBO+5Mun
/g7WygT3f6zpmiEge3OTo1r6+zkx2mmo05r1/mgFjYxiMQJpUoB7KpQjVXTivgJzQpygS/49+jEo
kte2oqwj5PdHtumWmsm7PeaC3XVKyBOoeLambbpOTTykj5sswRSXQJdfPAYd2N/qJbkheKExezxi
AvzdCE0P80NJN8cFKMPguh00eW8FuKycOzigPR//ItP5PJ2lv+XvTgX9x1Qf3g/Q26FPo3SAxINF
QVBoIMYGSJCJoh59RNv3IkQaUIcfs5XcdS404OGVJglPJLvrz6JAUL8MN7auJZ1g9LQ3oJUZepxL
5z+3CqPkUuZJmlRIfwDQFKKnI1NUWqKE0Ud7u4++sxbxWEzOH2rnp/7SbVurqptlN14IJUOIK7B+
4Xv513J1p17yv5aMJxI6t882op9duLkJ7rFz8B+D7AEbDIMIGwOjcQIiOXY4OS7hM73bymOncgoj
dns54u29y/Pjb4TFjlHbLVxJaWrkxUmQO3yOL8U/WcBKtZwAWflAQMcz3OS8zb+sCXwACGhkR4v5
LWQLnV/UMFPhplyyMO3glnLbovAwTjVq2Amnbu1jsn1MYvfElWMiv682Cvt763irIjJlIndycEtO
6AIFKDC9D6uA69l9Qw7Rv1oXalZmoFAYWcoDl0AqGLcrGSHohjo5VVSrx/F/WG7147L2ztctnehs
QNss9j7oJ64yEXeHkUZR6ZD4Qb6yNFetkiVuaHB26tGS+gBzZIUO3xamaTlXy4nVfZpjbuYMNbyi
L505Gqv00Ef15ShE1cc+TzT668KgClCuBEt9qxSCif9EPoTstdUAzyEDYn052xrcy9P7JJkpAXVI
vKt9++p3je7tLCcIvUqdEn2XPgVpwzqryn+Mihu7JSHxpAR9DLcUjZhA0QoEumqSKHjJEpEbpS9k
JbWy5aTKp1W4KtWEz8IIH4gjQLje62Voot6s5LlXjETXD5xwbaOnnFcWKH8HU7ZDbKhSzgTlhH1u
M8C7Bq35vc7sa7WzQOneOL4bGFGdcfVOp7murc4NL2ud7GHFsJ4K72dC0PaKRHYQLRA+3DpeNGh2
vNSz/mWrPH+jKiABeviY6tt9zOfSZvz8NAl92IH+k11OliYuowTLvdNb1xTFIuaKQzyST05jAzK+
mXWkyFeHabi3eWoVhksvTyafOs+rvuBP1CInxb3j7EQZk0D57Whfz3Jsq298XPPK5IlueLQ84n2y
5+3p6utQvyuhsBgxbuLfYaYCZeKvVwMJdHgd4oC2X07HF9z3M4u645q08GRUuCei0vkcoocPfZsZ
UaKsY1yvf1z1QeSTBZD3w2Hqjj8PsCPnKzbJdwDUJYT/Myh77o12MVILsyKM1AQYP+8eAUWOjo9Q
EGiQXwYNH4PRFVkxs6oin82xlOngKzcJbDz+/fqdA0CBgon+apn0XCC40e8Debw1NedPb3zAHu0r
p7LYvGLlbvMJO6t7zc0HWyj+pHjABRjnAuxCk3LIzw5xZTraZDI7MVGDIpVVz7Y+cx3j/xv+69YD
kuDvgL/JVk/p7WQCgAtuOnMjcDZQ0fSDqAZ24My6dk8itcGqSczhFJ4vKH14qrBuBd+CoFLlX2Q1
AF0GLrCa0U0sDS/iGGPwhj5z7Wo0KTqkOJEyw32KldTufyKLpTcAPfOUP+vuQdOAUYdW+dJG11Uq
Vh+TJhmPD3lQuVWsl/3imKUWW5bHW2OzcIXYWJFkQ/NcCBisiqAXEWNXCdqf18ePiMEFkrC+iqcW
YdGh8tYUh2IGdf3cD3iAZ/oCNoRqViraro65eudQf0wQTTJi3VZillhsBUDYoeawHrNRapd1GRk9
NCDqTjS3Ud6enbGNWl9OQCynilD6wvlK3ys2OKyp1mQHQgqpHsxfSuBBerdH+L/N8G/fW4TUW/gM
OkRbZpB0QRtSybu/fyPAvIy5N+B1NLcOs1B4qdNg2lh5HUTA5zxQoKa0BNQ2uUh6/ilMOupMQoqQ
qcl30rPsXMMLvciwyZk8ZpTA8dplCFiJIPzHgEmkCPJSHOz7DHVzv8Xg0RaGX7NIr4WYMu329g2j
Un8lhc330p2E8DS1op5sjTUDwPa7vXk+z8uCTJK2gQvMea1/EwBeZfbYbul2lFOSKb0AqG9zaX4S
tYdbpjIUGcUzMhYqisOcqwf7Ke1olLrG5eq83aBKk1HvMiQt81DKw1uMtEGVFfr45QxhkcNcZd5R
SKjq1aKVbthqZzGTTRO/e2ml5bs7HA/LU34ch4A8gPPDbrcNdWQblcKAQdb1F6mR7hstFkTzKn4w
dGdvA9/7TwqMOAirlmFnTSJmXBtaJGyPhCWZYrRHe7DHuUXFDEm35NN/12oR2MfAN0uhf940z0F6
SxEjKnikdxzlvrltamTF6pElhKZzMMLFWHTACmP8W++VT6FfVEhOsHgfZIsPTuEO/j1NRZRNHeRo
GR5T0tWLIe1KQoIZlaMFXdl80F9ZO3WfXoJcWfOdgQ8lTqdj3csiVw7s2Qy2E8cYo7uIhuZS6F7x
Vs2GaCWLGJJOUb1C9z4LByS6NwFBg7R+sF6hKhSmrGAi4xA5M+nSIO6y1aSdAp76b7XeeDwKmbV2
OUQLcGJFWiIaGzLZ1Kn562ZsFKlOH1lFiCdMrIF+KAk7RTTwrIiLyWlezwV81kBaxfS8WSskcFcA
G1rVa9yceEcf8tu2hnbOz9eHHo0uchTQUDADWCFd1r2a+kRUS0dYV93PX9Jr2mOgor7bia+1YzO1
/QNmQVE89igNhuqqRjNnUTXYP9vgqpHoAUPFLxRZWvLHWewi1VHCh3OxTCE6Ykgqomjm9K8LRVmv
ibkxyFYQADs9ySoyUOJaUxxMwf2zNEp2ElpAkXRss4p5lSNpLv3ZGRZ4fJgxSlQTbjbhiyx7O7on
ljy6c63Yy8MOcx3mXXkwvdfj1QLXQitT2uIKtb2QTzeZXwEUy1B/qfN7FgmCBWR+bhYr7L5dxeNr
WLp4EbO5ExQw/87tQy9QaRMvepzU8bRXI1a2HxRGz7nZgmKwptMPd+ivrTb/nDsuV6jRv/YTFZOH
S5jlBYDtR2NHTcvncSIyOqH4x5/cvJ4DwM5XGd2C9jlD9bZrHuk6epWwx9gPyfvs+L+65UHWxdzF
tHxYqztaISK9g7XYRvVllhZ/ewZLOx8XguO9OG40Pm4TxT6tHQ7/mqGEcJJwrNujKwhD8Ndpmvo6
miT/QSF7JMW2qrqJ5wdV9/Tc88cXpR4tW7USynXncMsAYbMNuLkzhvVlZtvgYTtVbqqE8cZp8ozH
YCjaM1aprMwrEdGJzlaTvS68sP2xmBL1z1lhjqoim6Axgu+Sfg2no4xzxEIVEuhadHMBFk0pt3j8
f3pp/0y1A1/h6H9SchgNDbvWzhpN2fG8c3aYbIVnciLFLF4rgCsHc4fjHN1/LEfWMaB8rff88Mpl
vWbq17KCzUIxbdOr9J+IyV8EDGML2Y2TppfQqG5EJpSp41ObwaW0Mghp2t7DqxI5kMnAhggm/Wbj
Wz9cmqvTn30Q13IIEI2ZJIU86gTc11c6fdHqqyvSvYyPXqBgou+HyUz62XStVdjpTZN0kTtmr+39
HXhC6Bku/cJEQC4nIJy1y8UAMa2BZ7L8E9Cu/zTi5IwH2x8+dsLeOinnyDMY/5wqKcpWPfxPnsxF
wwx7rUPUpH0unUE/lXdzgsjdbRtcXvf262dfpBMXuaZ2Jm6EwlA6v2nhGjqocmp4MA01M+76/mnK
SVZxohIq3JN75o+hSMJKO1zH5k1tF1Yds/HQfDs+CAlx24UFVXOc7E5joOI29OPb6Ho9YhXLg9YP
ypkJnq8JScLr9TkTsGT/fWf+kJ8jHzkcavIF6e8TIxgRrQh5QRYv2gEs8WEv4lF2rQaBtxHSQUcR
en52dykPA5EbMFfaldf63gx4ypKLgkg78gu+EPGMy6Od3vgnlQOGu4Rbhb3MWqIMMs/zE9SvfoIY
CR4/SLQQInMj6OMQs7TStdxBmYygUCSvFtCJPQz4VhJNliDS9fyx9RGgET2QieyEmVW9y/mwB+Xg
r0QgcepRHc5bfS2dR5R5XYrumFRm6j3izrj5Em1iAc4Z8jlEHvdG8gGL3WH+vq96zVbF1b0nE7x9
/EZS16ptp78cwEesUH0PpxsS0xnHxrbCeuTDWew0+96md91Rs8HZSv70EBCiZn9YVByclXPCxEXo
ibAXsW2tkeaJVfWJw2ysxLj1iFqHcCtA1hdQwgVERWD4EKVppZlLYwd4M+kjpUvIqJbp9LC7Mmwq
MPGtXpi3WVBzHo9iiOpVHUTZTnglVpNHsXLOR/jO4BVOasXoYdt68mxViRZwrjlAa/dv/jfAXJLC
UC3PrC5Hc41c/pz+PsJu8cHLhheRyfIxkGYkBWEuTHqKohTMTOBfVpBbXH2CbiGWBshgDOrjTnT/
5VUO0zkKzNUnKhchpNBNuTaf6ulPZhQbTqjljJkAK6HM1FA8m3TyVxMtMMDG068EjIm1aorNvxeD
Vs/29Cclmah3wW6IH7rrBdV+IgQK4geyi2v0uke1ToEAPvPAfXZOvrhtug1irUItpueVAu0nT2d8
/n7AVFZZLpaCimkAvUpigahf/lyH4sndQT2CwR718RWr1xJkUQ/yP0WD6Q0icpTwDPe8MY++JAud
7+mQ6nHtypDcccAoRfdi7QXm9t+kaJYyeG16pkGXx5QLF84Yb2gJKt8sa5mF0kfNnw2MqryTr56n
Mkg00Jq6TEN8QshVknBh14wnfWvSDm2hAToQo63hhNznGrKfZB5UcldJsHCBgjA8FhF8Sj/RlEbv
PATg5ssyT5aQNlez9NZ8GEbU31lo4E577GxH6zxhGVmCYuRQoTlSwLizdxH02GF2CsHnmAFzeX7O
kKSwCP/EXW6Osnul59EneTzj+8y/ZtS/NqC6YqgMqA4EzE9we5PMNqONIqCdZVVW9+Taf0QJuK0X
akmZIbZ3CbX4SsSfGA2jgHXsKNhq2njxt2FX16KdlT6jN0sW+rfABq/XI9pR6o9a1Tp4c3fpQ+ol
Bs1PFBea3xxlBoBwycum5Pe8ZD1coCiW9MqFiG50eY+DSK1HMQBO6u/qHmKwPgpze/UDRk5VepdY
XmjUyGEprHC9g1W8sIDwuDPn0b0ObeXTp8f/H+1h8BIdNbOmLhDB9rKDvY9rWP/cT79FquuqBfdQ
ufpkbMoWL3Gd0AHZVrSEbBtqFsgUHr/xsTy4vjxZ+tkKSVlSRMKXPhAB+oPxOhvIabvxIAlSLhh9
sCskJ8gqYRVDzEtR2EtD3YvAQIUzksekvQQncmzpVc5+yAypv7l9zt0cQQbeQrxsoaO5xTcgzog+
ajAUdXzLrftxLpz6HGCK9bDiBuiPgURFJDKGSTJRgxNRBSbFCHQPjkzv5Yzv7hmi1wZUCEttAmQ0
+YmKd1rGOyHCDRmLfZ1CneXSxUlyMbjpv/i7nUWMXZttrzwbM1IRT0qxzUYIUzSjAp77tMb8txhB
bQaWU7TN1uQtzG7MpvNbVXGlkB9yusEmFIX2n8cYHD+ivp0vu7RdNxN5JI1mDZ9vAwt4V4gBjzGF
85xM0BmviqFplY1Kw1pMgC5qvRypXRC4XJ/7uLfs6G3VmtXGRdL6zdmBMqH0CIuTE18FMBXELf1F
hU9LZv2E8fbSkyqkRG0E9SXY4oqTJjsFO8uesNCpE4l8I6iFqiwAgL/5dcTefD3qDwg2/e52Wydv
jU8A+w7EST2JNow/dgMxmlaY8w7N67Ps+59bo1Eq1ivxXAAzGHJK5N5t3B+lbNaGXbi1Puk/yZFz
vq2Rn5p7izRTNONtj8lK0BZkNlNNlh6S7OEiBIu0GoCeJgQaGeGxZLJAjKq2K1VYzyG+MfImEfTF
pCnSr60NQgD/Wh83PFt0cmNvSew/g3An1/YjLWrrvt/O3vn2p6BFqayqPZCAu6XJSlzrFc9OmZzL
jFSk3oAppYofU0hSeKvU560Ab34UhPy7R7uXj8E1kobnjyxQ77c2iGjQrL2U+Tv5Kz2tXh/SHRHW
IAB009Rj00ufIpubggKSCVA7UXDCngS9wmzFfFnVPxePMVFY+mrJFLRxwBUT7IicpKC0daUP2f2Z
G/xpk2A0TVN/3o1/ifuXr/9XXapaDMc+eERWLh1HfOoxwoxOiTbwTh5B2Gg1O8r2Q5vL2xPrconf
kaoKjpi0DWSiuLR4V+umMesIZ62L8kJPuAaf007UGTvJErVwMOioaLZWMDNQu5vvK1zZdxVuGdN9
Q02T4za8IqFukYa03GYagNzZxvpXONQkeF06ivs0xqQy17TyYI3Xoeogj85GqHZnOWU0FUSCH3f7
3ATiLRRsPzgvd4CZjLoJIN9xO3cAgKvGP+F9/h752JRoGKmVuKYqS+AL9ojNkjtxNgleuKbVKX5w
MuUS1athZ6THp3mkltQ/n9CYtBnZk9crVpyZ7AQyw4/A1ULDOrOH0//O54HYTvRhrKqlZ7iIE/9o
Eo1820CJNYz3Efxqz7poG1w5wAS6at7WFxVrXMcwpJQLztKj1UvBHS6+jFdFuTrWQE2m3pMbIYRz
CfLhA4KIFoHnUo8jr8MBscTWKuQ8k9cAEtqtlhX1bp5k5Rj9ONKoiADwJnUiS1bfKPTRdvpo+8II
qc5O4zDWSt97fIYd2K9HVfq3vhIPQ3r5Gd3lYZF7LaiKLOjoQ+Ju7ztAeqjuhh+Gg3Rg5lbPdUBh
9WEmnnL/uCRdC0NpTpB4RD4IDp9WQMsWXUEHj/8Z1bdrui6v7cgA3Jw/lvK5KqMae1KlLcqvQlfZ
rly2mILV76odrgLODrdP7ags+hVUrVs0gFsfyFLUOEjY60CT5CfpCU3JXzso7JE5IiKrT/Xj/XyR
w26i4+oXfk+C1k2SkfCofcWk2H5uZb9nM2OLS4U1yeMhy8tBXbWteZUZYMlsZ7k+sg4BtNUPae4a
VUHrBfaFoQ+ZzI0NQ9xkDrHZx17d33IiAzVojtn+FYty1LWXQTTLm9M+95fX0iMIRTg7/5FsJWvm
EGVykN2OyyOdvu/XmMK4rXMFv5aaDABXEmazrbZEAgV31sRnCGmPFFEUGP6JS579jqfuxbuE4Dgx
tKB6QjDU0GwSvrG0MrwXVmFpVOevWYwsMu0MTsekEiRQ8ov4H4Q+6FvXVv5TYjv253rf/R+lcAQ3
MWyn9/kY7PhTqSllznAorzsEYtPZTPNKFA3jNnQai1nFt37Tpi+xR1mYCW6fRHAg4w21H5oYkxTH
MuYSB1r9etambLYFHoKxgDB00tnZFViLiyCPpttCb/6U1EB9eSskwlWWsM1tj4+DsEt31cZ9ioom
Yey4/0HCj0ZT2s+B+chfUpjLq+TKSXcJqvZx6paSeiy5x1LcdOs79nb3G+gPRcAge3xLLNfNg9Qj
mqpeaXcerV8RGxgcAsWQsMb7CPi61LxGALRtdgewM/gKdBQ2OxuMgOMutkZgb6B0WKlMBitJtYWY
ZKxY3bFAaDF+1DaK+OqUQKdzoWgvdiAfNUWRNbo9eVJayzV2RM5S+snjZJMXqBY9w8akG7Nb4H0D
BvOMAQPw249VMrj9fZvHiExpZON9TKpJdsHSXjiHabmSB9QYiSiinMXqHcI43ex5nQfSwvZaNUdd
g+JOA5Psu7LyvF5csW5VguMSPG27dlz3osk44vJXmq7Qr4mL2BpFEf5Ephng6jFN+yLzGLDzKttJ
0jQohxIjNj8Z7Tbp5j3KszMzj6DN9qp295QSNmCm0d+gBOmzcrpbWIxtbmAJabfrMCB8UpTZPeZz
uhpPYZ5HSH/oCcO4gXnK89C7flHludNsCBGdXeM8BbWEaXZtJWH2cwfExqTpEZGDK5B8Q5VTPKWd
6u7yEB5yLqd6s+AA93sv7IXiwfnbHvG1vQjFDvlACucm0WfrX6ca9C6qUgqrzRGBCCVocMdoyQXG
LtCoCx190ne5MT9lhcbN8TmJQYBlTDOcz/AJhyAwt2zA72J676xFwGC2LfIwGVhIjuO4ekYdbcIi
brEFjn8ZQPkVgrYFnQChgef6KSek5WxiOtrRgfSjvojDOGF1TDbrF0cmA5aqgBl23PYUgE3YCGPO
RfqrW2P+SdSR9AeisacstbftAnsXsZnh1pWvc6fWb2YUwrE7Yu9oVXzaQlUMToyCoNu1RUjAJB0b
X4NmIwbkUiLn7sNlFKbAop+virK4D2yu+zEL5j1SKsCABBI0REkyYteR2du6K1O1fBJmw0v0pOvh
0NV55FI6dYD5RgVpyM5m7xxgSOr9smX/XlFEBe5MMpxRLiMBaS6JzHlNyeVnfQXc9ceW0Kox/4rT
s4iMwesYw9oJbQBBYJN5+83w4nR77U5/4lPwPejCJO+7+o0V/Sc7UOoo6sM9bJ8ujkhlTfnQEBNJ
jEFLZVN5/sH4zScDBdXEjVqFqt9nCWFcY6ynodzQa6uOpsZHXc7QV0yH2Zd29ThSdNAiOj5iBlS3
Hf+SWQxJ44LN6Q/I7ve8eddFKvrS4DsbLhReacOe2yzJMjODWy4fg20bsc9FnwU+yZgx04465CD9
XzaFquEWWSDmMbA5tHDO2c852eTjyK3+pcgHstwH4SAlP6tP7ICUlqhuLFPYleaADqz1uzG7Fldv
e/ZASHGOainFJweuc5LB9rUj5roUnxnsXOVOG/dJ9ZKEyrD19dSD22Nuui1PYtiriwr81mXK9oX1
UzYbqRW6FjJEZy9p3O++4YXLyIUbYVXqEPJTwEHs7FnsgM4fRR/6VhJYgDmrHus0JNsppiW5pxgN
7iMrqlpS6w5iRPeEFy2jnpaPp0VOu8TJJCVSPRTqG27G7cYtDIfJurFPCCjvRmD3XfZLovSu4Swo
KoBECJFo1PvlexpHAy82UwVtp+K7ZYj17LNVHL7NC3Tp1Pi0soHT/xwQ5gsPjcBvM8PFVndhycSB
r0k0MApJpEgXUD7lED0sYdzbhvXzZdtKEFisfk20tzDDWZkEux050jt158mE+JtZJ/gZdaoW6esD
u+/kACz1FP1iSlWZXjxKKJx8dYSxCFnJajoIwMX5eqkkYoLfkt81sMts3+UYVJDWlLXZYaPhaZXn
jZxKDU4ZExPay9/FPKAj8QM4WR0jYGCf3g2yccPrPXzLxQaal9+F56fbaNE8BDb1O40sb5FA1JOU
P0Do831WrK9gvou1NaByki1U+Yjdmam/dDmgCpnPUKHM4Vzci/VCCWN2xlB70+ZpDgoXzLhjnMFW
LCdPAJ7xUbHaBcZbLBZeQAM7cFd9arbUVDwS+VSlLd2LuYW6wJUdOFmg2Ec+dqu6q2Kjg7lilMk3
SiYoS7iD88KzoevlkuON826WEKem+TPFh1NGDJbh5yRWH1Cx+p+olMxiZqD62sUWDqiLU+SYEab2
Mn+X8onyhEnPrybPchSvNAhkXjYeroRx7O3A+xkWIEm8amRxM8LrDUb11lo0Qhoy4NYQQmfT0SCZ
Ou188cGpH0UwJLED5BwtIl79sA1xFa+22eGbVGRWso1Z3+Q3DPuQm21wACCD1QfYKGVluJFO0TTF
z5RSnqGkbOT2tqmLLwr2JzJd+ofSxm6k/s70HRhPW/wC3PCBDppi3Fga+FuqACwvzkXu01UMKsX3
beMtF9wa+1W0ZrwmFKti2u3ZTrK5nMimcTCxTDl61Wt0Wavb10nAEfUE95js+iR+NkOZ0+I/CXKI
Mk2nNfmOJ1A1oUyCUjzAG/sI7jI4zTLYXe+G3VzV/Gg18sx9mgBirjgDjJNfwzaSuUXjR1hShg3X
s/tZygPpZ5ofRPYZ0LXFU8P5XYj8C0iJWaPWa3vEUWUoNGpo+QbB7ZxWoSFDi/k4nXYNyWMrF+5n
Cj8xEXybKRRh18OhAJaJS0oKK6ho0BwwTNuTGnwwpyIwKjscmMauluEgdlzEKZm5uw9HOMlYgc8k
Y+NZBtTC1Fs34GEe0+QQ8pJ7wB9PFK43J5HhTh0eFFpUVWJcGfhm8oDcqazNVcD92V0S3ezdCznq
SP/AM5DXknn5bkPZK3/JrqeyE6cwhmaW6qsTSPvqlmH+2WuTjOAypgrVqc739NCxm2EuHXXwWD5W
BbKA3uKuwZCVrYoLGH97BirOljhaWa5z6d+UtHBhZFhnUDixmmsepou3GgLD9Uy5P6+im6BXLvmB
n4J3xOzJOhl/GU2WHiIpn2r8pBh/9l9w0EGDVGJ7xYnZP/8XwjuGU1Q0YpRWScRX6WtHqR09plip
3bDzf0aRoP/XAH1VOERqCsMj5Zlid25YRvQwLisLa4OAcYvMUGpkdYoRGCa8JeWP3Pbl4joJj6b/
VvnP9lgmFl2MKi3oHVbgtzgVZIDYhmhWcAWakFNx8bQnOqof9yGpMvxk3KU51ORuYVeG0Q7G0HV7
X22cUatr8L1jEEnAq1tCINaxseVpVZ+gTe525Tx0MkYXkoZ//sgYq1GP9buZlNbf+jXtIIpiOC1S
CCcdChlrlDXyD8wde0TCLyQBZ3knYsgDJ+ToOxVAQRh2sDRfkI3l5LSsD0+zfq8THHH92fjGjemZ
0fTDMI5X6KY9PXP/d51TADWrU2mI0gur+LjxoRHUDxsoC4bz3j9xkxJCmb8/h/QTgLEFxS8fvjSK
PYNb+/TKRf4T8GbTM7Rt0vu+qUJK47aFLm2ko2MYMLQsGABIeADIn8oREX4fqx3vCWBRD3v5ngcg
WQ97gDi7Tt9UIw7CyplN/eLhBfw+W5+ZVL19B0arTOOtwIE0rUirEIOLEe5UArtkiu9CPaAaIzOf
68aq6zgifKoAbYnKTHoSvh6X9ZIL8lK2oV89PmottRcOgKDYeRrx+sOr7vx2WSu4mlSZ9PB3Czfx
OSakurFO/uk1poXHRYtLEthjKCIkk6uDCZOdKR1ETLpF9Hu6b6eFLdNW2rnHwgaN/y3PyXOcSZVx
kd7GLiiyHfM3+yTcml95uBddPxU6SC5DEQ9sYr4wofBIjvRPj2YeYFCVyscOWrOzmH8fYt0ndmim
59WbRtCxijrcjPvqg9NcQSf5oNTBmoavz/5Yv9MUVZ4O0NUnFuBU/8o/5SlTEFryIz93QbZRfD5g
J+LzMKzGbsArhda9UR1emO30OedUkQtcCmR9efnGuo0P/ruDzCDpalRvD8mlFAQ49P4USoSDss/6
1b5ewq/cAY5vffPb0IAuWh8l0shs5FvYM+G1iz9JC7luC1Bcc82juBXISfb29j2S0rWg6feP96jB
mGFtU7mopq3M0Ly7tYXnuonuaZG8PqESIsn+Pj/Q55IZoMpotKou80uPyFQlXrA7XB2rXhEayZ2r
eOVn/IX6yl9TQ4mHuL9UmzdN+cktqnoPtaueG1imuRdtS3I1AIwwv1+eopzgp3/19cuis/JByDh3
ZmhNbHgagluVp+WP0bgpA7sfhB5lGuU4P7xIE54JCjDjWpq0vJYxY8U27SdJKJczkXFPak8s7fhM
CjwRO2MFtaov4aKs681qdifLsAHkeF5V6NARktEZzDVbiCEpLIcgVONULkrgU5e5e2FJekHdI09Z
6gXYaBesbRlJQPfFEbk7F4JM+rhacwtpjmmBF1hq845Vq1HuoSCsobsh7xDyj5uOk12m05RqeP4t
Tq1KMyi01mo3V+JVNcp348MKWCSNBQ09rStU5KdX96v1+cSVbg+1wE00Q/CBhNOuW9X3g1rgnhDU
+nMos5xyL3pzx98mGCczBXGQ0IgpgECnzYv9XOi69Y5krbVYCpC4gwdjVP9vTCSIrz/lOLYAYP7d
Ldl1ZNAFiIAR8kcrWRtqZ6JgcIyO40tZFXdInaPOzPS3vhqYwob9naNLt1NME2ufa9k2vY6PZf8W
LHgTkSyb6maoyjhkn+llCuSdk8Dz5s9JVfjTAF8WV6oYwN1O8yZ+qda4DhwI6mgSHUcabDNkgkC4
ddweJ0sxfvZGNihxa5hkS5Dd5E4QTuh6Ka5U6If66yEfG+/vcNq4d27+wvRv9oIXHEi895khDCQS
6tO0upvR1WjvUzjJ04qVaDIIuoUenofy566tgx01+/SMIVGAn2L88SmwH8jeJ1XBWtJuxrq06CMT
B0FjmoBAtlTjzrd8517yPumaU1pNUcm/CfQxL9xI4eP0x22wb3aauOOKBRUzcfsgj2jyKJ52UrSY
o8Q0Z8Rvp0h9iU8LP/47qOTkI40Fmtir3rLuROFwXWkb144IDgBQDXAQLiuTmfB/b8JHNjrk5eDu
XNUsc/rTZpdx63PijQNCQqZlOjQWroHeQhJXpmu9xzl0PoSRLT0MKwqAZ0Yicl9aR54f98VVjB2F
3qjcXZjRe/H5ZD0RgKpkv/3DTyFjREWGjGYzVeF+OKbUVbam/U9cSlimR+Oq72l2v0AaJ5NbVW5l
1tXzyeFaX3SeLR6GJh6U3Mdxc2oyELt78kDg85tc3yb0kCurMgXNirQf2TtIEzTrPOES5w9Y0R9p
jzLQM02i3nUXgNNkyWmj/cqPYwWanhdVB9gozya3BktEjibVQcZQdRQBusq82pZKesBqs63cRgFm
KgFuSzAM9SzmpHTkc+KiBcHKU9f1KHlynEjgncGtvwXd22V2wqauZLhyk9Ns5fxr3sRZUrxVzEUf
aP9KD4vzw3z1S5u6BWGAUrKkf/LOiZsDUDmZxvc/5FXzBUkiUxQ9TI6sXaTyjwkMGDhqCDvP/Mkx
BiQmdpZVFjtxUZDHuYdQyPHJI7vAWHauCZvS8THXLlUxA6xab56NcjTRqadmaskZDBLtdT4t2yZX
A+suK9z64pBp/zEBkia4LK0F22KZBk0H0ipG8sS3PvIAYNAfT4HA14lqvTBa722JsaKF9okr0WpS
aNPXvyp/7iwwgwqODH2Idq4yx0TR3Ll2hG855xjwRLZ/FDMbkQ1yNI1gXiiRlQIixFRNYuHBI/QD
TDsr7eYTcJ7MrIUB+2SVmlrVa7rod/ZqgnWeLCmgFn/yE+L3CdMcDUqj2Vp2H0LsZ7drMdLxh5Y8
7exNOrzTS9XPUDofiLnOTn+dqLkgwd/TQ9X2fuG/88qhj5EjTvjDgaypqkXlFHW8sf3xRqS7q6JZ
0AZ2Na8+frPPhnlpm4QXZ5lln3wsmp0HooZ7oT99w4dp0H7mnrbPLZsroDHB7dUv1sjmOeYMJO7Z
RBNsSSbJaM9OozLjt9p9O2/qQC73U0B8yT9vkEr55JwqfZB8sKzxLx1sTOxsDFFc18FkD0UjHMtj
txZUQ2aBu5MOamdZBcKBYdOUjxu+LHQCthkDuC63A1DM83ThK/XjIZxnWx0KwJsQqVLIocJ2LBQ3
aSkM9IO9H8HsDweSOiranQ6I1TfccPpvkqKgW87wxKHdXFa+ICn/X++vDs9jNIFSBSCjkAVPpXtD
D/UgTi0b9Y3W6v7pkJup4/4G69V5i6Yp8r1jFIGNa9fppQy2pFmvsIuRkEnOAj/MdamOShvSU6tX
49siJjxnNSNSq3gnF0MAVdn5zkU+2cIdZYlu8lC2jiqdk4ceeDgGPCBvLvTQpPUPhq1smGZmXHd1
PqBEBCV0DsBVLpn/t7HQlRFQOYgltGP/5bqEpnVAfYJP8q0NrbqMHWllWCM8JhRZXd002rTjibSE
r0WODuKgSH2jIuUVg2Qwb2dy5sKoYMRgVkFKdJz/Cn48lHucebt7M17qFzWMa6xaIw7K8hf2Agdz
wyWFIRDQ6MORADSvrHqDp6RJN4LZwECz/8ozBJFHZRjS0uOPZSUpHk/KpBYrA/08YLmj4kYAgm7Q
e+2ngrp3Ebda4Rq4zDmhRGT50PfUJM5O6PRCZA7mn1Etbv9knER5YoqoVcl3fAYFyLJgYXHxod50
Te/ohDVc7dqMOoK4GyfPUMWSMbVeFLYkqawmydRSedCNmqFypx9sm2jA7t8aZi/sYH2qoW65qX9F
kVd11/FwQOb6BR6ph7dG1ldLYg1gHMer6zHaqNNYEDz22SynhS7Pa+TOdqIC/njE5Nq7Ij+/mFPd
hG70iTY7V5B+uC5dZlYNEt+IM1WZNHpXpHeEB8+3MUkoRHOOmOZyq7piGvOoFX84qOU8k1xxJtIM
u0Q1FD9e0UCW7VgyaogfKpOqsEIhmql9YPq4YXt/aSDFM77KpuammZoJEo3arP1LZB3DmCUccwCs
TsxMTTyEUQYh2wbtbPeWkU4JumMS4QQ6Bb77qrP2RYuXiBKcSm/g6m8+winfx3h8CvTQ/FG7LyOb
5uYcmBXUp8KDm0jNoh6Kq8qwHR9wsaQq+xedF54uLGidUf7u5NPfRVt04PCEHYhwScLaJ9G8iUlC
O2BXsCBMYkV4+xtuXWuPssu4TmPS0yHzKEzYd6tgdtSILcF8jhs97bVs/2AmVuXTRBywCyCqDAOC
rqkWdXsl/UmG/je1RDZ5QUtcHR0olPwjI/PPEFceFxfycXFsEha2cvzpEPfl1CfXSebOdS+JM3JV
cR57H/86a0HSPCoa6f/eijy0uColHjv0VW3CfjH22hG+3btiWxKsmNxiMCB8lfe2BB9u6oDx9zY/
cVzDy5ZimhsffSqHpoGQ2kXZKcA0nPSCLXuKoZD6kxgKQrmXUt/jR47QlwahrUxRSaPzWfDL4D2V
abIESqgFM/V8kSfkuwT5iPBc9K4U4uV2yECldmse8IgnZ/qdXKnvJvJrqW7ITG+20o763J5bWmYh
YAWjMZQpa+fO0tz6L9jCRmoP3tENonxkQGmCMaA00S0REbK/Q0VcJZx9tz3Smckk4rvzEda4KT/m
nBiBThOFSlS6wzf55j2QX+k5R7hUn6gEUf7OwS4K5NFZEHZWSEAYGaPSR1tlLTP9+vhOmZZqEF+y
YSeNE5y5lZJr60jWDr2Hj3tD6y/3Jm47PIg88Fe7wjR7l/GT4JAKyoK300AJfxeIOdwM2nfIsiDj
RCXaiN7V69tvo5oBtHOdZW4OfDD6XJyHkk5W7eZPO4nKMWuyD/6AXiCYwyAk/tXVsj0nNtzCWUX3
yk+qeqZJmAD6ytg4qhgM7DFYCq2jb60r2xV/ER6soSiovRn3YdtROGikCwEmsNlQbhlLUnGDaqf+
txJ8nXDXeg0juEIRYKi8LQli+ytMTAo8qHfdGqvY8mpb0y9hvSgWYRrscqhPX/C0RffAkGItHgr8
B7MSaF63CaYMxKO5k7/FaX9jAptnO+Y+z1fCm1TSjLyfAaDIShlFdFp3v1jDgbl8QdZFQ9L6k923
tOaQqsFnpIJmP8buGSH4XEuEjv6KXfr6dRj8QXgGBRa6RFs1eAFpNHf9ruDHQrln2GqDBKgtCUSh
KLD8ruQY5tyVeCSktj9S5yHUlm7GcYJTLxr+VyTiu8IBAraJEKdTOwikGGmWprQCgS4RrSoKwAVo
N4w1bMP4EWh3TipDUUYqXO8nTNIOjXARibZ0vbS8Q0Pkse+r4DVBydl3HuirJGRgPKoEg8O2VU/N
jsoAyMIUEKISv7tfRa804fTslpGcBcmkkio1PaduIDput/ZAKMKL4rh4iV5KsB1kPSTpfnYP7SAA
/2aFtGfabzg7MY67gQiijjYo0RaeewwOdbWTdNeax6abClQe/lzCs2J4lvW9iUraPMApEvbgTf3P
tyFJavZpSsFrWdCN7/dvqKMbhkdB6pZA3UGU3tJMjD79PxfitbyIr2o0qrVjhLOjP3bhe5ftYJB9
swL9PcUualqhrO5LzS0jqoXGJ6CiL0HLtGxFrODJZU3QwCC3Foncw15hf8SHEBrzdL5OfetX9/pU
Z5ZHvVELQjovGzD974ZBzEPFr9Dx00aZoNGz0M99v3n/+bEt5ZYR8rAsFHvuhezHg8UW8PY90WOy
1ROknI/xgGZRmB+EC6UgTdS3Vxo+o1ojeZPLAOF1PFau9YxR30xKlN4doDzECCQAcGzzsR2iQO3o
xjJZkueiyehrH0hetgOKJj91nPfHOdE/dbPUvQIX6TB511JGR/Ezd5EhUqDXPL3OdNymAeYOdyGX
iWJOidZ5NWOxLJOzOW1SCet7wnxi5ljCYIdvjxYt/o5/CvCnu7uqzixERXD9AaxMUUN9rb+38vWn
vz83Zg51utQUZnI/+tPU/N4Pqauk7HlNdmb1oBluxLjws5OtZWW2gh1jbjQU/LKSjiv4V0+mYFNc
o9NBUAPW7cKl7Ec4MkvUjEkdyMs0AYW1hmfbr2ZsmS3NnXFJL1cwQKRqkCD7HRx43N0qI90ZICxl
tKT6wqkK/KsQFmidpvF0K+lvqP9g4M6AaVpyuc4hJMq/ytV5PI3CDLuITHvbr/zl0W5nctgcfFfC
f+u6CmT1XIASnLdW3kMUiVJY4wdsfZoD1MybV1uRSbEU//JWJQbEhv7tFWnHkz9QNereAnaWzLcH
IovL60hJOkqpF/Vzc75feFEH9VYoo/s1oyipQjF5hKMWZupjys3kxLVAscJmdOTzl9wDK0eAUYEs
UKFY1q96Ui62tNCbetD8nwx/LKYOS9hl+nfXgaWQI+wg7A17ygHffTTybqefFqLlJ0SrREDBzlJV
2f6E7+I491JIukW9Z81Ni/F+cvUrVATn1GjN0g5/WP6qkEtRof4ilmQcubL1QJv08jsPpzQMMqeF
LAObzS651kpBuF4HRexeEJ3JJHH9MlBJN1Yd67M/jbGLcbIVbaeoN4nlJER5hNbPaBNQ5ylgawuo
DJJiIt9oFRUf71ZcMr6ACei3t4lTSAx8oZxa2Kv1+dXfG+W3TRuByaT1LDFcNcNyROQBQ9bNOeQr
6Lf0jw0FX/GjLpaHUHeGR5wP7fKboeij+PDXdhTU7ytyqFIUiESJJ6urlzk36Zxaq5GVpxoUk1b6
+3+ZQPRaSbpHsvHsh3NvdbKMI5rvuLEIEV0TDnpu27JtkSMkdax4YztmLe7nyWYhykZZ96OnoGTq
lfwLz3mFpRXxwaLRIoAH6m5U0Dq8NK0uA/FpXEL1ytzNJi08aQW1Cwozgsb0wUkxl5yvKY19G93o
N5ySBbW19V3oYBkNKvxwW/ZfMI1mGacOQDDklDlEzABzeLW2dktLaGf4XreHtx7G6NsUpS68gyvU
qOlm3fABGstHAj66olRtLrkQnFRggXfL4F3xrnnLdvXmS/ZYJaSGASnBAscgUkPCMMDDRDS3y6tV
nu5f1L4osuhgpjiPrrK2gEpYJWsG4F7bigj7rYTpjKtJKMsjkvrxYZjTaToscjRqGPWh7IEQt6go
lTms4bmhP+ODg47uwzibN0vjjDhYcR1weRvYw9GTQXUv4yGOa2mqK+t6EI+IsemuC36MwWYKG9Z1
mBXsss1HDsN3JKuycRiw1gt3+Kw/LE49IIYuvr40TU1qvKSaG0wQflbx+SKEUYtvR1jktCw8Hgzd
2IvG0oHUpc8u6ocMyUXy5NYEkdWxR07iLhGwgcSIqIpwloPCUveVflbnkiLCHco0Ckzh2ZOuLi1Y
2+aFR8F9t7tAoSQHDBqYUHaDhJbVii3lJ1/Sgwjr90ItczNvFVdnn86XTJxEy5Jvnl+xQ3ogZXXv
oVtRABPd9bIbs2LEzFoE1uajU0bKjbUDThFR9fkfXX3kxoYgRUzblYJSyLysWFW4C9lFWif7SiFV
XPViQQSw2leL1aEA6+mALEGSY8nEcLGEVgZxE5XshQx2KDyCiphQf1A55qZKFgwt82bgBn47jMsj
n/+gIYVFd/o9jydpTzusvLe+xTZ5GjSa85o+iIE7dtAau/YoTMuTnbXmvyydUpcfHk4ZOMEwCiml
5DqvPZ0rHf3ZbhXBO3mh0Z9GPcOnne7Kq/eis17rjZ7iMM0llZ1p/oL/EEzF1RzhXsC6zbid8atx
/GegOQAq4r4n1nEv+XcYVp4OkB2lDqcY+krA7BnLx8ZQgiwZ31z0Q6GQ3niO6XpXf2GLJr7AXjgT
NJ58oJHWAsAdogF9mG6Rqudk6drbqCGPSSZbs+l+8PF/lXQGHIYj4G4HtLGbMBLvtG2DIla9OBeX
w9xC9dUnxU7Mv8KBJt8/rMkGQEyBxmYG7zOxNGGFyg2MeLfiT4gIcPwp8ta0LIVVKsjOLqhQHejg
yTeDmGQaha5A6BHs40gibr6Aq05gZFHw8Sno6n/I1AAtk/xEV6ITtie3SMD24ZHq8xRYV7nmoG3U
uXOf6k/za3uDGYxx+Ssqdr7St4A8Q+ZEjQIlZu1kGlLZ2C64f1IctR2JXuDN9P8lkrRcF/x+pEkC
bR9n5PDs5a5JlvNPuEFURgxP5/OkkkdlmMVfbLkEsDJJW4dX/xtWFcCU7F0jJXX12ifzvyj47TVh
L7TCqkUwwOKmRMXWX4s0WFjt4IRSfHLPVhag61jsyJOLCdQxvWPyk+JZYW04x2AvTRG1sToPYw48
uujVwExlfhDMu4NKhTxeUjY1bOdlbpq1NZTzYlvUaZvRSPXc15h8YBiHXDB4lNiZ/blsxwok/uzf
zFne2NkjfXpMK7Fkfly/QbYUvuD7fF8ouxKMgRvqk+IfAoVe0cQkYmBB4JY09nOzgw1ayArdQa52
An1K0two26ln9nmzi6WlL61YTiSEXUjlELwHhbuxMA3dGUtIXJ7pgzP866AmttdOhRP22Mdh1zJ5
tyJsPy0GSYwwwpWwKReQfaU2gIxoE8r/vFevcmkS9RusipPckb0+cmWdxFKsraW9yN5m51poqxDH
YbtHngoTiwPmVlawIDn4FMnWD2c+feRXHb3qC/0TfVhgreMusW1VSxTurQIfYEeEjt3AYSSHd1E4
06zynpk3n3qvsubgn+aphOvSvZJI3Xhxf6AbbDxFQeQ2sylMxL2kUMISr3Kc7zkLWz0405WL5+Pb
FEyzu6zevVeaXbGAzVgRkWxz7Ql4sOJW4ZLm5QItUv1Z+HcvuMX3K3DViV5Uu9v2VOPt8P1ozGvM
6jNkF9sZvhocaJ5wyUk3yRru1QdQn4YFYa/hX5+Fe36olVnOJxtMqfhXg4uBciAq7vN0JCW9KSKL
wmlwzoitOShUzkO7Efdmm0KmvojqP0/O5KT7wAKVVQy6PpKtD2eACeDHVMCSrpT5Y311kUllDzd1
niqCemMd7yhSdf5wmTKYnKdupnl86bFLzuZaOXAJs2Eiu9IRmisbiAm6dSfpYoCcwq0PbOB1z1PT
geX28R/1hkRraV6y0yGDtYMNPg0g2T8QnAy2AEqGs3Y5J8qvjeprK1jD/S9xrosfGdXa6ukaoMFi
ViSkMBLOuJ3SPVkoj/JhW67W0pFPv9phr1wxGWF0jwx3GCBDdgmdEwipoIEhjeCAa5CIffbGwBT3
QBmgMsPi4YZ3iDRnnN5tSmBhv/O4k/MnW9m/yZQlF0Vz6kDRUoVR7tGexxoi+A2hJM7RMAwj+6S3
A1v+lcKYCMbz63ZlZaS1X5WtA2To4aG7oUvj8tzLCKa5MWzopZXLhcdC5jA/uYhzRhvquhMvUUt6
Uq4c9NqUrKNGlfIyWj2lC8m17kOaORxG4NEhXJckuEJ1ZtPLNA8bhPQpLf7fxIQLYOgyRH6ISOc6
ruNAQSoQwyU0MeU4ZbeDXXgH1jyB5et+777WsFUz9zswkjIhu53XVic1n7IozFRIYyw6Ezshlqkb
SNjEvaxzYsW0WnKoKxXLLwv4bdSxVfGVw1T+M2x19H63tOoTJMW0j2IdEXy0XApQYTpfZPIU03fC
Wp852aJbvfgnXxebWv8otc+b8jHvEhEoapiy7iJ+uQf41X2KirSPs5Natdhj2SBFT1jozmG7YVCY
lHdC3j921h13llxHm/q/3It4eoVjsmf3FtaX0/oDW+ZGo2pmyOx2Z8SGmpX4VGlD+nB5qZm1WGFc
O9zjv3IkedBHjoac+KyIEG9j/han81ehpDgYpKs+8bKAKuaolwdgNKclVCRc6z2lD1H9fGaELZ+O
NjeeZBnYVHb3cRz5YKy9Jd5u8o44hlILXLFBs29GaeThFpzvwmY4vVrUNYzdZorUxsK4LgqlqvtW
cB0N1hHXSDd6jan4IJ711AD+geFi/WW2OelI9aXKnH64oAq5lkBey/AilORZ9b7FWlE2e/I4bWJ7
GLzaU837KAWJRfPwWFZOPJrtqlTK+Nq9qvXP8WwPAa8OrCnCyS4OzYmFbNEQzfOkocxPCHQOtGbm
pW4jUOw23U9oLxdM1I/QiSxQ7+EH/mheryaqbtjRBzCDDg3ojSxF8KhMyZd6iytVH6svpcMyB4Cj
hec0piUyP0DkhDu0bHyXxEPkTvTu/4LwdCzN1RQ+SiNCyubvcSUo6hKQNMxl/l+7MV+lUB+qqIEh
nHthXVmuAnz1sWftwZb6UwN6O9By0ksgJb9oUMkXFQqC8nkXAGpltMf0NE3+p/GW/bub3WuA1gfW
AAuP7wW4y/GVD5cdyPqFcFYclgRYNpK2nPUd9ZKkr64OwKYu9qLM++zN2G0zsxl77oeYrGoUAWH7
LqM45GryzXDbyJre/AxFUg6VU+tpZoXEKUSgjyEHjJmUg0VBr7b51HVyXKPAftCpnsLoBDWDcUsd
WpXPDdY9FslIFlgFPnSuCthP8yY8oBvDqyYJ3nhPSfYDkFFqS/xRjAXsdjw9kr7VV+VkfXDIHxjo
SpKU6qS8xhYaDb8OyVuQB6UX1/3VE96DcKAgSXjA+L+qCpCT5vqkZ6nROmROm8H7eMp5O8vn1ZIH
8M8O16IoHQK5Ewk+dcgrcAsKFGsE4WcQ9qqCtGYvARmhjhlIzuZLDOXKmaGnIvhL6TOSr8qiPyhe
k/Fw8Z3jT6UA78WEsgYYCFT/ZXZcewdACzPMv6C8FmTYiIHQwCspJjx+gS27FodHMpv/BPbIviwf
38qmQhC9am5HwOnd7HWvlsXfGbK0XtvRQiqkyo0m521OfnmBfUqcWKvRKkUC79UL599EeGgigTq0
gq7HksNOIv/xXr+56o6J9jIEgDywrJCHlqGnQTYU0un4o7KN5GgxzUjS2zTmudF2AtqLbUwwVjBh
C5G05szGUfaxPsN/e6S2zpPYI09bYOAZaVLGvisyecyjONKH/FHOqO+BHEniMr6tbfONmumcTmSw
fjJu17f8dA8PjD6Q1bDpPXTIcFnK3fM10QzXzUQCgXWdcCtq9js944i1N5bdsSoJNUZppSudDIEs
EDASHrWWx2J14wx+qCUjtFjTO9bHLOZdGrAMwQGGWXzRISzpSThyJ6BPC5GeG6K8izGD2fSPAkwB
xIIhYEczaXGn7F8H4hgIvkyTXpWUKaUQ1fVbTZykTDE+1JEqANTBp6PllQaLXF+epzcbtNjMdXfL
EAOdGVigGYSo4hcA8Ae56ILlTxIAyDp7nCkl47nOZj/rwBKD08cInqSVu4rMaIT/JCF+1hiFGuEW
keM7pqWuBfu8lDDhGSchGVR5dahHMiagW3J5HftJpcyPUAUAe9IUQi6UIXAsY95AxZjthva5mgpF
LrTSUNrlE1Pn8QHXaU3o3xSKkwpfGbFfVqhmR5LJZ3WnuPI+VaefhA1sAj9xBy1XTFXZ35QCGdeQ
tZOnBnApQ9hMcvG9xA2o95gDOmh9PL74jvOKuDYGuQEM/UYMAKbT5c8+C0FpmU3PEU68fIAhudLl
Io6Y1za87lOJdQ1FN7yj9vlhYpM5MXwoy/Wrb7G/K0QbcNZP4irOxgV5euBu5tVTbXvEcu6jULn8
EZWDhE8I/wAlNG9Uj/gqKkkzsHZuy95zSreOTx+J3SSJOohgy1c12zOV0wp1HEV0JyZmq3ew/Rv+
22LmCh5AP/oVqjegg/v+RmHhtefWr7BHB737jbI46hKeR+8ZgtEzCHYAYIQ9OG/ZRBX0UsT4pkcA
spIjJAtEnNkzgdLLxqR91ZG7uNp/1MOXNf0Xdllfv+xdE+h15IER/W+VKAICZTJ5vw7BV79JFNl2
aUQEOxVoECWvqklVUc0h+6zRjsRaUTfMdkvtOeTZxyN/FQHiHwtFxfdqnIoi/oaV+uSbzS6RJX3v
DPRH2anY0c9P8+2VUfQc6KPrsOzQdSE+KPidBgooWTsMTAfgRHLpump643iFj6RTZVILGi8kj4Gx
jQXVITfgZbDKqyOkBvwXcpZ8UJvoOY9WGaEt5LtYQWLYYf7bTVo84kZBU//47jykx0K9MFf9+y82
uNG0xL7w4+X3ovcnQZJgPYMe7QhxCJXW+oMX7ydvVm0/HXdyPzDiToW/eBOdfLrzkECnFim0Ze7M
c6dWLuH8Yl+TMrvMqiLYzzBtSuxPTfLuFmuvundNswtWIWwlqaPYKKdRJfefSkQARVdeITEpB4w9
NbhI76Fh6He5jzFIn7LidbLD4VjT5ZzS2Akio2BozSHKYc1ZyOq29qk1NY10zRAiEMC6DuaFWQZj
8/q+4oPJEKnO921BbQWgHHX7fI7K4crvhQNL+Ow8Mtr7BR/1GRpfcPMO8PNvR7ZFB+WsE7hbTMWe
wgAhxhXM6qqfk9XNn5Rax6gZSSL0kAqz4Ugr0pY/6eZNwDX2nZVrg09dxsQgsjcdh0qFcFTrJS4l
CJgmxcjGcdNsvce0L6g83mcjOVvcmcG8POVdO5ghLh+OS5ZOLNGW49WqCKG72lsS92ZFJooO5sZG
2uIdhzHXn57wpyfgmmbJx5SIdbjidffSPitFGysfgNE37pnfuAKtwsFJ//38upA7lMpXxPz3CPVl
DjySqfn/ZJw23wwCR4vvTI43tezv0n8Y7VDB6YkfYGTSi6cwuzmcihF4JYgtPwkYlDho2dxm5Bgm
e6UPV79bTqfJNVr5EkGdyCDJy0EXNuTPYTMSkcADKh4wGUZru3pHWQK9UXTSCW5WGgEVRQ4yR5sr
6eJ52euqta1guJVwBM7eVBZZYKwB6IfUhfeXZydZSGyWrCDi/34r6B4GaMrySJD/oo9aDEasxAyt
i5an4oVcjiyvvkb6yUgC5Zh6UGlqEwSOLl1OTLNoE7Yh2aIqU5/JPSdB/8pI7SSI6hGtKE6BpTaq
TY7rgbyO7uwD4quy6mLZY95Go2n4YSLdzFijWaiWh4/zDXaxHw3KIm+Ag8os/bEKRszDa3BGghVG
4HRULclEyOlqaRG6+fDfB0RinX0CW4VrOMPgOtlExRGTXUvWHlQP/42MDjB3UppJVAnQT6BFfucL
AJRys/H9w0fl0aWBYYNzDes8C2Yonu10BkrQZ0iibIGXAnug+rveg5Gj2ZcIKaVTLQ3fpx8amEvM
7kHWl+EOWk1qHkHk7hg0BybK0HcPvbNl53fP8xbaMc+7AycLzvAcMWlqmqBbWlFAcxwrEd+Z27Gr
MXm1qBoZGIMDttqWGUj8m4zmu7zOvfRI1T4Bb7i3/cBycS5qPMDcqejp8EWW9ujeZnUs9Ws4lsnf
2td1fXNr0T0W0OpkGSs4/lHW2jB+FJFL2sRc3t2z2WG2vTveL2zJhIpHMCfhQ8r5mI5/qgfuDnYr
nXU/A90ql54LwC6gIr276ThJaYlkmoQzaBESVy4CplYZiEiWJwwTHwvDcD8fF6uAPosOhLvs9lzH
k1z8Taw0k6zKS+LRkrbpoDv8g2HgopUAphLKnUX45MxLbeFunMRG0mdNQmkrga4jnE8hx1yhmkNp
vaxH1AcweHLW0MORdPpbJmCwDCckFwMVcP00ssuh1pb0dkkQ4pAxagxT6tXapGpN+yH9CXTzfSrJ
Pf4VMhmP+x2aIIiCBejbcHG1veq3Ka3NvUBCvxYEH+eZw+jXpWXd0Ove44j9WkN022cXCizUg9Or
m3DgpDMrkrfube3EKDNodiFgJdZL5RMlUmwbma28UoMilxvnaKhnE0QRBWMte44IWvvcquREqHqQ
cF1C1aDspEpDjRSt1vLI5j37Ch3gOTkHgBruTbKy+YbFkwxRx1xk/PAXuPMQsAa6EU//unRVdRPP
pXTLPg0WA+NR6mJ0LL2hOOSCPUkrtxFMFAkeZHVsfpwFVfe7Yl7p0Lis3lZF0vBVMlps2D3i0Ihf
hDPnw3m+Lw2BV/LGQa0MFP3U4OWlpv6bJPlCDAX4ImF3qEw1E/V3odSmfJfrlN6CMnYE6cFW+8bd
kUxkUj1muMhNOJEEoJKeDt3XEMmzlybtF+mdhIyKMiEX2Cifa8oyr2m53i2zjz4vqK+uE2YjNxd8
Zf3vbRbFUH3Snzje58tSRuYDVvnnujXohKeS2bL6a5J/iuuF5vMg4wRov+vz3nY3mZ8JxOx68v4j
v2BwbOrAAXsVmLdX84eiR0BixxrPr4/jAZ8gAdjayLau4cdIxHr/Dgdv+Hh0o34rRKX+TXy2BQ1m
4Bb+Cm+G4EWNbBW8l5oISu24vvPmEfsBMuN5A+SDADGYzM/qY58fi91V/lIjDPmU6IMig3Ve6sLF
GbSZ6j0Ht2d852VPrxP30EmzwdxoVfPvBQTxQ55efJ3AYaFWBtT3x+i41MIWdOCA/Cv9eZ7pAL4J
4utPxo3/bbpRQhoXeGtIwtGl/aJ8+HFK1HDSp3toKlzuL6SretsbwGt91SQBLDmIUuoPGpMcq0xB
AXsKsxKoQlcIJB/Ug7VOm5d0mOhR9pudkuIHfRHJ9Neg3IxRfAqsElt15IKm/xf5IpkUwUfInLRK
QBZUEiLSR7oBHFBqeY0yCaCGrfYb6KqhgVW6uvJSR5lrN2joOPf+syB2cs283sVKZWTj+tbsyHfu
BGwMIqSY4fqKiTTMCB4tJxoAGOmwXQnxh8g+nGpHyYSxghvEcgOnK8qVJJD9wzJoHW7VibAPdnf3
4ughsnPw3DialNHnatnt5/FUE/YlnKkEfuBbV7FF98xtXJP68rJY7OZpjfsUyogVH/gNdhrYcgJ6
xjTyYGjS9UCPVeeeYXInRUoi2LNOEX8JLV+9RBaOOb0aZJcDA5qD2A98BSH/JoqaB/Jk1dIjheqV
sASS7S42qk2ib/K9Fu+JsYMSTbGt8ksxVRqt9JKEt6toiEHAuHoOWI323Bg/T3/hje8r+U5O7Oks
bNST750WsKJ0wx+UUOisuct+Vfm5OF2PXpymsdJ5j2biEvorohjFKEgY7n0HVpC1zNmDvE88JuHJ
9vrZ5rfls5UWaeq4OZN/GSicMsHpxQQ/00uk5fQ6+n8bKPuWYSnxFs2vegkQC9BxeqFNsprjeYbR
GXRV1Pmc3IuUCWkKKGubirOYx092jgg4CuXxutcfBBbyEI70UkakFXLpOvkTVMh7UD/YwsD5wtuu
3PGjfgpA8Aj4DJjbBSmJId1fbhyDiNKPSI3C3X9uPBHOsIuM7OH6O2VpMO2FbvWnHQnO394AbcrY
SJZHZ5mVnxkLfJXkJUGN5MwqwCWHelIJh6+42M3610bzJHvma+kRt/hxPVtiP0F31XqR1ePE/0bW
o16jVN2yIP5ChBqreiwT24k1zcL4CQ8i6yogEx3Yy2nZYNeHPvmKo3i4Neobb4F2Ro/LHpK8CMsp
rvp8t16aKmITywp/joJgODLKU9/xVVWa5lYqOEtKt7nixasycLzkTFhEDGO/32cHQJ4noFOFg3xV
i+nioHjPXsm33pbILiW1EXGYG6pwqFpBBw+KcNKxwsA6Qef0n9ewCr+YCS1iziZSO0uav4vqZG7d
teKfceZQwqAnl1nmrHKVPN/TN98x2yC+jLZGEalzVMBzJ0TAo3QO7lfrX1pu95AuAR+oaDQYM7FO
6F77X5GGwclnaEIj+iqse+SE9aeNq/unC6oE9ewmDYvh2XWivEAt4dPuOQJfbmTXcTcKJRrm6NCV
22cw3XkHMDbyxBWMi8G6/Ph8pGunFyL5axN3A4yA/Rc10YXuONza/8fTjcDw5lOI9hp5jZbcQm7I
lFOvTAMR91dEkZ/I66LZ7IFgz8XJSY4yjLL+zmhglzaidFYZ2lNi4uU7SlyaIz/xlErBgfOd247P
FQeMTvnClwDZxc872Xy7liEsrP2AQyN+9lDWZD9dyUPkobS6byp4b68GYM6h/VoeYpVophDjEtiH
B9xmob+T21by4L4op5GTSYIvvQFkAPgfZS2FH2noGMWbOg9qkl2aM/Vq/gDv06WJOynBRIlRmMsq
huXHIxvX+BCHsxsUBHbUVSnYwIlMQkS7BHvdd5xctefqzVIwVoKwx0wNQZUbxV7gIrmEqJPi3Rq2
Nu39WEWj/hujnBedTSF40aEMj+Xeq/hT5Wyn/XFPBdYwithwLI59SMezF+BNPvFTSbvsr/WF2HA4
AwZWJFc/D70NZvPjJecX+cYOXq6F+kgJKxs8EZaHYtjC2tEx00h82WuSjKg8xV1I9E78miCMmCln
ZHeOtIgV/EyOcYfr2wlHfMvzH3Q/2jBnWBTdKGP6LW5wVfZODPuQZZOtmKNwDivFJkJaswXtkx6R
AAnf4QObcMPDd2xo7mxjntUgebr6Df1hYDosWsC+KPcwspzm348ShbUc+YYPvu52VUzprwPoYZ2e
WgOhjvILAoidwhJWNW56vxMH+tduE/YT7rouLuc0VNJh3uNEujqFdUN/4AmierDDZ0r5AKahDhAI
y6fhoPR9nrhJVaboMD3gIP9qWJFaiWbmxMN0WCSJuDOFvp2kT+H4PYuiXl3h2lUidzJD8OVsJ8JH
YjaKlBzA7AK3BxUEzjcT8Mk4iaFDrI0fSyi1Iyw2qUlNcaVH/jw4RK0UxkENIuUs2IpQ54kfR6eL
aQauR5Saks+zKQuMa6WOm/XYCXRgw7q5dHn1PmMuhlb4nFvd7lzfS7qLJi4F3VvEP20hpQaDKrUU
JUHxyZnPQefXjLSkWrXGqn//rsttRKnv1EJIdqZNcRaI9aJTvF6W511eI5S0jYg9v2TAwrP7ftnt
hafXt4M0DNIvM+Ax0FHmHRDUpmza26hqcqUOb/AFmKF+w1sXEpzE73hUj/C+Eo/q4tLnegrJ6cep
cIfV+HCS/+i/a7POtxZgmYICOmbi8DlsOhvk7XjmiNp/mXdBtlugqYJkoO7xC8fBaKwINRe2ZT2k
qVpWtlX4Eo6f7vdtQZMRjgZWoFj9hhZ0QhUQBAljPh7CG26upxdPUozTOdBOJutj77FWrGYeggtI
CIk7C7KWEMtQNBB0vdBMuo7YSPo61voVBq//X9wNe0HuECNzM/0ScnDa3LmPmEJbWQ1osRP6kFRc
Z5s6N2tPxgKYuwhTDbDXnvSVXEzjP9q9GVq5ZZ4QYKxouw092962HAFagLBns0CCB8kZQ1dFVJip
UP4lPLOcef138JyAtF5W0OvcAS/H7PNN+HuRwhzImOmh3iz19uhHGyneF0PQ8Zt5hDYZHeu19kYS
E0L9xTeTP/iWrPlnlopcWDuaR5MnX/dXMmPuDg1zPEfwsKPGXzbmr3kJPKfpspc6U3ZEKAs3Dh//
W2usIr3a9CYdeIHL+jGTAp/1Qhbv0YVEA1w1d1azrz3A/mT8Tzm6DRiF4Z4nbgICrWV316jaGWom
KobkWn/5Al3ffLYxllfs6QDHvQqDLI4ZGgJOxaPmey3fbQt2HWB8I/S7GLaCNha0eS05UFfsA5qT
SnEHqhYpqkIuKBu0Wjs2oBtSMmpFVkMHbodd+KSNuGqRXXnvGy46mNyGqUu3kzC39CHPhh8CQWkv
HJbbGE35V9yhi2GaoER2ov+oGqOoLCXzRqUPu680HOnJkDVUCllx5/muqmNwbe14OxWqZeZv3Jyq
gId5ayLpXzF8SDbmPywEXp7FsbnvY9sG+A1w7N/mnuIi4AEEEX/5QvsVsnTEMNFRqi0EE52xIDPp
BzcqngGMGgDQmV3vVI3MKE256ENDRpD5BpT1zHAnWB7S6BOURZhakvBC9Ewi/qAwbRXgcOyl37zh
dI6iBBhyOtmJbdnkhSFxFQIhUP7PZl2Mr3C9hr6DXm55VO9j7lqwBuDWjHKztmFciVRam88MNu13
Kbq9bSCDQk/TnpXn2DJPq0rmMDlmSMH4oPrYuzqcLXdrD7JVXPSy4CxNERtImbK36LBV2axf8OUi
LllYsvoBPsWyXx9Z38tULqTu3Ub3kEv/6/KJ3V2eUuAceI6dctbqAhfyG5nK63w1tVxbHRzI5HxY
07jRdvHGPqEFyseDxz8mFdtgt9jvdCRyz42hZBAKiLQVy5PV2DGTzg9o2DNSp2k2JIZSsVWxNEb5
36cSixX6lKhkNGzSp8uurVY6u38lFTcwazd+izg9TA0I+Fnp7/TryXSovhLww7yuccekYZD563nC
juCti+yC3NwwRdyRA3pHu3vYyXptC298CX6Raa4uIhE/Sl7PuhM3KnUd00KFPvCRbN+txUUjGfJj
FyotiPfysJLXAJ6uI8UW39r5otWwawW+9t3bMiNl3SQnmYfIiLXIqpA3DiS2lrwxFnK3oPx+qusx
5EqZjVFgPabfPne81p8pe7wYbPgI8T66MjUX3DcUiRnaDIGdGx7tHPZ6xP4MvbfWojNhkTuJ6BzK
Nrt/wS1TjGNsTTwOhU+rcw1hLTTfSiv4WnU8y+s4gN8Kk0fa+29prwhfRbJTvL0QE6dRZBzKbFU1
JfZljcFzd6K8uXP10uUGxUktSVtCtYIT5eRYlP3i+qlNKzihYZbExeQBrrHQD9E65AfoxC+h55MI
32ZZPfeo1laRPEdpOSNjtaGJNNZYH9nUefsQdt3xe1L8ZTDXbyslevfSBGTEbJ4tln5W32GfBiuY
U+Kem0NQe8RdTi+IoJj2t2tHaLaxa+H9xbFp1NkrheK19FdfcEzwcQgkB1MottmFPAN2mBNzNhCz
lb19Rc8jaltzj19NQAC8uqyXn0gAeYIIJSjiuGD8pnUGzN0I2AmZ3u7qOMQhkhCmzCqNZpDC27nV
5AA6Efp5TpcOuI1FB0V004U5PQFmWZVwEdlPgRaq2WUCQZDcFu5A8A5M6FtYVxRbAEDntMLtClv3
9mr3yO0YEEM0shdvx1Re/iguFq4FJ3dkgh3zUqJNVctswTgwTwJcBbJfb3nP+wnlZmGm5r627Fy3
jMk78zDHzuBt99Hjix4HU1N0cIKI4S4c4LRzCWohN/N6LlYA+3bSqSaQwynKDIA0KwVBaznBES6q
rYNHpWKdKXA3ra5v50XYt79xHyrJyK60zjXbDVPtQEHU5X/3vRxY/QnACuKWkW5pX+sGSB/mARjg
JAUnkE+yXRVj2l4mMdR7qzybafRkDnJ6qkxIZ0BatbxfrqQ1dzSC1wQS7W4bwsWPImt1D2MJG5xO
Y1+wUX+PtiuTi1UVgwZGgXKXR5abwF5NeaL6cRoDuCcZmLxvl+xTXAguyLT7ABVUzF8Ib/EjocpB
Cxx4f4S0huZeRf5DUq4HSY/1KJ4dUNnAVm1uQ6yHQAexRx4W/ZJDzO/aDaAuVvO06sEAYb6fnfUv
zb+Kce9zMZMsqMM6AfTaTDE7cNKcDkyxRISZYoI37GZJTF30ug7r4t1VIR7cmXoT8ajLr3l0Df9S
YyfdlnC0fgevHYcEv7hMuglTjsSHeIAdE00o9cCeL7sM35LhN6fTzl18iKMiBxtkbOqFj2sn/caV
omZWXh0k16APk2DYHuAKAcc0736J1sKScPBD6e+oaiXN7Fy68WQ5Pmodo1XHDgCxj/EcnWPURJn8
mhSGyu8X9HK4CAfjVx6DIgQc40IHPVfddqQa0WU+W8IIDy7jlrOvkuIkt3hNcShg+JVtzlgSNHIb
D0nseRjxy1Qb25bN0Gy1oNWohdpAPZOons6fPHX4zJWxDB3StTG4yd3yL5B7d5l5IqCJJXWBc4tj
dcZ+PojAHX0yXsBq84p7QalCsKMDgVAM6ent3Xe+wlfjOqyibTCZCbONJGO6Cer2fEO4fiUjL2is
sUeLIfG/iJvhQ0YyTVlKor7uPNtRLAD87oYX+Gg4lrwMh8h/emTbmkqLDbrBX0g6kqMlXI3YFGpB
9pkOBCiiqbdS00DE2Mvq9cMHn0idaCRkuM13T5SwklMvXGDEXTN2gs18YFSSu1FgUAxOqnaBnlQM
c0MSaEYQZZscei1YZ1/m8cuXoZbKhKFnvrYsrbu5dJb5q/qGC04qVpdWb8HNiZZhzbySCQEQ0ECY
iCrT+R7iFt73YTLqvvUCnbHcytB65neoWb+B3aIrbniopjGXps6E4j7twYLpHY1mpre0waLQN3Y2
G4HPf+7t7zBaRD3bITnzCQyTfflbKbd/G0LRCOD4QHTOmpGZuMBrWQ2oAJrry9aGvB82PL3beIK5
kLLSYYW7U9/PeyTvBTbIX0LtrqB3NYAIz4INUl8I7Zo8AgLsSbRcWfKgFzoVm8K9QCBmvDpOMM90
+anlRCOYqpJroTkmOjkbEzC2GXQiXMbSo2/HrXadf1sVrCU4nDnLDSR/xzscCfUli4AKubRV+yVQ
Gj5oJS1wqoPC9LB07j82hDXI4qUB/E5/XtBWbSD3YvEwtnYk83eTxV2C7njJGZnGw9OMr/9Hcs5q
3L0qe1F0MHUxLvIymP/n8gVyY1l0weFR7TgAaR1AVdMW8LjsjA8C36k2ws+41EVwNrNFtfCfEZ4t
uiwT1GM1qejj7B61f1UnmrJ5Sgeyeg/CyjDoWvDGatqdJyFwVOnvCNjDuEYwJBr8jSDGE23OULNa
Um9wCiL7wt2YXn0nuSSP7fH7wobp9H7jZwj5uwwt83G3TvkrI+JjNkV2S6QKwv8F7tolJmYQ3xaa
NS6snQSAgaQ3U5RxCUIEF5L7UjVQ6QAXq/iXZY6OIdfD0xk6fJBECtLS3wFUMhCErHlDUVBqUgJc
VjMJ7Q5/gKbgAelXXbnWAmTetMEbq7TBybdDrwM8nYdSumeDaw/58DebcN0Nz1aIuFCV/8sZfgw8
+rFm3SkSN1WywZ5gSsCCA9igS3vf8UHGJlBdCgizueX6vYOUJrZTI/h4OfM577QHkS/azM21RLjT
rwG+4+CGNMK1oYuGrkemdAGZ0eFcAsUDZBRxCwO/iKVVk1DDdYhMI8TJy/DYJOpk0cqsJZrtJxnq
7a0jCp5qHq9w3WLeRzeK3YP+k8F2cBmFMjhv9vRHRNk0gG8uEqCsZVnQ9iuOpEQzPeyV6g3Bv9Zn
egPaYFOO2GmGAka8mBfUC3c/0G0ouQo2TSR/YY0nnRmn5ZFtITQLyWG4HVO6rF5GHdQeQosswrjd
jgnRWhMd8CtEE5J4HitPlPPoS6Cy+TIQ85L0UGMZYIInhM7nWWAqDQr4DVFAMUFjgZWQ8ZZIYRtj
S//Dg0UfG3k1lO9+M0/AueflFV3JCjhGPZ2SfUdagPg4+Z1Cx/JRZs2cHLsBT7hNVfk1o4Xgt+q7
Ma2GMaAt8T053K2pf1Y1NSgrrPhOPbOMEzGym7gMe9c5KeJ0/nQ/yC4OHoqCcK/kcC5MaofY9h/G
0e8JdBi9m6pU8k1CEXWIriuIndn7WGe8vP2sLCB4bJw+WFhR20CbBG5RG8EuctITKZqnus+nFeX9
kEBJZ6/7wfBD2zpK9xfOOsAa3zbChwscIb1MtNtYZc4BQOes9ZITnTgkcveMstbztSr4AhdiXXQr
jxE84SZwL8QTULfZq/0Ek9xgrwic7XyeVhdur9k4iMW/25WsXqeWMR9D8doGOXAoP+OscaCU2CBX
PeTpfPRBOK/t0KgQCXWP2cxw1jOAyvPP/EwmGS/FfU8iNYH7woi8SZzWvnZQ9Pb/g/VBliZ0OZ+G
DtuyZCb1MgwHCrNCY+dwRioc7LdkSCdiAmxkx7afiT3vYY0FBJKnyjCVssYvFxTod0liTHR/PxGm
wPqA+ioNmFfb5eqJcRi+0N041Yhkv2wleo6Os+xUM21W/MYWAF+OIqtmZny7yz5PZNrQ3Yhpm2jW
E7HTYenso2ota4xRxK4UKQFu57KQoHIjXEwVrwOTil/kxSSco7soRjhj+XyE+IvdnrgRn0nFZrDi
6BFvM59bi40DRGJ+gMzbRfKEAlCMwEn0kBq0ZoudhY1QhbXohKG0QAQLg1umAJr0Lv6d6lt4uHPl
lWh1QJKiWm+VSOO4+G0Kr/aq0BTP7sirNfSPwWzW4nC+CVI2Lokt9CDbh5NnKhhS4kMcx96K3Lb8
wap1Axykcvoeu8PM2ofmXGq3nYts7fzsX4hE3EXHcV4/PxORMdM4XXqloviX4/3A53pC0HVxWeL3
IaxLYK5H+emFNk/4BmNbYMXAlVbAfFUT/HiEgIgrNAF64js6CbsZIRLf7ezwxhu6fXiLYipuWMmE
07qi3FMIsf0HhabR9l0H/Udy1JnmJdV1TJl34ucmCrSl21nq+lf1hGL8TTUV8aXH169wnz1mh7jm
+TiH0IkYZJqgu0m3Kq6Fd2jmeeFsI6FLQCxuvKbYyj5h94UhkSqPHpkNgqyilsU1B6mSB5TJCkal
1pp51XIzx2/woevYQAwXKGNa5wnVEmjeAuZgy7S2eQ6iebwR7IQYX+BPgSfAk28C0a/vxt2KDYbk
kZFx1scRWBH5N5hzYHfyX8R7KqZv/xqMrojw8imUkomfLjOA3yF35w/jRMQdLPUGhFKV8abOXxWt
uxI6kXRRzGpx1+oTT+Osr0DDu+/lDxDm/7EgX2DLr/LXTZWEhjQrDv60SNTgGoZzBT/RS2o3i5J0
alFgnGla400pU8p8QR4aOuhvXO0m3zOLZhxzNjh3TbWyA4zCzZRrkLQF/d/tELzWMFaKPM9tNtjo
ht/7s4qKczVOoyqKXoQsdhoAP3qya8X8TEtypP2Wk3FEBX+RNjZIvLBlLT7nxnryrVJ4keMpyspE
NNrxqq1Xe/F7+Dj7y2fb0ZNdgA/jhUiukGowNHCFOVJS/A3mqQc7PNfo1AkxVqNGQj5my47iJG5z
VKfl9qP3CCO2IsL29YX+eKWBHlIEWvO6I6G35czKdOu1eEe791WdrmEu9ckoaqkEdOa/2t9hoiAW
6jamfODOjM0ifhRCnTJFbSacGAdUBYKwJgqdK/3XEb+bSOGHAv3+HgQY6IYm7oZhuftM9QBdzMnl
8l2tB2OqdmbyP5srh5c5cAoTgG3Aw5ddJ1OJuJE4Qpa8HCLeLsoBZNq7jgrIFclmcNaqjAux29h+
b5fOLQyfuI9/Hv9HZfuB6QsOt0UHBESGqm29WcgyCaEo6oR6yziLtcksU1Jt4nekOZo4U0KdNAF/
gazPpFRELcIPM5s2uGwNtUoSidlXitgq2SHt8CT5H+WXFZ7kvnIGOKlig1IPmtH8IvkAGpEIdGAH
YXqq7tFZt0WifmPju74nzPtvWR8EDGsfV2f5yf9cV1IdZ1GZdBfvKqBmrc70zQssL4OR/PkCrUKm
tQHP8rXX+OJBhrEXFKzUFpNVty+uLyUoVICXgFf1N7q7e0xzKKDRQmUcfkA5Ctaica9dtupxmHTn
gDT3J5E7oUWNsJoydUU8eRirl0PQDup2YK1DnmbZqHzkeocdrYVQEE7gyReGCSh7HToBuQwKRflF
uwUeDIj092iKWa8mKzabnYFsGuiTs4if7kcCZYkpb7IB4tWPylq/zJSIHEp50DRIug1YwJxcWh4v
T7Ep9zUMjoMBSBI3cnU+CxcUvQ+GWNV993nwu5CCjhy5IN1k2wGB7O+LU9HS+N/PwbSFobuGvqC4
tPnVDwsUdRmfNFMhSQNGBrT04wXgPshiFq96rWACI9J5wpkkc5U5IebfS8/b38puNQQa/2n45TQG
x38w8nwX7M5e0cIKbBZB5kmWms2To2Na75fiTgOtxfw7n/iHphBaVyR3QGgTqS1ZFSML4xULGYka
pEwY3t9PUOgPBDj+6pTKeNKSPJlVIHfFs9NuSKJt2oy2izI98QGhZEGubzLqDXgEVTooguGrUN1p
/me9kzT1Az6Ea8fcS9D7MkDipllexx0HP48zigQB4Z5L50dF4BsP0g3Qnck8QvnKFkWGR8yPccXW
so1CHmus2jV9KTbafTRNEu84z8FMsAA4RLDjpBVhi0zyL70FEe2hhNEkxOshSlL74wOhMdqLMRtk
IrBaN5paKFvnaTmnlzjdGFdbIEMpDLo2BJRJWwgkw1xbBgvo5iC8l/4YBEMOlPv6Nc9j8ONQeNTF
YsvYiek0N4bHe4hXXAVN3L67GLywCAhXENm8ChC8Y+BfNnzLsDIi1ghoi0cuxbZ16R899/Lz9ygh
bIHurY8bMM/gzctM4SQNf1m5YX68XvQkm2s4K9qeoKVMHZbPpxsiuaMBpK6ocFwzh0HUuKJu0mTk
HIKRLUwN+xUYm3FAGem3i0j2hAJhd47EXvCE2w6nexuqPlzk4FuSdELaafeQQPRmsqersFB/7SJf
Dq+dCos7Tgezo6uvq6N/hGWGIWBYx+9w9vsqtJTflu5IAsiMsh0LOI1+tOTkiS83MXJoyPWH8CvE
DwigBMBuAJf2G+DMatMyQk532VycpA71fb89kY8iPgawzCipJTuE6dZMqzyzkif7tqLSEeYJj1K4
EZRaZWmZotsv7/5EumCSYqB3CSzdvngPXVFh4Mc8Exa4Tfc/7B1dQs5fFc2gKzhJbImpL3JKh/MU
sjXfX8MfyV1mI6MB4HFTT4ZtXZVQsiBk4WYDMVDOMloeDHCF37mdZqWVTBjuRAK9hvmO54hqQ/1i
eFi+oR4sTOkis30XfgRBwqZ21RCJgiP6sQa/ayt3gp5+vHiO+3xvenbPbqruyYR9Z4s0C1ZJYDSW
FtNYmG3qjxCphElvlDCbKuQxWNwqPaC6YZe20A3ewzojYZdObcDUdNTJ4lce9dWa+L1BWEjO6nCo
klp7w1aRDiULbtu/jwpNeseS+JIQXbpclmsCdwFv7T4dKfV7T5M/FdUhap4YVSh3MLf2ZPIkcWBu
Eledp+dJ/cnFAMupketU+WOIMm5FmvMBjNWSmKnEs9Ac+h4mlSUpH+TESjvSHRF54LD6sEIim0Et
WYwQBlTEjryzfic5iDQNvcZlF1kBszPIOZm/Dz6RJOlBvSIjyjggq9XcZeAPyRw1OuQB1xITpXJy
ghDMlhojEPvch28ZCXKHUV+gS8iwKhwW7vVDTGI6WkLJ3HNbaUNY1DyntpswAvwntuIhnkDjboc/
R82Nml361ywH3FvN7pUvf4O2VlYCBfEf+1wHPANSPNisap7Nh/cN+BNCg+FYvymwoLolpuqGsU8G
Yvk3RmrSC4uO5oHNEmhcDhynVsczxtkUWSCRQpQkwZz63P8LGE88sTgRW8x2hUmtIzVBEXDEaDa8
xn9HuY23Nv7CkrHDjImf2nNaqm/uMARngHfgbK+sKptbdkzhsKyIdaYg1hHwcLdbt8HmBOcbfDbG
9z9aS2uTtwDTuBjd3R7JN88rE+qZ6jmfekF1JBN1RXK8+3CQspnkDd8ZBQOdQyBn7+z7SGh3kjFS
PMeo2jGSOtg/0M1ww6W9sYyTqLRqI0z1cli3eXIvTfp3YoWNGJ9NzXbhexXBIuCIaCU0uZmC5yOr
LzK1RmK4rF8MVHb/8Jen+kzF3WhjvgMHYpXjTBpyCOaYQPkkqVpmKqaPyuBl9vnCnvSPsUXblZPi
V8DPHzOCwgFu3LkXoYRRy/GOtf9D88MlNBwwUrJkgnRGxmCwkF0pE687sj6sXUSsI/OJAfGxCz+d
5YbW20rirBO7qGdVwpnIpAa2Axwk/ZvblRcs6Z7gIE0uAVieynIrkcrnKxVQKx+0ZBvsYtlNtfmw
/5RZsTfUhP/OlWbFB+l84ozSStDn3jnXYSVUWPPfKVDDDJCVmOoHGZgtGGNIqQ8ntUQeflMyaCg7
Btef+7s/SFUk16UNsfSvBOoQ17e4WzTz5eEEV7n1RDZliNlFP03fd11DNOMqaw7sjC6AMQefCaOB
7a6mzRTWq/spSRLiTVxAOVXQE7p0+KW1JgpI0aEiYhYyvJgEQz16LGo9FSSijFaCM5JtEPSxaqLP
BNgLwQ2YHLVld+K3tUzPGBRb69d/tc7TQ4QOdK74FJodV88R6+UOAWN0VJDUqeL3oFZVlav5VxEH
hqwXh+g8026EkD6Rl4yOl8sPCmy5qTsrlfBGFBsmUJKAlSvLsJ/ZK2xdBFSZGOyz7u3CUeKbT5jZ
FRuhVs6d84kqtC+QfIYmwFMWUHhDoapdAoKw4uf3niq2Byr+b5Vp3b7YuU8uULWD+161bYW4R/C8
ex3Bu4Fg4YWxRU/tTWohJ72CRyvTzbStEQhO5pnFzyp1KaIPBNl4q0EZXN22CXMvHaMdkYx4rEJ2
+OH6+pYWPQvzWvtBxy8pUtmyNNxbLQCp5UzDymPyVpnjpHxPTOILLo2m5THo/08hwlpI784qPm03
RrCjWzEPhJnNm11EaBS7DpaLRCtIZcoCcijvXFq4lAohRhvlBsV07PB40zNHxga8gnqU9zN+KpZI
6ufW3/J9YmkUdlegp2os6MDTHTqN0H6sVPe5qfVabpTsl/5Xt3S/0xc8lRDU8zOMNF8liBZ1iKHk
k3sDPlk5S3t6bVozajtJzbwulS+i9qqQxuKntSUWG5IUvTcucyN7fElxBv5DyRK20LBIY9tlOgQu
urOf3+qxsobVGtdcE1T+KixpV5+9pb8RhH8cgoslGdY0VrXb6IOTP9TEaNFozojO1JUAAh1kfHq2
mgJR/DeVokMWyy5jMp1t00I8cB0bBd7NFAyWjzwBXuwnt8N2aX0S2pKRdUlTfQ/Fy3TSmivuarU9
1byiiZ8WEyAGeDIZ4htE+MwjUy3yc376lpuTVLewiTZ0rQRc+7GNHth/J1DWjLq8qJ3CBkTmbrIS
8/FEFPZG6tnwcmeFVijEJNTSJlsV/AAljWfm+Hc1fUAgVBEe9AW+1GKmJfFCk1zZ9BdI6cqXn8fe
Y8MALpU628QDPXEt5k8U+5OOz8BBct7n059d2wjnrUnMJB++28PAVYGPnrxSOuN6yKCTd+dt3vHU
FmDWHzI/SVKlwuFwgb/frXUb5kt5iFtolH96PBrEwjV6Wc21JgEsOtNdfwVVk+QzeyJjpBBZTTBB
B0KeQf6bBidbqlqJDL1ZH7fy6xPeu44WfkcRS/fhZa6P26n2sWPN6vfaxNjrY+jk7RdptsGOYsHb
0cQf/5MH28MxRr7asSstw0UHpdvGLJ1Q0nf/QrDd94KhFFSuOueZXxl2zN6QwExlvuM8qgM2e9L4
p/Y1vpp9t1mxODn+HGlO72HOIEy3V0+vrNwfL8j7SEurD1LIFWvVdtHhywG6gB+p0rjEWTyRHI9A
8vtGcVTGmbZ4LsXyk56sxDiar52FruZmBF7pZW7wyQ+A0gVFG7oXdBhG5Njichkj3FdC5awQmLqs
4pyIU2o7dFaWK5acjgW4LKU1atk785H8iED9DrOCLKP7RMCNIIVXKFiCzAlThOXDdKLQEoUUU6tT
JrGt6jx+ce+Ul5nw0BwSQ8aTbdWINYIhDAjUP7VIjUOMupwc51/7xd+FthxREkTnGLu+IWNVfPmY
NsblMwKDVQQ3NrC/TDgCVwSLlxpwvVFyZaipsXv1MZa2Zju9acNAfMKu3+YepKfl1WUmjIO7gbB5
JH68NimpOidPb34gOh2IH9mEyrdvoNO2t7b3ShZ90sK1oXbAytGXQeZIRVMh39wLCk007y/OLc6h
2kZZF7Lvzc1bR9zPGbEFsK17JWfmKELdHCSB1sprqhNdA2O15y4iT42foqeG/NW7tLQyG6XHrSnk
VF6UhvAdbr2cSZ3hhFgGDr7bFxJfkRh0pvzUWu2AWWtdsuTVVrCD9/Rt3wwlGg0NVlXSBvD4df/x
cOaqxtkZiUfAJWza0ODnl2cfU5d3WUHhslj1lM2Y4xCDp6d1j7smfXpRcweZ+zESRjSHylQ/hH2T
9hIW6m5cxi5yRWNtnCK12U46CfkKKQJgILMLtU4IIM9urxMdVzdxsZ+pWP9iediu6gaEWM9A46LU
mifA20htyOIwgU62dbx+x1vDyL+FhbWf4yov2Y41hO2k9AeSVOSkD/ZL/GNiov4d8kJhYyFXZu6p
CqXW7thj8GKgoDlcz65Ne+KDyKHwfgHD0U9MTsXuB+QOdkF1S58mHw5gkeGWJyHqV9UnpO0kVr0t
e+YOl4u3IpeVD7RDFn1p98HxAXzv9oIC/L+3x8O1rbJASpNBAex8C7U2EtyZXpHauqNmMzh+et0g
zQH+60TxZlIMc/Lkvni4nXji77iGRmp1PeQZoYjFLoTSK7RKSHPid6UIBx8kNkUyKWfWCvvRnwRm
Q0j+KcJmAsuvg+9q5sSDnjiqgfGSxC3kjjWAPSd1uKGqf1bUHFSSsD1IZDLNGOdvmOcHrNXqbCvx
QSNdDVIo9TCp3RBEjTYFAfFE6C0P3Rqv1UmnmhkhSM/OJVBayQ3pNHcvCpsakVMgtLgau8m+FubP
f/Ja56EF57rbtCKOVN4zs3CG0RrkW9dkSDlL+NTpq33tihSJp3ZTVdwdBSz3Q8a2noRdHFF4pcf3
BFDIrwZWikXTemtkHP1hmI1pF4Oz5x8e6e/3ce/Z04TpyE8h6W6rn2FTkrSiqmM04k2kQXtu/mbS
j2cmLOCLENfWNPeUp0301M3MW3CjlzufSsWAOe8gCkZs98HnNiT6zJqu6MdK7G0/FJKB2L6K16QD
IU09Jn03cZaJVmtQJYiNlFhnUK/ew5HiYPsIG1sG5pumVu0icibIej1TgvtdtBq7WVhRXteySq7c
cA4l+keDajj4VeWvtLYHpsoEjXQupmpXh1KLvcb2oa+QS7WH1MgcOog+VIUHrbto8lveD/dSIWuJ
OWAGHReMWWErTu3ET5h+EajoRTK/x8Zf5b91HNfjgfkkqSa6LXtX8moVJaOwn1OhqZ5kIMlx5TWb
8uOO1Lsmqc+rjmWXoIR4J/dlZKj+QZnyvO/8qINpk76LL86i5LdwJ+5RJmtM2NUBWaP/OS3DhhtG
NDI6qSGWFI5yGk49kk4TqswI/NwHha3YodRvIXqSxiLeOKKw10pqqiefKri65CfPGrDDcH7hgXfN
HLbH80ZDuiYg1k2DrgG2jjP4x1aMCatKfzPkhXBhIFA1jbOpOMofSdNJQsKdeGqCyIcvbPeWBcy8
A/OWutjJlobC7J5ICma2/vZ2hQfHeo6LBZi8mnS0So/OiXFPtmj6abkmqlCek1vVrvWpbXgzSD+7
7y1wJKydOsFHXI9g0q+ZrrDPSmYLOfXWN3ubT25K4YxtYxPfP43p/peOAhjk6FOkZ0rttYVnkRSG
JxzBYspn54FG7km0/opXOqUXSwmcVHNMqt0EvpU/ie2gJurP0j7wQAD0xr3xShxStjgod8uUx1hD
PntS57JwJNpzNzT07n84yY35zY7bWaITkixqnK/j/iSGZyb6teE1pVFHlze/MBxJ7ZICRjk0WtvN
K4Jf3z7WocPS/Fyr2eEvXpfpmrXg6TI4LR6UgFl2Tma1M+oSJQlA1MY9w9X9v636mazk25o/XSbP
ndo/3CFvQqjCMoz1jdRzUH61Hnr4hN8StBYKLC0ULcIXBiRP6YHrquuUa+wU9zVOIiHiVd6htzJS
wYPg1LsYEM/VHm9XakZdp5qHlJQLqLy1Xqh2kJZNdARZ+UBnfM0CeO2nErlwafMmvMhHkQKFGijb
GkmMccPDWk8bO4ic/rxUCp2uGdmnO8MBMpJHgK9Y0pfYcnEFFYOv+e0ju84emRNQGpmRwOlc/ZXU
+dhmm7nT8yXOq0XQ6m4p4K0+JrdJHUiMoNum3fpmHgCugiyyldlZ2NvV4CXCStzZWLbz8vv9/GBI
1AajxzrckOZqz199V1m2+xfnFi4G7MSTc8Ud0TtU0Sy99srnqBEqFo93JBODTKsLlZs8OjdlURYt
Y9PMv8Xt+t4mxLHEfgsrmD0KlSI2BRRHkCvQrGj0HQl31JOzwbotp65ORj03qrMqIl6NHpHRKKXR
wgNRrq7RMHUO1EJJ6OWDZuhiFlFi+MEJajHnU0V9dm/MskOij1xVj6VTmv8ySMpCx4WLTvFOW53K
0aUfDn2hzvoCPoUTcFRNvNO6PoIABQu3ddFg3PQvZH5nGBTnzefeU3LyUS5mJJw2IAZ+xY0kmQfC
3JaUWd+2cu98cOmRXV03yZAAQB9bB33uqiPg3XGJ2j1T5mJlGy8nEb56Zfnj1F/xky/vc9wPJh2U
HCuKETAzphYuM3NjxegNAc5nLnQEYM+14PY4jiUSFp0Y97cUU0kx8kQ7dj8Mh+7shx0rA7Ib0tyQ
reKgRXf85/knorgcMKW+ocvAUaLdUMgBltA+d4mjD2QIsDJ5pAefYvHrk9V1rrpHVvigA3lEgHKH
goICp6nBjCuUZl1Os0NhbZpoUDbNc7nFHMuuvnkItScnOwWjbVWlufAdZ7uM/gZPggqAnA+ycwRP
ASzvPe+Ij+y0btfP5Qmvf5LlvDDsophaVrU80XP8c4vmBFaC1YvT/VGc0FsGZcUCjt+m6iLlXHIA
8aKFRoAranhG3kZtkWqhTSinQhEKQdAXGlmG18Znnqf10rnImNrZOUGizGo+XVBj+SvXsYzf4r11
wK/RRZKi4wbtMHQ3O3Sq4+2yRgC61K/74oHMF6SoLIpKwn6Vd2qIvTsQLyD1Vuzu8d0Pc2oBhCQ8
NglqK1uauAKwfimJWpNDiUAK4tPsdb+kANPD+NhiczYVjH8oiehF7sdCa4mygwRs5q7C9E+k+Hlq
21dTL0XTBkrkXC/v7DNRpZCU9dHsPKx47lGaShvy0eLw00IQro6HW1ryCJcuPhzPdfdPapbEl/fj
YUN/mr/YaUFFJ+OC5PFIaYH8oBDYGGHx3QLUiqACGszBfkpNjDyIDkMmzF05l10gq4TVhaq8UNoZ
KkzDdwitPdwh8sDYbNpXANwDYEBzgoicuvDGVJ8XjUw4gJZpjwCST1klL2X/alZBecVuGt5G/6CZ
IMu0GzyO8F8q+QE9v73IcOj0JalYWd4v5a8xwsSYzHAFVpkR1eeRXistT+kmBpvaLw3LLD9fDla4
gbGdH19TdHrQ5YRxolewAdt0fZiTpsuljGcqIPOT0UQoD63RHcKdzfvyQCy0baiOnBFK4rQjPouC
jYAVPIyyxrFFl2WEjNF2U7EykOWnd6j7n4P5oRJhzqwsIyvzjtv6ZGQiwZ3mdMIG6rcK6TfY0Zw3
nv73KlG8WOCOMRzrL649HLFQqKE4D++YKGZtqOw89iowZgNiO6e926v6QUb3hWDob+sYoj6AY0wX
3KiDarevFrf1Is9OfDLMxJmOMfx6SxSlMIkZfuVDhEE90evy98WJtWppkoNDTl/jMVGstsgAsAi7
C+kgEyvB8cCYyjEzLSBK2sGuj3rbRADkIwwpdqshgM/TUQ5kJb/Ho89BAw3+p15NCvM6T96QkHB0
zxn9IfL5/EIRoPzWehN+Hq8pbupOVlvv3CZA+ZjZGNq/IPuG5aufkJKwh23uqRxmV6maY4N+pwI2
jRdIDOl35qOfO/5w+ZH6x3aZCxEGP48BoOd6ywK6Ai3Bxq9BwNbTrI5wJQWXoloY3AMSV+yFcO+n
Zn+OR+4nBLlXXIwVbkYw9l0fRprZE5969TOe1DtJa2ZkQqBQ3pOGm9qkwcDWgOBGwbB0XcFisf56
UBsdJntpbb980Wc7NWWwSKh6bYTNTs07Y3L9ecFINiQlNHRtm4SbIAjiWMKZ53/iLoLtO7XUaOFE
dlc2ReXGkTB6AsHbWcdy+luovCkHtWaanp5yghpsFy02qxlQl7gp9nSjn3y4xfOTq/MCR7bjfmnP
mg31axeh7N4GuFqVsqbl2vSsMNGgQmnJb3RL6rnedV8HTwnYPUfBjBBoUgY7vUcNaXG5EldY2Wa8
kfanUzlf7NbOebVOu81veJghV6jWPxn2rUBkD3uohBPewXruUS5HUIDP4XhruKDMgc66NT2gAoAg
cM4ccxbPhdeVTtUXEWrz4DKD7TCisHk9sCSHeHL09wDlHPJxUObeZB20RjU3WxgGwBS7+IGwaebp
w1pWUIZID1ZOKooC9+Q0msaVBm8ty9xMlMTwPpsnOd2m5e751bTZdn8y9GQ0/BTV57S99TO7dh5w
GPoaNFYBEUQIIFJ5pcCDB2Ucw6JQd/V9mKT1EyY1GIdaNMEVgGyynr6CAOkJ7TesboFp+Wjp1Z0r
NugczpbO0ZY9Wkw37U2br7hYLN65r8Q6E+YIZ3pUmwKHzdiLV5b+3cHEaQPB6tixe0xyug6RCeZk
1dMMivTh489UGdu/kWyE8VfP+mcfPgx3hRGQ8HtTAW3BdJhpjGPDt24BThISYOJT4sscek5wkvmK
YI3NfpNmi0kDRj6+OZ6sxjtTyq220kmXpMYoKL9EWvOwOCA/7dKAkjsDvlBKre20CKDo8bSyNX+S
S1aUe/1gZ81AQyIDZ9QIGP6F7O5UsgdDjCkyE4nrxoggiSTKbT04Gor6SI1oNEw/jGXSe7hpmWGH
Qs588/zQfO1ZLuzB3Mk2LmGh6OmwaK9uVy+EBHh0rEYIgv8ZqEfZsFGMUN2YcNOU/TwcQPtvmxfW
YBEK2vJfuAbNLMhfVVev4oSyfTQcY5+51WGK6RfIbygWc2aSJx5j6AgriwyNCkK6NclkVZNxR69v
+p5pCI2iVigPdofUT6KJWf6tPvMBkmXeAXSobirY5HKaV84Ilhi/GcXhlGlFZXJ1j/ZfmLYxkUEF
wfBmGucKqosfBmAY7blDNRA8FSlRzhTKfrCAmIHvBN0k9g5olXml+3u8sd5G2um+j7hHMf2elzTW
7Ekc7WIk5Kz76TXUH20i/w0AGZiyDf/TQqhkJD1BTXUUUKEJ376/a6FIhz1RsLZs3kwl6HHxzD9J
+wcge1k3/dzjJMDfpPaCeZ1FIATAsX+j2cQ8TRAz8XRoEv86D/aJS34RYIrKjM74nWfi1BOmH6Bx
QANMwUtyAKTsVOnpfoV1ZIUgo62Sw3LMmI20Lerttd15WwhoE0sRmDDR1vKYAvxhSxIw4edDurAe
HnBTZIcljVpXnhQUlHNxv+wr3pi3RnI5tylXthlBU2iBZ802Ct+n68pStlXk7aq8UKVTbU0SEo7W
0a3DW7O1L7UkFBYKkcrM1XPZgZkwPJDFPUHR3CFBQ0uXz6Sez09Gc8UjhpkAn1+MmIN6m4ZAm4wW
8pQqusoo1radj8P/N6GG/FSVkBahplKM4JgPaSIf0uO2Mdjm2MWJeD2Cs1/oJPZltH3v5BeMlLvh
WnPWs4y71U2N1b4DD0zCN7zzmobEOGJiWyjwOUJQwlsRiTMY3FnXOUqneEDJ5+NGf2wAy9Z2p7nm
BDZhEEhYphIEhrUs5P0kCtoRlWZAfCXPrR+Rt0bTnOGvgbFr38xZt7hWyZip04a7oUTWCCTzh2xO
1i+8GTh9a6yjghGNb6VQPM1jwJxEvpzN7ZseCAMemHGfbK+UIYu/astxHEWX7GyOrJwzx60vkVl/
Zrs9rtXth7hqyF7Nn+97HFLOIAIMKcqtvKgeFJ9wZdFPB6AOQRHrM0zqbqrBicT2rouFtKkb+uwV
J5DlMs6NVAAWv5Nqs3U7a3aFRfT/imWj10cqc8D1rRVGGjogcHpjoB6XXAiWta25AzCqAKjtuTcQ
lt3o+D+N1WtUF5uayA5ylVO3y23sBBZmUUEN7Nhu2U+xk1zjS7ZRvVBpTBMu7GVYZM1g9EvfudZ1
v/iNn6UC5ZE2/KJrmHkACu12L7algQOykFVroF67VFGlu8dR952kRR1J+PpSS7yiBMMHXUFEtADa
rDj9GqURddBKBeDfg/0SS8K70Pg6deLytF4WV8ESLj78NpZY9ryHTlHvW1lP/kq248szXP2zbUlx
KiZMmczeDZdsazMuhdjlVNx67pYWYPXIlSI9ehfVhDApji30/gfANGLTqdOj1C38wE15Sylsl4h8
/uR6kHIZJQgD5IIFYHvrtLOw0KA4+v5vbcrVt56E9zuCHeL2/mHCwx91eUQMOOgg1qkpP+bEcSw+
iXazjUn6/o9g/i7cNKJcjPGN8hloJeW+awseJ1VATwo77MH2N/y9yJJRPixbbqylW0e3i/U/yVdT
ry7FemRJmyj+/zhA8Icn4nYYCF+A3YPcFlcp7Nku3WhdQH1queBjzFGAJaHJXMJiGStUfh8XYG+p
5GATGncX+63kGoOlP4XQfu4I9aqoUUVJJou1ssxEoMS5DZnVV66VlYFi9tcK3W8BWUHmg1f5QhSM
eN1reB+ACXaTo1goDyq5Vaad1siTmHrXC0G5SUU07XYLYT1fkB6WgN6FhwkY5iLLM/r8csAERMHF
2/FiYSc2dPseIU2r93pObor707VLxINzYrlo57i/z12lyTgwUWyntrP2K7AtDK2HiFj7dmFGgvfb
+6ULnOd2fW0wyKdU4yNLBFX9Nqd+H3FQqet88t138aILCj3jQ+rOfEHpzDGULuFAdK8j+WJWsEf1
WWNpbg5DPsiWd3dYoNGa9yHlbB1jQEsoQ0ryIhzVHN0w3onU3sLJDZP9xO8d8D+4zGCCCp1Ro86h
DEzOilHyx0mNGR14Al0FqE97fojBgHcVJ1dedmKdSDAWnV1+KDooVNoMK07fyarmx8Xe6hCREH7t
8pbpAMhYGeidOnCOYWJauNQ4rkRM9/OSNZbpiaGwfBFMA6mkMCa/XenCk5WQrwsxQ0tshGR14til
rzBepYfNmqYMQZNixBHJ1HFQOjS8CZjFiN11c7mUKJDZOqTQ/1vG0yFPAbMJYkRbtK7W2bKmcgdg
1PlW63nlNhVjQqx8U8vMwt+fET7EaGv7jN3StgDeYokP29faP+lvNkOys0c++8rnHv13GHS9Lfhv
5OeNTDHGJ2L9N8pOPaqioSeZlTQNBi3hWmywC5sr8tkKs2mbKibxj79c0GKKAT7F4myL/alDX82w
58LoAkSpt42ee43I7ykLZkGAb/Jt05VDUTtjvtzCVShnsO8vJ0m6tqhSvGV50aTAsZWq0JUVZS2d
8IE9UMpdt17wgtJSxrj9RKHxeA3jlliCsNK94p8i2h6JULRYusV08D8cw5mEU7FMzSlHof4pggyd
/aodCtM1nb8FUjiShub5PS/6XzwjPBJDVH/All2G1XlZP3U6mRYx9UFTNqEv/Rum2xHmiQd0cBvi
vk+IjDb6/fosSZdwVao7OHbja0257A8x6NNwajvWfcHNm5OChTc7SsvPG39MdtNewERIHWe7pHlq
WFC+cUFGxESQrqMMpNdx/j0yIeaBMkdJrdUvbzNctcSu38ifqv9w80PkWgvIOBxlLzMYh2OhFXvp
1eNvU4WsSjQhIkcZUk09t7us5aNACkLYIHtDCCtgiqpWS3c0boZoMeAuECIfHuQOdQwNPPGGJnU+
TDgn9Z0zIhnrCYCUM807ESAtteP7s6WERwdxwVLy2Zn2DGJ8IZI1VcaBq6w/rdUfjTJCuJ3ByDVM
WuUqU/AGuYPdN2bf6S71UVZ9E/nqyF0P1uSn6tfu4/ZMUqGc7j/6OXC90AEJreSAAKjVLF0RGfjm
st1ZKg+dnniJZBDgI0Wt2fD4+on62AYSe6u6HI3bu1j20/HUAk5TRVdTkK+d4YP5PEOU+4gYlKCE
9vv9LKDRkCK8GN/l8tmLU2YUxmVTZFIzs7sZwJBhcp77OHSqqjaH1DoKzZvF/d7MRA5gFwUdBDzv
v7X2MFVfbjwagwmXDclrZ7MUhGwO2Aq3NfJb3hu7gM/W/z9QmQUTx8vOF6ILL+5sNtc0jJGEPci4
SS2OIDiE2Bo24ZNEzqitMDI29RNV+G5XE2cpKJTevV5lgRpEcKt+5s4UPV/IzEz5OqzQzWcjkcVv
7Nztry1cnb5zb7nA1LdxtgRBnS7n1N27prVpeI0DZHQPKzZooZb4Ekue/qxdXtSeQ86Cko29irGO
f48pjtvSuqahfk4ww28D14jkKjNsONLRfUJ2GiWlub5v37pLSOq2SSKn7BS+QcqTk0CzvNz96hI0
kR3o0+Tg2MHYgqVq/XbDhYSjj84wY0ibynfgiY7EXx6zHcgzAvA1OO7k+LkYziIy/ORLqE2fx4/d
hwZWPDBwX7TYYAeOma4k/BVozjTjz/tdDz2dF5YEFbQq74LH0nW6j0tHYtpjTzAmMYfYZmUXPHjc
N3z2jAdLni0RAVao133xzoeqs132Nx+jsRo5/Z34pdZgz2yBf2JKMEQuJDolSCxZQ3R9b4Y4Q+vp
x8rVUFfhetmGprIcWst7L9mrb2u7EPdeNSRJEmzp5Q6EqxgAl3lLRwvoe5Vps0oxkiPGc72Gsbrs
aMW0O4fTDqXTeQihgYHR5B7BCgJv5KtZ2VpW5+IOkaogJXyYgphRyjtAogwGIcPFtcII/ei5zQli
3aQ75eGBRPnJoyTREwE4oLFjWXQPpu3PyqfysLKgSBoxCthuwbEOJPXgsxivZaTz3KErkt5Elqm8
exaBZuNwjz7OTa5EVS+O41v6DkvwJk3qFiUlivcpAcZuqEDidlOPvE3CKtxZi7bjQ9wP/xRCRm4O
dukhTXSTbgkNJDt/g7T++eJvBAdjWBgonpIXPPS01w/ZfpOPCVnB4veMomTKhVaXKroZLfu3fEw+
aRhfUKuw4vMHfrXUQj1lx95LDm17nce8tZ6lx1ad0lDweLnlgmWr0wfAHTeALvVY+EVoqqaS3+CA
hZxwRd4CmnzDPdYPJi1rTr979L6/JaMkU5z4rj0fSMVw9RhP3eWYryj+7/Be8C2gvrTrln44nagn
64RKSl3qL7O9f7bS24vV8eTO5wIuB2bd48uOs7l/U+r+HusFrtQWVbOHN1Ce1jNW0wL1/qA7DFDS
embAYKPcKod4wS9KCB6bnnoe/636nQjp+7zA8TZ9UwbxDqwJp/JjTPWC967kfNNGpcgus+Yo13a1
ChY5+sTnhKpnIP18E6PFfkchnI6SNePiB6cZL5sohPhlcDO1rOsC9sva4nyqSrBq3eEoHlGqL+fn
y8a4B/iLggtJXxnZu9D7XXD2mH9V/w78uiu1mDLNuJu7rUyerfwV5HjfvKyDZGD7OCMEXoodd8qu
P5WRqlDO4yhzjXrcnAO6vDjy/aPW3sP1+55Ep94kpqGqFPjw9Wq7aKda3QP7AoMsDmxG23bYEqEy
/Oy6kLM6duud6Ue6mFAMt1JlCLStbgBK5mZ17akOp4R2DczCcM7XTmnxwtnqIsuzt7ZtmU4uSwOb
4GigcYorSO8M01uZXGIig1v/PeWB8wzPo/epR0CLgj0ianebJhQu2DRGA9HSUBH1OeVAFTuBVB0J
N6/ADg9NogftKOp1EgL9omV8AS/CER7eRNkqTrgNrjrhlx1aluyNSr9ugnNZsDigcivFrW25r8t6
89cV1NpMgGXoUiCVd9TzzKOBlipzv0PZxt6UklVR+MaXJ2ThgcTTOQBMS0kEGK2WAR4LWwUx7e66
NyLy81i4vpWYwU5tDWB6QUo+6EcBmDT4YMikfJHcS4M5VsqlLoGuLvMG1fR8te/k3vDGiGObWbEk
xlrY+BSKU+GB7GbEo/I7tzVJBGkl8fJThLkbHWbuA0UGPz8dfDbDhtmkg0Cl+XMCI1Tkp0291lRo
E/CZCnMYCO5DMVmdiQxdvJh5cyeyqut+RAMZkIyFmeR9eWMCwxJwneg8RBTl/QCi59hbsj67QNWd
xPclEiEmQbn4zvB6eQRT8Oywc5oETvD4xF5SQoOHAFqyo1HSZ0ZZO8D4DSGy/drNALd5nIDpF1ec
RmlYW8YhHaJ0mMUEGsHaOdOr33ly+mXR39M8R7W5v2noL51ZYsou5RFTcMTDx+vrrQ94WW7z6vWR
uPo2O6B2mRo95TH8ubvLxNlnTVTbG5iq9YzijiQJc7eh5z04ZZlFInv0Gan1W/OqqOtOWrkKUfXQ
XPqaANildSs3U/PY2ZavVsKWu7M8gC0BgYuSXTnKc7IYA0Xi6ujIygaz5c2lTeqOrERbmBC+Lnfe
cZIkWJf7sbzgeJAkuGSKoA8DECundAKD6tXOWRVpEFcZlDlwyOEai9JdQY7I5hp00qEL0J2mnMFB
pc7f6/mzf6NqNsFqavZbuBUEZScboAi0dt1bGsxSvH8/CESyL1Mi84uzmOUWNy4Xj9CBHdken3uM
nU7oFjIoQHLtzMGfZrzMqk8sN7NuJiYzpc2ExAhVi99FrQRkgP1xHks7PK12JnbxoWdrpJEpK/XW
X0r+kgRHjYAaiyY7ON9+kUVS0AirHz1wJdYItPc7le1UKaPM5zarR9+dUVmJXu0eijUULc2IRDLX
kNLVxlgefPCyxZAKjw+4XPhvWSNmvwhmdXWPQeOM0ZWaxsNkeFlYmkCKXYOfNl49vtbaAMn39tEi
CEA7ja6cLiszrFNGn1Wb249PzyV/bEG1rQJ56PIYdR2/TbDg29AG3Nlo+M2O/NtgTpcZ+bB0VfV+
pL5VTqzxnLcluUIVjoFNgRAJH+3OmeTRoo4sPzcCq0c3tPayWwnNrPwD23JPSHtWctgpORZU+1ng
KMkUmQW0dJsqGT12MXrsSMbS75wEqR2m2ofsaBBwPHIvcPnnxY8r2I3zJXg/6MoyQqK8WxmEiS0G
e5kUIduLnhqRssRpU/1NUDtyPwJsGTCVZdhjB7eGl+r/aFzM0JgMogXJMTGpJ1MxjtSAajuywWVe
cCJQr2uEIm2159zjsArybHxSCD6ZWT0tdVBX7l8zeiJQB82Fffya3iysZuV5AeeQ0drkOvwEgwM1
A27NQ4XmasEgcGrO0DN14rGb6bMhhwVmekbwLGCSLsx/+y31HijenBQHG0RJMaGSzrFPVb/isHeu
yDIZeQNkovJ2MALH+q3oNb2rdo1lw8UwchdENzJnRYvVfHZzqh9mK1RsSldoh1SNoCDQ2k7j067E
pXXoBlZKC+YdNBR/ZMeroqPTMDry3T2YMiBkyGj9UvB2hr+qSpSQbsm5N8JdtxWDbx/gp84pYt2J
0r0xDULGh+47rM8YsyfQYesAJ6DaXCTt3+q1cxz4E3KuLbwc0RSx0r+5PUl3RGKdkK46Eq6bF8QB
nyIoW6DgAZb3qzGwIP1L6ca9ViP/cFmzsyJD4pQxoxMZIvij7g0mQQRBptFVzQJF7qwCUtWL9SNX
CXlirVsVYxfLBlMpmPfaxQeQVFfdrjaPf0CQ3yIKgTpxGUs6SZJOkDL7gHIqnmdwGbPOZxYB6tlp
2oA/zdyAqxaeoDs6gRzPmPMPVzQdeI8bM7DX2DuflBZU/WQ4jCzInl7z98e69jKx15H0+rppBI+8
ThDRZtZZCSFwW5CchZsXbN5ooFo7IJmedo+rwsRivDI4zDizl7mzryrshTgs6A9ZhtYPLt0m+7N5
9ZU02P4cdUd5RZTO4M3Rv/ScaMdM9nQCXPBWv1/A6yH1WlTc9fGda5rHTS0c1BcE0sKUFm8yebYa
Ujcus2BoYpPZIDLheY18voQPgBU2YWkQsxXTLWRzvhp7wl2yslWeH6iGqy/YeHjFlYt7jmq7UYf0
JkLe0TO4Y1CtEBKqly4R39Nt1GXXPXUoH9G1ryiPGp16Yya3LsqxU9bu4JcQ2GahhxitAgr5LEZ6
ecExTWCKQHUz5h61bOwfed0fB2bSqfJt/mz8bTgEArc2yixc4nRyP0/4iLl0zsUMGonS+dbKqaTy
Fka5SSAOAcjrD4AmjoHKypTY5VR862tMa2CdOScu/C7ktOuPy6XK7wJFmM1mgP46BJoH/eufO0PV
ymgmlQ6KtW1/G1lHmirbrnL/U5mx6B6MNpmoPv9nGfAr0C1WCXuftLZH73O7WteWx24HQqfASL76
CEnx5TcpiCVXnoKHBnqIHfTY3nszIQJHDBRJBT7RR7+zBRDkHD+hkOVsZdXA0f+cYllw0ND0A+Th
bh7q8rJ3i7Hk8i+zECxBthsw06BESWc6VLxr/TgnCx2xpueCPJeb+Z8TW2+cy+xIKfXrfBE4CIso
XGpIXcrL+MYucwSKN6/EYyqLwI4dL4nqDeX2kp5O10egJHwkiYGa8zRSWHquPejfeDqmvb5ycLQ2
NdprmH4LFBbeb78oI0c95w7q5byHZLC/wrfADwFa8CdS6QvJtzVvExCi6j9u+p0+oKsFeFlFwRSj
G2JFhcwfsCDMU4y/y0jt/RQIzG91G312h6huPjy4pR9tuSderTLfo4SMG++kb8QOoX4WUU731f0c
UGVGVymYJGAImvXv/MsVsHJAjKJa2pHk2bhjPRSAlplK6VGRKXWcTUkKR3VWjsc0LPdLfbyEdR4V
61YjNe7p9Npsm/JqBXH/e8P/iRv7v+CWAXZRCfGZ00v4XC2fvtsjLhSsxdBWNmGkx7NU8+VuewGx
TQVdQGirSthvYnIs2pDQ2whyUbhMVXNJ99l4h8/9hWUN1UxhrXxKA8/1Y+LdMOyAuNOUGGa7CHfL
QJ6S/85c7VheutHLMx/RtqZPI16WwSN5g3jCtZfTj/skbNYtLVhtuy7KTlSCxoeq8o+TmUAbC3yn
0Hg2PqCk8rPWHwNgrk9+/6P6PfH9S5qqsYk6tu41dFo/zm+Al99P90tg78V8KD1kdaAgqKRait6M
dcpJzzu5s22R/jJxWjJYV79/KHzSYyxjfAttkSKaBlUhEB7i5fNkR7eoFPOt7Y0QsMnX3ohC/vwC
yq6ICyRWTSOTPtkf9fHVfn1Ze+ciZSebBCn9efjk1sz6BIk+y9LhUXa+bVeRlcPuSr/aDeN9X7VH
cxzdRN8Y723dXlzTj0e7iaK/NKwMxKn8oJSKl2IVIjw9AaCiN2qizdyMT9WcA6qQOMG22Py9cR1k
FchVcYFWS2UKub62ShdLmkQ0lJw6U6oi8v/tl5/Kq4775UF/21moGWWy5dfK4f+ETSbQwcSxZVvq
kvO9GOp6eKXh8rKosueTU9jmd+Kn4hOTML30/eAoAs184gqIKY7Dt91CxtT1xydWFV4KvvKKB5Dx
pKA29GZvZ26IbsE+5hp8oVDBVm1BNoYpVIX6PNUb7YBiyqdzftOsr/A5RxZB7ka9v3xJYfxk2iOb
IKoFCD5B+h8wTBQxhY5lJGcycAmvWDPs/ocg7VU55NyjZcBCpBKAMSDv0NfnAKFEdf7EBS/LrrEy
jZ1CWtNf/xTl6wQNRKka/RaNBnK50aDKMG9ML5L6X/0J2yerdsaCb4FaSpV2XmhDhRjv5OftDiiy
NC834mY/olK/n8gA/FhjgehbKPi+D3cczQzMwTOQJ3bGJ+gEZOnzf2YgY40peEYs7jW8Xfiu1v84
x4Vz1uu1wucyH7rP/0CMaoixTw4bkj3S28Etd87l1TSiYte6vNBQnkxCWPYdJ1fNJLFlZYO8jDH6
+A02GzWnWAMRHHeOtEAEtpr39uOhkRLnLbnHjDhc0UvUP0WuI/XTX+55uN5iHOTCugMKXn4AYwc4
GKlxvTkLnQ/GGIJ3Hc9AEbF1v/Oph5toa8uH37ATMQusr0HeN26WpzO4SUQhAXQC+ivpotUbTE7O
mN1kz8P85xpSCPH5p03OQwN2Yka9CoJRqlHPL8zIY22rStni4ZD2HycZDKdSEv0NutG6305PeEud
J2l/ZqKpErgDwNLGm406NXJYqRwTvBjc+d7p0CzI43/y+XW7rNVBMU4DlydpNdR2RbTUUdVUhaze
Aa8iugT2wXdUePo36bYk3dGyhp8HsgJ8ZXHnB/XxgQPrApK7hhZOyW1bQIuqUiqik+gmu3RsOvEj
RrUJAUxDksH8SLJUigmOPMthQ8cwIU7Xx3Os0tpSnRmcOwfuGflVf7+l/48xx+sZaROHMSUzS/Xr
7OrJxEWYaIEZcCRGve4sNIMMPSwRVfhu9YN2tMFRQvdCWjxPyQgBwbEYWbqIpwUC3wBLxbLi7dFV
JqP4FiU3vVj76804L9sbyJ8u6yLuMHU4JKMfFnPTCystP74b8o1Qo6XvUZQ+PT4a5oKTIn2Qm5y/
CbRZHK34t7ADyCMGXv75ZZQKSLvfVdjVgLcAkDxMkhejfJw7hFmBVPwWxwASA5Bwq7419h4eoD/K
qZSLeB7WFO2RJ4/wwTM3D8lKIV2ZU8aS8OeupS9dNH3sfjnKGrUxZ6gQUO9pCzto9u1G0bPpX4Hc
sFaWV6iXWcDaYhSt2YL58WHdtVwpqIA2Mse+PkiEOWwZJLApuq13rnZoTIB4c5o4iwdkOJtsmysK
wANxGGPctc71rXmyy5KvkF6DQNv/AiXkTtJW9eoLBxQShDW7WOkPxUZY2U4hfMmQ0sooWG6IF0el
gOByLpeuF6uAjC1vMTtACi5ROplvAk57vs5jH/CdH16X1OuYP1a+hAvOE8l//e8JmQnRMFJircvs
h2Nc/2sRyhyl2cIW5437gDRcGGeUo+Bagx7XZnYGK4iubacIzRyPFmZPy8WPkQu46wF8duevuwDa
bSzoDMrcO5m/bad88IT4VmOgz8e//0279PlsfoDefMdSyiDRc8au5zTB/cuOk2UNXhbU7xyz8B7t
sQYhgYjXgnv3yP/cqtgCEl8j4k3lGkmtVyidNMcmYu/p3yGBJeEcQtRIPyTpvEeEq2PKfStCFgHf
VOx2AV/Z9VbfgoGUlvoPJIe0QgIgt2+npvY2isbHx9IEdWViWbxK/9ed0KVEJcQSh44msg+Ph5Fg
drFSRDd+42nwfZlo4O84VJm54qkKsYVw2cW/h5CFyNenXqBtVW3rfHRfu76vgol7gAKyYPG75Vat
Q73ZDxE4WGJ46J8RQ1r6zfbKgMq9iB1gQZL87iGF3RhodUSfz2kgm2pVyccQDsZfhKpA6JLMI6XO
d7p+Tmoqy2KOr6/GsDDxqeI4AzY9bAqjKFQc+NTYJZMviPbfD0aCvNiNYFoAX7ApLuqS586gNtoN
/2JZtG7LW5a2jZAVgwt9KeigJJWB6oLD0qS3xRvYJ3N/GETuQP7jR38a9WMp7ut7+Ol8dmBWukeb
KX26IFOVEdis2h0Md6AB/0wpS9XMtoX5u9m+S8HcVcyKVGFd31hO+0oc+C49K34Bp6TNdk+kXs3h
YWexHYfd2GyM/xeAER0nYOADztVj1xJEMs5zgALoOQz0ekA+i6q8Kiu4VfyRGoqVzbTS2QVTN57d
Sw7X5t9FsZ3MZj39O+ZjwUFKX8MV8IPQ2N9CkglrgxYNr6jOPqtbs9UKADSnWfwzrvoDO/2zZw7S
5qwdcaA8VTelLNDe7jIRQIkAfIY7iOzjnGxboS0lFfCiwaEVZcSP708IY69y+Fw7/WQ0efgBDBWs
jYUKI+01kWbJwFBXlhC7A7d4gXH+odd7Yw+A0jGtZOjxlXWR8oXeHGxexn+Ccs7qVpJtpz9ARqJg
yaukGSrjfkHBu8mDurhsYdnoQw6lP22wltRWFxbHE8QkrnsDw8fqYseDj/hNHces6yh3ZjR0V720
UbAK/n2BlsbFNnBrBmpX9cB8ACSZy9rA9pCklewQk6/l1nHjLkQhbqDTaMq1xRNb2zKF5JR5zgHl
vk41E3tffc9TatUPlF3gpMwbM82Y7UXkWkiR7UDGv9uaoDMTsrOrHks5I0Dy1G3Om+t+tcYKOXxa
c99YEYVr2V38ABNBXcc6TeSzYpwYf7gt/gxITU+nBwOJ/aTa/Vkn6h2IKW/r7IZmpwglPQETRzSF
S+gHSqVyoErjj3WiRQWAd5+2nCMxDME2vLVVw5TJ9AuzELujupqSFsQKYWCNikNS7RVmYS62D5U+
alA4gBiuGfCjKcjOV6KKeOVeeEa2GRcUZ3jcA31w/DGmZtF2urjh78qXTngS4yy4LALMOXNxbtX1
MlL2YepQfhRevfUHKxWR1O2n1tC1BArDpUhvaeph+wtssI0YlTipCljMBSRTj1kLEGj1jOGz+LPN
vqjtgRg8y1zis1GeV0HiTQuuUTWZ9bGLc4q8y/Eya9Z/zmd8P/QJ2+0+Bjra0rqe/AoZ5i8rb7XJ
LFtMIULPWUW3HoiauhDa/RJtBjRvyIqT3e+wLsSsPruwcSOV8Edj+KeW0adhjfoMT7gbaYtcUANC
VSXWEHSbobuEmBAu1/4pOLnzc8yKufNVXO+rUBctHvtYTA9t175QZn3ICu/nYQ6sOG4RY0+byYTe
uYX0uELeEnfNg4/1UNU0vgq3lVGTz8QKnrt1IGTtpSmVDJWE1oXYwir0X6aujTKqtE0hpXqWRaSl
3gCGOvb127OKFpDxPIZyXgomNBcN9bHCpRXGescURApYvpeuA9ecbBY6eVjEBZhiUarQVs+/dMR8
WuMOIJ/RuRtf9ioP6AsKYCufuuEEtRDR/gmnHUkBH5Pa1YV/7Vy8Nl6HSuUdpEqCLES1v4l6YLd5
6qVkfEeJunoMHv2CxRShTrv06iLiut0v1f26nUX+j6pa6sYktRuHgVERGNsxN0dxQ2vCIoYyYglZ
AJQ2dnSgdpA7iy5ktl8YGsLOrLrySwffA+MYas0eyG5t+QHUkRPOhkZzbaGFTkmsTuZxSUM6gYYx
PrJpR5davmzbbjFFi+Ik3ZBb6VMzVXIj1cdfHU6ntUgKO+IGdfuM6LF3MQ6n6/QODFz2kDKv+Om8
8mD/4+bO3McQzXagEmQDAaAmysUHq+FGGEXMVLw0EUrMitANWwA4oBvmNbdOfRNwPEslgfMKVaVR
T9GTetu8eFU49cbAkR6A1RvV0RTMH6maAUFPVdMhKDCnROmydLasAIM8PYVIfo1GkJ6kEaSJ+RiB
QSq6C9avST63afd7k0z2+QHjL7NwmkJX4OQ3vDTnq+g09gFhNz3A4lpMniw2utmpCeqnclR3O1+2
QbUE4YAUgZzPmhY2mH5hEr0D6yzKqlcxcRB2tzpR6PHU4uVMWHpJymajLivmeCKgSzjCStJB8lLi
bbnIl0gKs7nRcnRQhrUff0nQSTiSgk1YNpv8ZqXLX+wwYhw+JrLRP6xm0UJFxFg+ca5buLIkQ+4u
MYFF0zRkz+hJvl6blyCqNKUoRVfxfu20rROHeYXpTnJU/vOpPMVPN1ZvoIsXKiyY2Li0eM57A2g+
z9kkVkoprQIRlhZIhaOHMO8zLib+GMzxmWtCYqDuPX37XELSwOFGxKxN3UmiDRjbVmFJPvbEn1am
EBToQlrNPYJTF4rOMJu/U+hcnpVumo0fz5ScgKhOCtEFthZ5vqXMpR0nvOqHdqe8ElB/6RpJau0S
ua5l8EuOBI5I4S+PNRjC0VtQOVQeldnVSEDAYG1CwJnX54hL7+tSnQoHhD/ptWSYk11I93IRIv7K
+jpnjEItXQv9y8aL2XvjBsRAMO72H9sP35scjXnHNtYFEUFhCRruxmbRX0AimnSq3ewp4nuS9TFo
VuwtwzRdLFwSRrPqYbGMsQjL9l+68iGANjPaLQP2kMFy9ehVpvzcDkaZKsc7w9romp/a7DIirUVn
az5NCRcXnGCwb1rNul9jMeNOTDx0pcdGl4NsFkVuvJviXe5BQl78Xhq5D6KWSvMQ3x7Of6RaD/b+
ANdBy8FmCDfeV727XEowvnZvYF6Dkrva6q/NU0T9vFlpJ8DRZRP99/3vuTscdmHomoq6w/09ULSs
OzMlWw2XLNQmNndaS0Yf/FK54vL+j5OBkEVJVi/YI6dy+c0iVSLXXwRfbX3v77/qqdvr2nNU9GZG
43ztajZwb2jUB2jTwK4QDtudLWWzPdMZjUQk41OideKKQKYySvtPdqybrKUW+cCn0j/IqYnmATBh
YrwZiUwEuT/Du2oN2QKa2sTsTAHjc0jjkSYzymmIaCbnmNHaxm8pkFesco3gCCg9hgbttHPoHcZw
hVl/fZDP+w39NDD7pHMwOEs3Dko0REcvSMQeoPFbXhJPNthrAtekub4mTziPvD6kao1pSeJzL5tG
tb+fN/9AtUOnCzNgyzBfvuOPLzcsd34Jl4lnrEaq/QRs9B16HS8Fz4k6q5HhkTuRkUMaMnMRzw4e
ZNtzyHV/3s3fPQCHlqUpjDm9XVOCNWFFz9Djj8mqe4U4tMH+lKb8qGgPTYsq+kqKUQunm8ZS2Ny+
SJ+iJr1guPoSWL+TSPB71bpysdajZBOedQfkbQGuzKrev44a8hC64p/yMx7qQ8ry4TM1gIdGpbVK
ELBP6AOBAKKQK1XRgLx47d77ZPbXoKZF3CMjxFkBfhO24XUsuUWgU9VRcg/18gqU9FoXB9CFVhlH
Pki6sx7FbLK/Y37l2/l10KAXfaP8VSkVJr9E9eUBzhVNgEhL9QGM06E0/CPwZ8n5WU8Sb0oOFgHn
g3J9v2XKKuOgzSsc0nxa3Tfw89fJgWY5XY3WmHKwTWm/KfniRDXFL2tZX/HW7Q1yJcqlSaJN1pji
lWChxgYc/YxuBXaZDP/ARE+AyAuZwWFJ7bjlizY0rJ/Y1Ato57t0i8cLKTGjpxiH8vmSWzcuoAZu
2Crxygsn8h5VzQCtFHOsU0Sc33lt24knyrRd3xYfcmOhNry9vXmI1BNzoX/3vuhaJOzbOqxjozsJ
zfaYrfmNoEtOzwAxCVkSnaYICq70kjAAOisu5uFyNmmywJRGqJqyJtDVw4azjmrqvaS5m9Z1fNlh
lKHfbsGpszOnZTvk4S37T34QDQbTIS+gnoWRUP7yhAwPRsSIiSRkEVqj3wuPvdzinKz/FOeV9V43
v82N6FCcIu8QsJkb0GKh9dYYauAnEoTqYZFt09pei+NTDSsEuskHULxRBBU2IIiB3nkbp3E++uuG
7IYSykz6KPOO7XsDK/NTBUGzFX+WWMwXjZp0m6/rRwf1R7L5Byy4uKp0dwJJucEovTmjrnNM3gqs
YZ+RnUYduMQ+8HUCeS4JT5h2rG1bvAHOBMyGu2X0c1Ick4qlmZ8V4T+7/t0uvfhEwir9t9z/lbej
ZWi2y5R+P4WVR5cPk6KBk5SbQsDQKaDUxDYvR4vWpDxFy5EKXrYMN/yZli638BXY1UhqkLp+3LVN
wYVRxpFKwCv5PSpl7LsW/KRT+ekrfrb+f+FFyecYBAyCqdJsQ1MPJP/Y20RtmnedOgjo1UEGdIVQ
hxbWnysPzbPalB1OfATezQVMvk4G1795+kKsiFupb6caAQ4UJpPuqoJeFQGFP6X0h3JShBg9NLkz
Z1e1odydTZ/7dZE9+f32/c12Zlaq/DO690vn3DkDiQyE7XTWmHusQLM/LXXArMXYTVvKNk6c4tyh
QMcagghzUKemWbt7m0s04nKg9QcydT/rdLwfHwrUol59OLJf0I3DrVA5NxrlImjDQL7KtpdAFH3e
5kYp1eOCZ6qwGxHVr77t1gkvF+AgxK8j5SfzcZr307lfIwt5xu+zsFIdV2tLu0EvRIkzv1tZqTOM
zQvI9fKVUKJdGdqWVTLSzRaI6Qe/no50CHCUtexvdO+hXwcHgsQzbUevk/EeKmL6yVB7xvm8GDXT
LLxpaqxL6YHgSoQ7nCxoV6bLB78hCOlVyURagevdjivl4vL+yzqlTDo9HF16/4vtIIoOnEWxkgae
NWTbF+jgcJ9A3WlbmRfI2q/XEX40u2l4Hjl+R+DkW5stLa3zVIPOrRFamoW/fQgQDkq3471NlOYI
37iXVhj1+6cFQsSC9xIEy+4Xh38SGnfsuFyRMNgTTwPa3aiefHCr0CPHKL/m7NOOMYUz2YMj1PF6
M+4oxEazFHJoVt6su1NoE4FJXkw9giSmbCGvmjiviFlgyGiUAtBdFRsglsJQcTmQa/0//cli3XH0
6Y90D+HieIT4ua6AXQ4r1MUsSDaXV9HjQMkw+j9PmTL+0SwoKStUF/WnfdGxsAF3ocFJuCUw06Jo
GSd+QWKbZSNKIj9SY5nHVgLamSKMafbjXCGxVzLYzXhETR6NBx9YfdGY+CX0nlf9/yzqxj+9TKeO
0BZKBEg8FctLwARrGTR9T+q8TzwOE31QsOBElCrKR3V6nfl0n6DB9dQYTuY8HTeIwl1zGZWrNjox
2HDLOES2U+hsqkUVuVYovfJGf+kD1wG6XI2YmT7VOgDcSELdZLV3gio3Tse58Kz5uNVwwA7Rkv1Y
7R5MzP8KysFH1FlfYL/YcVQHInMljters6rHg7MQwHKqUwNUmamgBSg1Hc3EK49x+yzCplUiYIwh
nwDItU1o9ItL2IvZNWlu32t38be1AxRFtFnEcM5OEUCeSuINgx/wlE2DvN/y+q+AUmGm4ecu1j74
byXimDQBUzGWSvwy4l4t5q9azY+dea2M/ZAL4WIe85lG477KHBSyqsNcfKHl9JkKArkebWRmTKmk
JlwRtwGqLRLchSHZ9kPbPs3SdE1JNceroYe8pQGAEYWWW3X8xYYQLJyuTJJyzRc7nrmrmWPe1ZBF
ThffcFAIY6OzdbqdDBdaInYxKstHFe1nfSOPIF1L1MChadi2OevZsdNrysbVnEbOLRHAve1GEVUy
FrhWwn51BhZT35FhE0x7BSTTvUwoUytSBBcFfp+41pxhiinyRNToMoXjgqc6wszpc1f97vOSTTLD
1ZA3QJFZEE8xbfJrJtfEDl/eMeqBr9Z/MuSR8ENtSBXOf3hpncbHSNNlW+MYw7QUlQhd879xLSJi
tjnqIOyWkMdcszPzQWeKcfDER43JUYaP408zKMoguUrZSGgQ1tME0Z8pwH/eNeuH4R7vT8uDP900
NnsAT043QmJupCL+X7twwktEr1MVk317iyPplvsaINx7Yd3wBSn5S84wIRnp+4eDlbHBI6zodTmZ
0TmJpOwNX0kz/AgHBEf5SEfNQ6EjsevUNIkinvqmXcR8GRBzlcrbiCQIUoHpnqhLywZ1Ch6wCwQe
QdORrNYm/x0WBZbRsSXoSDYhkWP/1jwdXwcl48pGHslEjv2Kx30EAdTtW+zcWeQW/bXhfzkOBXII
3w+2zdXaBllS0RTxueaTtewevLFqY+F8kzTuh9ji2Dsjv4uvmoQipbhRNDGdpiSGQdiu28GyuIG0
zhh9EzEACYif508vKJZfykdQrYLCenCqCqYzQhYFXdb6cpXLRiF3VerVzlZEHO5wBlLazYwBYtBF
gby3gD/3oOR98TLSHLksNMKSFpWriugvvFSJqMGkNORuF52N+U9rhw48wuqgfBmGSv93Gdu4Ir5W
ifmSI3qZHqwCVpOeNT9Dm4izgS9qqMnEpV3FbBsF0+jTFpplS0iUyXKX6j86KUU32yi4yC577QR3
fPH35FpESANzLBJXFebM8zq4XDDmrXTZwifnmEdaUpKnZ3KiP0Br8tL86YPRvOrHAnQdqXhrgVqN
4k5eJxNtgOlxHCQUby20nTfPa/A3T2knsdrAHqd2G8A0mafm8yM1Mn6ziMtg7ERb3WJPn3jrCuu0
oQp8AWIrBWfajXIbkRbOk+w4060u0OGvvMGm/NLUHjHYXQIjvtrMe0SJJWIoefXsba0Sj6kMBVsv
fYYuLgEkK6zaH1Ki7X59IRYPQ7MotQ+PeMiJRiyKMtEcBatyWIqNPBeA97WPv//dWPVXf3rSlH1+
Jm2RirZ+t63Yuq3BuIr+dQrgPb5wxAQztS5uJPwYJJCxfXMj70/uw33EadDcHji14EEmq8LrHVst
bQFlUOqCcu0jpH3zt0PKWhnLGLEXQbSaoWdzrdHNy4xsIsLXStS3VWA6y8XNeO/OOdj9FE4yCVMu
C1RpRYqc2fhzPqGu/A4ssikXl8Q0bE2eJfJzyul0xEWxAevcN/n3nVumEtv6kjpR+gqV/RqMVJb4
OI9PqIpn9X7Q5KsnLHq+hrRh9QS9MDCXLNKcrjH16YYMyRNiXwffpiAkHKEWWxi0o+kkyy82iV9T
iEPjtJjHAMUGbnA/eApA1Uqvir9Lfg6ebpp059zrLowFfe72LJSpwABrNTT7vWCWS46TkVLwaSRp
tMYrp5gMofqnw+HyhXDicPkOM5Vtguw7Un5WLRuFkuBQeuUBW25I9SkVt+99Z+uNl703duFv5f31
pMboCl5ugiaIB9Uw41PYyVk4YhQcIi3Tm2Wg+BdVMpDx6PYBoWlZGxw3rRKpDK266iTYIwHe+GhP
Bp9vNsW8gUrBFFYutb+MtxjZAq5L3vxuN2MhqNWgN0iJ6Wpd5U2cR4SvYxLvHWPp2kPJRiXoZZeq
dzyxEIBRJUpXIkc9zoK/gsvVSPxd+Lp99KvWg+hBQPvW2iiFF6di74Ko8EdbwIAIt3tRXkidHxQC
VYRbmqVYFiZpqKx9iLdOZAjF1HnWXzHgaaQg2oTLgRahCJQ3yfrmoof/zQs3CC18h2HFgSD4cOZe
NOiYhP6GQZkCEfPJoIvd0jL9BQJxGjtCDWWNMERC9i7PcOej3B/B7l/CfnrJ6HPupPFJxkP1/XT9
glFicYifW96KSicSudC/X8vqngvwRUTAWJvzmfDLYMKtkGtacKt8MBi09WrpSpI+aDYZODKzU+46
yRC1UiEeicHjZqqUzPoTcunrB0kS1akM6EzQvFr00G0QdTFOGY+vrSCZPW3o+ktmjjyFMapXBD+p
A27nOUMlz2Zxf7OmCdjr4b6CsD3ZCLIqzd/obxiDEenpGXUIsq/vPNcsOPGX3jrWJx4IdnM3MpuR
Q5upNZnMuErFTykvL0382au/8Y+h2XtXSJsNUHo2oWtHw1Z7XgdELgfBD5KSmsArgQpKPRDCBr1i
L6x4vZgP6rFvb1vWq7YYXjSpRo/x4QyDnkQk/WIX1+JSitoX6dVO590uVkSkvkVLEiWPNQbZpkAD
F3jwxBX/7hMgWnyWDUkTO0D0PosEK+bIbJgjAGk1WrROYE8EBH6pEFepZsijo/rkukGMC4UisQ0o
+ccvAJV48MZoOcqzl0QzTRmfZfmLMc5vBNzLWoTBYmiN0PmlMyYxlc8K7eK566Qh5M7EY/xdsaUB
DJodcTcM4urAFVrtjCsCroyVI8hXRKHO6YPQWaU167yFj1zrfPZTUFdnzMKDH+W+Suax/L9/F87k
whXZ3wW1TNFP3ekM8zjBkkc5qZSUkpC8OGhVdgMVGZlreY0Ted1UCwncuFBCL6CUp0FR7FniE7Nv
GEcrsOXE2x+17pArpcBzoi4CBNSCu1JgfXXL861d5RhLv2jQHit9BbyXMFqjF4uzamFzHd4/8KvL
BKOsols0QbAaA2QdqtaCHaLiISQYzcxuUy61ATa8q2WKbW434TTs/AFBgBAOkeOagG5MX4Gmwa8j
4BLTSsr0uBix0QsocfdWYBzBOHOgAnxz0tRmfNF6JDrdavKHZHpQTiH5u4EJAB0Ilf1yYZH+vKXU
OoWXZ3Bzi2Fhce6pcCxLyt9ilUWAGmvZ07l2AqfabJ4tEpcctFDX61UT9Q3HgTeRaA2QKWUbxI/l
asrv5MYoe7LCJ7HTIpI0ZwMCbo/WG/yagxo6mpLetsvG5P0jaDiW9SIREm5bvGRP/sZxJs88+F1N
2WaJPeCAFn4YFgUwkkBMA3UqiwR67e1UiUlZ8khwupRaWabZOXMnClia+dTtEzF7FNjqzz7xSSYG
u1hBiA93TW78db7SNWdQCpxvnAHBnEQrcf0euwusp/TP48nsgXpvVoyecZV+eCv/0CfpcNu9cbk/
4r6Q7ZGcXO8bfw3DiW/KJgw/iIWyJRDoEQiYqbvmtoQxpDLGK6qWDdtcHBPBGEC8ov+O04gFdiLZ
69sljthDjnTpnr4m5UEY1ewAaGYo66bt+AI3CaE+i0HooeiSfs+FIa8RK1RtI+Jh+xJgWuUgCOHZ
j3lWaPFqNEJ9x8cywBIYJy7uKN9mB3sKG+dKUwo6d3hJTfOaCp4pRRe6+w5NVJeZaWaUBXUPlmLy
Srwj9FbCaC/wqA1uHcL7KMTIquXEP2vp7nyOAG0LS4rfvsNkirQxKNg0Hee0YJPQVb2nQav5j95y
EEOYOpj4i8JShjo0a18MQzOGwI8efzYB0RgyFlXpQl+OLXuYMUdZyNkZrYR9h7m0ZAZ3j0fLJE+V
7dcQlJVXdcQQziLijeeKQAh+BxM30kSbvxqDS9l41hJl2CfYamt8RSClMf+O3jKrcz4kHDdou8Iq
ejlUQVbaPVi641ZOZ+QW33iP2UFru7vrYycCwYSzCM08m0DPcwy1l2mApn/7Kqu1Kwx8dDTfHrB6
x26kgazHune7kTlaAjtFlLS4+nBc484lGjqO7Sxmp+l0hOL2FIXQ8C9bTuTl/fAt+5cvkMIijkLO
kvpPNYh2/jzkFmqyGFt7F8mocTa1Ja5r9g1WBYvXbcta4g5C5yxuKFbYPc5QJ3xqN3W8M+kVkfqL
Sm4tYxqi52BiL19bNyZf2NG6Z5k1Ll8zqsuFr8WcmPFauYwGzOoLUaaDAYZWqjaWR61M62eOq64E
8ZoZuqUXd/V2jH7Ufa7jj4q2JdbISLiFW6sa6c0+hY/+V1DlREeoO7aneg7+/tUByb4nlljUCBl9
3j4ZeOKGNXPSYaBgxZ5hAEJWUOpLH3H7rx6CE2B3n8gfkUvFS1H4XTGk9mqXkt98RXLYSW4f6Moh
RWz2l0/pKNVnvNZkjh4de39MfSAznGsEXBBt8keov2MN+lsckqba1MGNQg2HkEcVRu7tRJIvJt8j
j45lbAZA/rsN68axqf7pR0IsT16m/1R929WIKUW3zY34C+9Jn/tC/6/NZuZXMT5FYeM5+2Re4VSP
EuT6mohAw9pPpuFXOuxraSo2oWvjpbabyf2UFAkMAUvTpX0VbExmd0BkPFTcWpzfEEiUg2PISFGf
iw3up852J67hsQ6I/3AlZpEPy9SGZ/5vuW1RqzVXERrKZhPfAM+YXWpmBIuv63VThtQWVVJw4OoD
x+z4XqpbKiIOUdhCCzjPwB/uAK7ecyB+X7l1nCqz+qujzDzAUEFcLiogSwDbzVQY9RjgPxgrnEeQ
keishvk0qG+hV5YhRz364HQQycM78Zuf14OG+e6mpksx7Mkx0EyCkqjJGHYvc2O6l4gsDMtR5L/I
15/4UKtaYakmeop9/n0c7iObjlbmh53rw51KhYbo+F9vSGr4bRBXmqkTR37d60D/ruy+Zt3NBW7T
qWo9gQJgNpwhUyqV8rneFyQdO7dgQlI+ZT21qp9J0o8yWRY/euUnVJdST/9Q13eElMmFYx6KHjN6
apqq8OgaJnQpPKQeXpdymhRsDeYRGaYouRmJNby5FZdCguOv0iOPBDN0lWp5jjMpdWV3hhWzRvqs
sIvwnFaHsSnwzdSASwYbxLrLig1tfaHUvHjiPlC6cvDvH7J1WdYLcPfd3bo0RXwngIAsE+MvPWKJ
XeEVHF94Ee4TepgDQ1Av7mRAoTuVDd+bsF19Z/FJO8cemN5cleYl/vi/RVu/MBxFqECzAEnubVMD
SxUJ78eRrgByKG4r9oZfLkkeiv4Je3Vr7JP0bcrh7J/uCo3r81GF7q3g3sgRZki6uZ6GoFFizgoM
XjaG0ycoxLzo5iegdhEVzF7Q9Bf4A+mh7/9zyIhbx/u8ej2pK+RPFCjrz5Z1cjlpImmlu/VPen94
b2T6pzhZPsJowPWR3rVN4xumk9GIjQlnEKQT4jT3BEWAdA7YtLU6r6O8iEZKrtGNQN4PhBjVqOJQ
yZTIVCvNHwGsNFtma4tUB4XivWOURSzb1Qbn4AjRLzDIbp4zVYDCsLvQTB1J7nMDLY5vWojFZ6mJ
NCiPfaA/8nGWnPsiihjsK5K9TjZEIzIJ8nNgG6Yy6M/1C3jEKFhRCiLzL4z2O0kqobAdeVGb9ROw
UjY8mHW/uUeGBAbAqGm1sBLmoPOVUOSVzp+lZMsMh70HFbpFXIhLJsU4fuP7ZClC0zRXqSKT2bsS
YFbyR/LLJ0FJB07gFN+b5dly9mfaMx5dDwXrWAUuJ3mOnMjmzX+xU606Meji//c3p0Z/dcv/BdX/
Pud9Opg9bBsSs7V18Towe1FFGb2WLk0jTm9X3Um1C1uvBGlcaq4kavj8xjNpPla2D+OkZyXaP37R
jhDDthKw7GSwmkYbXMrWEAlS1M3SL8/04fUjSKZ1xr9l5nPrTeLpCnwbISolpTrqmIW3T4ezdS2c
6jbfcBU7PJgWc+TJZlFtfJFEYi/8lmOfKMUDo2iDkOhjySoOQ8cB/13ELxYShN/dot5NQs9Rv526
IMliOkDK3dnGTibL0YLTg7QA3JippYLoombrTSa8GfBOValRQ/L+QOWLZrQ1tQKhU4XMtMQ0dyqS
fat+CFV4b/p7X45s1V4DGolM6QrVzaqtBeevMWiFtY6DjGlMturS0XXNUI6AF58IWoBp9VHfCxli
qQQWaimi4eB3g2rsY4rQX2BP4Ec5mrIvQskmZ9vQ/lDACeVlcOhJTqtjeJAWsQ2QyIHDdYAR1ktq
tP6DRZMEDy4JbqtVnHZiOk6VnR4ZLIM1P68Vz59bZ3XH3Yq7Plkr521x0dFULXpe9iHF3usJW9xR
Aopm6lC7p2c9tnYEPzX4abKtR6FoCiny8FZuHJlNb03NM2cryYUUeHpNAjzvu/BZ2uQapa6GvDdQ
2kEZSKHUKxH2msNXaUWuA+hv6Kk0o9iX85sBZefaG7VLratpNBa+pDPCd6ssp9wKRfK+N3TVNUfZ
SE0x5VxP9y166/jBuITsA7/FMUwfJVvnaFYN4G6Ciqam122lDZAC/oDMLc1O30xBR7BUSrX1Dbx3
bxO5qWby8FsQ3F4S5oHhUsMRO1vmgvVq5OY2fmcT+YT1LrlqHBTJ+GA9itLYAtlvACCq094lwucB
LbR3b+icbgBx+kZ1KSY+1UU/rbmqqhRlqlajls5pFV8n3xcZP0ijbBT0C32+OnZlrgsRlwrT/kwI
4fuaCg+uhoEXtwC5hT7x6gW3kxlc9bf3f0PJyJ3KmFKebMqyLwBVOyBvRLAltIBTUp70gM4BJ9Pd
1Mn1+YxLuFtNFkoSi9br7RxzIaWrlYULCbjw4yi60mYg9L8+RHNWu1erhEydPUtuYzh8hd4sfK/d
09Z3Hn9o/fe/sojCnZtQkMIFxPvC12cl1QmN6omZ34rAydedqqZcB+H3bcOBH9HNUTmCr2uQyrlS
yLn/slSiz1OJ9kG9EGV04B4ae4+sqfHZZvAUd/qmUkWv6KgTzp8MN1p7kI6OAUjwP0JOBoL/FLbl
YhDd+jZ0XuyIbUTbWRnGbimjQcvUIPAl4FbG/IPT5irgfGhVHuzRikkhn4KGdIS0Nb5ZtM9KEgMD
LEGvZPxgvEaYGXGGaShIVjk2u3HpGT2Mv4NbXdBAhFqgy3jNSbWXFTE2uJK+cM7LiIlhFpMiqBxM
FKff+oqkp+JKO6a236rQ2W3xRC01jwMvEwr4a/1dazUvbkNwS1XSM3AbxSDiNscqZLupIeN66+ma
AOz3KtAofQ0YA/BqVDz/7uDqQk8/miEbAPWbH0sYuoXoPipSmsII3Ly9vHU/BiDB0vbJXJqGAVA6
ZItsP688kvz+ZRfwRzcHKp/qqYeP9JrsTC0Vj5HtzbNogX/A6snD5ZyjBmqH3S9VfKMYrNm9hwmX
lRhlAgjvxuZo/IJM7RKP1X9XSGHOcVXdZav2TWklTXIYY21IUwpk4icGgZy/5rUwGBrdLmIFNYhq
uTD7mkeSzhuEiiWCdONCZYXpk6XqvgngpV3d/gtIH1I83jHFJ7RaMO9/2unW7UPJmYnSFxkfV7us
CPntp1vDAPdoquqE3xfaHw4g3CZrpki+GmPjtyiQnDc3M+cV+mcNu9uTWame1pImjQI49f8Oa8Pu
VBVHhEDK4wYSD2aRbGwJq9BnoxlI8rQ63CDmksCfAZvyOdEk2EK2C5VeLOplsaPSb48UJko2U3M6
Zr5lXq8QYTCfgk2YGdz4WI0iTfV5RQdXVkDiGtsFr1C2O+YQpzYV/6T6XjAoDDSr6FF3rZM/CK20
jZef7AAch7Ab1cOtieyT38k6MpUrR65KVZX77IlpwFHZNX82a3++iCyVKwWe1A9JMCommdupfyO4
dLMjCftq/r/5vBnLYY/Q5hIR4O0ga3sCNGXCexBYQNL9HJCRxYLzzKeID64aL0Ze+8FB6b96C+hr
H0VypX/H1saAqPFRhbp0LSFWV0LwBDNye5EQfWI7YmHgK1K2y85QeMBUfMnPMM9VDGMKeWfvOsqP
fqr4EfWXjL2DmGrh+cDuObVVRGru9SPAL8F8OzkcrBXEJJX/+dYVAXdLxAI4u9c3X9jp7pBfYusx
+SMfXZlYnKdmv80vc3wHTqcQGLcech0GQFXK34vCi96ALUbJzI/l6aNoMXa6aXxQVaqkzj5pU5K9
jYIapBw1vTohza1z7KWS4OG8YNwpZmgpU5CqgHwpsBv+VgjjPqMrf17pL3IdH31i5bGHqVNtx37h
vt/Fdx1ZNf3K/BixLvO0Rgt6GpmlUwwftl/Sx1a0tXRapKd/gq5ucqz+SrLjLZGq+W4smyXmOjSS
U2MXBv9ute5nD6J2LvBml/LEJaKv2PUjKxO0XdBiMfiqcNyccScBnA/ZBS56UKHfloxBefEkMOWE
7toeRuEdNGtxv3sdVYs4Hm28UZGN0SKK02fsw0nXohF25mGFSwqyPAc3OZGHQkBB7oPKThewErle
mHBuSnHxTLq3oNFR7GbNl5FXAav4bfRjEyGASQ8VnECC7n/zqWEaDb4nA9MCAdUdYQr9+IqCmTaZ
ppf6nzVrg6UrHd2AMFrgt9+iIcPRE7uS3KrBFlkvdBzbivdhxGQj3S0hT/e14RNhyuc9ix6ynFVO
LMQ0Oh1Il6ERwBwChFk20oVFfcVxQ8vMmv76LOHuQxXLZ5l5dc/9PFLEGjjvJt+Vco8OfiDokM0g
X0FihX4se9Wj0c6BjtY3fvJ+MJguEUV5GgJpAoIRwm4iEJbffBa84a6EJsW0LauPQk2zqQR8UoJM
LIV8sL3Xs0sgYz8LLb7VrLyLMhF6AsfzP4l6jtV9QVpzuYtNEcm1b3735NJS/+HGyHP13BEYdbuD
sy+Rn+TzVaX7Lw1E7IumKMIOdRdeBG6fTrTir/UUo5omEiSJerrICZN0r3YPo0c8HvsttZ3CA1nN
qgL7coXUAiIq9Y+YRJArIkWb5Hs0Isct0jC/F/Wo2u1D5W4FDXD//ooSDfSClz1wKv3ZlJ2Fxdnt
UitD/eyj9T5T04I88y6gNzN5xJBArniMvAlorTpXB6j10ups68gieHrAoMAqFTd00BhSRhAuMt2a
ry5ssc2hnKHr++qCVUnq50ISpLl6IsvvTIL6eaCeC1yz0OCjiq/7yVdXSMLI2Mq0jDLN7UK1IpCr
6FsAR+cS00G7JIycLKniWnVpryMx7LRTKjIoRAGo3Pr2NZwajh6Tl4wPRVt8dF6JJsMZ5Y8HQElH
W3Ej4wsHDGB5XEJiQttJ18FkdIV0xs4sxdjc1fEp5OLA3KGhvjZe6y2Me+7uZpLaSBx0A8vxdoNh
9ilxG1+sYMMAPiN8TczFWiYbCjsZsBFkR5wnlaCgmHOO6d92nUibYXCs7IWy7beJhOYgU5Qfm5yi
2QMp6Kc9b0nSm1oRwmaQVKZ9TP1lQdLzKegcoIa2C73JywfyfH1bGEC7m0WUxA6/UHlnvbLfsTd+
nTJD0ceBgD2u12ae9dIy1VX10FUEPFnZ/9aySNp9+e0xeN2NiFqyzsnzaril0eHytp3PhqA/URBT
2+FRMtZg/diBnedzllrtHdIWn75R/z7j4tfAwlKPPwcYVlXDj47DfJ6p5lw8xbxTyZDunipwPbrT
q2jTgU7zS6lh8Ujf81T1q61GvXNGTf7Uc/0MFLvufoW4fHwcC8TUClvXSZ6j7p7uF8SmNVqQLdKz
Y4y42urxQEIxbfEhCeFdgz/BXM3E8ig+H1hUs9UiWzI/us0avig1XpG1/VAjLX+LBbP/hB/Ln8RA
2tMsNMaAwqy8zYj/quBFyF7UPnDVLJe1MLfX+n38RRZiRb41oJun9xpWI3TYqC+FFjPkYx5YVtQ7
sy6sPmdd6O8WGEUtohjjYejVRg2Vwp5Q47HbkHbG+o0M1WD4vJcLHVY/TrxOWwJ00lFS7IApmkpr
tXA7ulikrIQAujQ2LX27Z9sKRQLmz09dLFetoDknhCb/I4fXLMtlgxQ/N1+NhwdqBzkU4lSVVtZI
JtqHscxoeq1PDIVFHjUCSTao6b0hVkf9UN+BLLs7BOknS/BwhaDTwGZ3OQrS0mROKaZULtWPMaEM
8QSmnOORXkQjm0yy/zo0zEL/DV7bYwPO6Qhmu+XSTW3wus4jFuidDjuRQ/+sNZ+SPXKFYhlkdhNw
ZH17K4lZm/Kj6ujSufir+1gGsdDiPkmBs74oqF9qbqyS16xDZNJHWQ8v8fsjz8mPKmn0ZwD+naFz
iK8wZkq+YXgo/hcK+JTdyqaKXpe3SgPiItvHc9ugXWcu7OlUuweArobBHZhIJqDObnnZ03/SErjJ
tNB2UN/nfptl4umSFx5zpbtLVWEiFNlgncOu/P2GNmaqplUBudB/DnEw/H03O2/N5XXRH8wiFH3O
jxtDhX4ISf1+dhoSIS810aC6SpmEIdXsNeWr4FW/vFg8X2uQ8PhkVIJkk+oyIbYb+I71zZGv8jRM
qHO+h0SN2JX3AgSh8mkPyuH1Hl+EQEDW3d0d9KPwOEJyXrR44c0tG0+IMIlC6+H1NtNsJqcwylYo
I2rzEfHhZCrOFCODOHply/BZdcPyWyhomX1eovZRnjUUO76rddI+fvsvrBAoFds5u8CVSLBYt4vo
D4vYLSQhMnYafUM4Y044Qf8RqnV7OHS4kswpqLLnd0agmot76AM8/yIB/Qqh+TZVLPkPIZWA3ny1
phnO6AeWs7o+USJMMOPTOJ2Pp+QnsOtwBYYC2Ugb5T/zmy+uTiuf951sW1czwZqQ1qBnEVg/GvkX
8JvF8vj9fWg2TuiLz8KpwS3kz+V6bO3TfupjeC/RdXcQ3u6lEAJdLnJ2XchV3AlC++6HZYjKWAlF
naS3kc6LqGqvr6Iydhp+anLKprKR7gMtk8oE5kKYMScIKGZdILnitcJim3V3m5qaqjptG3ULzMxJ
D8dGueA86kMBjIeouPgJ8N5eBUPXHjKB+n65caH+pX2tKExnpWnILTAGAjtCfXoFGsd2R7RpwB7u
4Iw/N9Ev5pYiBJPfaCK+bJV4jnCTwqRcI+gW5pQ4WgZcgHXr/cMTWA8xDSbseTkr6A/yN8XXKP92
WvhdNFdNVzJq0hFoW8FC6AMOIOy59btwj+3FgkcZ5grH42F1ePzbKI5+lsB2EeDkiUW95F30TLWs
/Af3q5uwLbmRLMYGwFbv0EbZISidDky+G9lU293z+dHaAX/xX+kes1nDfgQ5wd854BV4RpJq80qW
s+8P3PtWrhvy3QcyLHCwLnlzGl47lUal+8L9TmNiK3nqEwb9joeY5CUvh+YOVAfaGNz+arhYuho5
+wPeqqRJl5h3gWCCbd8Tir3h3tNvPi/8ZxJjnZkYm9Cs2jzqfzvME+ypOy7zpdMmxOo1zkRDlHui
9USxUuH0TV+RUICXy9BJ/7vXJV7dYyLk3QoSpsK5wod8Yjm8CFKjAooZasORpzWL4TRw46xZcPaJ
8EhJjA424GXn1QnwQe5VyKl5MbdQepcjZNneegVviosBvwxsFWuPfirfQiTwKN9AwXQu71cHT/XI
qzaNU0Ke+4GDLpiBoUMuUAg+WOThf4uCVsFTXMak+T2TY6l6YTJT4xbjbt0CL+2TcNFEjBEltLwE
aAVLvA4DLHvV4m0kSfmRIqPFQa16sWX6R8gLKFD1Qc6CzgvjBfzoEkHLtS6lSGSFbocdXHs00Mi1
ldsG/NjjWEevfCFaL+UikqjCB8MvGwSaj2uA9t+rNPjsVZtb15Qoa54iKHhcQIoTijlLXT5mRSiz
H3Bk4mMJmYhP3ePLusSPgoEedkRuv8fZEDce8lFCXytXLFyUK4ulFbOhXxwn19yQkTwYxQ6Ka1yj
xy09vRKqlx4ptSo3HSEbVnliyZP9KcKwQyk+CO6bI72iuP4ULc+XxGjon/MbBYRluK3AfAsy1T4x
jEQEsOaEHGwZWgOw3W8bRTKGMzKUY2/xuKYJVSOuCJ5GXSvqz7YzWbiVmP8PiCLgjq9ByveX9iS4
3atJ1zIoDOh2/s2GSIHfzrXgG8jYVQ4P3wpy9vKMDrVVCYmZLWEgRF6oQaCb6kAJSscUc/RqS6r6
It7CH7QaSt6GPJeLgtBmahzgI8z+eYmmKtpCFSykCg623BZEP4vvYAYEaMGlFEvGqAVjDxWKk+u8
dhwo5yGjoqMRO+Z6I0ngVa0EnHyX6gawgh0Zdwc9WypBAc3cZRspVPeL1nc0Ihtr2b8mAHO+Lbgl
CMUGDKq08ShtX6zFTq7BZQz1i9E1Exm1W5z3ANi/W9V6p55pfyBlrssw/3ZlAMW0OqJOuNHJF2nd
iFisjXgF/PUIUVg7SQAj/aVe4vKf/G/09+re26qYybGpCmt2x9rPLO3XiFIpdeDoK8/WyQpY+/xp
waSpjI2N0MeXs9yTEgqivNLfQwm5fs9o3x4qq4EBFNiJ+tgjQE/+Ab3OlWCawFVHXVGth/PEEUpF
qFAm3oylq8TcuhmiG8mzGkNHigTcW8sWgIbx2nxovPXV8haiclDK/adK5RnA+zTnKHvpaxApLUak
D7/SM7Py26UOUv5lSiNZKIYVcyTjFskgarpl5yRpABVkPT6WvAoUMC3SF1ZA6v6lv501G08IIoYa
+jwMjt6lF86w7l+YO3ZAD8fQ+yopwsSYfpb6Fx5RmwVp6NXPjH2PSxQbrPMFmbQi9Sm4EWHPh4qc
ZBlNSiWbHLpxXkw5NQC+BSBwkTWC3aXoqPmQ7V23y0bzLze8Jmeb67mriQbDcDQgxIfU48YQs60s
ptykXy8UFXTGQk69Ibt3bprlPImDbEv6BOH2nw6QhhQv4saCdUrYKonWLFhSvX0s1wupUZAnh+OH
8Zu66tV0W2FqpkEjToCtlDtRetE3wNWSfGZ4rzSpnKYd6cTBqgVyuKon/jBuWZeb0LfNzxV5oI+k
o4+JTC9BWBjR5+k8fUrBcUau9dS3DjPZt3Gvjaps6QG3q9gCVClh+5CnH4+LF8N8PoJA5eacxcUD
kE5B/XPkPG5eYoG+uQpb/L05biw2kTVD7P0AN89GALaPwRvGmE7cf50mXEpMP+ijxUDTybEbslAi
kUfWI58sgeTLnAlu4xONp8WcvaJ+o7zvNRbVpaYw3m4YBrLL7rMxuEB69CPuZKfSvKLnON1y2iNA
3d7O0c7grpo06hCTQz4bSqBiqBbiPOVS0q8gV1qRByMo5PDLtwTOU+lRtbiKR9LOrXm/FkYooZum
p1xcFf8lLNs1SZImp3GoreFSE9+Pbd+r6yPySoUGns6tRLp1uKSWy1A7dNB/aFNInFR1+J97gMd9
XnYZ9OMCNiZtV7IwyS2vXkCk2BKkg8XoG7giP2HqkKrJMuAAnRARIAgAreh7hMmHXZ3Dj0CC7YH1
NoWO8nBTPGxkUDvKucTD4GyK9CoBeFyq+rnSrDvC9liis1NBt32RrfYhm7VhVghuDDPHwNmRy8W7
5QTNVnt29NFfPq4258ACHrgYJmaYe2Aw+8btIv2EoW1yDsUQ2YKwIaC342XTbtURJHftY0Kcdx4y
sUih4GGHgs+/86vhjSmd1+zIy1N8VvfOkAFNtk9mIPGvGzuSEre0yXe2cesiNow64ch5rrjEhIfO
k4DJ4Xe7+8wPr+nTWtoTRh9W9QvAR5e4Vcm9GmzUJWdYzgks8sDqgnj4dVidvngjosrj0LaBFJTR
v61q5ixxIUJWZ3piezeImT6sn8tw24+ltutVE6vCFncQLKzW2N3LrpfQqoQZTjWJFL44LreuxxQs
WqrQkKTL46ZC+8XRxLwXSXSq6KDbd5x1WIVpR4e1F/qVysJUNsrEcupFeCGkrs6rybYugNnFZnfZ
iKnezMiOGqAL41zE//cejMQKafwjhdjsQIHiliKKAHnDIcisOYgXCUG4FA84qDAaLbd8Xh5JQc/B
Qc8TEpo/vOA4fkuMXEuGZCGU29/+ZA3D9mGF9vUWcTWcmRSJkQuWojtLWE23ziwivxIIp0ZEukVc
MCJh6wH06CH4DA8lMegqNyQmIv/KeE2ClUUIBBn7pIwWY2lWzovSHwrgexyTwd9XR2Bd0mglJeNx
62TAM38519bGuySZylgvFS/dElY578GQrAw6te407S8JD0TYwzPgadfwSnGxLmZejSmZ2zOOc4sP
AvQQu4lRfKstmaNf1vtuoD42ryjpF0MR0qEUoOhADnCbmlzAdw3bBWWU1q02IVbyiiXFt5RnoU6u
Q9qu1Dkh2kQsf83i9orGUFhRZUD2RbZmLpn5ACd2C+C0UW8OM9ylgmnonjqmikC9Y+k6lV5VoUUP
nl+RYLIKWSBiLr5QOYvF+6DQ6rcNQLaXnXTGL20UUxUyOZ3+5sIi8/4sigLoEUFHxnUYqqecMSL7
0Xg0W12YatzGfk0uNimHODUT0/k9Lwi6LPUFq8VIYkobmMqS4uE/qqXnFoeoj/26I5GcnrR1R1G4
VbYuMfc2m45cNOmu+qIVFvPWPUOf2kZcSyyHiY33DAwcoX+thi2tmEjcYwn8QXBI95R/wbF9SMvM
g/7z4R/jznBR/arQFjCEX4VYAOUqNzpafj4xProSXrPv9rYTsPlAbusmb1JpjeKugFsnK2bu1rKp
Aqw6C8IksA4Fy9uxG8B4weojUy3rYnX+Gn22NNrKfv09G+ZPR+7sRi7nIRaZgnLDApLvZlTaDHB5
8MG7bg2TkKGwLs43pSqHC3n2U5zh6v7Tbsnx21f85Z0dvhAvFB0DpofR9nsTlDxivOjjQpH/XYTI
IFF51Cfye7wMnT9VkxeG0QvyXvH41ffLuZ8wu36Fo2umvVmokNjHwt6O+DIWZpTJEIMEtlwZRMwV
K+J2R82zVYwLXxCTLPsal9alY7jm22edd61uHQWWec+IGf7W8GfsKy/cv8rzfSuP0F97AWmPIjni
CAnQsrwXL1lEG35PqxDSUxYCYjtlZkW7MWiNpN4x4ZwTHRkz9uAjFCxYftHNwlA1+PYTEHRYfcFW
TfjJ9KFLwxTZFzC0EmNA4sMcK4zF0q8b3lEkfqwCJUEWzTPAVt92GAgQN2iWx+E8PJa9bRGaR3fm
eq6VZU53uCuHXE8ZxxSRQoh8FTvHo1BzMDBfF932NRZ9fkW+rziKen3E1AfMFV811yg6FGrrW6w3
IZM3FmUjgY3bbGiG7qH/MVV/TffU7LGqwsu6H/n9a1jXzCyNS4DkdHJS9j1KwOOglfE8NAmpmvcE
0+3pEgYkS2kG5Bag8eE3UtvT68InLT6T6C3Im6+HveKHiTwpp/oypgXA9HWSj8qyObBZzvIigYK4
ounRUkuCuqdnbXweRtNzB0aN9rhcBbxh16wVq2v85P1JP1/cZhsLlKLtLO395EGmggTldYvXf9GK
GxcS/WJTUUV5NvSZmvklO7GThbWXXrBHaU1CGzlNcHgdMpyXc7M4rSU2Vc8hq8uOdNpdTwRBSKjQ
lc8KnYmMPCzP6L284qoP3068zUs/COYaE4v0SpUYGvGfB1YIhQ0fGDCIjBmqO6F9AttK0JrYUuCF
v+kf/YSI5LZQyTYPa4KNJGLpxSmnz+wqqg418X1q3USN99JhLcSrr87QhE7wmX673EZmEOXnD6HT
EfglLmx3uArY3u938pra67ZsOMue4HPKGIPfrV/fmn5ls8XcvUY3QfE8w/y4GT0ZYh3x9glRZyF/
yq6VLoSaCMwu1aoheoFbuGUA2cdhKEFoU+X3Oy85oBJZEUxBlBJfF4JQP2YAk31XZgOmZXXNmZE0
cG7m6kMSTlamsPYkSyHj5NVlqN05+a5hMVRV1RE80WELw3HoXMiD+01AOLMbzw6pHdNiHLXUDyHI
Z66tVhg8dT5XaEYgkIIbhfl9SwrGN7nmz2k1mIuqlypRgPEGgfiCwKoj/0ypGXmao06Z2J+hbj17
QTqvGF1NhOdCzdlg+JwzI9dJZmZvlNIfPKNUNndOaL+0rWEdwxjbBHqbRE3WWj1YRSOk676bHbiO
Mc649fPy7lDLs2alzqOshLD1dKqzhYi8s9yLqEck2rKMnaH93zD71z2Gt5rDhNo1BrnqP9/L20d8
3Yhkz9DYj5aakyu2/tqeDoETRStdm1otKouT18glbvDdFN1yUhYNSdq8EicyWf/1oDT9zZ7wt3dU
DeH1inTLGlcwPGBnU6FYB80v2+2dVmvfxgcSgV+XPmNFMacLybkJ2ebapXcJeUNV29uqRR0KzJOF
Pri8JdN2Bv8jWmqm58RNbqF4VFoYp5PsLn6iTDef8F9HiKLlucdkWh+eH+F94dBTN3Ddxt3rbs2b
df8O0ALIgi60HLs2M8LQfylFXaxgRDOnYaf+OnXlleS0nIxawuuw3NcVFg3oS1wILudSLKQb77Us
cdAFlWqNSRWg42Zm6I+ISa0fo/MgQVbKpuFBaR8wjM4R6ngGhCNXdHP0Pg2NeyTww+rCPdCFI6+3
ynaibGBmHG+HP8r9Y0N2vEowCz5Io9JdokCebny4qJ9hrj8MsPmXVFzQh+ITBULAfmlDdmuZonKP
4Qc0JLLrmI/eNdbQK+oQQOMVN62aIQ4s1glfJTkmnnA/PMnKecSjejwrcEWRLvxPQEbaO5RqyyY3
mx7svm3BiW7cFhc5uw1uSg5oXJ2rFaVurBfw0nxGxKFMHb9WuY9pwoBi8KZe9kBsDd1jZHrfhSx1
AHOie+Uq47kWnETjB9Eo44PiVeUc8T2RU4M4g1Ch+kEBZ0tDnYTiQ2ocFy7EP3AXn0OjAr/BtCqz
+50RprrPk2+eD0RijQNo0Qnbmf+xgFpmqGVgC/1HHIwELjlaJ0C3PkqB6DB8A9bBpfQPn9+eBDHd
FOyCx3/pkhHjh+OTffAlGrAY+PY6g8YY2r69MRn3qjh8xEFJ33qnHyKEUa6ics/zx04RcKKetdmQ
1INF+HOMCcY2gBwbCllF5bAds/wl6t3wH4KmIasKd7ipBSgQ6HSbHJdXPBpZk0S11ov2aiOnbqpm
yxoT3SJSfFZ8w8B3TOt/+F6C9jJqn6HTEQAGiJfM8ceKn/BhJPin+pb68R4UKHUOz+8DIjgMA/8d
oeIz2r0MgvWycNG1yLW2hUQ/qL7arRmf0HrRG1U92vafzIHUR6tEBW9ibKWFPmY6agGWec6INGBs
QWKtTO/63KdSAGR7jPn43z0zEr7/3Z34E5P43vFP27GlAzSlETAOGh+9qsYP6JUn1vzt36tYHSBD
md/pw8pD4X0IWmezptzsrmp7bcabgguVMugUWpppiX2l09w58KyM33peLLvKjbcDTPew80+8fwss
r0KcO4Nos7C+RrePtir7sAPVaV2790ehVcGnh530OO4g1qkE9cr9igEkJJvYc7hnq7Mrd4kKX7ou
7RbnurmL5/Rb5gzCYUJYj6/2+XY1GfzbZGxLTvYrIRujZW033p8SapsHD6sqVUQuK6Y8V/0DYNtK
0MeTGRNSeLN9+8wIvLIIJFviGH8Pj8SAnLFGxbMby1Uht5X4XS3QcnPvaFe9Qbd0bz3WgB2BEQke
ywWMH2DHnQYJOiPm8/KCaM+bjsNr/qpSTdpXoJD40P+DCodKRGVLuXCpnNqW/n9f71BaFRvanOYM
37vaiuJfxkKIxNZWduvouJiz8Er+XVa1VziCrxqTIm1Ah7u+89ty/KzvuuF8o9oVQ4fIkIZ+XR8V
PRGA+R4SiQrBflqc22a9Yyn0/ROXh32Ileu8hqVn9dINTeuNGhCawUnXiedhtjMEJhZ1FDOc+dqK
RX9bPZLvL/mxuCNGCSIJBGLNFFHKXOiVSG1ZtwoUXKhvFNJouFads6KIV+FZPuiD5TCGtSamVSXb
b5JIDq/I95hecWOL7Lc64XHVIFOXF+tWxMDH44vfq424+ksVRUIHYy9OmWKgh/ksldVrwl5L8oxm
1zn2s+5fjnmCKAAdiWET+RjSLcu49CCakdTvYPi8g2CHDhCze43/rq7X27YxCZwP+vQkB2CzQ575
D0SPoyXCTtt9YSvCVXAmZJfcG+l5t6sU1OL/BKRVnE8jQePNQbuOngRfrEHr0KUjos6o1HhLHJoZ
MP7Ww56iKb+LXhjGGC6GdZ5jfkKcQFC4ymI4J/+txYg8HoRpomHLBwcxrIUO9s3GnBwYq2HW3NQR
9AYPmi2aHd9otKCneipwJB3ysL+J2dwgGlDwR+NfGRyE+Fo8Tt+7Hlq/tNV/xPug4Mo5hQyncekP
OIUMWyXUNYnU6PL8kwI//oChPaE4jXV8iaTnZWGBTCxwyFINFPypaq7LQPlnpNztV3y+ckrXZ2am
oCxfcKwm6hWZVoa/DJt6joT5fJGmVRz7S8A2jooo9duKd1f/TaThRUQo7r+ME9T7IhXWKqJdV0xy
y0Ia3XHH4GjeE2thSxYrIkD2L73Dv2lhJf3kaiGMeBia3IMMppwFiu4ucje/j8xH53Ke0IICf7dZ
NUxPOqrs7jaghb15kOU0wMHRH+mdWDzArgXWgwirYNz6N1y1B8OofUqxCdGGB9uWjK3+n96RaAhh
3EpojiBJ8jRhfuX2rIZHW9lbkbOQxGqX4Jdcf0K6SQyD0DGDEYXdNJk09f9PdcDMFh+R1GcJlNq7
6WAs/OYc8Avptk4p8+u0Augqr3bZL0Kqq20IMcX+RD2NiUQedLVDgSPVxA0dgLs2veAjkm+FxBHC
FfaLw6SP6XBnnr7thuo/ZQwgwS/17meS/BBI1ZkJURZ4TzyxHUYknwNO33xDAwlgZCuCWguilAOF
ntnlkzvBxzpO+IDr50Nr4fSQTt04EFMDPt+dvxAB8q4vQVtA7TIKcv39HrM5lOXvoA5WQi9aCzZZ
1UXv3EnTZuS3qcPuG/TpnQJkM+PIzoHlT8ze7Wc+4pjIe1mGCxdGrb4pFzdB5J9eask8px5L3A+v
59RJhJRWS0VjOz06sLZZgg2biKDeV4y3tfMnwq92vaHWc2Ltf4VAdWKAi6rU2Zf1AOjOFERKyUCS
1xvfqFgSJEN2S3BNtWFDtsO355kSTJQWJuhIw7r1A+RQ/7U/hogJV1SbppK6j841OIB7vJMOYT5Z
GJkIwTORn2Cr47htVzPFfdtKzWNHLSmdrlZnwbu8T+wcn/4umqKkx0B07NG6eOLx2P6rnUbLMz5S
G2rruWxgEYexLsyE28rHamdF4txInhNWBeFgkivlyjcS3N6BHc5m94fmtDdG1ACXDh2na82Ffe75
bH1JEochQtN7qeCGlwjMPqZM6baUu3vFiaq6JtLezNDzk6keyTPr0b7JMZ9HNHocfhdnYFaZrLsr
DVLsMZlXGEKNXW6umHO7mVcrlmlkN7jYDbhrrRMOmyphIGGWzyfdAakvR956B6j0PM3fGN3nuf87
l1U1UwiJtIFjrjXk5wlQVz/gAcAmO6DCecZ/szlbtIa8t3hK+O2EhrjxS6Zcc22g1rpzrJMC9gm3
Akcv960vgi1anSklxlrwG6/nYM/LVMrDe8tc5H2EHmV01XAWWcm5sY8L5zLvvRfKXaZpqSC6NTi+
6ss5XWa9fflkeWKT7DkVkjIs91NeJG34n40CcVZL+2xbdt2Ea9dpC9nvVENgp+vdr8jjDxk4q6QQ
tJuXFtISRW6Ll+WsblByxP97IvOFPbiHlmmKmDPtEwIimuLqEEjg1VjWy78euoO8FDcWCiakuHwr
1UOKvohNFT5SHUlfUlTWkgre4+dupbMQGgJyqTXy6wcW8DmWfBFSCTNPeXKY9EM/EOwPPx3yW21l
V6X8zUdtD0rB49K7hgswRFX3rY2pj8YGtvumfjstsZeGCYbW6Ng967bJzGLy5pvnbXNvvfnJEcLR
/5GZfFTa7GvHMK0wssTI2yTr928LelrQ+C4nnEy1psAQoEtpZthWMImtA4gjTpf2YhNqQz/5OQN7
snyydXp2pqZ1uM9uqylW+UZcEMt8KkDi4QKPuj8U+/3wZyV4t96bBLO/JOXPvu7o6N//kRyCfTu6
BCfAoz6tk4RIWqvkBGVKXWcGqpIKxx6RbIkQlGt3Vh+HmSR7vZyYDR7Np9uDEeg/2S2U7lZhVDV1
o1rv/MHPtH3WMDkzr1ZNOc/m8fyT6VCF01nBL3jLXy0+OPt9oZRm9yDbNkoc496evTArNdGHoL7h
8UzUSpLbRgv25sHDPFY1x/DE8yAx0N6e1ddHiK3DUsh3cEdYhPgKPBg3a22sfAN0kjadDnSrcTvQ
5L+vZjW+5xScstCFPj0Z78W2RaausSizcU91f89vSVm6FAcHM7qRpoiAMLnmJysqzZ2KAL6wq1Xb
6FpTrOkzIB4usNX2opS29tNThdb3Dgr2dhW53IS/rWTYaxqEapSdLtrkK2bl44lrbpsnRaIEgIqD
nHj9VHSdsXwlfP3rpKJbvHH53JU8vud49P928cujcAT6XC3h2BQm/ePZUx/bRK3lQiNXo5Id+a9u
e1Tkmh4q07Z9paKsZ72TPiOmmzts+ElUq2+qgKA/braUGpRGOVXN5r1NiQtO0nJoJQuv8ZKdcKww
W9g6aVnzpEXXduj5wOFYWVKSovHvsfGDV5MWTqmfb6CQqBppYn8HnFPS2d7+IfUTP5uRUGlV0Wyu
L7U+SjrZ4zE1opMKdPNka3PhpkEGMN4AC78PQyyXcCK94kXs012tKrSaGNIvANfY4+ftuAk/Wvrm
NM7sztdm4vqj/MYcPujnwy7MLJjEU8k0zkgVySoTXmDg/hW+P5eiIukGsBaP0uNuKX0LVPsCfhxv
Ib746QEQKH8oWtgmo1M/NdanPfqWsgPEpGXCY9B9RBELiFAVQFDgO9Gey75xbYgv847HsYB6Ho5Z
NDMmycFdtsMcby0rY9q7MK8LldlcrXEAIc1JNjkyRoKpKFkdoDKg34aDlIKgax3BMcHEFew3pNEJ
twyCWuyIJy5nUDHyWFGoAvJfVXUFqy+a2FOkH7oMBMC1ExxP+YoTK7IaliDZKm9hfp0C+zIpLNK3
qxejGMY6Q7Ft0YqzKqqqjBd6IfaJI0pKgceRJiqXjW0MU5fBIP/2kIZ0zda6DFo6c4bTFYIcoiGm
NFlHh8KpnlxLnzHcjo4ZLRnQBeKJJcxdHvCeYhG+4AreWpTwc+JlUkf3SV/L179g/GjhfLJ+/skx
lXR+hnFMcDvF6u0K1m4aWaMk/KiGGqmd+dfK15IktJC+JlnRU9TE2lUoDcHnxqzZRuBFZmZtNS8Y
FOzW5/ixNs7SPNxYAssOKyEwgm0InZ9ytzq28MgGSzxcqFcg3ArqtZilupg7Dh8F3SPiq49au2RH
chKaOX0GGJSIs4hr3pym0gEm4Ybk5dyN5EZuDneeWMSnJ4ry+7YnWDpKX/N3e7+SXwcnr7lpQOwK
Sjc7YSkeQ40PXBrBSSM0rvezYidSe/vU4SxZT9MNvJOv8iPT50/K+fzsnCaAXlkA3fIRlewk7Et6
6fPR3X5SQWGJlkaMLQFJ8LywNsozjXy0dfr6egZXiYhcaH1v3C50f4TqNJq4b0zvYEoE2Fl30Cy9
nuKbkj7yOd2VqUNg/1fpOc5tt3K4bMSvdaArMpQufOsVQ1Du4xGGkUsMmtMKVLNjHTJxg3ak3l81
Nc/qXcPplDmvtBc3U7nt4U3j8So3rArjedUaOfzX5QPJKkHGbFBzWSEz4NL+JbaY1WL2x0t3c7L5
T/cCebeM7o29Bn+W9ckjFq0I7M2aq3PYx2TzJ9RNLV1leJtiwI6DVTvnZlhi2UDJyAd3JYA72uHQ
J7+tBDXNt9FSdNrByPo46ysLz6abNdR5YAcbQFCMwTpgUwuPdlv2u2YQ30mN97pvQWt0OPgQHgbI
eo+EA3d5PLAiJllVWNT3BzkFXjejw1m/awjlzeQoD6w0avYkjKwXrQxWd7X/hL7SzFgaWKsUrmxT
UM4CHr1n/jglRy41Pc4OVOibNW9Occ3aE5oSNtlud59bPKQmDJBbKPHIW+eGOdFNV8AsW1BScQcM
K1eOjT/5yfCVhUwCTZXjMRkyB6HM6RtC5dNiSbOonhWmSQv5t7QBg6hVtcBe5Uw/5dnhCpIXF1EO
8Kcin/cOePOlgDEYRlamw3Lcnox02r9hJlWWiackWl9I45F4U6hwEoj9pQBp+UfSm1CTpgHTqbY6
qXUx7SpfKOpG5hi66LLIdT00Eu03hCwS8sqauu2/flk4VODXYZ67ghSgQlWsN5yZhlDWVUL+SezY
vT+EGpJt07TQBl0catC5QUcg5Yh/Kpo3rCkpe3+5q047WCIO4z5w5+7SKDqrTpCHscsz1BsqVlzk
EVgogLdu9CdxrFI8C+mLhlSS1nHnzYlDFoVIlu/XUJMDmbhtrz7uZBIqH7xZTCXQUVo32lkak0qR
pLXLJUQC5ygkgdbDEOt/j5HxsorPn3F0pEAr05HzEELMQ1hUZ5xPKME/0UJIICr1MR8VqO3brsxR
FlGQ1tSdd8KG3jM4jeoYzcwNJkrEr32LHUXcJ+jm1opbdRMJLx2cM9eam65PJG5RzLH8vAgL/X6p
Mlr2tlIGisr1pDzq+KjpGoDG/WkoZt6TuUxpLmi+G+DHN48hSvNZJLle57WmKtB8wIIyFbDFMob/
0sbmuEcV8w7K4zEJ0vSDmRn0kx8Bk+RhXTsAjz8/IbVdQG0mLflrsWwGXECW16UK+9p8CCw6JCVE
YgU98g2MbXPk9qwfPvAHnGjHutzZgajMxf6proAL1MzKrw80vVPyf4hVcib5A1X9ZvXPvB7NZTDI
WouS6ZZulSX0j+1ehCN93HSznQQsSUwRYwIySOyfgfKSom3vFq+j0VTO27uVL8zgWdGz7bIjh9pm
WtVdEYVL3GXKxku2cg7o+DUP+TpJ8UZppQ32jnS26LsfqhYZn9tA4PKzxB9YaBKehdjOZdOgDoAk
105SRg9yo623/e+FKiqnMHA8C+UHxLqX/uvu+fOoVb8nUp3xQ8ymA3fNNXNdd1eFx/V1n3+HtOFp
upx9h34MvwsSET8UkF20RPd/8EZqU9Y28DpBOlc50QbS/dHXIwZgKDP8bQMyEQ3RdWxXo+B9Ed5V
iNfAm32xUaN/1BcZ0vX49FLXZc8fCMWYLDADjGiYvgz7vGWTOryZY3BctWptxQd4HY3kCzoRZO4O
eCOcNGYT11BcI2h0OybIJg13E2nwPJroNzz/V+uek8l92+24OPLF08ss0tkEjTEF7+itZrtj6Jju
vTvatvTXoHnifpgpQ57liv9fpAEX/8niIxDpa8IkIKQNiQZ/YwSlo8xdmdsMo69M7z+DLzPyF0mH
RV9xzXeIFAGUWtm+FNJviniYAYc1As+ejyrfJeOhnsp6aPB/fI/TJRww5JE5HgaBEEy/VtnubuiP
w82jdJnrxPJ3xvgy1XGoMtSbMopwMO9f1oww7/K3oEFx2NyZdVtqL6aDJ8o81xFzH9O5ECsoZ/M3
hO1v3FnoxkiiWiYdUx4R9+G2isk07KFk1YPblO1bJ7ltfYvYNZHNB5vfB0L9KcERFZznaU7pmLSw
mk4WSUc0+PxU3bNC79JLl6V0VYtoABIwcxLTfMVjuIJ9EmYr9H+HcrLDmutEOyT0o6sWQeNmg1cs
SncQls1AU6HwpZzgAAFagxZJ407xNYhwpc/unYt2gfQRGxrCce3NRlXCS2hD1NUBzmZJO+GSyNPE
gONLackMme2s07Ff2JpqLhuXYFG7TnbVEXrUf6ttylGSku3yZLTT9G6m24qTzXM5tzd/bY+6usof
7ScDde+faTap7abWPYqDjE5MpeFSRIYYp/NOauNv7hveq7htjOgI1EizI1w0k9O/S1yBDblaweM9
bs78hbgbHZNQhArI57THepFGIDvrOoNJjSDum3e2QRYRI+nUm4p/USJ9Nuk5swD2s44n7Sn946Bj
lroqY4MUjDgEA+oXsa9NBn2h9MMtQ1LOZvWRNInmX/N4BZB1ZfRCronfOlFN2mM0s3WhCYlmtyxi
FoQVFPmKuElZ59OrfnpRaNwf6T6KMtWRUIbUoKwZFht6oR7CFMGe6APqP5BR691Fw14aVqWFf8GZ
qyIgeb/AY5POWV5Y+ajSbsaD6Zh/BkGTLerUEsPA4CQm9xir5HLJwP8Mw6fXtZdu8FStY8HF0Cjt
3g8qrq0hhnpRC9F0sxFAFfjPBnqs6Lok9KrLTnV2IJvNE0Je3vkYMSKGTe5zBAx+OVDms+XxtNsX
EhFInxFzJkg6XoQivH7nNgnNLW4QhqbN0x5M1sfTyb1EsuS+nt4OTG0Yv2CsBDilRx71Y+dHdawn
14gJIIWPjTmW/jSgRoMXdWTQWXMmOxPCclD6x/LrXk1+0wuOLAFqaMjAQWIA9ZEvQQCyJuNWsUVz
zGJlT4w2tp4uZhEhNeohOkt2MI87IwfsO5sr6pbUMHuYlC1CQBGr5YvbW2kio15jrQm4GosLdwYE
v6x0SU75KSmnAw2beuabZ5PwLGDRlBcLVWcxXGp82mtT/J47Wd5/NesAFT6tKJ9gPePIZiWk+6t1
DTHBaSRJQ2f2t1tBlFcFOyHIhnR08axv6fzgTtJSq6hzEY2g6OFKHLAuhsWXzczQz/ju3o8nxUeK
YTdTB5eFqAxb+obuEA28bYc05cyYvnnzYGVXmVx24QuZEZ2siiE22P96ydKLdf91r4pALZc62Lut
TcLpSAnfW6cx4UtbK+3fFmrNUJdnli01zR4ZFA5g2x/K9FdRxc8v7RpYVZJxpSgVdolbaoc+NQsE
twXQyzwtlKQwEXzQEOyxmD6ps4EMVK8CnxxU8qtlIY4poEjfLzeSpAC8VVPwNCteoeTij5HDqNn4
i6y3BzOCsEMUscdIYyPkde7XBhbR513+TjDAlodUcT9IF+hjlSulQ64vtXJmRi/wuI2vllquZFFM
cBguXYLRefF0kpfHV0sHU7Q3grN/bcazRP/DJI9QXATAs30+97F0/ZbH+Hu22hK6G2fMg4XGdiN4
sdr7KE1RYKwRZUQUfpjH+NqCMdVxUJIvJYm+trtyMaROvf9mAGEYX40BN/aIV6ILmes0MJWmzW86
kpgj+ejswKXjpkcphu6Q9UnIuTIN05Ixp5E3OjebHW2hvOUhFc7ed6skFvyHcHpswpW5heQobzeM
LHBiZIJopPKTfBT3YtpNifKOoQ95JMrmVLCX4pydddx2tQxjsIGvhnpeUluaaJFtoO1FsZf2Ioz6
RdjuIr4I1Ipr5v1cvyy0Wv9l8kSkPH23Sf6uLKfNH3zsOvzPSsc1memx8xW3Yb0I6cC0+tyaq/2O
1ai2hoQtZJBDrxJyNx+cY3g2KmyEK5pI2G0TRqTjgF/cT7Qa13pXHZXNYjCW/KlJWSVKljGIHeFi
GemtKfSskMG5x3PN3WI0J3AD6d4umpr/nbHGOxRIMnFuARHKsRopnyrNjw64o2oFSXEf9D9F1Pus
M8JAsEHeIIUywialj+3vaYPrzfZNAOMJ8skBVZOxZRj8ppAcmxpAEj0fDIiMjkrg7Q+TjAYwR9Gh
kqNdDAjWvbHpy7OiTR5Gz6C0OXFpPNFc9w2Fpc4nhPjwXlDVuDs7b3/uLa35plEH8Rx5E4pihu70
lFoX5t667bjVZdmLsWdr5SC7zvSWpg0g6yeBTZmqnkQGDCkBe7DOeQpgqo+uS7cMV2oIe1YhcRCY
Cu6cw+YgTXVCstkOenTp/M/rmLa5r3KVf+ql1l5iIIBF8elNMWq5MEjGQ0K01NSxPY9mU9VMwDe7
HkUilTu2VHUrlLd8VOOJqFw4P+RbrME6s67yM0ynLJ5dE/FQ2Kr1tzUgDBgG48noHP6fNR18a48h
im4W1tVMx3SMGAybRpuirqsdhQExbt4sJVRaYWIbLzDJH97v+3AeNWHImLYceP+sgWGEFefeVJa7
uvcrip4Gl5IcfNmCjFSWlqUGGPn3HSTnCo/2j9hKN0VWRZ8+xPZHAbRkmFfXjrRhifgdsuQN5mMm
x9kEEuRlxRle7zCi5h4A9RRtivHkje6VcOhFSAk5tlVV91AnnC4FpciqvYhLvwzzhIvpVbWUAF93
/InurnOXXdlLUHeTaW+Pz11f4ZaLgDvrZCPHAHQ5C8u+3l4Qw/fxKqZjrpF0NF1qJpVsLHC3/HVN
ELtbwH57urDFEfgr6NkKePQsliEVedK+RgB1uKM2S3h6De8SO/CuH/Pj+t3/VNiXQcDrX+UOmUZK
oqkL/NaRxhwj1LEZzs7efe2NMyzRrbi9AYZ5Ccmh28jZqxmT/P4AUgRg82co9PS/l86zIuGXLHvT
16Eqt2dQ/YeirzNiTrR/3xzFwE8sYj9VUdStilWZojuUi0vbsrugUStLhEPJw5sN4YQSKXqnRoMz
TEibVcNuz8cn0qbL8SAPS2/bodiMIxV4s5fHVfezQi6lIBmaqyzD9yGjDy9MRw9osijd163p5Ow5
FiM2bPCPyMuf/Rx2RQ8WVnbNWj3I9fTWkjEqHyjZf8BnvjpglMqVPLCgwPOJ9KqH4sV6EdyvyTJ4
+kapsGTXjvg5Xv4BLTpJkWfg2mT+uwzRa+oRHUpRI9L38MtZQUzc4ndNOUNwD3VppOaIp+dZk4Kt
hVAWc11qAINHnVUgBD+uDH4g7CLV2uQaIyYxM1xULg1YWhuT8jOIy+DJxUpktizEzWrigN5l6j5a
f4kdOVjEgo37G013J2TBBBXtpLkyt3A0HSd3kyDM+niXaTxKskDva4WL2LtE4707Fhqi+sjcScnQ
g0aW5z+FQ+BS1/prVlfzU+0i3+l/S7ntG8xyQAjIoFIig3gRtMRst/8YPfE7prZbZDgg4QengVo9
Ic/lBTr+qmSsaoevGOBF6HbHGdEfZOKl4/YcRnmxqybV2NaQQervg+D6DVydQh64cNG9klrvGTeW
mvNCTH3S7GlS59V85TIhvCsfS9acTn0YskvhLke0CHdWVRRdGxsXV7og0q4UVN9Lg3/2OIs45MBj
XQYqDlwKaK56gmqbKkHTcRelo357/fxilnzda1wTDyiwNH1CwAs++JvfK/jnfvfA6GVZD6bUGkIz
wO4XIGMP0/m2dVQpaZzt0rhaJctfIUdw8HT2+e3wRvzTzryLiVjM95b71ao9zRpMv2Il8SuAsWg8
77elUwJN4uD7vu3hn2FtffvnflXCRFlBbgfFKsu5IjK8rggCDjDc9CZ1VAlgM0PZw4+Beh7KkB6d
XKovwZ5YAA51B8tWGI0fdvNwnEcu23PHwlv6mmOD1dYuU0R6hzCjmEtpQXb2fAgcPdsgLHSAU+tU
MNALSUO7XZxRJpK+Cp7Xw1Y9ayjmF272oVA7+q1ShjJx4jWp6TCmRCJBsKyA3E6n7PD9kK60XDB6
mM09Wou43grIX96R2GqRh0pneAGmEqu5wgCYChAeV6ufCIFRWl9OGqRang7xK1lU2TlKxdoOCvH2
e+q6YoJH72tyc5g5YZiL/G24ExqwkvR3U1J5IernHuWr/LCfmXl8yyE3yeneGDgMlIgfy0c6b1ZH
t9NCT6CA6AwJujaUfyS2glM0yZTz7flwm6RoRa1OohiGn0r6tVfRSb6k0W94rC/sw07JsPqSHmOQ
Q5GmQh8nooswsXKgLtiLfOyRUMuzhj/kpOJae/efe78mU5xstBv9Bb0TYBJRjI3n0lDSiCn1DHCv
HW4IxQ7SLWLKUXiajn734bgla6qu95+rjzu0WBBOjaTvTy45gO38BvP5Yfq3mCj5NiCfOLbvp/HN
s/SllQawO/M8X1JYrtQP0zshrjn/RDofvN7oF/DLvWd/vRfL247D2sBfz8TOyuNnaZfMMCangHIQ
kzaXy1Tx19SxCfFMybQvwCVQtsQFY1GOiNt8JExMjfuImOe/t0lYKNKCALDrtxV571UL4+BynC3m
hUeEmnYnq6CwTW3Avsq9mURClqVUIYHtO+7CAxZU0WNt3i4j4P6aDIgpn4PvMmc7fLnmXvjOF1aX
1KYJ1aC/B17UpogkdaNwO/GfzZfleGUiygLuWQEv5SLedlULM+b166exuTrNztFk4HodwPO5CuF/
ANMaIc5+fBe2hAwRfMVMSd7a0pIbozvA7JgHPF6XRc2G3Mtbq4zFXz0fP6uh87WnjDokBxzY18PW
+iSMzxvcylGnvSwJErLUHEfQ0KcxLPk1CTdG+rdwgdqD8pNoR/c1LNV9wsIb5tMG5z2jToZzCJHH
sQ9ksTa76ZpBKbPCA4btX27aGKp9UunxGmUps8Mh2Og0GdVwIBTSNEQ+BWzMPVVYTG0/PJACqNS3
BwIZ3SpIPp77MtkKtbgXDGHOku5E5qNAi0o2P3gh93TS3xCAMkf81F5kiernzVJJ3I0ZKNBspTP4
m4RUmMBrHBERIUBLC1B+VrwXt9spRiAvj3gJafOv3cmv7MSmaPaWLDiY1fqnbcBuIMQtI/XemivY
vFzNoSbuPrS7QTTq6z75QGbJD2ZF7vrZa1t3t/xACOskE27rip71IeHAKh2fXkcR7ZCOVnOMhwzA
zDdxvpv8HLdzdt3lynNmFwBxNlCrze6NJph6WMaankvZJx+ZdFaZ6oevq5OZh06e+fczGFIRZFTb
GG6L6IPHELi1rwX6k5BtxPK9x/7buvCyPf6AFlz0u0BxorPXwjNSj9+aFiS6zvEoTAW+1AKva/m/
ijRs3/x8NWcqQmlURp+FZKoYwzudZksXembm5cVx+KO+ceRJYg4aqC9HGEJSa2HjfCnckLzeQhSA
8WxdykrqFXal42R3avWyp4nsh2QSwud+q3aeVLE9XJwY1ctuY/Qlmv2+wlH3Gaw1a44tKS/lqdIC
FmdWfNkdzzzuODYzbnBgkuC5qOP676waeO0wY+rPKdyzNuylT9vDGAYwdTK4CbDwLQ5xFtAiRZn4
Rvq7wKQkHvyiYt2dZ6Mc6FxozMObLnYmIzux6H44y33BTK/Ybzpti7zVibvhRudAWS+uCK6CACGl
rp7WTcZ4hEieGBqLAMrp/DXdCLTfVPFFcuSJcafw3sOiwojoM707VpRDY0biWzYE2/i0ypavEf3H
zOKR3POFt2iUI6bkQGo/FQAtgSUwY91l+0G1F+BAHqUL3X9MTNBx382xMeEE8eUAUuhT/Og6+Dvj
VnrJDUnzrOHpkUbIk6X5ndhOZW5/iNjskL9R4cUuzDNEnxRgsuEFQkCx+MrXgpQHqtAKUeuI56h0
R/N/EFxiU33vTgR7IWwCHqFUycmXEZivbQPT3okKkLBk0KI7buhhVkiUUHrPn12dJgmGegmed+Mi
Kj1X8u6ofX4ummZtv852jBuD4QKH4yDuUxdIZH5Jh/gwUIkL/SxVLwXKApVsEgcI7anzcOhdT1ZU
KqYcd0al9jnB/2OxERcIaZWuxmAiyPjcMxqCedq0/oSa8V4tddBdy83aHH//PolmHmyUnDhgRJFz
f2pM7ZKtLPxBgNH2rIxdMJj06Qvg59odegRcXMSrvF9vbvEGaXLzH7sx7V/30hsGMUYPyD2LqaVB
i1Py4tyz7o50K0cALnwBazJoDcCCYZ9TuuiD8LfDGvOddoPZ1nbmySODUH308jL4Ly+E0bwnIAeb
BnoeJowS7PtT4t+bKTAoPuoAs7q+LPrGEElQ2qzhro7MbPO2OXtwM7DCgfXk4lw7dQhHT8y61fxg
dZtIf/xHnapleKYpRGmf7Hslr8+ndF6abcb9sPifzYM+zIFPYxkvYhvCAa6ceHnnQZrSej018UrK
OOsesTKbmQtjUCnTb/rxxWrIJeiFMJWlmZeRxWnDmpU5INyhXGLaug7T+wHmgBiZek+Os8VkosyR
FRQNyBodmsnWQlKHAI5aoNO01ynVjEFEFCq9A6wJ8LIoW2IicE9FcUHCwnjsDy7ES7DIeh7flnMC
mXwZIfwDWo+A1/sLltbjRO0e3qXUdIc6TBjrs++F/UqBwN/WyivMCkSxSY2FczrCoLtrGI13j3Qb
S07AKZcKMp1DMkp5DYMeogazKpucJNpTC69TwdAcHkOBbHfhAxTP8blvn4CeStOGkzIeI24pUUBJ
wWCSkzqlcchW56i/esk1AI1uCpubgTEqzgNj4Ul+OTlBmCFMTHtvWoWknAKvZ3UGFGIxwXVw7FU/
8K1HDvOWNkxsg0boFqNmfTm3nqB8fqi/0JuybuBy1W2Sfua70Y/ElQBq/WlnB+uICLzqe48kulew
jkbHPKQb8TDfDGrU4vQVoCuajntVUPJhVRKMbFGF00etoM6TCjaPdjxqy1gDTJFpWaM+dYhy8B2o
9zPQ88P3RODCsUs4/Udk8fA2q+g180gsW47tW+fMWkohyVVQ3uQsyct+Ys1cK3yGraYwNrq9RJMc
aMJkbTOTm79fwvk3KhZQ2J8bBXnBzOoeef2IqmLeVCd7r5/atRBMgd06s0RphWUOwBOI2laOo2Se
CKrtSkPX8WwbhwA4jNvBSXxWoNepe1MFN+6vHXhWHuAZcLmHnCakOOPPhZbwsSx7dR4tdPlbDoPN
gTalxwk/KgTE4K8Nol80C0Yxc2NwnlYwtZeEke+jdMHps66lXItX7T5VWR+nNQCxoSpVF9SEbk3W
/frYORuwQeZK/cf75cRtW9LLl8TTcpcYBHrTAMcXTeaiyElv8/5A1ATDv8L56JsItc6mjPJpOgPq
FkpBVrpUmCo/5VfOhvHQAxJhmNlMsV9A7BFMduXBDdotUjor1IkkEq8eQzmdnDoBT5RlY83XCGAG
e9GQYM4TGJ1c72gccsnA01jBSvwiJMCIcogcfRZ6Nwxnl1N0tJIB4AskRbKmjt+GPOEu9tDC2hiM
fIFhwf8dqsGSupOp/oZwJjb9vXRtzPA/KNWs8xznpK+VSe+77RDs9kiQEoL68pvhg89QpoUJtT0v
0uNml74DtUmEGvsdacnlH9Hrud0GQ3oZBo69WPxiqksn5QBfcKs/p0Jm2cdh2KlYxess0Aurz4wj
GKRvTxE6vpjPiBrh+l00md0T0GslHZ0BLuf9pLUC6/d3jjmPWnPMgwMGhwNwDtcm2mWY/hueaUZF
+NQyKilH77OmZq+1zj81KUvDXTwzuKeqUTmkJXauMgMoDp9aTA0wCtDoYmEZMNAlfNoyxXuyGMgR
NTVLT1bbaRD968kalbk8Qq94Ro2YH6vZ5TC3m8lgJmML5AG0kBIEqDs06/42TlwHiw6Jw8OB0GEG
HSr5pjz9zkvf9Yaax9OlW8Teq7PE2DEwgFPFsvQazWjz7Zzezpe7/JZ8Gasi4AzP96qdQkhvdCRA
ovTfl8CR3OC6RISr7jbaPGAJCqcC7Kadbv9z3ej/PmSyWPo7P38tYZF9mKywsCsZMlyW7iLVj2OB
Uas4csF1eCn6vV5TDoA6YhqDkCrF+BMbZALB4FTPt6pS0ZV5Byi7aLKjcyx8JkbJpRZCVabRDPqd
ptYqkRqu29eRc4ZqCOEU/MdXin1uiLc2WAy5jEGRd+blUj//Q2oFOtYtF2tarGva6GDyf9B9lvTo
z0sQyHeUXscjva7B+VihWkMlMSQgJFrOGKIu1E5mhkbrYekOrNK7zrF/aJNjReUGNdgkQ6LkJ87m
dC5sUxakLOyex/nIaQ7/FwMOjenpPBpEprdGgaK5dP4yKv8095vo3RR6lFqkYUTOFwUtYJAm2PdE
r/nmnww1epMFjt21b57kSiplciF6mKY6KvDYg8DfOf7hKOamKiGfqLkPiQz+M1yXvqpDpTFRGw2x
gZ2rRTHJmQjZImrRjQz9xCA0+gfoKEpC6CNsnzP60ZUGyAcscgxoW5elzlb+GSj7sL0qCDcMYGiA
Xh2wXTksDnLkE3jw0KfyllosniQlHtmG3yvVHE8wyEpcTlXTUfGQmhaiIGymPXGm+tCgK7iXoUOx
hMe9TGWY4WmKHOsLwASWQEe015e8l7Upy96hqYGrdVYdy8prHdG5L8l5zu2OixDIVoAb6uAJpAFA
DiSkwmoOtHiQfhazN6HUXnNVHH0dvxL0lKtvTVGnbIRgvCYN+/frCTujU3lalgq5Wt2l+0fJIckj
GhvR0Y1nIvXbuU2RL+SXL88AF1VRIw7e2btNLGIZ3oOzJn427U2SJKoNfMqD8WGx6IJwEF3ll1xS
NvasKAs7xP5TPqw5EOdAB6heLaB+vhj5T/va/RptZ+ZXhf/gDEZ3IAHBQab+9mxEVig2lqbaghWE
2ARr19FO0OxBxpOQVLZ7YLeqXk0mc8t4di29OMklrOcOePH8d6+jZlz51DRWNdFxqnG0n/TWMt7N
GjY+Yaq3MRW3945a0CqEB2kZfdXqge28d8375Hof7MTscg1ch3T3zzvwmKURCbrmsGnRbsDfkSGm
StKyGd0PseJ9iKQRTWPg7r6vH6nkvFBYKbthnq/u6uqpcFLQC+W3OZR9yAja4T80j7W+piH5Cnx7
DyABlcYG965E1XG4C3YCEwl5A2CqNWFgjelG7tthJPP14aa3D8BeVAgwxqGA+WL8R2hEzP4zQYUb
dK4k2YWIkU7tE7iQYgo/FC2VI0R14VaPHOicRkmMhZspKyVyRvf3sWCMP4jKfONltkmpOOeBkW1t
23r7tcHEcXB7Q9ne4ulg7mBfTuUoeVH/hspZXasJbh1nQ/Brem/7PO7WS12QFXX/Lm+uNybTmS14
xoKv/aEkDC7cwnxv9A1XUyxhdgOK9iX0a3/HguM7Udo6HBda8gfIjwfwfZ1chfNVPxbmtlyWX7Hy
KidISJlrHvbNLmH0zfPjmn8f5WxpRFP0YUnSuFs+C7BOLX3kZcu74cWQBiQnXKakQy1Sr3m06709
f6xIKLAn4B9quVIV+F7tJBQezIKjR8VPRpXIH5AHSySkxwQBdiI8SyBM4XEB108j38vJprvFcDUw
eWfGom8EtPIIFYp6jhsm/iq4HTGOWkCUhrqINahqSDmkHvEzNzWAkqN4e7VNiScWLGrg5U4ttfxm
GbCRSz+KBCdTtDtk9r6iV2hgrwPxa0DO1kfeVHzZCIN4LPLOvdcsV35Gf9AG8vG4VIuRetq7dQG2
GZ/B17fUwqoKekd3pzrQ0UyP4P1qeHLQbDjqmoShGXvVrpsczFaV8K0ntmDoiNX7vzp2R4oPpEbz
PcREQlzCHTxbX/3TqgiSJm8zQkbeQPSgX6e7nIlZyo1Yr6pGNl1vuvc/xl/vlfm3m3JRCtD9Mp5G
MdBBCN/nil5xb1CIHr1fJM7LCuPJ4pKzdcS7QD5Od5ZhldvWrT9kqb2ieYJ2CHJe8Z4ojP7v4dEs
6ex43DgDrWC0hXwS44MnphD4IL3fdFjJ44GSCaMwvzGhTDp+QrfJyHVBryBLc5vh/aJKCRbvNfZT
dPfUhT2v60hXbJHzSwdLkDIzABCgF+z4SExCN1JON35ebzZU/4yIY6bJ8/kKH+VNd5AFcz539vtb
hrRoTZadytGQalnD/ax9RI/5SYu274OmnfiujUgvxhEvCDkHQZ/s5srRWzL+LO1K3Ok1nCFvGzFU
9ZqaonBy2Pj+ZBevE7/tklR2i5wkh/wdbOqYEdbXzaCrEKF9FZsiA7JlvLFy3kCGdTp8E3YVDmnP
el88MMIBD/POnAPj58VGoG/7+596MPH85U4L6uE9ZwODHGnBH4LT1BylixfRLsU3R3qVHgMDocXH
BJ/1z1z5+aNpjKIo9Jgs/S+Mrd+rMMxEqNB8PqF1kYR3GAfxON4kYv0lPNIJKGZFmBl1/IyWGeAb
qf4u1psD85nelqwKz7gDodJXlqsjGTEO67QYYIWa4PnZAYWCERkFWjmvBsEXZTjndwUyf1C1SYsI
SAxAYHeuGXREa2sAnP2DkqOmz9QU7XS+aMIQz4O0wGCHQoZChfQB8Z7t9jCSQol5AhpdKHYE18YG
98/Jws4LvIj30xKhhgGN2uOHEfRel6Q0fw9X4+cRPBIR/J9YQB84OnSARDG7ehUOlHTZj3KtVQQB
NflQ7wddNaWQc9cbPDbFxMEnhZqoD/zNEnh0VSQoVQ6Wpja6zhyykRbm99H8bPg2yXhf01uc9tZ9
0rEWF2u4vEQ35BpAUq8vCz7LiO1tpiAF+lqTkU8gGwpltjwzAWjr+WGKcJgTtGGBrngrwcDuSVge
jNvyzCFKzF+PS16XUUlylpBBZg84so8XlsWLxATkQ9ytSsIfyT/UB70PG6zxmrxvg4lNRsXGXBwt
lA4LwSIMhXqg/NCUxOZE7JQcAYp0P6fFDk5wMY2vWnZZv2Vk7nGj8p/6WU9ycylxN3xPVbz6b9sb
RmhPmjF2yt5eVhw+e4wzj9iWCESq03BU1hixMzjLcOy3CvZ3rGvFOc8XxuVnwX5Nz6OhZE1OVRNq
GnLJzuSW/lh6cZF3sp22rp3+Zi/GcPTTjf6cFTMf53uAB+YanRhI6HTo/ww/jCrSHduoahrb7B1C
T2Zj4q3XdwVMbHlsiWVDIEj96Vt3fvAsB7b3NprIYbhBl7GWfBxIgqCg5tqFiT+fLssp+MC+dt2g
3h6PGW7s1oyEdVJtn8fz6Cy50MTvlFaIb2YJyt5WCFErSQH/CarZ0rQ4ph3YA6d2kR80kCC2udeG
Kmlwb6DxjV1iW4Vjsa/ExnCeuF44CIoFULoTboQGM/n0xatWv0+PuC88/d8FmkWVzl1NaqqcjfFu
GYCkkPNBdSek9j2okHgV2mNcP51dVVnP3iUzcGan0sd0AV760iKjsBbMqmqlM783UocaOeaf4v4m
xOyddCgPPymDcsq/fLiZeCJNB1k9sYO1gMAh6MKk4hIXOlHSmvP/cbLAA+bXAK+gfvgJSsF8XX0x
LztieXaZW6rsVvhXpZogq8m6Ju9/n7UuA5k5K+2Z2TPNLRZf3SZ8WzpZ/vR2f50G1f3t/XgJaO9h
gp1QeggjCS8FXjLK/s4kO3H25poIMfM7sKcGNfiZRSMQd/isfu2rvo9pH7FdR7qby0yLEPyNP6SC
RWHY4NBY5K0f8gf/JaeQPMTCdyGSuxZyt4EPLCD/M/Ps/WHWN7OvioYFW4yHwMbipGr7CGYciG10
CRXXnfBFWpBeEOqBpz+Ry1NCKoCaEeYsPGZKMSydGkLDT+sfY7OpoNX4L3T5gwGVZps3aB0vRlmh
P6ZAOQ9+cXkH4kFX6YKMpEqgyvzGRnvY1gseiGbAcAc/rHrRgRPpi90HrhlcDmm/Cr70nwaU7tWq
hDai14GveoNO6m/XS4WCjYCur/iO+0MIh2OROW+NEnWQUD1aHsJOmRWxuagMnz3vtqOpoWNYM5XD
rxgxICWyGlKdeVjHgZB3Th4iK5CbM4MrD3UQykFIc3QnkaCYK7Gk5PAjbYVJdKfIwf9msPwhHrks
6hI6tNX5IREWmora8haU7yXhm5/1u8PfylBPDNb03nnjuKmhocCYj0d1dQ3dAYMG2bN8GUOqXzRi
OkeY+b+m8StRI5XIK10xBZtJLIv7k6EPcWo65Q6YgIhl9/exKSF5oROCjM9pGMitex+A5CD+nxCn
dC8xLVfe8yyEyw71tKLd6kxa1fNH0CriEMMeBa1tqqmv9JkyPrVxuQGhZsBE5yNcfQfIPdIh2Okl
BdN05u6FiYCUQK36oDw6nKJVeDcFo1ybyOGCPF1+cdBMb67xuJoPsNQYbpyK0XNMKj35LQjs3Ztf
1rcwtISyTmqRZz+tS4SZusS+hZFNoIhbd6Ud0MvoMDWNrk7ClkOfr8QqVzyd9kSrVda8QkchMNuR
jRYEEkC53R33yj/aLzb+duTZY6Z2LHxU130WKjpxupWQfZSfTibjvCs0jnlajGSJn0KHEIVNG6CY
hmoSzK2QSB/+9j0gPD7H45fw2poWlb0h/N5XdIdui2n9PBb5TNxGex9Es0p734u6hlv68Fx+QmN0
NW9Vp2VF97uv0D20je6atgV9ARnZ26KqzRTL0b+0AVIaSPmHqWweIsLyZIoWtVUzEAoXQ1NnW+aD
JU0w0CxmsMiJkhltq5T/6rVdtfhCuMQsBReyLhDUD670Y/+z+6ygFj3bLu9bKOCymXBc7v7h5YBA
GsU1658biW8JD5zouLSDLjOBCs4JuXcQNxrNzakYrUz2w3MA9DIJ2TbWe0V2R/94rpcRkCNjbebH
O7JgeyuVrlpxSVtJIoYw2oFj/ww1IEP61UjopLUiCsDWefW63DAxefBzy2gysALLyFl1bflf0xQy
FV9+ea9L61ONtGiN5xxI6954MQZjVJm+SO3MygB3Q7BLE/ClTgu2myvYa/4gb9iln61hgPm5Y2ag
QqJLRRTZLPY10R8sbb8azj/Uu/aQjZycL6Ij/GdtezO/GaC57zy+CsD1vAp7A66AILYvRzLz24/O
4ddxQUlJKYDJ17/be8upHSdno8f2J0qjjYfHnTwbDMbkhit4N7LXWqVHmhahUvKpUo8BDbv57ffA
CJvlQTMAZfdFUXmlxICv+TZuCJB57KQ1QbEQ7WSiFADx7jQrK2TNytdqRWrOS5+AecrUA07EA6jL
igr4UldzKSKOESSygSO04HyKFW3DvEJTcGZfnBKN26EzL8HhDXwUqvKLkHlKMhCUIe09Z+th+XCv
YnMaQPALwPIqj7xm3JcIYUTBjoxoLmOcQW6Ba77Umu+HvZZog/QLDVXrTnVH+uHDYW/X4IoCTW3Y
8J8MaI7XCRRM4BpzmKi+Ljezp3Hq7wL9+uElBQp6P7LMZ6JlFXnMcySZXx7YDprzNxLdQFk4nJR7
4LC+wfkJNOLcuto3wnhebWYWjSpD+hMVlm45ZOmJ7rs2dNsFP+hMZRRIlN2pk1EC3ZzIk2cmgpF7
cu93VmBNs4wRY9y5Gkmg4B7WbtudtVZ5Ef9KxXDqQN8IrvU6J5xsMb4TIQChoIk87Ur+mIUPrsnx
4ElycxKEU0Vx4JjupRdYLdXylHWOINB/6GfnL/L0PtjQO6mabXxg0MsoxOSDmt4dNP9OSxd28KXO
ETJ/4tLyU3ZqZeLJUNCkWU9m0f0WF9pZpbMzglJZBSjTIMHI7OWzJx8KX6yn2B3bqf3thIKvqclx
8rGQk6ymC64waz7y6/+tFIPeZyr9EfH6mWetRtiaxMIbO1OAgEAR0wua3sBn81RGoMI3D/Seuz2L
CK6Qva8Hy1O0+Q6a8yf6tvOMsVXlwSymLQ/lxYuA0c+S82GeE5jI3roXIgyvuFHSSB09hWz1u5I7
1KKon6nUiYxP5+kpzTY6Ih4EeSQzz/frC6yCzLbyQ7q/aJCUpuXuTSI9uMH9C8I6TzGythlFFbKu
8FPCk8oc/Mb2NRhcLGGicHUeGJsGL6U3FB5bkB0pZ2JhimcDFNSW3x/eSIDgsVKfQPN8DpAHtX+Y
0FKKeMJv9YPDwu++p5F/ja3rIt/FmiuUo1vQfqbq1RpVXdLtDr2D6SMUWYD7ArtgyVf4gzc9vm5U
4Yju738YMuku1ZqF156vQLtL5BsqWfTnYHNoaS3VoYys4TdSyqA3tZWJ8CUlIZvZlAeGSmEj+5nW
8ON68UgZRrgGyQySoPVZlsKC08idbZyNbTnaNMWAczDwL4on69ZFlkzecUz8W1eyGJ+v8szlyKwe
0tveFGI+8GuijuvXnF/c1DTfoICrnFhErSJ9n4UykdtUFGGIv4QunCrv7jZgp2un7OGcwx68KlNn
BOsQYrbYkEVSKZ50LmkUeTd7ZGUno4lFFO7NRjFGSMS0fST02oNcO5MUvb/Ws7AMBcwr87dJ6zoJ
FIbqqwFp3hbUZM6ptQwZu5tiRN0ztIokzoUjyy3qCq7q09DriqpaaQFnGOKLsMgHCtFh2qhp1XZu
Ln4NFuECLgJmgW5QMfhTydw6YrhoPvRQ4vuj1Nt7mTg5lFdCDbabxtMlCyHThGPwQCJhhaXYGHoP
RfuuA2C1J8ZZI7IyKH9O1Fvpe+Qjjh6ZT+d1zTUKU2RCvtrxjYRydwLyMLJB45iM2EgsFYsy5+cE
nlGNck6AhFaGPqrz6FVB+D9v7fLTGIMA+iJLptpzhme5zjb/UI+Sn4xtlno2CvDDLtgNMqrSTFFX
oj+C9iOEbiTCr6CJlcZQRo8l3n1v5A7lCdqWXhDzpXiPYk2zkhVDASSMU1DMkJtnhtbD1VBQRrmV
nHV5yrZqlfUJHD7fb3IvSTtkyFwprrObH7gyi1PDasxEJjUuDOeI2xzC0DywQ0XCFnggb7zGC0w0
W2IpaSRFkrEJam/tVVL4yGqImM2XhjbCmcwv5rINAQDKboqrsM+6aQV+r0tCQuDb7+z6Bs02w3V8
nHDyDl8fGtAB/VCIwnlQCb0/G8P8+mkjU1xoi8mhhCbvjNA19dDxgtcclPIvev4ERXx2ZoJ6zrtv
iCur+sxTeXcg5ILRFRwMxUTh8kmlp8eMAtuBdON6GvPLT5qS/vKd1vSBUZV3+gGDhgsOZRNGS/7X
DTh0oBFWkEoqULgEyY34LcDLaI0R93Z+NWgvT3W6U5qifj0dAqnhON3KeFArb/8+Hv0//NEyDR5s
WryHZTEX7HqhrGpQmm7G0T3PrBV1w22f5WS/CGt2k6YJSYn3MqlVdVtx3atAWX8Vu5OdTt064MA6
JQcMi07etwGjmdiPoJfgxMPQYJSrrZQxRrtMUwNMePaHm4h+D19Aa4rrBfNv1q1z5SThQglGVolk
Zy+4MIz1QTaDw//eXvd2marQ6siWFSWU07rCflrJfXmPcWjgq3Mzrq3dTvz7IUaVTiFeD/5S2R9g
5vcErGzgDr0dCDfaDeovprYh8Pe33Bp1EUitLAhUkikCDFZe3JYZq06Y79itlMofNavqDcvN2dyM
B7q/F6MqrFXE3H/+ZztMHa0/SY0lwjq+/ey6ip2hVnO+yEHGJ32G0zwwLDlb6DhIlb9JXsVonx7R
FKgPDuLy7DbV2d2B+Z8GyHyf1zEOg6vGGLDodyTb/dcgdMFzVv32X2ZO1xS21O+o1EuzyVwwI0Q/
wAP/TDk5zvvs2Sx85d96KN3HeC5KCbBYTA59sRxfQvPFtXUFjpypQQ54RQ3NpDKrZUQy1BCcND3b
nxWdHS0omGDfum5FO7KZ40fb/TCinIXELxVA+kqsvZ/de13Od8LrsnT5M8rQX1SZEV/5JTozPHV4
BigcmS4rdqOqC9LVXDMB2pw7whj0kNOKvDJLka9Bw1xxOfBLGQJ4aySIPR6SKMmNDFE7Zaubo4BV
Z4afzLqqlCW2bdb5GNNOQq6OFN8KaT6XFdEgxNKbfz4JInR6LWxkMsbPJauqyrmClZEuNOm0SHP0
79LqXTD+uJXiehcR/DCd2s6+r+UyrCFV46lMWJAcNhMq9vqC2Q3C1llDT5Bf3VH8Th69BushPCZb
yUv0PG7mrWS89rIy12iPQlIMRof1by4jviAK1eVMd10krCllkKgQzGbOJi5t0kA0q2le7uKP3gYa
Zd0uaLOeBG2rK3d5+ivmMgf2evdyaye+i53SA5H4bFk7Rc5cRw+InCTz8TxOmdk8aQCVHhZutTZo
I1fQGk6b/kOtk+K0Yqp3TuS6E1QE71WQdto7RbZV0zTFehZ434Up1IEg+8Jgb4hDX6l+ug2eUpsO
NNsfcTt0qC0Rnh6S7lfgA1t62MkMwIXPumr7Z+iBszOoGAfPRl6mPe7L0HyqUjiIIqcChdEZl96m
zqb5m3eEEj0SSfAXDjjor4MyufGMrRhaofqG45eC3IJaYb6dwOZW1lTU3lw0kSl7y/tE0BsW5EeH
kmVx6Q2960V74F+xBS7SVZYGIClw4jGBsHxouUZftMVxSUCzLyilzieVW8bIdV3UFXTohklaGCEs
dTQRXTr0yLQQVePAYPIh9sFXoWPbWAjKaHxwzuwXulzviU2zKuiqHpnOzwOGuoXvGXn+PblI2is0
oGhI8TQwyyf6/OaBJ5G52vLBUadGwFxY6t2XbnMzYFM9Gslfd0/banGAv+3sJW6ANlzxrUTDL4f6
Q/Rtz9YoFUC2QMEedd3tpOtxekfn0e/6IKOWvjiu2V4DVIFWxYIfLJLTkICwfFh5tseuMf8d4oLW
yNrIPwSEIhANSt7FuMs7/Jpul463TXV23L5CVfHEcmMYwEq07YayMKUi5XY3C2fr7mWFVJU91gjw
MlJKj7eBfZ0hJp6CyMn93ImL0JgobWGrj2KebOLSHRi2UsuWAp0wNf37NzuJ3Z767t8FbI/ibcKt
tsF+ZFZeWcxhnrLoKyH/I2W4yXo6uGRVc7gCISlPmDLHoBCsIPPnKsE12p5gbfJWrjk3QFBoNi35
HKU68/8IrtytzyNo8abmHzytqIO+HAguJ/nIOBcp7b87igoDs/xX4PC1aie0cLLRn9kFErdMoRFA
O/rMuWKObtbYD6W0eEHL5KBe0rrvJOTTUMwyBXDrJARtuQMP2rc7MftLze+gamKr+FLCbjLmT/nW
dghBYw76dvIyFleNEqUXAu7CBVmrEunRyx1vKlCJWeTFWhrkhYFAR7zhkpR1vneSSS5XHRwXXXGo
yK4KNgJYf6BCpQsg1STpbVlkAp6hFLDkibz4xdup9S1THmjN9E9vWEGruWXiXzi88rvxOD4e/6R/
l52dnH7+rqXNcD1nfw0+QDNcBkDqtL2eIw+2jg+LRjyY2QQn3cOOTWDUkNk3Nk6RCXnmjqkTa2ZH
zXTPEMp797TtDWEuYnHjT92W2cRQ8Rsn0pPR8rXYS1t38mkxlepMWHzh4XyuDqJxz6l3SXoqYkNJ
8q6dV8NVCcQ4W5ApHVcCyTNDcZFa/+90DWKQ67o/hHl9ijt/eRWFBgbGYz1ePUbYTIsNW5ZyU5EQ
BwFCToSXuQctDRdEcWjtDBydrWwJYVYfbqo9KbGjIKB5DScLi9WDl4IIXGTMYNCp+QL2APhWviU3
XFh6W/AbJjHPXywv/80r7q6n2JoMPG4Wqc40n5/F+oupaBFMW0dyrnaLesSQZR9AnM8eO/CeuCK9
JLEBoUvJ+IzwnFT+CFMWkFf/vBMwC582zOdMO+VL1wTBZF62EySe+xHDuXhhtfcihDs9NcSachlQ
IkZichXH0YlLemzDQfRoj7deUic1O3btpBUGTar5RGUlo1IY4kjcFqomEIUedMftafN18mZ6KFNI
dijrYZNlpTiMW9K3n9D9WKE5p0t+3591Cb1hvd9HRgBKCumD/DgWsqJTeXaPsv5mkpW+fwmEZwiT
CkgguBFlnP2/AfAS3/Q07ssfbqOZvl0gOH0nKyl9SrOv4Vrw6IWLyzb1fkBEeiMyFxA+lVCFywWC
BFJ+4sDWg0mr1Nit7nWTIJV2st4nxV5KeKxQCKwuLyRrfPYvn24u/3n0zzOgWcrZ1z2AuIlMH7/L
QJg/D+KrXCDbI14KFPuFULW2pRlbUDka1j+IpEojzCb9OliGqZx78U3kBM53na7ijYhgYaq1N+l+
8szF3WKoeJ5Ae0cEQlqprEPckU5iQpFG0BaJzbM18Bv4V5hkByz3tDaMQIh89+Bj/4Va1pe+cSTD
fjJSV7P2kgR0KpcrQHPiP6wBaGbDuAJiW0I+1mpOCnYxQ9u8UNzU1F70aZuWKO5hTLUUEWiUtWFj
05we76GRpDdMhGBPKCR7YKdkGDjsDvmEqxBcQZi/bI/IPejMQcfWs9UoebcG+8AywqOrIHHtCzvP
H0HkFDxAgfOVZX0eI+pVL1L0bNM9YKVjrATFxV6EskAZ1RR6fejLEysWqJ39kcitgYverGAZN6gs
MRQNDppqduxhoECQJObhmC8JrXsfAgI95NDoWR/r5VIaIIzMGYmvlMQY52PG86Pw0HAL5VFMm2ZK
KbezQOaJ2rpKCfkOcDCLPh6T4KWDAwY5vyy/pVpwLQFu5RKpT4f+jkqzGOy1DjS2KPmKefkETIo7
qMuhMgwUSuHXpPxUIFH3ypcNPdADjmLwhH+VGSwNu3lAYcpNFbQRhM+3uVKgK5iaj6PyzkrSMi5p
mGx3svAuPnLbZ3t3ceBJy1DZU7L7YoR5eBrAYaT9RF7fjlVGemY7HQlh+8QOweVjsGgraTHxH6Ob
pyXC/Z/mmVzQMFPBPGJTMJxawnFGLcZR/dF+rDTCPd8Bkn5XdwMzd7kXj9mTaMFats7qaOSOX5VJ
ygux1qoyZjxFT7n5er9WJGCVjiY6pskDv7FJr1dgFS8ijn94NjDFdyA1SR0SRhjoFa/a3AaF/sok
BIBZIFMlq7/glFNkqphHnaF9PcDp/iOYzf0Y9Phs4NuwA15jz9quTIlOAxPerIYwfSn5zqJolnj/
eN0qShM0hg16ByApmKJ/0SOdifb9lHlQP7M+CCKCVz9z9poOnSR8NmHGRGbVO4IDDyLVmu7bEL/g
y1r7/OQY7kZHdnSpP89+FNDim2hobeK0DWjr+sah7b9eW3QYHiBeBwACwAdiC4lLiKmQ52t5T/jt
1P6Krk1VFdbAK1Ch+ToHYVLxTTIwQrt7EshdTtSH4/5hVyBuIjn1RvWnWz9XlqOhDv480QzIQ9K6
9EY/s3f83IXBVObFb0bu72EKTkNNurTL55MZ4nN3otu3l+sSfH+nD7mkScB4s63OamciVqdEmth/
RYE2A8RHgI5Vh73EcNOt/CM17N5G1Rz4euUhppKYQAdVF7SmE9+12S+TEiSDy1yshDE9HHXAXjIO
9O9UtBBo6JXjvunnyRaOps9W+km410G1YKRDC7zeX/nB3803mpwTkKfvF5alTq5j79WE4M+MFzDv
UiEDaG0z3hkRUlgqXVMb4Sgfy0GcTKpYnodT0gdWb6A+VlYVBCESdhsV8rIFW44C3A7c1tM2y4Rs
ToOvkUo0QVv1AaeNxp25hs1vsb9EJ33lGXzJvQw4lsfUsBB3hEX6nY40jwTYarGLxaGvgrNjNtWM
Shr6vJqD7uMGwBXWHsj22ijfZiwO+UckxgYT3guxGn07Lv/lV2//80V7hZ95IsdlwS9Jon1pOzZ9
yzJ4LQ2LZhfEJSBLKEYnSIHOqkzYwrHQb1xJNbVZYbANIQuAOQ0G6JWjL8ev0SdZuvGn7PLqe2uq
48umqLFIxK56hMryJZMVs0GnOVGvge+gxf3ezyg10nmNw7TNvy0CUQDmP2LXARArB5BSLFXXVnkL
JBeYJI8ML+3dxpW4dLs2z+/3LMmExOiAQdTVGE75k9xBH5C+/tzpPYaiVIFX6swQeG5l+Qe4fJ0s
7Cgot24d2gh5lF/tfAK3dPVxkGYOPKoAYP8UUwnVkkaqz2pK/rraEpmRznRXRP9EjeUQvgJHgYjp
1yWchR6IvtsrFgQtLCwMYSbxfsg1u/hbZfwjDKrpNmJSNQBl4qpKcjCIRu9mXakOklD5e5jbovzM
xShMgI1J/vISK22gBmkSmBGGJfjvMqcOmusVMdySI+R9aE8SwajM/KOkQ2kL6Tgl0gFvMASBiLYZ
I8rNQr7aj9+VGMjr8gj2LjjX7c7x2u0Hay7YIs42IwzPhBlzGGt5/pjADAtkaAnmfnqLRQJUsxTr
DndfFhul7ei7uofpFOk7okHtw+1BJkvwNMCnHksLHJWlIo3zh0GMsSG5LSQCJ7ccBPW8knpp2tA2
pFH+7oCZLpKFPp6sSDerGsDBirUPypqWbsmWdjIJItOBxHFnXIa67Tm7F2K0s9y+QmuXxK43wsCE
SD/WzOURPy44YofcAUOYn8D2W5bK6ZJrENIQU28UyisxA5f+Fv0drXHDY/H4GZP5KxEDmdj0M+Xn
7VTmon5lNTdeOi83r3GYuy3KvVoeyK42yGRYFb4gWoVhR3hLbOEn/rg+Pnk49M9fes1Y3ktFZP0k
gxi8azIAem6LdtaVdCpnXbIEVYQgVmcjICGr4s6LRjfqqrndlCTPokiNQDMR2PolL/fcdHbJRQpo
cKvLA74hNsU/2P6JW4zCtje1eOyvFZup7bJ5CiwqjZo3OYE9J4rZHjmRmAsRijTAyveLslPKCN4A
Q45137OgQnXMal+Iq712P3pdVz8jEF9Sz8TSgL+mJiAQwaJoUeT8hFV5tB9cJE1AaDrFl/cwwbKr
gUSuTA8myQYvYOwruCxuYVfnjpyq3dstQKFrFBIP8liCrus7T3ZA8zRXPq5MwD24ehwkeM3mojdw
n7CAZdNxLHUiyIsH5n0FPU1PPe89urZ/JNsQs/b5KqrqPtZhImU8YFc2MynCwjhlTRGNorb0w2I+
k+Hi/MzfisfFPeljyCev862iSUkqA9TTxhrgdUDyyt+yNAO1ouG/p7nTQ7MnG3iUDVU1RC9b1Z2n
1eEbLAj63zs+qor6sMdG5a594jgJMdPz6FIx15EGxXuuRil+IarpXXWsmhuSsITN9AJbr+5UEatV
8qhmtieF0PHwjdNDEpnijJuo3huklwHqfNWCirmksCFZsrZL7n/6TaJKJs7tB0jFIxJvnrvWB/Bq
1Nik40LdyCVRDBBxoUQtb4DnoLk5ANuXFFip4/4CeV56bwPV+cDLIJX93lZn5GEM799SDP/23wo/
d+yXYz/zZfqfLKqCj1TMbVUz6Z5dXCI9MVxVtfjXrGy9bBTZaD9OQDQOtjuDDIjKDYEDrDBBGw7+
NdAq58j02qAuvRxYIpjN66sojGQYIxURXQxGBxwYEmvYmgkHwIee/JZIkQEo8CXTNiA7I+0YXRFx
cfYbpdRqB4bwm5TV8TaI8zvBpmFo88oF7kwHIriEGRR/TT/ZuT8c9ipxsdO+Kv++Ml/okTFDHSjC
KdhtLL4NgjS5k7kRZYaqRx1DK7NYJVzP65x6iepZtUZK56P/Jgog1+e/alKSdxEKdcCgtLmzTsLZ
fjQRMHvWwxA8RjlEowEuyMSIvUKuJgZR4qEvFnhszMMLwKDnsBCI4R+9lpjPwG3gVTAnZL/8JK7c
9g4bCinjD01SdBMCbllisYLgE0cBvVyRH5A4Zz9gKdJcqfg9TAy3fprfqkoWugJOyXKZaFEQ2kcg
ajLorw1J+ACOtRYpjSBfbTvws+R9xapVorSGe+GAsiYdAcqC+MGrxx3Ko1kuci2SZoNH6i3Q6ZLQ
K2iem9QK8WgNhShx0Wf8u8KSX4IVlpqj6r51iVYNB2tjdtvtdVOPXOq0j1DH1qt4AUQV5aLdO5AD
3iJNmGlQ48gXLIagGmY9iNFakqOhFSKY0QoFXgJA0eio6Au18c3OVPUZkuvPC2sJRT+zpwce+20X
L+CW66b9SYAiyJF6/NC1QW8WekHlMkvD66WruSXmq3R1b2ZFU2DtKcJmNLJ8DCe8cW1KYs0I5ESC
+cVMsRicoox1rygNQdr6zC+D95QTvN1yOQhEygBrutOMP1f48SZ9vAD404qshcIWVHKMrVBD+BVd
x+al25wMey6475JuJUfku7dY3iNk22zmjqOja/sV15D4KC8JLHvNVDhWKWf4T/JSQEEAzw0lbgIu
mZwIrDbiKPWTardLu9tltyO/ZoUXC0Ul9Uv+B3p3WD/0xvwr7uFdMsZkKFa0od21kdRlmGEM5yr3
B0U/ky7iNzp/z/hZkObM99LgwlicdrvlULeV2+01J70sek1EpaBUtULj8SpLGaHwV6P/8kOqZpYy
NK6U22f0bKvOP7xDtxu6uS+KF0xcJEHzdwYWJ85Ov6xyzIwo5hAdN12D6yXrnMsybGuhdOzAM1lB
BecHZlTgRl1/y70NXjI9t69jJnlnIDgxzylhERndYKF7KqHadAjzeeRckU1lI6cK1dO4tuTVxNSV
E1veKuLWUsbkVM5a1EXl1/tZbf4e01XC2htek+EBbrSOTzaH4Qd7SknvuSC2Q/0NhB36wQ9257Y9
M0O5xhwnvOguc6lJFPjnB9e5y8D/05IZ0HSa6Xw/dbOih7JHL2SBH1o3QDgQ67pW029tq3eeSd0E
g2LEi4ZTQzw2LpvaI94MtLcIqWGcZGnvJ9ChLkwjoG3SSMIyIujBCNMtXh0RceYkqRFOTqipnOKJ
WItvsV+h9brFRaCbfNwwnDpVgODqhMOtN6x3fK2OGspFv71uEuEPzlOfqAS9N0uJdLREtUS/X7qh
7nbjHaCg7LS8IMAyVUnEsNb7o9mgah9YFw4Ypyzq+wMYF1vX6945C7v+4eu586TU+ZuckDFFnKoZ
8BGnXEVb0UQ4POUA6Ym7OU9177nLReIZWZBtCo4s1T++v52kvCZlwmOTgIeBJnMWuq/OyjrBRtRR
1BLUbD8UCWCci5IqCtv3Tm3C0LAEUyDACsPAcosBnO1SkdSaLJolTyMHIh9izM7Eglacurky7KHW
P8TVxYAtliZTZi/5XuO1DUJASiqtqoFR0JPTlQdhPSJvh/JgHCtiuon4OL5tgn0ry37D1o5uqiHc
Oip9g7O+f8ovslR/jZ7Sf2julC+XKS8DScol7sRvZBNu1PlX4GOy1K19sImHQMwJstFken12oxVC
ss4scLJNdTOD5dLNZo3pUMlcP0/XyN+HBRBuIwKQFBb7KAcpNAAhyqpTlBIr+slkbnxP1DT49Yqn
SM8kNOk3pjWW2jmjDDBH8rADS20Eias2KILyZQMbwBX/ecyjdArzaDT0eBZfOKLj9kvz5VEQ/N9B
0X70d7/3B2EDIRoMySduNPTE7CXimxMJlCFJZuS3VacQq+dE3PFiasikhFN1oEVg2tZnSX/CYfm9
slICL+TrBihOjUBrQKK4Y6AJAXUhwoEKdnW8DGsiTYnDXtPbR3LZhOSPhghpiaXXnp3+gkSSpnS2
DAFEoK5qQpF4ob6eKZ+ipF/ILOBADoKYQDBTcfzJv6H+eQAGKKC1kHrY4Ugj2hCQNHPTI+HaWac0
Ves0SrYsOAtumdVDG0mOUWx/vc7xAHFrxrifVPlmnH/gPZ6Lc0+o3aaxtAwqMeI8UqODk1mgJZNN
a1F/MFqktOM2ctAnxBUKISFKcC2RSZwDhdImHhZVpvk8DTMs5VA5CqpBVVF97AdcMGQulvaGcAUT
clj1hh9zbrZdqyM1yjN4zDUDplCgL/hsZdgf09EdzVukFb9aGLGplDJLeWvpijhAKb2QAOAIzn/H
yEvkz5+IDU6oSHrMqBajoocHSGUJulXRUmg4o0lDX1ICsFXRNziMUJ7MGdpuV4hfNGfke8e26hFY
qsJ9OsTfkpbaFRuKayVTBMGSMYn+N7rHZLZd9me2l/E7meqTsy03hAiyWSpcv2I2VJR0p41s7t4c
8y8dYUS/AXej2NGyFD/DSH1z9M2Pk3ChZ9cYFXE1p1gfXN9Anbgfe1Yn249zmAYycdRvZcYWhA/N
dSBunZ3h9MNKLeEUB9p4FJZNEH7ws8FgfR+z8T9vQUs+dp6y4GMLN94SuEo872+/5kLQNcnnOhSg
qQ4x2oLfiAYxluXUmq+8vlp2GepB+DPwVbH5qATdTgRy1S8cRAWeDTdSJLSPGDysJA0DlxkvOhho
4XAKCoUJ10cT+fn9spfSqkoe9yHjxkZ5Uw+1KboX/C167QCnvMVdyqtVnv7QFPsOUDZYgWKfqfCP
yGpg+P9+ypqoap1pJc+Mxt/nf4Ru18evVs+YLLWRIdfHRKxWT34I9q8qVvRGyqK9nZvgMjHcVJJr
K1X+mUpZOtMJEzjbI1KeXR6XX8iMMv8IlbuaKuoBQxYPVIGzfyxbDXcmaX1GMtGudBauhrzaU78c
rJgQ+QEB7u0FFavWqfuWQHkHeuacagoxBujPytgL5ba8o7jSMq0jguWklQWwhw2XlfWZD7bfsCCv
VebYKBjVWHxzNMp9RjcyWWis2+sgdr49swPsYo3op4yRrj4O4Y+F87IgEFbpZQLhLN0u/JXaL+Om
Owb/buB0X9FFz8HRZRJwDhfDZO5dZX7TSCOIDIm2mAs9X7IIueuDPqo8EiEPHJnj3kBi+Dutpdvz
IBZqpk4dHWfk810UVRuTn5CLKfO9GLLPC+dByeCrGPVdJvHYOplLtBJeFcrrg2Tu5aqBSIDNUuXV
v2bUgpOXDbmrSXuBPwjsw8VYkMCVhAiVJ16CcoOznvh9zzaYV+H/fwUYgvOSQW8ObIlk/dxb33+F
cc83IyxQgkw4F6tyFimB3aGMGkzw3yaGfdWUZUOO8CnvnUBYqyxnSYq57n++aLoYLjBLpEDoh1yH
8wdggukrFOgVONLL6/qz0QuB1wlhdfBzw4+rUUBLeMtM4NYtmkWIaxmjJuyKfWA2BYnUOC8KP//7
atmUNA2wy/A1BbsC8wyXGnt17d0uSIrz5XToejpMYeqMf+RrA52z+W+AEvkcsvUQq6+CAwR05eTi
lNNhR6kTCKnLCJBu9exMsi5YT2wYifdcW6wna8Rm44pWDAqIUkecqnnfWOCEepzQCVf/DeZ9Q8GF
QXW73NigDv4Hji3MQ9niGqRYF+HpQMoLvMdCePPGBXSiVyw8hJ5sWwNvZKW2iac4W24s/o5Mdlfx
VZij4O2ltfAepfB5HHuyZm8Yi5PLurEblNrCTCVYiVxoi7Oc3tkw2cf1mXkVUuEiUD6ZfvuKiNEZ
Nu/KuzGeOKbBwWXuuLU006bZQXRywh5qT9uHFvjHz8Xh5vSjdqDF5UpZuNGNlWLcIFavoOj8DJh9
DEyV54KiH/G3RB5hgdhyFfk1QAmMxpJFJ3bLTLfSJAigU3HCdmN5IYaBL1/RnrXd05H73MSVV6ug
XhQHTI56q7AjOgaMdOYePfZOInqri3AERw9jcZ2zt5pufWrrCMk2oeaaTUSGBhe15p0Rop0RHO6G
sRnCYucNVosAN+B0kphHae5OwO4/YOw65junI+fXiD2h8pyfLiBJgGS9OAW7oXMi7Lsxz2pyThBV
oua/VZulApDt+ysTjhUYCPWWLQ6970VYYQAljYqeXts9pGPJ7Jlp51EY7kt9qAoAzmeE+zaQxXEA
3X0YH6jcP8YbwH03sKXFMO9aKlPlsxkP7sw4IE2YUOK8TiVGZ0WpaR9B/r8kNxUpiGPYkOvil/XJ
PjCHIkW2qZuI42kGq5ViJATINFhd5JeuCqxBdjUUv2rluH/HQXag0ctlJ/T1RC52CFxZVXRg8QPx
cwolmw5XY+wcNOXe157QgeejEZKnFV/E065wk/lBkUsQ7985QFq7SIaZv5cbElOxecMsK3sEjwvO
1uQfrGPWp3Hd92yTPs2Loo38jv1p5+MQdb43OMdsyM3xAvggkEJdMCWtojikA7CbdKLAvozhCjAq
GXZvjpG8qs6aOXckCmiIJSqWjbSYUsBnYjDwtbgPiQPn8VD/1capmu92v52+K3OpNbRYGcn/9Wa/
fbh93od2Sgte2Evw2AEcM/dsu2rhUyuW9ZM5LZvukQo0dw1Mey0FgVxFZQgeeg8WiNX8b2fQhwIk
d+ptbmPEfJdegV+BUh7+i9AIXhARU36lrb50k/h42vMVFBtujaYCZd4rBE1HeBTj0jBrgiEQKKuf
vyXDq+X8UAjOkp+ZTP2oQQQBOYD5cdofMlQ+r6jE2KL+cV0VCJJL1JIAWJvNX9+guXWu2Ts8hBup
e2rUbJDlvXI1X5t0gX1m8S8YsXdjhNGfrLXpp1FmVVUe/DPg/bGg7sdYYArakGPE7nFe3IIu/Qqt
mlxiJ56MpDmlZLwUZkrOPJpH/kUj8c+tBKc9Ci0qh+eNX2c2iQbScks2L0tERRHMNi7UOU32gOlE
p49F9ugUek90QwDCX9loxQIMwGNYtnIwJlNwCu7hVabYOCiDfAYZUFou3emlZMb+0CofQYOqDeKd
MZhJkhzgr1yUIYLcw3Gb+ueAqr+0FAfxAIsQFr607CkhSf0fYOXgb+QPIPZ+9IZQvMWMJ5t3d/T8
oTefi6TEqq2mSBxnFOrhEwR3xTX2zHhGcEIS1ZDEaWcAhPReTtPiWUip7fsog6nL0OosCqXbsr6u
AIisepkIRQHxyFTBFaSa+KYxecOcRtEyUB6Jiez015D2P+SOyPTkBOb1ay6wg6NIKCtIQ5vCALXf
HyMsJc9CP4Y6yDbLkvDnJV+ftOj53ZKa8wOmGl/73oC5MoGMNvbtGwdD1FEt1q5U1i3Z5SOu3dVw
uYg3wcTlUZ7J8ssgSo9gbGv9fSq4drR8PsPqDMhJY03ENW1dSMz1vBk6TXjgGHCa0FqLGdK6GRF5
x8J7IIWhDcDrcjzkP6IDXTp1HhrY13LcggMrlFhDdiivdPgxXRlGgWRWpbdZN/YAA7kjae/rANBg
3N5wJhKh0tP7xAfg7M9FSZlSpXKp5UBV533d6bBX4CX2n1ZpQWurKmxufMs3vYz6rtpggKG5uide
Hk0dZ3j86odwP9P8sIKSi8SZVsOaXvtL5J4elkIkCvGyEVKXAy5KePAavmMfAewGbcqbD18Mhy1x
Ewkt4iJtN5329knILQOKGfRJWgeC5ds7FL63FthWqm3Heq0p5MbhfbXJwD+uLdptMlM8qPhAxBOt
eW60pFu/zfvRxYOK9P/09no3i1Lbyivjlkywy+reldrn8geJ5ocPFQlye2QQ0ETr/HVbXvNL7awh
Sa3COpzASCVXu6qHqZTLJ9DyEu55jaxj6bEhBaQQM1mZw9RMvToDyO9WL2qdYHo/wlQxIAMOCh03
M0fqEAD7KKZeIzrzgBMiv7u9fqpFw0U3t4pzdwe5delmNmtLpMOpxv/Df7Ynbv4tMhhVDOCiwWmL
EUtZHW1XMwQylkXVcldP8B/JAqVRkmi6rI9mirkAukrIbnFEZNk2qYaZAZu0oPCqMdfvjrG7tmWo
hChTVPSj04UW79JKG/7A5cEhl6hYFZXtpQnfLUlKOPM+3SdiH75FhpUhsi77pubq2008SDPSzRrL
fwBl4xlH8akpWP8sw/+OZnMkgYBy411wtM+GikvItBxwBxyPhdOxjMS87l5x1aRNCEGBKPV8Lisw
DFmXB4wiTUWbVgv6OHSHkL4fG8n+9pCRPHqiHuybbV0eH1seWoNCSAV4DXoDF/UyEdTZq4Hmxj5h
OKGDoG5TGocr1iNdbTRawHemtrV5SrW2alaMM+Epxr6dX83ASQQ0Sfj2YS1RhqT/hk6LQAqLWM2m
214dfbLU81wharA4poebU1GU29tMZlv4V/Qw8eV61YCltWF8wyu+A+97pxH02NdAjfOATN7bZUVl
QFGTM8jRpPxdgEP+irsNKtWjyfDaJTn/k1GIlIu5MCmw+Lvj43TJh+3ZQp04xGHCLEjeD4HfcP8H
vaY2Ndxz2Aet1QT8Z3xoyN5Wp0pe9mp04jh2kSyk9i10Seq9e4Y5sDxY9FHQXHJZNUKD+1HpsU2p
H6RlKc5Jo44n/jKaqGiAqtFILxJ1oi7oBL44PPozCe/pXWbVVqnV/ckM2nTCa0+Y0lVESGwTvSwZ
WNfJXjiUlOnnW+PEkeO/VNh29k44FgADfP2XPkXCELKI6v8OEGvHzIbS6PAjR3m2bs+bGImx9ONl
uNDJSQqixl6olOtag2yvb2HKAYNLp1BbleKA28Eco5pwcChP/FAzdeCjr2oIVV4i+yGt55C/TzHt
dearRpZRvAELwwqqTQ8a0mpgMdk/Y4rSDhz/bTW+23cTTlJYA6JqFEbEGbHIxRdwic/vcTYE/Uil
E6psfUQ3vhMTw28arWLPsTTEb2X5nb7xH+HoT1vZzIfBPYyJDn1zwT2KlvK9jCOQmdYAzIUWYGM7
BZ8fj5YaDT9MtwEUHHels7Z0jPWVOTNijjua518Ely/c/GW45TOSP/g6EhR7M2XyTXc4T897dlnA
yE92gsbIh32uVWM5GzXZ8353ouXpJO9gjve8f5S4KZcJbbB3L+8RWCPg4DZ7+4/uHgc1EPFzjOdI
l1D7A8h4aO3tioq/GOdIwuSsSfzMRoEEwXRn/C9mDZqKAVVqUuu+O29nogVKJeWiLNBt/ykXOfIo
MUs0W8bmOM/aS9b5b7zIELt4XtdcJFiJBvnM0OY+z1ZU5HuUPMBdUXWMwe6sjc2bXG83Z2o7JiG3
lC8BeX936fZhrrMwNHNugnPdHup5E1aKtwbAVCSxg40dZOo4KFB75yoDmvwDsV93nev+Aiubv7EM
cvlrn7S7l+UO7ugZaMAwcixmHRYXpSQrH0fCmYWfC8XEgXbIpRR12aTSMnlN8wnn6CxXF8Sx0eTt
2e/lCxl5fD01lsZFkLExUTJ+bm5r17TfFDWi26sUop0aK4Eq0D1jn5MEkgfKoRPPNGn2Ctk4qMm9
KnH9FmWZlx7J+m6ZI5y5k4Y84SwKClCceSVIx/aexKdtY7XmsPVdpZHWM11ikQWu8tDdngDpSisH
eutcQwUv01PB1wIo1oTFxa+7gCRl/eKtrky29afKM8dnTnX5VdhlnFh0KH5aZWfTP5hV2CvhTVtH
GxQktmREPSg9qGOpdGRt0W19G/hdLqkTCiNu3su+LhB83UViQDzUy8EerAyCKUSna1UnXiq3SDNc
ItviOHNanchp5H2R0gz4AsVEqLjvLmfdoNPonxOzTaOzNeXsHNVCpVCxaOuTZ+eOFwE6NJzzcf5v
Bk/29AqXIH0x0Ep+/tvAJspZg+6IB6sNiUywenkiM3a37uBs3iIhxWLXg9kl2GNVMsMqCA035uMy
qXB0gWWHs6x+NkbDYx6+B5DMnj7NhKAf8OWGBP6lIHmyX1MEZJbwAAtfpEzot52mPOMGSkJ7TV6e
oBV7qWxoRgl2Zco+vA7+7my8RG3AbAsdMYUOPk+fhGLYPC96EIuF9hi8mlLK/7ClE+AQ8mX20w9v
PAKcqZ9sdKjGVoi9hOOkdHuOk9DHVvKW+5RHUaS23oCkW4gilQNSfjL2O8j29PKgoeiIJXN9YAmD
WPC6vX1QEZDfP2dGMQ9I8snghytmOJAbgyQaz2ZbJFe1KyoB1NddKgCsGmuGuOfWG9w1pVJ8F7aE
XgsBtTMi3uZTB+B1HZpsprGHJmCuztir2Si7S2dFiqpBVF0eiqceTggC5QeFYFqemtFMrmw44A4J
s0UWlxiQuXKlDe5kQb1wg70OX0USwmT/00+tTl3b2gvVtAuYaW4TOoW5jnLO9UcaLzKD3+NbWXR6
I9yL5f2/ojGSfVKkjctxnX9BTo2J/9puPUEysqxmm/GbZd7pfVMrl33rHLnTGZtneUZuJnG49/b+
pfAglNcRIAqyHPFxbb3ryCs1l1vWU2NSI4FdYYMNzlj4qv2QzSbcqCp1lJNALQliN1MeqMWVWKqt
W3e/mAISsssmuM0xfrgu+p4u5KzKoPCRwrpkjyJDnFSwaKnYvPUnPer+P83pL8TgZlf7J+KtB3+3
ddmJt3vs2TgtJbyD0YhZsPKALPdwdwza7LMhtcx6W1vcDs6cWhja6mDtmmxRkIUZKKfd4X+caBZ1
XCzas+k9RCuKfRoghPnsHFEeU6Vju5WbNAD9a5kTUipy4uVWgf/hH8C7ok+7o7XHJ7ElT9Tz8551
ahrzKDxTbp8722WvOS0NC+nmZtsxAY3nBaS7U78hrBUMHZha262Z82526DUVtpeyutmuodoYtN1B
hZJr3r4JOkJ2r0rKD+zameoJbrrphPcOzoqLnZc2zHPhxw0RDV+0Eo5OsW08m6PAPhbsKJd149P8
3QfdfrSH0H2aQijys1JT2N6v1XschI8hwEYFNSC39bI0CHqJtTyHI+M5WKgWutm2RsmC1KALC4AD
9foWToVrkpd++huF1fF+QpUichh5ci/LrONi+n76GGvWWkHTi0Xqup3nCp90u8VKzsc3/78hzvy/
6SG15iWDEg/iw+cjITSeXnhPngnqihLqcFDjJdj1BXf6Nlo2xHvI2YoKzzm3XZxLNQfJv465dDCz
deUlh2SoMUBOEsBcDHOwi1N6EkD5FNAOJCT0or2qXpL9ZJ/cacTunNKvWx1PTyjW7++XPx+BatVD
ajGfi/PZd2L425MvmyABuu4k0Ve3GN3Nigw4K/Zua8bbLj6YWRMgPxS/eRI9c3JfRCUMqmxmS4Rw
tl+DVuY97aiaKS10rs+b7MCxn0j+LnJ+oRqNoaqVuxYninwd+v7uS9aFANZsM7Wl+jXwKc5bmzdR
SEcfWCLVXl6tNa3hTcmMkrvOeLtpTQrH093BKOEtrUbAwQfWJgRFWwnum1w6KBLW+pkJTMKI31ns
DTggJAuDMhZiqQb3E1KSnURj3lQKfQq0WMTcoCA4tMmVApuD1kf2692G1igXhybjnAMIP/vz8F+o
jzuFsj/vqauQrRFaB80MX7DSjjMrm+OZlSqslCX9ttXN+yqbr48WeMjwRt+8Kk+lOiC41Onsc8q+
vDfDK36Bq38Qz68/FZavMUxeDDQrdT/+A/tJz8WGtVG+mlAxtRd7MBqXm/+1V2b0x2ykfb6CQtbv
exz9WcYkO/KL944b/Kz4obheLwoB6RbyWP9MbKPQ4qIginrZfQJZoSe1Qf3tirubOUYcirlm8WiU
CNSVnZItuaL3qHr3t/hOnbHb5aJN50NRq/pHCh0bS2/57kezf9S8Ob0Q3N1IHsKQvA8aImug5IpO
sc9jsJiUoZIW50e2PHscaXTDg8TG+6x7q/8SY7AmrZHHNPZMEk4Wlb+ybSRAOSOOTrR9W+Rfd2eD
bgKrWBBeZmDRmFc2Fv6kWaU1DzB2zBYEC2OrpPtCm46VxbOpkpSoL8kTo0NaQaBh9yAQ31cPNUIs
BU3xD+mwGwo3++ym3xrgEBHjMIiYbhP3SogCdiXa5Jyw+38rPCslOhMDUcjNRGLsNLKCLaJYWNwi
9TdQK+AgRVu1iSeLUWOqcp07g7lAavp4UK/bwPSGBuEIvXjA6m2UrY2e5dm7rhBKVkCTzeO1c6lH
DXsH5P93EKDZiFeq3ChjmjRVJ0ymss9BHxwwRrCPovep6F4pgBvQ35c4jdpJYCSA6dy0rBHn2G80
zUdgThXYKJ3pG475oHPChl9JBPEl/NW9/+6QaE9zuZ2RBrOZbtSJudhaHuqDn/neHMK98aVbgozP
UczrhrJAjBCLMasZJoTGRT0JRVP4PLAsEuuOQw/YZpOTxF71HKG8Rsrqg+7PnEhuQeymZCWiYXAM
NOKeSOLpeTbhaDtpBMJOaAJfOGt8gaKtjHMnSgOvGltcI0OITyzLr51I7kS+tIFPx3vK93N9bCDZ
uXA2BxQg128Csego4pVnMg2zZW/srqnzwrq2/iseC36mnL4Nya02QPZ2viMLBfm2Z2Z8WqMdCkku
0t9ZukGZTAAWM8ULcsWUvPgtsQH7A02fsWk8pe9Oo46GAhcnSJJUa2ZCWygB3Yj5v9RtM1FO83NL
oPTxvdTyW9g0k6rleM1UDUYKiTugLIpBbroy97kl8KY7Lknlk8QDqZGp4MozlJCv9cVXiQ11Macd
/bQ9tr+mAH53LOxmj5VfkP6ul5tVjvnb6FOiCo/OINR95JwTMzhhzEAUSPMS4CkbOMfPC7P5nST2
snBhx4HpbY9iHggaOnMg3+dr4zvgEChjIK784nexLztSs2e3lD0v/MM3NanSOF2UD7gsisDwTWlv
jvCdC6SSvWFs8Ei2i2VtyKx9Gz+0BLYuxMgWEIdSuysoimGxH0SYz9TpOh4sT7aDVGDse1RiQmQY
tDH0FfhdV0aI2ud75hxPz02ez192lCWUWQctiCHlPuxI+q6HAYF5jbKrrDoDFpjeQAQvE1PMGsSZ
VgmxwJBItERnQdOvxMe1UWIjpFowAbqgsUtSZAgNNcXYgSIlH+CJbJo1iFzCLPOVUa3lZXfDhBc9
oRou78V04kcIoT3wKvmEdtXD8YE1Ll06K+WMgbPB79h7E9w75kp9uwnUTqj6PlKXDpxuISyKIh+J
JMf8DKuqvCvIeMSxTn7pYRQF7jSP920DHR1nO9lNlfcnjieKkEH7iHu9i1bWJa5KxhfBh6qU7lOU
Pqd1gBDKz9AqloP0svcrN+sdx9QNlQagJSD74j6tvQ1JItm4glksF1QzjYyj3I2TRLBfShRARosk
I5MoyH3nYqpxr2jrhSk/w16134fyNDDKHPDr22b8wLQdHLCdkr5p+2RXN9zecRgALjgNpJG2ZdWg
hqAqjxs027Kq7wYLWY09vwdAt6iYtCB7T5PZEG0MVkcqmYphbE5A4aZ7NBWIGduntviNv67m4uPe
rq5dmQtLq94yq0plXklAMUb0glQ/LpikVyHIVzlmEGXc3FZq4s+LuOQTV9CnwxtR1YCOF3pRrxQS
65jNNFijmpJp9lWFzx1Jm7A7I/EJrGThJF7WLE7hBNX/bVdmTiYf+T+37YhJx+o/bR9qbBKh/TWU
jbrHW0yp0uM8q6A5k0hAJjd+aEQ+AUclXlmbzDBCCoHaFlYZCvP64Ts1abI95LxosNGroIHVEPeF
fg+aTpEp9n/HUzKyINwmtVu/8svqjjhHMmZ5fDuU+F3SsDyMK/yw+dtN1H1OYt9FcsHljsWG4FVR
ZpUKFE0i+QdN0J1pFakItimKSeJGUh3Rd/i9N+Ro4l74p/NceIzTCd5h2GjP8FGT9kRHVbYZNjEx
mezTNzxdc42M2mkRKexenJubnErcEG9hhs/yidjTJ79UpRATNudnuhkzrcIeZE60mhOHisd3EGqK
3GQoCRhzG3Yp80q8xjGbMDab5uwx4r9MOD8bcdaVl6h0NiURnN+EB8zKdZopd8I3OxDYYyesIUPC
/xDdhcwr0ELp1tC/5qsjI5arcjyA7R1Fg5msiq2AVCgEsFkaYjAcUyFCcWqJism53FM05n6DbbJ3
fgWJ2X64GVhZOj8SUcFqk7xMqcYwCAi95Nz0FZHx7eVboL1LRUE0GEM6YGAMrs4pY9jxcSzFL64Z
Rc26HjYXPSjDI7Q77hAAijOeEFvdm5PQyEtwpnvHS/rS3IolOp5TPxVnhzL7vx9hP+lKjG68igV/
kDbNfcuk3sBBAzrKGVL+FjjQdIzwv8u4G0K3yqD3GK72cBBkSyE2bH7PdaAxfApQ+nBvp3SH28Ta
QsqU0RzBmX8brWxraGu8BXveKMIVB+Ouyc4d1lrUESsnaTP/KnxALyR/UglxCOAlHuAvD41OXKvy
SG8atCJ/VuoBgM0qv9Mz34I7WXZbMKQqQghi4sRrNl2OgJfe6OMl84zQrPkc+FGIHeB6bUh/SRGh
sTHCAdAKGP8+HVF/KxgnZDYdNj5V6rUBYKqNoTARgheOjUbOgM8d8A0HUOIqMkQVUIbw8ag24rpr
FBsi0/9Ub8yB/U1d7I9dii14NpaV8T3QwBkX9zRl8XBQaNNxLOVYVFsitMOPKresOmcuwfKYH/+W
gEljbz9/3AG9IpH9IdlBIG8ZTckxMuEp6fLR8KEfD0CDxAf5zn4rJZW1+opDIXcfRwuaBP4rHzcr
ZXDFF3lwS06TmuB8vx2kCVUewh4CUPI/ZsEMF/zFO6MTH5gIyUXW7r1c6s8joLtUrZiX1bby86k0
Lv/s6zuX4IQ8Dw78x4kzep2JjSwF+7XNtLYUjlFXtXResCQOgYFzgePN5siAG2uiI2C+nbItJp+z
sloV1jUa7rzoDShhbXJsGztNQ4KgH08Jmtwqpw+qqqkc3nCOWDGB9lZiyku9KYgXRl4o59c9fzLp
qL+amWqPXjRjbqkSj2vzF2YhjcAF5a5Z4PhEuiewh0yNSU1ejzX7xF0fWlZA+A3w6IQYJ+7h4jhS
dO7iCRuue+YhvJbc7wUi19xdHk175rF5e8w2r4e8W+SNOAet0nCEUuc4UgBLp1QQ5qPaC1VLgUOu
oTyH4ix8cW7+WcURky4O958sEw52fKCdkllGStk7XuIdzPdUqQFfm5zXsflHGWktL7gfxv5TxXRu
Bh0Lq5WLSGsLQTJ1XwuhmYp4DTx4Fp1YNTwnVMG/hBqMPl8VKuJoexvYP/vrS8wzesh5Qx9CFJ62
4YKGHT0yWr1renuCk7STBfsbnc7OV5HLVEb1atPRHPYLmOVV6OkLgu5/AuUUVTS+bClof9ie2ocW
i/++G5GCr77rvuEHwUEOy+TwdsZBw2y3vrlFq/cgOHPlvTthemr/tGJsJrwrW1LKqLnabxRts8rM
lUGfB0ZPx/kJXqUBoHqI1lMBxAz1EeatCGhB6T6bMloQODA8R5wIfT17EeqJ99pQ7XRz4GLQ/HV4
ksCh2lAca4GrhWDcX6wJFwjWWGaTbu7BilXiCNGBBWoWsefrvl/p1Mf9OyKJeq9GYNov/Csup7bv
ZSuZJLQHHlzi/DNGwd4lxHENq+8VJiHNg4o5mgEa3mCZbQLRlSxE1ViZx+O6cdVx2OoZse0Qn9wE
fmaQGS14ko//J5+xXzOvIqqlI5rUT5UBkATDIwulaphHHf20tN+LbrlETFHo/W7NOs/9tAu1CZ9s
e5XT6WUOGf3P99w90yvy9m/x6ZClRZiJxBI+/ICz3yfkJWITFsQMCGdmmGWfF7YTJwUOA8a10EJl
zqRYFimd/EDVYqrBmdaMpCRO6FQUgnplEoKXHnwQj7TeWxj4Y3ZImekqblKJ5r4zP+c2v0vJpCaa
8gaehqXn2c71XQSrx4v6+nOCz7vixObo6NU1xscCt5ySnLv8w1fcfJkg+l6meNP1BmXpiHbaA/MN
KQDGYq9ZaRLHeyz/b233kImHU51DWQ+5G4yjCBzdyFJkPFi83YfNPPvsxZ2vJj+SUuJ9QFa7JgIc
jSGrYrr2+NCH8CKwyn63gUnccNniBsRG57Z8uCMpsuvO8aC5xXpBJjTWREpC8O9OPTX6wlEVb5ic
7kaYfgxVS54ljOKdO301IActjpdWPJKBkmBbDzNt/R/FycOXEay3V0SeCOJJAetv4Ky/KFd1owMa
8Fgk0z7Bh+r2S9T9sKV8uItx71Fg60+D88SJQOs5cmfY8CZQq/VRkDunCL37UoUZda83pZk+ZJcJ
3hkxDL2mug/QmH3TDo4Dp2Thsx9G2DRnvqoKbvMXmGLwu11/FLGxLT5MNd8TVGBCov9aCcDxQLmJ
zrd+cu8Lfev4LSxu5YKhCssYhJnqdpmD1ZjuQxueOJ1sqHRevHwTjEeyAKQ3MyV4Fq/fto/l2SYY
CrnA8rIIQpEUQqYWzq8GoLqxiLSixl5vh2STYXPmjMgJerWeqZf+tfQoWE3XNk+ppU1NK4fUi0QF
M7ewv4zp4ZmcetAvnAF+XzXVg05JI5grL010t07QRxtDtueIyAxPIuMbfqnWUlLTPVsgIZDr0igW
fEtSt93g/cVY3oAGku5ns2/UGVHkURYMVBbQK1I5qECKPZmAmIpf1vstwAVscLKHpIuvBAO9TXZn
caqMZQVSSETZJ3k0eyoixd8dOE2CobsWiPs1+FcSsJhXAZUJUSwrVO7/24xgYh9wk5b6RF8/QLjF
AjZJLhhCwxi4R8LRwQj+IpP7ENOMzMWYNWy8xN3N/BdTFBxPXS9dIRz/ZFPab9hgX0K1ZdFPnIYT
6bIGFFVhMzXA/H9sECADKaSqCznHL/VC2iDiCDbQjRCW46+wE2Ci37w/nwmxwgZBsYtO7ZCV+ZuU
LTQxF2Z1Bu/zVSXBLWHTFRJzZVq4lhzxmTN+hvpPy/JcU0G4ONWuGng1Tv/XdbXPxZ2DGt4tGBrg
IB0IjvMbEOGzW1EKlCJxcgaSu+KixvIykon2dfMysMzrZaWqEEKwzyBZqZePOR5Ky1uPH/YuLaVK
Py8TA3i/GM0cYDa89VvL6Lo2bUJx76tHNcwaJ71Y2HMDF1LJ2Xc+Tn36TQxNJyljNbhIFlU5FLA9
IM/Z4fsKCwEM7LujpvSSN8TyfZrG8M4KUjwU0g7M/crdsQJrejSwiKB9zem0Qg3Si9bTHGoaB23H
4pRmw/Pk7ebEYl84g4dzEsiqVJPpHcndsmJpFuHRW83/BfOBoVWMnvUXKv6PCrEb2E3+VInXCD9m
fPtKNmAcaiOAr/bBAZBjJDkvg+Fnb0tsT9JEVXSmql89mDQNUniVp8OnuiGJSzfkRjauyVZUKGkO
mVPY3i3cEIYt5YUtKAyzLL8qqBaovylDnAMnC/vEWbMwiMrjzOHY9V7ln6JRNsYE5dW/0LFN0rbp
MPZZXytg6+pQSkwNQirhITsAnhwj7cg6o6+Wg4g5rwJyWpq6my53F6oVuDcN+MlpSpT+7bLwxOYa
6U2TLF+DzlKqMON0O+ul6bgX6Jnd84eeLOxEiBMIymRYL82zRCpAq+mWp/TyTBGl/SiJg5Lj4C1r
MHqIQYPvnYj8f9SHOqpOdOJP+xRZzwE/OzR9QxY/dz5Hi4+E3zDLtTJzaRQvAx+03GZJzQAsoULq
jmG4Z32Sfxsfi3/dNezKz14tRhZnr1O2yJY6wmeTtilEOtsvet0hdN44xHBWrzEh4XVwLdDisjQN
ECCAIyHcjLOON3A0vTkh6yKcfDw3Hw1ZCu+5PXuL8JIXfe1zAhiI5Tmn4aCZeBm/+1bhwzyA/UyW
YUiKUV6sLINnRGSesyRyfCsrB9GFh8LWxv5FM87rAlVz7qk3L1cLsENeG064+q4h9QLbdZm/+T5q
NL3itJTHgHnLNG2Qogo9SyTEVgO4knr4KTSvht8VLPKs3qIty0JOp9C+5T/1s5UqEgSAfLvrXFx2
KIjQ3iDSum9pRrbOTtlsHGcdq7hvxnhXPIntWTeOMH0IHAXi8wQzgtdbZLj+hG4xtIWWecpo8yLY
TTYAIOYFkn+jF0GC057R/lSzjbtzrXOq1vtfeOIqUw2LPTLUXLJSnDqxAnoI14Ks8lLzLua82OTl
uD3Li0STzAJSletSZArpLzhAyVsgSrnlRlCwlVXyvqlj8HkWVijnz9zn+ER+ewtbp/jXj2M8qoiI
sKAxsZ63KJ7jTccdMtBvTLjEyRfXSYj9b2LD7YuGw1FP1o/QXvGb5SYPJHWW+394sa+FSlksi4aL
BAInQ7CCGxXXkBcQRnGs3BcFITtzRv5h40ZAbSuD6SUKPE5VJW4dSJtXEDwov7Cbm150QTAmDZdG
bq3kyoKUwJVTcTFrBmpf1CvDaR8F3uFh16v8TFUpNN2UQzrbciWriTYu7gPAFEne4omUCTZ1QOMb
kntxXMdnKLSSRAqYh/yj4RafHdrSGzve/4uifp9Pj/JlBG0DdlYc0SuIesOytZwsenupIc8rwGlK
8XEjqFbLpLjBVEI81H63qjC+7gzNda1al7IL4ozCpt5x6ji4WTfkBSRyunCb7JRQ5jn3SRRyMatZ
Z0F3PPLNkasE+5bGlglRHT4xPPbCkSOxEhZ1AEjmC6mhw97+baJHNK8hvebVzcPgJzqOaivLtVwn
R20eHsb1RRFBDXnWkODqnG0Ew2uE3F/Ha+hV3SFsBNEuZY1FqReEgANGvceOYNf47JmD6yAbvOjs
Pmk4UTnlddqcKCC/NPEqDYiIWZMVrcnprmtGf3+dEcaRAfTHa7OZRIjDhMJiFwgMtHIYoWlMkEJY
+B6OYbJd+RZlQigfUWNVV3ZyK8tCBxEXjsYgkNt9BFqJFRyJFrPoQlq9hEJWwQVfitKNH96MOz1c
JINrtnvrnz0MLjvxSnsE1Yu6aTzGYesybOIbCDAeUZOjf2M+JwvNlmovMLhFaMA5wlqpka9ngqCS
4iqOIubxTAKXyT/DzVo90tPd6NOm0+HDoi0xhekKH6hCXLLaZ59Ex3jKEGEP6B8UacBO0M1t9s7J
uasA4013HZPHRiJpx1EM0JuZjh+4oIryUgx3wM/jtPQlSZKqURMeu194FAnusLzDAbKrKTjjQEKv
sSXhARpz1EiZi6VDz/5h209pe27+iH6pzTHjCbnzTSLBwIVs0Sm1KRHyaxRmrlMH2IU6nQ3QlJKe
+r5nIs/Xr6ZewE84tSxr71FowE+t0N9leMZ26pz0Q9bls5RwWhs/KROrhXp3G86+MatMJp41bj+m
Kg2psiEAMjLcWYtFDgH+7trSd5L2g+NDlCDOcgwZ2ZoPBxrM81Ktkxnurr2sW2Eao+9zUym1sqW6
cD6YyGorF3Cg+HsYcUd6lLPR/0QPmPvrdvD3cwWc5av4w2jBSEimDvlAynzL6nV/9pvr2frOySRe
ZjqVD4D49DXQqjoEHwBX15AEFi4EdKilZEQmHlTJGZx9DJuEBOm2e1K9aYa3F3IZmmqYdb+e6BMq
xDNRA82lFQlkphq4P7i6aNp7vMJGHlxlDFUQwFyuayXS49+Gor28mHtQ4hf3074RYtGVPuc+L171
/frsKQlwRpQCHGmCa7Hm3rzRTFTQx1vYwW640rpJwH9+EEHtA1jIlMr3OPbUYiW1wyh+foBtVtEy
ZKPOdNrRg9rmMf6Po4Zu91cQHLBZMflVjxnGr8TckFzI4ZvSUqNyK+NwHB1SPHKfWbmER8fszjkh
qvzXb0elFvfJA0O6beX1zgxS3hTzQo179RQ8jfkjF3yhFAQgWSiPrEk/R9zrtVwTVHmNxVde8hkg
feIbZCoBCN0VLhcGAU8IXuTrbPqqGiYL8+jtyLmLRaFVFK2otLDvFeQ4LYEhXjRCfOFPSkkfOh26
zxwx9DHTYv5DwJKKjRvBnf3RX1EUyr4Cp+SidY5iO2A90bkZ9spf0c0bKjYKC40WPFQAudDvvUm5
W2HZKfbe16hH2eylda34wYYqOVn7oMDGXBlg1oTtjr5Ic3lLnLnkuUVM6+Am4ZQ6Mw1QyZ8WGQlG
EKC4Ogy9IJjrG4y34X61asOSSYLds3HeDJpwwbN/gD/KMF6tpIR1rJabRNfQqXa+fMsHNcG6EB1t
LPobTFWvOYfFuY9FA1A3Lmxo+aIz0ovajAq1EO/KvEPUTag2RYU3+5xfBwjBZYG+GeJqz3/WnzfG
jzbNIxu++bSFaWhBIDA+MX3mV2tDzOhuhVYBdxlHu/CAiqas5psIoOnylmPlBc76mVbHf8wb3+B+
oiHRP0fbXvK75r30dtK0/FYrp0d3Wrpqi0gO/kFcoq7cogG/z76n0u4xHuHlhk8yY3Wxzh3dxKxI
qLyUX7J/pLgrw5TiWyJZc1pPcWC92olVvBSodpGH60HZ9u4nJ9FzxuSREqhT2EBTJnYXdVRbTVcu
a0UMzcsvXnh63nTlEsyusS95FSZpdIxPdFoH8XUOUU3uzC4uqia5c/hX+tfTV0f78j48PPOEuqU3
gSrxxvZ8xy/o8lk4bNOOQ+8XO/VKNKu1P8InQbYiu4K7lDomgpK/aWQkRX6a+tWLvUqnz1rmOX4j
xkUALXIsRlEGK4aU7lL/fY446s0P6UvzGHkZa6DxlhkGRlWzkseKP1mIP4zRQA1bwiaf/cIlEPOj
z94uas/v3G2NvZJ1GtpC5WOS3rfY8rAMzx2XEKcOj5Av35ukogdM/xxqb4fywreXOJvQEdkWD8pu
CiJqMyPuYSUwuegD+e66yGwdEi9ZFjQeecGEoQLCG/QZEDVV1sptkEvf88kxfUMypVm8Bmypzu4J
0gii4dCQ3G4AvYqvaRHH7IUdmx1huD6j340IZ9Pz2kI4hFdz0DLlGHAIPU9X4u38okC7LjNJbpUx
AFT1XBatrdR2DdRH1eGIMWA4ukyQ4NFA9smtUEsQVkRSQV1D1RItl76izNmySxys1ViJUd53Grx5
fTVN+1n+TARA0XWn0Fp9SJ01Xjvrm3IsFdjqUrbyUbsrYckZBM8ou6li/kz7LRk01CavUdkOxOnl
wxkPPDAcUpihzP3w4i0o2+LRFj4rYQHNjlGXIw/XrEpvfVKm7+iiDBAz0U8EBX0aPEXpG8Q0rPBQ
tD1lAZcTx1YdsYQMI8Ydr5NnfG9/pXedP1dDVnUNcJ9Zpfk1ZVYpOPYDlCF3qSzFj8UjtBI/qr8d
U0wMOxa4HZedeWIVaa3+v34fzGcAdqtefJQ5gzB2hY3LtLz8Nm/zUnyDpKgaviyEpHhK/8QoQBDm
T6P742qw1YLrG+pUBvJeoXfdFbR7gtdRxe+7ZtSMF8o+lqnTzQBoAsAmCYolujsguPVTfIIVbQ/Y
i4UZPvjjdDPKcOoy0hGjMqAtPztKqhoaAfjFKStYeUb13SldPZC3L+w2mF9kv8phpaZOcoVvmuQc
CeFvv34+OJHn7G1KVwmPmx+1GVAK3jQCUUh+18sdXr/Cg7/6IxNQT0fU3RG44PcoA7TsYGpXITuQ
OUGflz0xUrwtQioPxXLujQej/ohncYzZ/9PZOfzt9vpTMxnAXnl19Bv6MHUIEZnrnhdhmq9o98yS
ARbGwmvyLKGa5wGz1tlORtMUu/RWO1AMlsg/EOuFmrJPrgxbS8UyPp470UnUjU8AepSYPdCjRnJs
q+/bLAPBvGQFZ5/HCLUMRa8rWCzwXMpHeRI8Iva6xlwFkJ4ZZYOoOKlei3ryCbgrtV305DHAyMX/
+lsF8R4fNZLd6qkfE8ieSVqbNq3oEkJcfkcwgf6tQu6xcSCK1u8zO6d5Mj+//3YWooSDiEByi6xe
yn7QICIYnDIUK3EKi6bSLXw0BiLURAbC1aBttIILOyXg4ltRgJnL3GkCGT1j14oAA8+4mPEMlb+A
x7c243GCWz1e6+O95eKwa410O0HObOqH6dlyZU+TPYxsQq+UMktX+x7/SmclAnr4B73HyQmBmTfl
h+xMI/VjjVt3OdrTw/vTKeeYDr5T8VNs0FRBF0dZZEAY3yeftulCyA1X9JIeey/WINK6+SsvRCEk
mr/froys6vfE1GbSPc0i4+Q6SGz5FfXZIEeKWA7baQSBeoTPixYOeSwqEq2WbyyGpMSpC0QEeVGs
TqWa2GCEttJQ7DE1RVoFETV/Mw2pSMPTtfl4y15X25g+y2I1ry61fI2OCOnVcMl1ql64l9EGMyk4
GTxKxDp/7Py0BTTwedSePJeV980/goCdOE+WfgbOQ9a4MPK3Kz+6e/08YUZciRf6k70XZn77KCS8
FY+6OOzC0+5iBknDwogAZzQBj7v64uqb1rPEBjRDPTxnWK149b3/YYf2nH9oJ0dPeXUQ9Rlmo1AQ
5hRzOlc1MPzPtYh06cv0KcxTpAfZ/87lL4trze0gmvySr7a6fMxqjAaMdwnL7wLdR6T+gtzdotd4
mU67dJAeFF+IQD8nR76vbgqZYlRuth7IosBY3oxfj4vCKKisTS1dcPfcRKwd7vO9xvT9s55bAgql
mB16p2bqXvc0hl+Sy9c3nMMrf58EBlE5kcgm6cy+r+8YXTsnsKrnPP/yGpTGxXGc1l7aZ+N5FO2C
Wwz+1aqhVZCwzsGhqap7jjjLc33ZEYvyHv4FVvupZYEGLT2RhIUulCzhfvzxbn3rJZVu7Apu2sWu
iYVYXwMY+rqPCGY3h4jkqxbeh2rMzFwJivJpAGq/b+gBj4waX872tmeslDBSsmuYpFDk148HqKB7
jQ5mY3doUy3+O/ZA9Mttf+8rbRFHhgCZ6GkUK9h9TZriYc5T21R786T2bP9UKuNwomZUHUTa1hyi
FHTdhN2BGYL6ZtqazSHA0Zo/wjNU3c36kdPaZTcGbibfhB83kSrpPwHOsUou1eDS6JOi5N3aTCcV
x+paF0cu+rvD1NCpeqrUpQPuwGSiIyORLYNbJfFspIzdg4BZXq2W5CQGIOrHaNdsti3z4hp7YzQ2
uSUpeud4T9O5HLouWcCTiTQYvFkFu70CmqMds6oWa3UNZFH6pSBjcQbXvJiroonDdvT8rpscxP7a
92lXIFyEEyCmkNk0Xh5nMUd+VkJ2s0iDqappLv/orqFAtHrfg+pzkyna67mav1qRbBDMV323q6sa
IgHOGQoOPJYpYz6g7OdQFzrpOquRzyPY2p3CrZnqKC9LE3zH1toHjhfQ0Odu265MbDdf+YOJNsZY
3u05FWfXlEG/6jOqlNgmzsS3pV+624btij8ljIhzhL0Dzhfxn90LSF5MXI4dxU1OEo23dAtEvCOy
ihpBiHkzd/iDv7quAvpg5qNJw6ZA5WVH4wp+wDCKQxL+KJgy0j9pbZBnq8/Gv3+83OmS6aJqoAPG
0BelR81vSR3/frlz951y+Vn73UxJ1cQ9h9XwPvdNaU9oqFaaKqIEeB+WMsWv6ZM6A0prceue2gWn
cALD5C9NIrUCMnhltuu9npx5jcfMlCFMoNvMvUIwXhD/HvmQUlHe3LzIMAK4tYslBWVUt00lazyc
QGniBSTLdJw4HyfeYeyf7xey1IeG6jxzwdjc8Ss7/MqFIfGsKHgax4JUoKEYqNrAwyueKFWwi5wW
ZkAh8dEWK2EmP4rFUJPaV3MHk+lC/zvoJeeiHtIceluKAvTjv1lSkK+BbpS2eJBr3LXLD6ZajEk0
psR3sefhYRfKeL3N/tqUlFEJArPmMT497LxgNiHiJAZoa6A9L9RlnzGcSP+pRJgSaWNvWARW6r6d
Px5YLTzUIbbh2piA+vDymzIW+HA+AtoGEeMfvfndlj18Jx/qx605oRmZh9iuKYm7bvNQ68qf6Bml
8DogoFRHrPB+UmRmhf9tO+N4rIYf9JutH0Bi6Ragf80J/LJpnTG6uxzvi+olSL0MGKtLOKfb8CLk
vpn7vEF+fmmGp4u2fjoapFi6FLfDBxZDRjJSyEcMzKH+N7ti3qHpIUA70MvITv/mAAiGlPkraVoi
ru30OaIvy5UGuK7FycJoKEHAWJGKKkOP06RwL8wLSWVDcZrzRIHEFLkKtpI7SLH6mcEHneGmxIMS
576vw98SmkKpFd6jNsxU7W8UQDSED45gRJCZJVsndgubnGSwmJobPQ5qA5yc73w+KPhDNvCw81Oq
SQmXQYh4yuvNs2Akt72F+ySM8p81WK2ZKi1gfJshssB0tBJFwywprhxCUtch00evohYgPUrV0eZZ
y41F7Dp/MeoEn+uyx0mzR2+DefWZbFkmog2Jmk+ZWM6zU+XQ6Sx3IawU2KO59SDFj729OkYiBcrP
UTHgaTH2oYl/YgkMw3o3IFZklp9xTEYx7WLP6ui8Xdo5yTTQ/aVblfrUAOG0KeS7HPKk7vHvSVJH
3TVkEU+c79Fpf+gpcdZHqwkGqIxLwFzDFbcwBMmEkyu9nXx3TQh50nF3AbZ9+Mb0B+RWFq1V8J6T
ps1sXeozjQ07f3ptgAGy9jR5iJ+2HJs+K2qn1f6pe5k4dlMxzoKH/h7sspxRcKPywdGoX8ciBwNS
TCDnnyCCec1sZ6M4cjqHvJVb9Imxorilumk+dREXfHTdhlFPSbU6Vg1YuJAVZih7wKwsdTc5veqT
ZoU0mjT0k+9RGa676AUleblr879PML+q1VTDYfs9TPzuk+h6RbhAUAo2B8eoZIf2Bc+bglb4jdak
jTScV/sbuALQ6ViQsjmExTw/fyEIcC6d+G5/ULutiTip40/ak9XUtUSvnF6J9uOcetlJMQENdxbU
+8GzUORSDlrb3YSMpjx/BbumUei9sHRpfRT1FAmngmWz5iT/VkNMY6t/zMZ2hlvIEEzZdyL0nUyD
qFZCoOwmR9cLCfhOlNOt49szsvjikF1Gr22PyePIMtyVPIRX5g5Q5RDR2IS9t+u28kk0HiApjdT2
hUCoWmkDE6Jn1xWvF7sXptBTRF9gllWobFHsW27nfqZVh2jGNt1CxYXsIcCXAq5kI0MrjU56tbLX
Y6yJPAgXbLkvDFj+XN5qjMtwXSDtpOM6Ha0iRclhuIhv/Kb+r5ISn5R/5Fk09mGtGLTf/c54d8Ju
+OZKTioVwxSoriuVzuwKH1nhY5DxZ59XitvsCzp32mEK/bdnUgDbnpOSu40hx0OsgCicwht1Sypy
VsJf0JsO7KCLlBESNQs8umMmtb8Rl2MCb8IgoyH9YZt3eES5tgRRLf2D9c4eO/562tDSFL5hLffp
NXy0F0+JJsPwnMzjaQgWF92BKnnXP58HZHYHO6IfZt5aVh+tGvBZsNFBGuLU1cNgHt+idGdl7gQC
eUy6c3ntfmpBZEEjye/ALesXyJ1+QyAZSRkNOsRCM8p/6RQMO/5CY+7+9mk8Po5UfX+UnmRuijpw
Xo7pMxgffsOxBkJCiIl4tGE5s80yCaXOsA2dCbzZxO8yHNimIG1i1KyTOBLlAh5wFu0zXc+QOvO9
Go3v/lz6i2R5/T0ijjZC3gywbNv3AwfTc8bYdHPOsj/01dOcGlLJGTUmhot7dVEl8J7lJAHR+ifj
cI8vJBiTbfDgHBJLbmZvHAnMMQz5MBR5d8Yi/JiGUC44ZXjUYDDNX6MkEpjphX7lNsfm+MyFdyEa
W4ig5FBzLuRhtxNQOv8DjSZ2VTlNJ5fezjghKRlxCpl8YQrTb5DRaGgXfx6ji/uc4Lpq5WyEdccO
a6NlGS/ydlt5RgbgNZ/c7Zxbf69iyMd0nmdNz61cR4qg2+OlOn3tldz7MVhpA71wUoASfe9pBSpH
z5SuTVpEjl3LTyhBkfra+WPZMn3O1pQGj5tUgdug3ciaKrJSPrOtiCkUsuwRGCzixPr8YvhQHWJa
0jo7trL5S/vSA24YVRemDMSH1Pj4j7DqlYtxHQvGLMky0MRt8M9PNCKwgUJb7+xFkGycQtXEF7uR
tWlntISNvQ+h7cdpoOZ73ehcx6F1GY+PmmMLEVC+U0TROZ+w45vZ6zXJZtw6fu7E81zv5LW0Frm/
1i8iXJzBS1hboLKnSxy3bA0jeFxFJ+A61hLOFm7oXmXp0LznwiPNHQdvbDWguwOdXsTZk5jrfh3W
zc6QA+81H6emCJeJe3Crk6Yu8a3lRPAEd5SDbynpsCLkPqvuvOwf7Eic2s/7Cxf3+3+BxF6BDeCf
db113Q/5k+n5PAdO1tFHjGhQ3UusMpQ3GtViL4/o6y1NtYbghXW4x2SjVYAzCzSYJpjzOQMUz7w4
Q5xaXvhghhXIDpz3a4BjMeOk5GBvoVxkQuuKKPgOQKmFEqWkQ+V1wmxZ6p4OQFy1WqwbvU9GhJVk
1keUd5o8aRTzCKAs4k7WMqZ6VVPkEdNGsk0sQvVCuybi4AEIwTnM3trtDBvbC5v6QKeHp/iqp8+l
tLW7mYbdFOn5T9nJRoL7NmA9sygoJs54QSHErY3pCfViUQquxKOxi3wmQm5H7/T5DNeAAtlGBHvk
KSAsokxkrBI9eySXQeTV5IDlNRv0SM9/9IyFmBXom9J1o+rmZAjc5e5uxZOQ33oHoaCY9MHLoLux
0r17qXeMa+3YNHZzVx8Uzd93PzVS4mLWZ6K7u0ADCIA08fsAQaAA3+T3Uu0w68ZTwehhSatUZbwp
VDuhFw9v+mO7LdrCQHMhCAHyEPZ2UCdcJVRszOfy1mZAnSZ6/op0+/BoXbf7db4BWhloD/+WqMx7
JnuOvurdApoJ/Gi5J2iJl6bVveFRHZm+bG7DN0aEzYL6UDxjNuqIplVR/k5KVVVdHlQqdyvwdqB0
FOmozBvfwl308UzhgWdIt+VzzYm9GhcXnJ+lplroFRZaNZeb/F0tlbVmviWbT8MSDaBR/MJbXyvb
vcIqq1Jrrq/absuLlQbO1fsW7IVQQNO6X/ZAtUBsz0UcShZVc/4NLEKm47DGFwwbVRycecI+PLV9
VhSZc4SjNnPJJRRQQ8phW1l+yySMfkAWK5UFsPnBNXJp1Y5Yh2ut4Ut/b7Vxv9dHChdMoa2JEqES
epGN+0L643W/wWBq5deO9KT2nL/5dvVfEN2ggryymZn4VXqUp+rJxyInPIqZ/GFdkOyltEkE4qHt
yL9NL1qEYUpTP9B17IzgAcdYWgAg/fxGi1v7NaL8G1qUQOzR74GQT48vXuNvvEYnDWKFHs51clHt
hQjlFYlFP5+gy/2wLucSXOBEqM9c+90jkphZqz+Amjaq2mpEtZcVyOch0YeFkt4ZZK7I5QRd3PA7
c5KcZ8yGjthyDD0C1YbRSwAVpMUXHH3xuGc5TjxCBu/zoAG6rGk58n6nvXe6RL/B3fZ9+Si66v8y
2Py2/glk76Ht+3Evh6gBuO6Vm4jhlfVeZ5V+2NuGvsrXC4JHywm55R22HT0hXZsse0kJY9BFR9Mm
LMI3M0EkQ3SUHNIUJI+p+wGkXq8gDoaYZxax/FhuKkJGv9e8aGDrDffynYbDkFcsNR2ERxlnCoDS
/jO+a1i70UINOenEtpe2TYVK2VHwIZfvwM4fxbN2JbKXsAdS8RzhfUsjz66n/BwmlipYOxWPEa7k
mMOnpcypB1p5Ci0New3jMvbAbO0hOVcK1WH/vVosQjojOrYn0lopqhltcmAF6B5fzrHBKK5+7MXX
dKDkYaPe4qcboujkpCBW70Eky9rBZt7+YO8T02wIKi7VP1HqZGQd+DmaAda1DLyX3h2OZmPj64Hm
ZL9d7ppY/tmVK+u0zGnGmzxBFAaeld8Wjpb9VoFOYKhRa1JZFhCSfsvh3szqWRPYGwgADnEnxAhW
hq8qrqfGraQtMWfMRtYKX4usHtIPqdjChvifYTMShLNHhTONa6cvhRYUn5oFUR3iZMPzby1RS5E1
8VqnviedvJ0b11Lr0DtuUtguBQkOkhp7xntcHVF7uN1J5xZU0XcWAF4Fsxc/vlOhmCqz88xd/3Qu
1IpgEW2tuEpWCKMdR+MA4iXnxu0IbGPVSRj+aD5I2hv8SmJXVPqMQTdf+SU7C2Hbc/+fvYcDZpxa
mdBZWg2shXA7jvEBT/etwvC1jqGAe9XWhBVXfPVZC9BoLPehGsO2qq+nxnQ2hvMFfb8smEyCP0u5
kcfavqb/Xv57uVwCYfqrQy2ZO2eV7JLNKNEnhiHDvV3EOuINjrOgYdoSVnD2NjKAaq+RZgGrneBx
jBoce554BI12jBvFgzTLq9IsB8KaceomEUdVAv/G/b6DXv6shD/z01GV75dprSbDmR7+ev+Aesdt
nBIY/IiHSoFLIP5wHeJIHbxaUMlYCsfUN0iRKtyUWQnx4gucsW+30dYFu9qpyuz4ayMkcuYE72jW
K6IMlrGwDwJOrYQjx5870s6FKvnxCIva2EJS5WAtvzX2anfI4aZ+GYXW831+QI71RptRD+hcm6Iw
z2m1p6xHmg3Jb4mxBMQeklSP9ji8svKTHPZ3X5Ao/89xbW3HXj7peBdSpDEUxfPWhcav3i9vDDFk
1I83brJsPxwDWwHbkVDSxRT8re9Dmue6tFtA2MYnquKdSPAbAQQODE/Cf6PxlzRRhAv5sbWm3EUO
bk2xD970ZW+mJZihrD2x4CQeiiQEzlwSDvbN5182GrpXKjdt0CqDzDS6/lERosrTMCjTKk/3jAVU
Apo/cq3PnCwCKCnTfb98f6QvZZSbCUEbn4iJhLlL6TuVj6rfc63r10z5yqToJ7c8ZV7xbE4Rh/qd
hn7JS3GuBHiy9xCdHG7vgzmSBf2HEUu5aw94C4Vz9tiaB9jHPLrQ96x+G/dA5cq+glPErnXIL413
Lfjfl08IYwYYuh+dzukAwXxwpeWPM9hHIVmP5SlxzVIoc+hyV33jh1NL6/9454AEgCl6AJWLJlBR
iChj/HXYSe+X1YQtzUOzjnZMHeJNHqhbtnWXDNn/8P2wwQ/QylA5sUth/hGW2BBoekKEAWXbi7Mw
4tssPH4kwWmJBg0Qp8bMII6JJWSlIXAk0kxuiq/p0vJgzfh8+MyfLodSBak6BDUoGbfWF0+z4aE3
pI7qJVsHD+Uwj9SAUL5JEhKO/W7C1tsklp3iFzNVj8P2aq9fotw7egqdaEl6hD5XuFviInu5jufU
kycbDwAJEErBt/1fP/M56BaOQmXtTOPaL1hEIN3ZWSifztExSXBBR2DIKrZB8PIUbP8BguGmoDSC
HwnNV21PabTJPSXvzlDBeSy6EWMLFIaBihQTNGLke2Kwy525EU1/B09PRGXSj5WVWaBM0Qe+oadK
5FkQwbx/Pba4s/Hr923l/Om1iqySZ80jWuAlnUsaAvevMVBeWARa0q8tVX+DL/vJ2gASfJ2o8XNc
r7FpetAdNLrW1W9hKHfnL0PcP5HaOvxvMUIeA5VQelQO2I2W3DUk07nNwje2pzMmV/slumf1fWfU
szW5jy64MD5Kw8KonWgLwZF9vhHlrkngr61hVA1YL/P1AU/oZj1AaJf8OkVziMWSAFFHH08rMyNP
MfOTlCtP2rXAhVgTa4JpWXYuYkRwF0vaGFpwzRF4TxNG1H9gFMplmfom1hcCN2JGi+ncmHjPpsdR
UaePTPWKHGNQZZgAAfP5U7UAfIAod816Lbv40c1jrZkR/DENWcJJrrtwIPM6Xuh6yFfYrhrbek+t
gsJAngRWPPsiZmbAF9tpUznWR7AtzbKgOn81hxKkRsxODXRcLHdFdwIF3rC3euPXsE7/lLwzl80z
l+l52GzQ4W0f60yyE+x5m3KNF5xOAoAsYDdcLfBjMllc9edCGY+Caqk4DBkDpiN50lC6quOIfaq+
tiPkG5UpQ795v+4S1YY1gghU5sYPSBMu+E4HO4bKHKkVZOWLDwEuk6WIxZwy45kfp3iIYC1Jhit0
s/nwKK5JqMgZnJNQYiEHAFxGT8zACDnp+UfnBzCjkQAQF5YyBTcy0NcVceFtKlu2+8pYuogoXi8v
9PEwavR7tXwJ9dEfWYOA8fmJEsmGYNCVgmZQ4u2qVOc7DXxUpguV0/wcAlXlNcObYzo11fpBb0L9
df9nc4kyyqaRje7h4pkRR2yW2tR7u+1O7W4JeCNh8bH0WXzQTua2kBLMCvV1ztioC5SI8EyY3WIS
ool20/bPDM22nWrahtH8w+u6IEwxs2bYTQqMcVyA5W0rbPfwiXfHeHw16Bkb0Q5ZH94itWJorVEi
TDu3yfQ3roR/U3UVfiIDStq08bR5DYrwjzWvS3QiM2tYIvUKafj5E816+B3J9sFe4m3x17Ps5WUF
conjSQ9r8Dk4ANynRP7nUEonhfuLCeYPI+EYAdHTCZF6p3BN+oDp+8UT+2m/IVhSIfd2I7jE6ekC
82JPqGpxWE3tBxHgmYD0Gewh4UPp9wg6GEbmMeFcFR4J9S1ApkEwIRWhbLFs0DSSgQptNxun3hrY
Z/WPaIPB8Oj67KQYHCOJ1JoCA82LyO2HQ0jnkgMy2Fh4NKCf+1Zy6wL2Q02UxoWuNdYQOMSXBXud
EXL1PPs2IVjpO5qbG2QlIugCXadm7Yg2Dpf5r+kKU+zdCVdc5V+uef6kTYQeVSGsOQ/k8CJsVLyF
zQue4PrHvvNRsAKVNIA0i/ZmwxxvST6xEJ4e8QP095/4V+beadi5HtFP/BqlMK3PCtyKMIscbXzo
Jghvvu8YB2FSUyuk011m8EUqLk8sE1s1sv4A/FMNTnIgSJ30V0DsFQSDcqde3si4PNNCci2acm8P
0mxmkwvSNeZLMyl10ruq0NDHqOE741IGZnQoJogP8ZykkABt4H59Lvx8RPIcJY4Fsu+9wO3FRso+
IHnDs7y3W716b2mdlzaxoKOg5cchPrDuO+Kelw2u97EoA2QYWDfAaqGhjoBuSiy3RkHk5mwhPFKK
LBGF1rV4hat1bkEpfKIRDa0wZLNthMSNLdzxS2kdQ5IVuj//xel1U5cGZvRdg84+mwo/nDvaRYni
Ok4Mu5umPkB/cvi28DeHlkTl9UwKesr2D9FMwShSollTtDCV6xbeOLUdSZyA+R3Id9KULAoidEtE
WKOxFf4a+xOvcoqCYU9rnr14S45Kn6ny4CbdLgxt65XinNCT+rML7rXYiRwKh29zVDZPDz3r+ZUE
kyYvzci5vwWomgJHQjAOFQkAwWidlGuKfhJZ4ukW2qi0ihUdpDBpj51PQY0b/v9zlTmaBJlqTm1/
7hYOtvmRuZ2Dr68pMQspXGcrGbkhIwXV1N0uXOQxZ70cKz8g4EhmSJzTKjFNdws1mLgfz7ZzAu7X
8Ni4WktmOIj+Jf5vlB8wfkqGihYZ4xU7vgKDSk56Y35Bc/m2rIp/kz+fwkwV3RZoeVpqKuQphVjr
bPn2bd9n4I7XtxIvOcCW5frxtY5EDCjFEh46y+EO3Kp/HNePZykqg5nAEVvVBSk00UspJip98gNG
TZYsAJby5xtQadt2xM6FmoO5kA0VibWGPiD5vIG+s0MYQAnsM1KZhRKKlPz3rMChs19bmmnri2by
Bn6nsSqgypZT6E1QHdCk/iwD1c1B4vY0gfYbqojeDqMFOE0+ACtRNYh7BrhmGJsoVo/NpHo6gQlY
WV+VuPPxknx4nCgZj4jKotxicdnpavcrQW68TeiFNZ1qEhg5vEgn+iH4wuNH56SUzP68U0/yrmr/
d99mTLuwflHt1cExRBFdEHK5ym5No05BdHga3+z6YILVnQD0S8Ab66eX3tOofbP15mXKp4gvtpfr
er1iHRnONgJOBHU538ye+XMszRranm8eHTNcsu0antq2Pmws9wdGuRkM8YVXZ3OSIkj4+VmuA4hD
ZPf7JNrIO8j3RcuOM+PCqwXwjF5VA7g8qa1Pp/PHeQmoS0iOKEsB1INTkNwbh4v6f8RFdxHHvHLn
9apY8IV4rOLsQr9jZRkk7EIOsU2XsTt3BgUIEGpkYRLrlHAh8nupBBoZVjPxaCB1LrdTUmmDaKzL
fDUEQFQSOseo1zREiiHYju41k6zGtpC889kOBYk+/HIItTPivtNlT7USykHiwH/RYV+VTXdvrdyZ
EruxxwnTQMegkaVCgFM9nBkG0SxeC2I5uz1CKxYyesjMUHZpSyFXaQJUrqPW1O0ltoQUA4i7tL+t
bBqaeLv7+84HWcHU/rhy3QpVUY05lEUaLqwDmSJ4ANckY9mbzaCGRPnfDEj6MYtkqTz3jAYJoXxv
tHqTPiLkvnkR7zo6fQNbG7O74UPQkm0IOwGORzlAs0rGnGBjVMpm6SEMPV9kfhNk+zNTRQKwEIs9
4rF0GpaW76OgEBk3CKHBz4nG5wC3G/F0EE2BEw/6Pdts/X0PVZgm2Hq5Q205lC5Z9EbnbgEyYvl5
i93CD457dG/DVdkAVv11k0gjTD/SVm6fS4FsVHYmxjJdSVVqO7/OeUF0y189IpQrNrGiM8PB1Qqw
uf9GqZk0HssSKGg8spm4kLKHFy9qNjoHsA9ucwV2sWNxxNnKu+YYgBg06n6iCnqOYPLkhDLKYptC
AGjH1OQ29CkDKeMXWTPYZaX+PP9FQgXVClz3P55dW3jprhQnW9x9SqXVqvCVX1w3Z6dJhTTJ/avc
wIDzSIHHOIjJB+wKBUKTdO//Eaa5j8vMLDdVz1Fy0B/AhT9jX884HfTYhgRE/PkZH5MXvXVwRYSA
XaQuoKYVJKZq6K/mO54rJ4WuZi7Y4melSlLmazQwEyH2eXSC5RDR4ILJse25MwqEGVHMOG/egQCt
MIMMo2Rg3NMPhMu7UmITUoCHNyMNFspAXSHUZ+QQgc1xg65BPDKX6OccZHyqLDCFAHHcz8WdkjTe
5JTf1Zw/oqBavUZKYiLCCfVkp64Zzu5k0kgFdKavQTWygUeSixSRoeEzZB2eQlvfiuVz805tsRVG
kLUZSa4tOi4hHjn8reg0717ZTcPwWh6/n4vEnJR20Bj+i+PAjJNppfCOj+yB0uoFIo3fIiLNjyeQ
UkKLQEC+g+xn311ZWzZqdiPDXxl7KUTPVYJHU0hgyFQ0jR7YKFDhmS0NKl6GSWm/zka+o8aAD+RX
QOOIA0OWYG+GVmDAu97ny1cQA8/iYlE6Hq7hDQpPqG55XOAk/9+qNjXjTJzFJaiaSKkvvegKazA8
DewSaZOn8QUV/9TZtaG4M1c9FON9YQICRgLCrS2vloh4UWKaUaQECFLlEcscsjj4tbh2wiP5vLsF
UYAEiIOEe3jJgQ08C1dMZ7h8Kpz5Dq4NDrGsiq+FiuNKkQ9Y03bOl8MeejnLuTE5E0qMfgMJ0UEA
gnGg0ngF8soNEab1EjFuMtxeutrSSQ0XgzDSw8c4GzZ9tdJU5cs5D+aq9uxTX8KnCwSe8pqKdP9i
763TSpsDqVYd72Sr5rJsLXEWIdulDnqTTrxBi5udCGpc8HSZYsC86nmozPyyOcXlxWg87eANVFJa
5r23/46AhnD39PCivui+fwDQoBZpmNW1iJnSgXL9WoYg91XFCrWWG/ca4/ANfZfziedxHyvfdLnL
veFEmN2R3u3dsemf1OS04e4V/U5Kw7c3vXYCOMmKSeQiOpVMPuRXp/WWdXnsbiXEPkM50+ig8uJv
SlmliR1UTBbCJFPtCQoYEQ1BCcBhSerqkqfy2/anG4IIA4Z0ozxkuXuTJ5sLiAU6AxGXUWnCxMcG
vm1UeV5W1//vfK+dlzeEo89YLR0ZBAd2oZVa5sL+sbO/KXJED7vr+ADfSckZ8MCrj1YSu1M5VlSH
aWO6d3gYF9XrYu/uXxFOFw5P0NblKmJx6BKmAxUaN3Gzz+/7romjMHZLQ+sTi4zbiEUdod1lvuKi
Tuw6frPML+L7sP27ogvmqAel7bYP9+TuEKAPByx8e6pcLfqUAqawazTEq1vdsW3U4oMcj6wICr2T
KItX+/Pw1hp9SIa8H20vQ3C/oWYIk2f81xdmvj5oWr0Eza4uX75ZVPZj2nYY6ort2LafrL0mK55V
GvBdyvAJd+L4K8XEqoAuvnRfyvkhgRYyxrmlN0QK+7CiIuTnpmhU0zzTHg0hmvNyvshxV3b6akah
a5XPIWy8ERV6gWfELRQygGf3k6mm75nkd5NPgn5uzMcW3t82jEV2X5281awO9I/N5/c4LQ4BpJAd
1wnoIS81nzyjL0CfMOxnnHZfp08GhG6xthPZ1DW1LClnW3cgEklkCLkGXrHigMXeyb9vTZuy9ofk
trCw+UHpcpkSDWXx9ejJvFH94y86QkuaaoKiQoOub2vsMku4aeAv63UqCzmowEGjgldE9ZO+vn/o
5Vt26gfEwfmn3AYuJUZ2EKw8dFWNGHfU9zXHfR5wXl0aaVZ8Ss572o39zK2K4+Xhby+pfl9YjyuI
b/tiQc2loBV1EdlCQ+eVRn2HERgisuV7O94IbSr4yMOVtB2b5T7R4uOfqihUVxuaQrgXPljDzYsc
FvkhUnqzNKye69H+7J2MQwtOMS5mWIkMO9MlpqWj1bTBiWLfuOxBFJWSN8VS4DUry+fczfFoI5tr
jPDcwyDuZb42Pac/Zhsv3uwV1W/1gJKFZs/HAuXXiAFbF48/sXzRo/BwCE1r7nrJdQGNYTvqcyqz
UVhA5plYP9od8bQnGq/fiVClWCUFS/iOS1KRj3pccfyZTQo1/29eB1/9alLUrUr0sJJsxK8GVxQo
PCkOFctr8Bl1DYt4M+0udcxPyMYBT+pxiHQfWWwaN4Kba2+SdTIukbfeurj/ZFfanRBlSawSo6E1
myf+WszZ7jCCsHmsOgfpztD+ltATvnBbb23d46v7DI/7RuyCtgUUJX8LQ7NOkxNd4saSsUCvzTUk
XBnyRmdLTo4CojnEbwBY0Es3fSIPL7BkNFUwFpLjGaKxJXLt/OIrYUc0JRq2raUqPzmwgeNNrpdu
h1XtY2j9aRrGiwCOB0HYKI4ga+Sn6Gajtkq4CylGMvuFl0nZ+CpmWCwonEiSkUbXch6upzUxauej
JDg6oSQkNDMd7VGpC8gumDxz2h3mbQaYZGWZcqHeGfdUBeFxZqy1eWfUO17k1SngrQQa/4qcII2X
TGtPzDw0pBAZOsftr6o4BUiU3YUWFeti6nE0HgKbl5bR3f82fYeeY4qoiqodaCdHth4QzIenq5Uv
rOZxxKogsiUgWUFkPzRTRXbaV5Imv/LMROQe60l8loDHh8Yh0tuwvPXm1WNHKGA45Lc0pRLN9dAQ
giQhFjaTUwone/bTfw0wO/Iu0aXjmPtvIOjh7zeAYVECqoXmHzo5wpYyKKUTOpivxTe9kWo7RdqD
TtTd/rc0C2bJkYH5czWbI98LcbInc4yE/lo8DHxN56+zHiykjYjduOKF9KxeZf+3K3YgYe4rIglN
OntpKOezh1wTbYRq1X0hXxaWNbvaNgbbt6ha8b42tnLP+aZzVo8pT/vMHhjvIYzuIEE+3WD5BUIc
gww31WpofePF37AySD15XzbvKBPUQno+e0cTrlIEpOENQdFrPSArux/cX7lEEnEt8CZ+KClfHgYq
KoPJP/iFApIJtS26mCsz26NFauPMzas2XQ9PGbf8DmwCplDhpSTwwsqkTpK1A6xtvAwe9DhGn6cJ
a6e9qF2/5G4lbJtga97zMyPf5jtm+qKgyOngz+90fcvZRBRQxasEov/oe6kdVlpmBQFUrrWJ8RQE
t803dqsXgrsVKbBEWrTjm9CAfmTVgTiWwBJe61KD+ut9dQgNVWjFTgn+a1twMwTlt149kQxCO+Bd
fi/OfOPdTzKSXXvkdaQkcHxGVOGB36oaxnib+JJV48DgviNu+AgzDt+Wb6cJjYckYT1yxsZs3Vd3
NAqRtOjgP22X6h+G5Gs1xBw+rllL4q1AarCXWKc20ZcQ5c38WLjJ2etYnNDqAKWLUnlZnY4pBPzT
/9h/4mK8zcdwJrXB+z8tPijxZbGYGignVZwcJDSREGnVQVZOZ8cMvKpkwq1FyUPOAimYNSSlyzMy
gHq2d81y/hJS8lyWzUEDtyJZBg5Md3hJp0qHFOkGUn65EDG6l4uFi5m6ymw1lVT7xeziC7x9L/ZR
oTpjnoRbEpQpNOadeMfVoBJmKdGDyC12hLduF/nD+zcA3+aDhLmgSzTQac8d6Vx81UyOw2oed9j7
OsaApfnjZ+9Wo22pTdnWkKz24AMDeyH+jB4rAXI8XZyiOVUA94ZkVJ1DeBjlXIDKE1YpHuwFTy84
hvSUiM95alDBOvhiImEHly6WCDZrsPZOBuVQaH1pPkulKXDYmCnX4Z9QH+ar/91O6qhUC0vUT0H6
LLRGZ1vuk2Z6YWCQiRW2E+7fdqLsLlc/0SajkuWkIeCQM+rLkkPbrfnyle5DQY76mH35aN8AXhaQ
vGcfEOjbkrr2hAOsYPkJtT2I49lA/zB40WL/c2p0k3dZEfXDx5oso4UvuKuE2xr65xpIgCpDIOcN
C9uSenIQOMYjn+V4DAOcITiymO6wBVvpw2i4iZcLkIiAYwvMjJ9JClvUlTCjqV0OOBBSo4+uNDlO
/JFOix+BssQP9gPu4ajt+mO9+u4t6yfgE5Chpq0Gc6edBaXhT9F5xpzXQu2u4/GFEvzU9Q7nIGrr
v2t8I/nBJTIrmiXdls5GHBiOBetS++iiT0hwBAzszjmj4yPnCsv9wfO6qhreUrf2aacBMtR/Zxwz
Ao5KIRiRshtZSbZQZbrEsMJWJDUX181fDb/6AyCR+FvoP05bjYqFqvGhOdGN/UNAgsNn+r5JGu67
vcv5kkEJPcIInBPLDkFLUkRFT18o4w/h+eZ+OmZOBaYkrBYvYmoZ+NUYT6LD1dtUclKnQbzmn82M
Gaib+mO8c2KWU3Z8/V/eIpJEZMOAYvicHloPBhh+nJBgv6ZSzT3bHoQ9jQoU6qu5OiivnImGRgul
N/LZnWOpUaBuufGWVZ2bR/aMYgnz/s1DG0hRgcu/R7RqN3R2cfCD/GzJmGnlg/aFT21SdGRr7/44
2avg75yCfDNTZA46fPNQY1STi2Y+lrMwcQFOS470D0u5Ou4YQj1GlJgBNzIvtcrROpDzg9pw7lni
zn3pJpwTLXG+cUeNRVT0jxVA/53zZrkoH2UchxOhy7SW5DqaFtrgex80gMCanoRBD1/SiyX7LIAE
ym+lZz0t+HgQhFU9M+uW45I/B53TMyjAbthPhdmh7zCDe+sznpQf5xJsz7otvQYNpznHrWa6v/en
2I+/lsxVWRPbRhGyBUa+iWgEjXxvdEnb2ViyoK8l0XoSTzLL+IC8cm3pZo4Y602O/aNAvUHc2KFJ
5QtKM7me/jMPUk5stGDchSLZZCadUNkdDXt2BN0TwBOQFeD0wtOFlHOMizZIagB5zO/bH5mDoaDN
HW/Mn/SLXsaYKELDclrP8uX0vPl+JNmFdT+knGQ7MXb8IhjoHf7AZ3hhvR34XfLQ9FPQXnihZWGd
Nv2b1Z4nmXtIdX/81mbewMy2eRbwxRHuQOb732sRjdyY021RHMD+fSYlmtQxBVcVRbV1IMHWW8T8
7qLUXanMKZMFDBjeKPkNHb3Mk+1BtpIV9EyKZqnyojuJx4wCpztKxOYEn0sH9grpCfo8JBFxj33f
NctSDlltU9wlSfBHMPpMi7UGzwkdH1Z9lh5W9EFQIn2x+m12zhR3YuLxbypFYgq6qc3SjtYAZIYP
BDvnP1IfY5b+uDerLkk/zjgTYyg4LQBqA6T3k8lHI3khMjPlnv++BSNN57wumQQchIfyHR6kAby7
r0TD5iP+dQDKq3QXNWoRvyJ7w16oOuK9+fCKStka5Bxe5zwSj/3hSDdEceFAwB34rtfQvPvwqB8d
8sZMjMvTioW5svwwUC4RmuvbwFcQc7hWenJF+kLfhHEaAb+U8ygLvy6WTlsLb4jd7U9xYOW2OOjz
Km4e3QOlxplVuf0cNwUZt+pgJJWgZSOTHJ1rUt/qg98AKTae9nNDtml1R+GYUbZ8e+Nd/xbbpDjF
qeTBrr6AMvpFMzrMcJMIxq1Ge0BcJVhsWZf/H2CSeTjZve/mYhX51JQjDkNzheMJnebRO06p+DBn
Us3MVhnAzHmH8p1Z4DmSZxCPDsv/MIjbwB1CMcyAW37fa8p2eWjTtRlFup5TX0JCC1F+q5j2H4dZ
o143sfod4Q4YP2Of4s+KsXF7WRERd5HlDprcDzJxfthrHTbU46lAILJb/K0Z2UybZvnXKeKLFSh8
sm1iBYxo8ZriczkWm0G7BUgBHBaCBvr9A+03hBH6zVnAonc+zLcgHijCmY4tSjunHKTEu1DPaUYu
kmc7nAX9Rt3b2LZMQ1o2E2emRJAhs6HxK+psQuTbnWL/UxQbW4WXAbn4R2yNx/zdwcQA+eJkmzrI
H3VY7XCe/9mqpa5Z1t9I99DFo3wAekcc8LYdQr6uIF9dcb8Tsga2DhcgCNlChh5lk1PmEk3Y715Z
cf4zJBT4G9dvkfLyungvj0j0Ibtbu8mVtzUoBEUvRwTFssPlQHpnwhurGjQICAQlutYGURGDBcd1
HpeJXbhtABD8Yx4HEQOPq/Dv/Nmv2ubpzMr7oeVrV1k5bn3SjTQ3gfqu8Pgrag63X3gW8dkdKMJC
gMqBFy60sFn4uRR6DFDI/mEc/PlpwGlzUJ2AM9aJgkptnghoQGbkvd2j5AzSZiI/oSKsPjGMUbEr
CrmDYHLXN4MeIpsr+1XOmO3y61+vggGvqtRa8kNgpnnv2TfsjQsDYgBawkrrUhlV/8xLKKoImffB
yGRIJrcD+usl2a769pUBeEPeVLWWgwqP/fFDdguy4/vRlu2ZSpoBy72Tf5ujZENsTep947giQ6io
y7XHXFh8mGccyqIl0Ssylj0aniNqbn6p4043xWZS209iDuqN0MtAhWfEAi/Fgc2xm0V1y2ndOTS7
Kkq16YAjh5+Qbbyn+BQxjGD4kydza7UaukHR8b+Sd0l75mxdaxwjuIwz0oVnSBfvw2UR+XzCvAAu
4rNXNSZUOdJpAuXwOnafLQ1KagUNbWQnlXQLT0nH3db3rMFBGlykpOqTZz5QI+N6pELKArfuWjf4
7DKxYcS2GMjZ99b4S4iTBt+JWZZ5g109AUd9j9GlrSmv9Q2gkvT9qFDvYPQEhTpVU40bcC2juuw3
ihYo5cq2yxoIibaBCmHwj46QVrhMmhyO4YG5kN+fFWLDdH1jywqRi7O0NFYxbWnCymrFAph04xNj
g0aEwzeF+JP7V9kfQTMzSEfj0k1DWOQbcd6WHyrQOxAKgtlKieaE7BXK3xjgv+SdbyVWe38b/EHi
lbWPuj8NIOzKnxCvWIVBXhbHA5gzFHeYJQCJtZcKzCNO3YrA7VStHHDt7wOcyqIVZsIWOghP8je0
QnQKyjCqoofL9/4hlk52nU8cBuWfHnlX1VtF5iaU9QYV/uE7+/mXVN0TsGPeiFvYbO8NCcMyiig5
MAnVqOOoJPM40/wDDzMIcz0eGbn7uEFVL5UDQAfwrcgYrdIQxeXhung3NCXf4oPnPmUKWbBVmDUI
gfjANktsQsIAe1padwBHeRmqjV4N8UNBIfMzYX8Juc7PUJFS0MK9y3PSOeaWqdLqh3RAPwPDqiKY
lU/LobyF/t0swaqP/FeSIjlUHECBkuV1oS7oosBvil+Ur3PpMNCAW452BDMv9HunG902jFQEDRej
wF0hNnDT/QiTgGsk3MSTqpGR7Q5+iSPh5rUiBKxU3MUyTaWhsaxt2JQv3+/Gk9F+Q89N37/4pIPT
8iqIUlRCGFcFWIrK2/A7zGDQFnqRFAzzeN0PNif9+4htJqx+31xK2mqsp+D9x6ERNwQSJrzfL/JR
7ytDumuS2NPDdphPxVpVYaGPBlc9y6dQkmsYsqz6z2JaBqy6VDEpcFXeqMeZiNaguy61Eta15Q8n
Lpb5oVe6jv4fPmHzKDX/uSreIZGLn3OiY5V5l+jT2YJs2Tp9SYiU2jWMlSp7E7KOl9+ORPPkIEFo
dqLi6SO2/RBhStPQYDrh4waPxuxd+E6+AYiXZwUoekqNrzIcONX+kmPGGyTVMyxf4PwuuePQIC2C
y4DxZQRt1t1hTXQjNwDfh+L/eL/Tv4wzYeuqksVwcqp63XiN5iyqHrNg11MjTV7VQD9BfGsNDRi6
OOpyFohmmlYZexL78I96yydGURxHuRmYXU7LHkeaAbFaBCXKIczjiZY00e0I3EdVkVFF7WtsGtmP
cdrDWo3XzMjBvccnEpAQBREamry23HPHIHLZxaDHR2ph+uRkdkwA0CaugRsm7N0I7/kf8ne/ZSIJ
gaYZmMc9eG0FtQVf9dsTzjGF2yQ3cQcTImOJEyZoU7j/aiUOaYJpkDyY3IKSRO93nUVZwUJWVO2n
yZeRpETxiaPtoQP2UNWTE8DHyz0HYdwZOYqmXug9ZaAB+N3R/69iVYmT8iOaRQNTbyZ4X5wEODfK
/L9n052iYDFRWXSSDGUJv1lWxT1pJFH49MBRSWkBL7EJbOhb1dL6sRFqfFdtc8wzhWHs42yHeHWm
80K+6QGCVrH85y8BOhXRmgYBgjkln0NzaYvmG/61UBsTO2Km++ChpzbV7naVXt1IXyLM6ihkHANT
EZ9EmPgEZwNLlB7yl51/JL0JGVxG4FV2otTcQXGzVu7h7pwZ09+uchatmol6vw3a+hLzui9ZKLdN
S14HEcOzHpGoM82wz649jecl29UZowY1praX1mgpMt3Z4fHc4IocOzO4gU5bWwaVHw4VXFcYh8YI
fRD6BI3j4P54bA4HUuXvPP/modqzlchxZD3gkm//ww3RIhTZ58sowJPSUJVIlFM4KWEKeOaU9GAI
H3NFcXeE6gTsIUBhjkdKMYpn6Qu5LNiWZBYnzy/Kp5203O6n0JWdOTYCoQ1zOGYuN9LL2uMYWtA0
U5nuHOO7N67P8acSIVbKU502gg/Otxr94KYldvvOP42jT2hFCj1aYru9BcIhnpHubwDEgBQXNFQB
OFmogBnWEVpCyyBmOn+GQRM1tVgL0DZOmHEqErUoPWuLF3dEc3x1eZECjXui0pNG9KMJ+m/tH66e
LjXczWY9xeV0USkas+6Tw/Z8U27IEgUeTEF4Rp8BrdSADpqnCtjGNnRBOZy+LCzvoVghRvGD2UAv
F/DI++kwmT0O3g1fA2Cw8OUtnlpAVf+jd7zNR3rbq+oPPm42MhQF2fkbdVIOQ0FBxjSI40ltHX9L
WRbNSqPDnFVQSssWLpEeeG8vzzQzAB9LWaaha8J2vTnVkKuTpXiwnO7cYutJmCd4rccPg6zE5Dot
BEHVYfvnaTt2hIuON2D5S5YMTNL5vTXasirLqdCQxgkOqPxde9gbbNrQwGd/v6bdOla67OBqbzaq
U3igPNp7n4I+vablSn6zlaKqjcRhnnCdnCL+mVogLPktbvsteArEDWGthmsS04rEaFdP6Vu1eeeZ
ySutlV4AWtQiLN3ow/2qpwf2dGCS6JMIBKpOYy99OF9eOw1cvt6/49kP7iD/2y68w3qhn44zPwOF
2X+0iDNh3KtDkIJekVMRRpD5fVtTJbaqGaIMxQYmSli8XfVih2EFixhBtNjBezdcxbwpwvKCfDji
us/tDs/Nh6vNbfOdMFEFVk+56IJZAnangc8Ud1z+8iGumuIte6T5BxtRiSHi98+X6te7xNrgXNdG
MKgdQWKyuIFDvCm/1mORjoKD/f+XjVquoEtgLiapQV4xGEUxqH1bq+nwiPOXcxQI559Y0cpCILfs
bm2YFJjKIIluL8JB2ytDWUDqvbjDJRpl4U44RfaBtSqOifix9D7KO4uVyDFnKFh8C0ygrrYyuy+D
jQ/PYHH1m1YNyhpFjQz8HIHuG2KxQOZiOJcRkY9/SrC4EQKVxvjGipzPE5f3u0D28FE2rKLDEaK9
fZ3QVDyxPv/RjmeA0WlIcMlea09N3PhpFcOdTo7YRcuIOgdDffmEcVyY8gjEOFBGKRU9R5gYGAWZ
1+rHrliM/g0uwP6lk57etQ69TnO5laE4/Xrtbf9ZfPvwQH2ciCKpHcoU1JikxNlssJ4zGZyryLzk
DNrCQ56daIKpxFBqVGTgaLnaqj+fhe6Hnc+FMmOKkOhnvFGEUQyxnplXH3/RBYgs6ooTfnXs6bGQ
G5NiWRNn/fJsz7WYDR2EIX0k5wOrjp1b4CLnRp0GFRyppjhDvLeC0ogUCen6ZkYeamgTRC/y8iof
enVQJGmdzaFUhlxQhzxeDPbx7ZBVx2aLcyP9zD/oKpi+EJG9UyOmr4IBQBCzvYHou9N06uxSyUcx
eymhMxYUzP9aEL5PQkAv0AyTvzLcBzGkvC7/VHX6HjrS6d+wtaAUeribP5cHDqA25HBywK3H8m51
cv0zkJLNRjgrssIJJA9PmO06dsrzTaZeOTx+1bc5lo+tAx2KE153fWzlhvEQNGGvWHDbdu+vfmhj
80yVpnYV54DzV0JWk7nbnO2h6fFRc2S5u23KFvIsA0n5XINgQPrkpdlAJ9x1WWDTsACZ7UwWClgn
UUQelbG/0UykEZS9ngW1VYeWXLIdZQ9e3iSEclmzb1oUSMJj/xKnWCcffog2XhXSmSLqmd2w5tnB
BFGUmETBYb+U0Le+qDao5GS0LUjjBbqxo0C1K+B6OA/rK6AQe5u8JaILkhO5pdZd2+bMQUudjyEj
mE22/lm3eG/FOCJPvskB3oSXcSCBrTA5tUbArGiiSNRP1PxENp5qqXzT04+iXbuIsBiJGA5hhtYx
MwZrhTXMb7VfX25yk5DT7dckcemF+cjUD6SAItCqlDpuJn6N2IS/caPpcB6GmM3YW230Hxa8KIAz
pELbsRbXG+wDpPdeZWsoqPpQD4Ppd4HAfqu3jly+grdeOqsv/rxQYaO1B4PfzBb3tIGr60xwh5rV
eNVMuqbMuT1JqIKZTLKUV+LNvTSqwOe1lRFOI/IAiZ6hAJyOCskQKlFbqLMUtO2mEC/ZWwNpY21k
kvaS064dNTSNcbcOwmZpywYHvX53e6isi6seRyJZVZhaK9RSferwEY7HUFChd2tK/UzJGOexrT4i
z5iiKdaQ5by0wBuMCBPkMIJ/Kpn5Larioka7hH96yNUt8afBNnU2VwjrEcu1LYng4UCH9uN/ma1Y
fmBusHz92UZ55Z4erP4Udj6vkUFdVa4BdxQbSVIN7Wufxfe4ei9CE+WLb53IH3oNIq3rZmsilC1o
zxOnzdFG7FDghzO7s+qSFJd52o68dKS/9+t0Ij3NVhHXBaTRXs4jfVouc4KdX8tNDy8A4CigojvF
OFm0laL51gT90B0UCC5zld+Kp66K6kXAloXyOuIijEYVr4nXF6/3nQJHYb3JZmOEwX4BafNWIjt0
1b+y1CzT+WStzVQOn2cdiU1aK5JUsZNVmyz99RWrTEESdKRMocpp5sZJ8cnBsJSFeAmo0SuSHg0e
aAmsK6eh9ruywRCXdYN1YcWZvQYO+MfFcVDuqkPOfC+7WC31AyeiuJjM67zhbZcC4urYZiYrfqAP
DR19u78NwRqiSUR2N5uL1W660IKG2SVE9oiBJ8Dy5ZNYbbDAOIoW6TOP6zgTidH1df98i9P84Fa8
CHP/UVNf68dqygxFpokupDbXCQr+iw+yQDz0znq1S6GJ0GYA326keP7uFuF33SNPtNcQzZ0UMFLt
R5EG8kTRxbCWq0ztoP5NEX0OSZCHZO5sRpHIYoEAL47a6H1sJeMYls/dQaVRKRJ9swCguHWSzNiF
cmmwVo6cdts0C9hYvIjQtiqfxrcula7B2ib8ETAc/EY+iWxtlVw2CbsIqxlrnqKVK/9uO8NXCsBX
s3kwxaArzNzUHBC/nNcwfpi3u79cBApMgU5P927KDosClzmimpSHYtpMvmk1gcq9FMMsbHHUq0sB
EwCHD+RcHGqL5pi4+I3rdfTTPvzX/K19QlDaC10ZGEQAmzPPRT6GxIzZK9fN5VJlJtDn+KfVnr5k
yaBECrpZjNqCOZy5Go7WGV8eR8yofxcuqWiWU7eI0zXpcM0cj1PrLk8cXErSyJS17JOY14lpEKjj
bCZWD9paffUAts+T2wIL+6RcBwTUanyeo2Ul1HPWlrgu4pcg/0Z3xsEhzozTTaPAsEO/aA9EUyPg
EWUyeaXAOagzSJ8nDApSQi5TTH8qHCoFiPOKBluTUFkXl19XPxUZJDwFXu2YoixnMd5U06dgp/8m
bl6EPGMnXB990lbUGSQ8SKSJnCOAIDpE3UIOrorHcGNwsUt5XGTGQE4t52sbnzcqEg6IMhA8HgG+
jk/e4EC+4o6CJsTOvUmmuIc9gtABFHCw5cyRITJnlDXE0bRw5TF88Wi6rmTkJCkHHqe8eu3Mf7Mu
TUrnPkzBzqX+OKFi+83eiyA6tDJlO1KSB/B/WnH+XZ+j7kjI1+Xwt6ssOlSDFxc5D4pRd8Q9ySD7
lk9un6CNTaxUZ67sIoVGKBAPGZM0R8J59we1GJyjoxKOeCue/XL5N3Yw3BZseQ4pxJy6gTQsnPhx
M8Ms41/5bm7+Q577vD+CpBFs0qspqPzt6bqHonYbb2s21x3rfOT3Mv5NVZDDRmeNvfHdKAahCK3x
GbAq5YEb7BWVj+QiY1LjaLO/Cj3biwqv6HnsgbCTx6Uvcou5g87M1uJuj1OXN46Lbp1QHTvhwJQG
nxO36tkR7uh2j1xhrcXJDOpZQXonIAFML3GcW4e5VLanuHcP54A5fXCDncUcCx1pB51trli5++Cv
I60ozhRr2ryVYkbKhSGnjLnhmG1+3Ca3M1WWIJhuNMjMaCkIyje5MuPbCwTyexlUG5qzTCdWfpA9
uDqYOe2mKLHCTwIwcbV+kskmM0xYtvMbtQs2PqFOA+GONkLSJTWI6nA42z9ZSh3c4Z/aD72Q+gOJ
Lp5l0VbBYeav/BSxiKA+TpOLyxCHiO0/60voG4Rgybo5p9JTlOYnuui0KLP6oj51GtNXajvIg8x3
Wnst/qA6lGebKzUZWwz5t1QiGnz9V3l2bRq8Xxh1NSy5ndrOuB0lDJV1AoFigVUhRJWMEUQJxYNT
GkEzv/Fy1Y7I6QwYCo0EcxkRPVcZAsoAiPwxtURMDpJwIdZpazQTXmCbm0pW7Ukp8OczxeXs6F5P
gduQbKoWr4Jd1U+X7dOB2cYEy8Lpvr0wZ94iFs9OTos774aZf8LvAj5Cbp6tXmklSiSHfDvziMlK
RqKRPgVhtHEU8OCxhglzS2XVy96eWw1A700U5LWrbQqLQhWhQ86dmPv20w/3yqjQ/hsE6fMHHM7F
pC0nC++ex8Q9HUW42XUnzD2avmbbfXMsO/jfmMGH07nj3QIIoPBly8EPEBLJ5wqcFGNw917N2wzu
1euL/mSLKuMKAqHdtrhpfmWxqrAJANRqbNOoU7viQ18h1R0RQbqrGvKjhetTLJMGWuPLpXKvbhYM
1Oi7F7HKnbTzqbGn+ye0bEWSG005GIRIWfMM6tVJWDcnzpkOLjI/jRwcDPWqvTkILKmPkHv0tAr4
WLVN70NOLGLVTQEU+3uDjweI4OWnXAyz2iN/9rnm6nAcpul5y7h7wuWh6dT0DvqmTqfRX31aLzng
VLVLkZrxutUl4BPHxMUeJI1d/j+l3s2FdLoOHwzo3aM4oNshmvcZAeylvAuN5yYUYjdYZt8j+JeX
BJZc3ASBBYZEya2zl3M0B3bzNIr13dUaWD0OxQW+9lRobpuuUlyNl+QQy2Pk2KGciF+nlxKg6Oxn
tcVOnfX2Buu6NQfLn8Zebpc4fjgkmHByw+DEURQ84jvTI/Dn4cB8gn7qcKdiecw7js9RRB8l0yLB
0pHxH3Jy2nxbi7ne/0uUsso9iYeWN+7AUzutRh27AmHpHO4jj4wG1ERzQd0+oVcmNfRYMbEXZAoX
lUM2uaPfZFV5R1jwaMI2agEuQ2BL4akTJQgbs3cjfvHFr9s7n7ZkmyZY2bb1cLMjORrWOf89sYlV
T7vS/8zLYHVlnG7WDWjuwXrQCntxZhEPfpkj8HBgdXKeMR9LdjceLQcgCb2AHMsAgZKpJNPycDVc
N2T6PnV+Sf76aknYzQm0bKiFrkttrkYK72Chwnw7jtSTxCGEWRKHVpWuHIFqZoLxPCrlDsr/+bc0
XkEUZYyWIuGfc3GipHuqecQR37LeDygSGIGen3sunY8r4DFShisVsWK3jKLnOFuubZkbUdqDIemz
jg5t076RpQOQV12AhsoKO1w9t4vSm2NP5wB1ZFeVu0Kc1/88Bb0yXovsSTLmCvttzFb+XZ1tnT9V
NUH790VeTp41Ij3yY/uOfLl2A9mMVb3YsZlCFYyihU4p+q4AHg9IXkH7yPzRVyuEYZjQIr2lhhiv
590kN4TQg3JUakXRPS8WXbjLxTj+fc18Gru24mhOufZ2mXGAeJw64fWHKQhvKB7Pf2XudnjhbHYI
DZgyk+ZfccPZ3tQvLCMgQHaMjxMvl9baAPWS+MAdcGsmE60clX3QDQQEOTF79rwFL/fmWvwXhqu4
qcmAmCA51AJAs7rfTfdgXDSeAKMmuT1wlTM+QQxq0cFRzzxKLU2JNIjHhEoD55KmIiKUFSzQHbBV
2eaa1ZaJZWIkwrhnyuKQIQmrDuWvouuW3kwkUZ+3u6fbfELkyU4VvBy7AwMfIsGo4YOJJp5vx9DD
HJx0bkCtlOVzK4VVH51WBbIidtpMqABWeUpF6vVshcXgxzRi9xvFb4TWy1T41jEcwRuGmXfLBy6K
ifwjABdPGZA5XT1fqtmvjlKRxSA5YdstyRJrwbEgs579FkXbVUInPQDY0BiznJOBSweC9QTriO84
/E8k6PWjQVre7A+7mRqIZD36LSo6jgKxSfnd4NpFtW0+hkBuQhhuHaPuAoi1VCQ2FRTWN2BQXt5U
D50P9qjaZmdEdFks0YkNNfnnfoF0yT2KNH9E6s+UTZwnnZpi8iNXVEU5hO/WYS6dthmoA/Hkuotv
Yqk1EVan2z5mX9ayW8TdA3UNPll5OX9QrEx0WqBuITg9yWrg2pmvShbmBknTj5aixEZrenTHwL42
a9TqVH/FujqJszyarkoptPIHNXfjiwPAwGLKoPx+LGD2nHsdTV8Hy4N1ljvSNwRC9yyO2iE2XYqH
HsmKrH8HC1dgGbOPtgiUzh1vLVPVP+xSYFs6hdOrlJw++5PIXVgRQpc7/1Ok0KctiDpx//dgbYNS
nWlLAIWMQkuDZtKi0WDutzppJTKBLKvi5ohuDgd9IufVyXP2b0IqH2hQRvB+oUtBpPBENVuMDeJq
H92cJ/KHDGNW/do3ekzOXxAqpr5EMKp2Z4BH62tfz3pB4Cel+Gg82n8U5BFTaMz+CGeQUytvqlzk
lRQuRjxuaG3acIK/OS018yi2rfj8YbJ06pZK25y+b10NohIpLexvfufFw+0NHvBYiHAfscPKlx83
MIEeUPLY2vd26OnG3EO9hyNLUtD2+WZGfXk97Ngc+K0C4NjucPKvnstERTZ/yp16LxnYs/1qPkkp
/A4Chi4XXw3v+PbqqKS7d+n1s+lPGB0Yob02v5dsHhVgYzEManSigVlbZnkXewl0z/llYBBIBhuF
HRBVRTdi/UhsxYonw0/xFnfFBNpDfqBry5EIMt7FdADtGa9ibCOXFNto3UDYXEeb2E/JjkTxCaC/
dk+EKwsnpAFY4BGXAOW70Jht6vRLd/xKz9UhbhykZzjW962ZX2wKmZjSXni97wwZtD/jlUakc64j
CD2mtzO5B2HXIjS20AxSR5sPJSExwHp8niIjQesklJo1YtxLP75pkErB76kuKsS+m77216nlzFM+
TN3IqvTH6baZL5OMLkWhM9jVESqwIQ051Au4NsLOjw148Y0niVj1pNRLtU+GllQO2icbCMutHS7F
1w5MQPMYqQo7MzWENUcT+DEpXsatdUV3JCRV25N6Jm++SikA5/F6QXHvYdEmdbT40nnJgWHPXXvq
Ze2bRo9CWPkswkwh9EqVB2h1p2JzrEMMnN5t30eg4Qap1FN/+n+Dk/3761jty42elQyr7YZFTyjL
1o4eRHutUV3bp9cyeq5iMw/IKZc/hJbvJiBZcuVzeZfLBRALgRNtdJq6sti972yHtXVrBS902X5D
QgFrVxbqIXAOWXeIwdcrQYasrKf/PshBDlvz5slVqeXLMxhAuqkTofTfK/QqjtRG3dA3KDyAFVrC
3A0X5gmSBeGC0wa+H7/RHuK63tXq+NJQFCGHPlxjUbl4Ar9ZViuKg2wFyz2orjIbecm2yj25dfGw
6dYw/S6dO8kiygvb9yuVCtT2ZstkOcNx4+h6T8AjSCUDgXa+EyhtBhnwLZDCJVCkyZkJrr/fVw09
1aiuEqZ7XuMjAbtZoSzvAKpLZXkRq0s6h3xSIKX0zbPU4LILOpGePqUomQPUGcphCzBmH/uP0vb9
BTCBxeG7l+OfDIIvkhQCw/fX/LVLsY2ZjVplJSdKVADEgXpaINwdTYOxuxAFgAy+Pe8zApvFctHE
9h+5DqeAYZt5qU1C1cqwhrLsLjev72ZtmvdPQq/DPSAeFYOiXilZN+lo/hHeJRI4BrsXlS5R0rPF
SHE6KRXBu1hlVFr4BmDwEyEJqMoUjF/AJefGf5RYH5O/rEfagUHhKPfBT8V1icpbcAvVG3lJPYtN
uySMUTa73/dSZjcQgC45JCzSL4Q/V/GrnIbop1yuhwWxs2Fu6EeBo6lMWrMHY2KE6O0Pak1t4dEz
OqBrQT4LY8nTWNoj1LKyzK+rJwY+Zny07sAtXVHXhOIYqILSeZAptLSOlWuZGwtqBxo/iISNDj3u
vHgVeVxen8j6UZ8bBFl71ZKSz71epEfJxPWbIe18EUP+yLYiLNuWuefBTuO1flb7SOy7AX1fvHS6
4p73qnJY9Mzgok4awplpKHySv2zNaRHaROY4lRasPlEaGyTfhcoQiMb58N1hJLakZ1uJrmh87K07
huUCIEB/wwE5g7m/+wENo+9t60bTIN55yGtkPJCcUrtj9+Vsska8c6KJZtf1NFP0r6OUMkHAAodq
LB4YReYGQ/955JNwlFCWYRHcglktUe+I++uV2b6xQnTHrYTPA4k4Mz/GXu+UARRPmV3C5BCyxlma
6GuD/CK7pDrlr44PP5/joCq9RIKgsjRZVX/z9elX2Dsgd73dDZEcFG4ZR9HdydPsdODQ52Y7VM7y
uFSpSTrri/YiOKbNzHJBp6yS1pkQorHxo01yIG04fN46xux76J4uKt5IKhgxy2e6jqHzuEgN1MfK
XzQg1Zdsqz6+cj8cxuLDKRoO1GPosQTpjSIAKNv+4Pw/g7K63Pp1Aj6IZdmJu9c7xt7yzXCGEWhx
tN5aTvON9bh0q+qO3TbHRpTUGWobuDJJPxcTHpWlmqK42K0j9dPO/nA1eK+shQAWMhrXtJZ5QtHs
WHlDJW2U0TVljFfhwRiCs3O59F8NOdz8BX0Vdiy2Rc4SU/AUOt00RjkbFJBq66mjbItrkdT9DH5Z
mku4aHGDaonM3cMdffoUZbkcfcjxurcjns5/8sRbDhuhXELMciuODPYszUTset5hK+ZxrQqz/Ce2
BkxAITEkDvU+sJczXd4OWauHaaRHSAoeCXxcwCaVwdBLCjx6RLdDtnslbjsXcJNS5cDm6Hu19yzo
8Rhahed4HOwWnxHVhhCM6zvwOay5vmFSwDlf4oIer8XD/eocYbGfWofu/Pb0XW2xZ3jwdXwlYFX1
DkJyuIA4JyM2OWvAnlUGuWgpuzW6AX7Unwhn0hUlf0PcKv11rcGlR7DNypZHvP8sZmfBpBXae2Lv
LI3kHR4hoRtRzo3s9+EdNDlXnCjjC/56eJKKH69X8PNSgcaB2w4mpoLfbZGS9sAZUHanRQP4cVaw
mTIu8+kV0UEzH1n2wfeNs0vm80jvMJNiIzrEyIhxughACPcwIvNFFyM1NGc0nlvCYyeF0ECZLNfm
0O5r51J2eZswWiM9VMsoZ14X/kqUjMf93w0k30xWMIxc7ESgV4NT9r2cgsJN6/0fzcY4vrvTAk1Y
IZRunYH8VCPA0rPGsPZdeB+TWURc4DDS6kp4Cexg07seRaCclFGXSDde23jrZEZUGDouVRZ7u7D0
f+lZhQjGbQdZI8Phd5HdZRIyXpU4w56RKz14qlyO8IiiTlelKOfwOEgqF0vPY40nOpSuoYYcdqRJ
mxlGQZyufMOqTJOIdJVW/xUhtONsXSDznAPhvw74nq7matj/84uNE3ETBZ4SMQ/xDJ704DVku4Dy
wq/8hoL/+knrTMiuyAyVMixjbiYVStnCpaVzVGnWUj7nTfBKWBZnTfo2u8YhAPN4IxyUK0ObkQG2
6O/ADfiEAk7WGNHs66Ws+7kaijBT6Ue9NSiuc4Ac2XKANt4ZJ6gyo4RIGoS5GN9z1gMbDO5RDFAU
IA76qApilBgoAShxx68aNnDH9JxDY4RUwbhjRkOh4ZGTfc8o2Za+m0ZNTvpkMNX4uWUQY62YizFq
8/SSgTnRrLaecKxUBAW14SOxXbklGxPcAc/AG6/H3+UyarImk3Jv/DNVvuoXlG1IJ1auYqAtDpoT
fFtjOOAgUhq6RUABewV3euKFn3xtEHHi3mU/QCxN1LlmptVKbPhA50e1U2tXW2J3rif4fRNemkGQ
+KZhBoNSW015d+msiih74nuj1ZAQO8IWddeccSb/wydOyUwsbB+aTt4CUn0jEtPIpS6Ua5YW8vdg
luiftYzwrd7tqBzvBB2mSSKMl6U9lhJKMWVGrbTlvj60jkunLbmjty2edrgNLRWGx5Im5VzNMBCZ
3vP7jtowWhlvhKK/PylgLPXhkR9Rvw18+aHDiY98gmvHLe0+hH0UbfDvi5m8OKTS/aJyxz2PXgan
kKZG6kzAnTrKv78HUV8UJVOATsqVG86HHFAX/bTIoW/TFhVXvRQ3HJYxUfVr+sHcABD/LQsLLVS7
iA0O1FL6am+sv/zjXvgtXdDvm/HAw4/LCdZJdpKP2IY05DFjxraH3t8tsG3GR/lWO5ImbwcLx5qx
Egr3hkT2lY75XUaKHO9Zc/jq9RrpWI5VGiR9AqLVIUK8kwqxYYGLU1ZgabyA4Km/LKkv3u1o05e+
2sz8WgfqBsGgyXaKGWgQ63k+xPVthf8hAsRJydZvXr5Xh3HsZwxRWnTGN+PA769HPZFTbfPOQLZ4
xmPRZh4UxkxjQvxbSxCn0Mcg5iQryf7EIu3YopBhXHWkZlCLI5JL8CYvuBuHvLg/GX66XpTLcDas
1jCYdgjeRUgSPxymSvjlOD53gGXJxEmRO0NEGsOq7zyf4dZYpPLrG9UvmDHMacszwh3zuJkAr/HD
vR8aGkKyAHl49r2/eiZfsMHLwFYGKUOtDQv2f86xSWerNa67nx+xAjdRfi52TSlMAkKmttibUqRr
rFzGxjJzzrNmzm1bs9Bnpg8NBCW8/NS5qZTzETpKpqmzCcliPgRbLS2YeVDrZAqx8UvAfKBCYkTR
HKWS2idMqpZYWSdfcBn6Er71rnUPFSgdOeeGEBblI24Z3lPpC1vGuA1Ta4DJlHF9N+8DNFQaB5yT
qnDN8pcEOxxovCOwdZ5eB476GRcwU7+FW4G9JdWmEm/qA83iI6m9HsYE4SmDmbGKMU3h4KfJ2x8L
kWa01sLtOrf78yVErjf3Ic3Qj1nMxvQUjL1M2MrXnruUTcnmQ16FMEb/p9e5Rj/pRs+yLAwvGJuM
7waOk1Pj6xB8TsdtNIOwxOSOhOeYL2Sh4Npup1GtzeKXWKn3at7NQtDJ6/vvv+3CpX3rpArZdllz
SSRAf1ZD/iBTfA4kC7hIjVDkkzLDTNUHjjm4GXkSgqj0o3zt7ozaJazSDES40fXOYwlSePpC1DvL
JAS5vcWa9PFf4+Tw5dsIvwpaM90sPdR+gB3JBSQkj8/kWy2Qcp1eaK8L1gdaq1m1Vy428doxN+cn
FPUFbdhBrq9H87lGG6xMPFEb4CNDelfj6yja2abbvCEmtAJcFO7AE3qcifK9ToId7iTh9iQR2+Dx
SXN+kpYpWdUQpCu+Gm5pGKT497ZOgBbEvlGCnHQ/sgCuw0GsCdRRR41zk7MWD1+lhgwKnCIoY/Ah
tJ0OcZ0731aMbO4Jo9Tpe3POIO/MYwOW6a7rDRCNdfx8BEivP7aSwK1a/I+XZr9BMDHdj9qjYxFE
k/0/cdviMM03rXNqfdJe0Cq6ikuEmL8TZeTYbsx7JyWEPbSVxqL4I1MhF+I9L2/DAI0pfruaI0TW
RxT4DoydvZF1ufw6x4DJLproYgO6fWaPEUUl/zb7vyKAavISgFD338sx74pRod343NV2BNaWkTgh
2nD/gKwQCPOJ4qkjLcvS3tElW/K9nSHXIf6yz/mcGBHvw1QXcEA3Cm7gC2x7owz7fd1agRT0WKQ2
umMT8Yj8otcTdsWmBIpZfVf//V+2WWSaB5CTPbKHiyBsBcn/za1V0qlVHk65A+e80Q+0PO4roz75
7j3yOUqdch0zH0mBM/2Duwos3yTaeiJLKw7wJT7S46le86AFB6bajNpfURT4xgMuDc+kRPzoNZEL
DIUnKmqNW9fBvzgDLMtXq13v22ZqFYQhVv4stkKcmpdDMKmiyF5LmQMFgJX0EiVp4eGI8TSEbJrF
X5yvvn/BLm+ztX1CVEAPr0UBD9vMKWDfedlA6fQ7MCFfoEMdgKnwJX6ngKNbAKLjFoZJK/5frIYY
v+nYoXWUqPLBTAAckQHqb3jaDtLYVSCC7lZpX13Yf2H9/8t731NC99Z84u1sF0LtjMuqj6paNWRs
Ggzy5G3Tknvs/WCqUUYFiTawEOXyNwdki1FYAPuXf2kBvXO+PRVErtIAd4XzrtR9xj9a6o3UowB0
lARh8nXYmTieoFWeFIDTFS8Ih1orz+hBp5FJL4z+c88jsudMdmDqf49pVMSA/uZpd0FWI4zgxTM9
VIiSqxUCZNtaiLKP5P4h8mLgmABLH6syIljKfkIzpRLlGuKM+qCYOhZ1H2xCN73PvBXs15faTy+r
IIE+7bY9f47KGF0d0PahmAeuUyGIrenezerFiOPujrKFJzD6qJmU1HhKIfI+0g5WlGE54i5Hpc8r
LNRBcYPp/4eculETk2OMvYXGblmMvlA1AeEnw9HRUG/vDZP+YtfWmuQ1F9VrgEaN9TvLGi940B6n
eIffT2lWNGv4TijcJrdIW676ZEAPNFNOXLkyyPBvrbSQ0aVpjnSyZ77Kl3O9WPz8KnGRiQxetRYA
XsAbUc43Uxq54BQK3GRhlmTKIYfvBoOt5rdPSAzBPl+DQAyd1e/M/+okG43jqWeRs04wUYx/nsMK
tP1v9QSMs+DxdAsY815klEXyKYtWCRWhrkHZKdcnVlpy+1yvNNV/GNAB9PCGAPXhIKfH43Ch88Vg
PHfLlzJruehspG3aKkFSVjU6rgB0i19kdJCrDKCR2O/2YvlTQR6aUFx1Z1Eqs2WFp2AG9UCvVXTR
0/ypAcHeJRwbZhFIU9PEsrHJppdki3Hl7pjoPoTX9/8T8JHD6m/IhpDO3Ee8sqAJW3TyhDDYq4K2
Q3esDt+3Ct7/0ImUsB4bg3yzEEsnvZBZFeFlsM2COAQohH+T6Kw8eO/rUbA2d96UNlFcMrNay66y
z8Y5/A9IzGmzOGkU3m2GDkpUPUx1DqXAiz/hu1hcJNKsAy51CqyI61BTIwN2RSrAlRlnWcv3LP78
frefOaVOQv1O2V6WGDTIuTMH7Qqf7E86G3Hf9BMJTGrzmO+D/Jm3+4e+J1pNvePOyG/cr6ioAm4l
iwehpxqCBTxSP3iOvW3sPipW04rwKVidrgnSrbA0Du4lcTiIfgBke9zakKGTQvQ9h1BLeMVsWfHY
Gx9dEs84w6EEufU0OQaEV8YZhW8aeda1JWSDvUhnWre4gNJPIEQiVbCP2S8zmweyrLgbmsXioe0P
jI7kbgu8QX2Ded89UPLvKbf/qRs8NEL0XHcKDwlRfeyg5UJ8wYXGPoSipYAfU8CNAlgiLTiDSkEV
9X2UtIuneyDKixZpU2lXu6Lp2B76LKU3HpBT4H4GUCkYrgG919nr0E6ekiEiT+A75ZcfyrUrsRMm
S7T8POlBffsfpUjcJQZQ3r9hyqoE9IXlrigopqk7rC5cRh5QI98kmm0Fwzg7S4ZRVHv+brRaDAkV
B7/VWn/UBdQtzWN7re9hEOK0pX6J7g7wLpxW9FBWrwk//YJBlMxF95hXiyEqpNs80UXxhUSpRaKW
x5ur7qExwODJycB8ukw/ZD4iKfWvq8FqPgzzIBCvuLNWpLCjopnQH68ANi++ZyHIwqKdb03TTU1N
vbozUB/Tctoa2GaYcNk8CcciB2Y3RPBMR9gHYatYbusnMa5Tr5TAgeJ67PX9t1wfUxyw8O4CdYHr
49rdXQNDuIAsIGVcW1rgKO85tnD50EmYSvXu0GC2A+RlGP6U4AXxvF1TsJhILYDea1E5juP3To9E
klhIncVCi7wKHmvUSP4fRTZFYpJ5M+3eyCQw4rbyeervVv4mgqGmf/6OkzBFwzyb9AMf6luxnrW5
n4+IzlpKpX4ha2r7QQNHLE1QW+u7g1qpyiZG6HVBeA0LrkGFMOMnZxCB+e+N6r1eloPrk5PSoOoo
jU3RL6B/jGpAen7YbnppQADRoqa9mNCETSlhGBoXtHVgQWedzGnYBEx+dnp2LM0Efoq0bSwqB/VW
Ra4u3lKBz2iz7CVjzKmG57TsUW598UaLG22plMGMRSZwrKeEBxyNHohGp5RLv/rTgUroWiuKZdDC
H9b5DelinTgG6ousUIfbzTGvW5e4/F2GVXCCpnNeUKi4IjCEG6VM9jfG8ko+/9iGb/sQYbYY6KB3
MQviO8QB4oYLpt3t37/28jxsaiVNiS9rFh+mYRP0kXXGGcN1jLL+YVsCh4dOALNqitr9F+ua9SeE
RSCqMM9KylYYYGwHJK/N6QFMrEN1IZXcaTzK6CdtXr/CRKIiRteY2EfU5YDMUFBkH8OrbZ06oKuj
WwXF1nV5k0nySg52p+7YRW6AyY0S8/+9uvnx8s8Uo/DHtDaHAYle6nJkYfXSkxN2Bk7Q53OuVRHe
rlG67KtyOobETvpBYU1/C018/ETZQh2+3w9Kp00hmLpgeDD3LJCVoCXiauxV0lAyf8rHDPbiR36n
OxGdcbVD6Q7gc6J6pP4yNE7T7dmnMv8B/aWUjB6uhKwcTCP7RD7ABoe1+tjAsnZJc3rFOy+atoiv
3ywAkgN2jfVlWuH/4dPbTvwMwE170AdWsBw0Yw0JeAc7m5exrkz/MKXX/cyUsfp2NFKIqWQ12e8G
hpKw4Nd5a8GiugrO/f4PyLpMzE6LO4+1y5rdGiurkpqBAU1GqnSiTuYim+5/8ocxpjQ6haGbij1Y
795tzGN58AlYq3tYKsCPSLYudwnFj3LqeGoxIP2We9yfr8b8LvWjjQ8QHG3OpoxyJj+4K/G2vyyf
X0Guy3MeOb4rkyaR0V67MTj/TZEtGdgEquv1S8rSgDGoZYauKSsnXc3r+9u1gkPuzRG/TGgsMQs/
TbrsJthP6OVJ9E8al8sGBJdP5OPdPBUIRKlxwWjpHpFdpuoTWvbQseOz14eIk+/YrC5Zg3DRjhjL
dT1YeVrT7CfDnFPCYHxGgnUKFYHkfHe3UT0W8Ouhpa8zqNLafFerEUAbi3aXxSVwo++K+FZPQPjB
gN27RJ5NyJNPUsAuIE8dR6pZBtTgplM6ic68QQBKVxgUzdiSiuSXs0wQ9a7k71wgjGXc5VLr42eL
VMYhC7fQBhfcVgUOWkvT4H8XtrrFwnMCFK7g4AKtEkzu7v7LT8kK2VPBY2k6FEsTYzCrtR9DmPqX
bxKuW9diacckECtJF6441EEfK4nGThwGPfPuSmrr5iXUgQQEfoiBEumKRT8RwVusrH1ic8PS1ekT
i8Ha50uvXxWXto8IHEHmIrJx7J0KHZ1EsrPROlfF/M3bS4xBzk7KeMoPcozmWOp5S7vuUSq0q+lP
mOhQjY3Jyfw1UoKeAKNJ0oXlwPOBRZmfZJ7QspK3/Ck4f5M0GBAXalZkyaV+Ew/zknz6FOXS2TEt
n9NIQvW/5oD7twkb9DGbHQinDzcPqNeTkR6687UeA2rkEwzD4oTWwGX0iie0lXo495VsjYZeqTqe
ab13oB2p2eQk62PfjZeGIl2vpeW5hEgQQ1WQkI5sutlEBCRW2bGGazEvgzp1PkTQXvPsO6NY2wv8
rS8LnMCm5mG1g+OZoAeMLGYfvfyuxPYPaBYK9ex1JsJDeA52dtaosUWiIHWqZZV7mbqqV3Q7f81w
cnz7woIKVnKBxqK1cgKieWozpRsQ85yjGni6DV6/YeVOz+Ewg+wWBLouD7NMmX64s9cWd/dLAug4
zCaCzVC4XF2uQI6AJeFpBCehchYenDLoGuhQWF9P/i/pld6U6rqTiQEoZFJO79HH3yo646Qt05JC
46jPngWYvWg1VBuMn9EhIFWhMzjqg9SvTWZzxcbtW1sEPJqwXHkqVN8uIdVi41XQI8mCpl/+RA1T
MlO7cHiRBX6kFpzDuH2peLRmiUOXFOzcQFqY6jiAz0UmV5ScoBoa+N2JTV+Jul44j06nRH99bbfe
/vA8eY130ZWuKrpf2rB1482P1j5/TIxtfDEjgTiA9KIc6fwjOk/lz8kTzFp21JomDOxnQYrIhIu/
WGuCAdAV5OqA9HYg46YVYwkqdsFbuZV3QQIrGtf3PJ3ov+hzbg0gvo5gIXWoTLLyncAcGBh6hNIo
EePcoiFrpMbclhPKcEsbi/jhHk0U0A/yFUPrUddm8FkeJlnKYe5V0N/vF2EgLnmduqS3p2vZc3ww
3G9I3OF2rTv0FjAEJkcYwbjG3irwVrrKk1eOMELQFfKm/xGIxjw6hSsWeApiSQRO+sZiQ0KATyWN
pKnnMLMs3SQKRPOvR0KjSmUHVtbKTY+6n6NLXu3OQNx41omNvDqOLQRuxjPZBpdhfcNr9Xq8vtuE
GjHOwqs4PWoa/QBbsQXxbXzVLSxLlxhNFUMVVpO4LDVKCHspCZ40RvcxCn2hqiq4lWBGV1dHGzCo
AjK+VJ2CWP3Lil79E9N4oz2hq1FEpaUIyCeX1ATdo9TrGuRfKLZmfnKb1ppp9W5ejv4BA4rIo8CX
8x1P2OCRd5GfjCr8ejm7Et1BmFdvWYgQfPtE5JI47rXn2WCbUyeV2vDuUh2FL/4BWzEHuuv2DXUf
0yl4uc6vbsJuoqKgnzRcE6C8xIF0kWFaPv5p1+7gpa+ln0+JIcIjXsv/q89eEls5pXlm7+PmDVje
9Sc1e23P3l6jeE0G5oesCDfW67tGdQRf/d3VA+6Pz9dMhaBN0uXBlh7Lwfr8vO4vzoZVx7rinYVA
FfHrFhGp2iTuabSEKyRHDN08hi8XnbvfU1v37Rx4vIFO9sYqQcJdsxAEEE39l5EXCToxcvIvfSOX
5io8BhWaHd+B6GaMtXbnbu3zb4dfn1r9cvHWg6ue7nnV0bxQKdFuhgYFA78wpEIUtM0CsmBJzUea
yaxaNweAIAgydonaqW8QjNUHhBtvFfmm98F95j95E6R5ABXQdc0TfPP2g3f5Gq/XZRjNaYSEc/ES
P79f5dY2vFUzQFIGDXaUEJAzw/hF8GS/RL6a/l8LrtbauGbxFyA440BFUojMSI9WRVjGvqyuinxs
XF/ruTomEwDmUmxFGrGrIY+UwHumVwVg56ubvFjKa8nCsOvq2sd5sQ7R1DzS0wn12rLpggnIRUs1
4yEr17ZZplyG3NPxk4eUGyfVnnjbrWakE7XfD8Tyw6FkuIqL3OaDKnVbAYWaMikL7WicdycPp33s
xlJauyv++HMXP8gq3ppIWI3GHioWkS3FscP+1cPqNtv9OXZfqfUrTIsWVOg+D6ZtaeRlTI6N/Tzo
f0GFmAcnwWv9e9VKry7/TLsl8fo3B2kG+ujSSed/Ygt1Uavr58z4gay8+gDcv8WCie9zVuackHZz
uLrlh0mlnpDine9raRUC988UDywxzwU1qLxJb3TtoEwLofsyafp6E84BnkhMbNBDHMWdVlC5Vgjg
RAn4aMdTQr6DfUBuicissIFfDKCL43BZReUoNpOtXgsTCDlDfVhsmvY9l7kIAqfajpmCWhL96FCL
EnDIe6dA8yAPsLUYD4Zpc/TaWH0L0FcKnB1KQeSxERJzxdpVnfXL2qD9CZjxKhnHgsjzgRLCla9M
KZt8GcaxA7S3Ous3G6JituEpmu7P6viwNljFxuod6dVWm1HusFAdXJUtLyVjEVCHnQsoLp79T0p5
Sa49Uwd4NSWSZLEzUEKrkxZJEEYU2YKIc4tsD2+eFYHRfXrxabb2qw75n+CN1PMJwERnkJ4IunOT
lbtj/zhZKjOOF1h8+MlElrVvBFacuWLFlS2ecI9KvdgHWeMeifeWyp4/BY8eZAj50cD9UKzI1F+D
/2T08EF7Hbm6mX06syHgDxIVups90CVgxrBl8UHapXnAQ8pZtswxewYZ8hn4fX1hLFkH1AnwfGZD
UnwGYlihyA8eAg91TnpTNXObOpHlS7mKnMW8KRnV5kJgua8kQOmIzfMld9qHBXODd7x56IFmr1wO
gVy30Iok467r05psG4Bell5yN6Y4criAcrq4zVRrGJa7rUt9yPwSLw8WP43qSYtJxEsQY+il4BwH
izC1fMiRLmlaZr9iIEnpLaZRm76sPthMa5esFTiU7j7W9zoufVRFg3hCnheoXUPFytDJ9du534/W
G75P0iHvxsKnVHGbBY110O959QuXeoD+2rOXQ6+q8GTMMJVfTy4jfAyapdzcWxRF0fou61xtj5pA
TQZGVyISo3TUpyz82Ktu0hN5fUvtTZVZjBzRm0VXKClBs5Hpe2EtnmYsg5Ol+0Wifk7qhx2rUuQA
6PZFO/KN9zqVeOEUsq8w0LX8RujDl0e3xZ+iDDsVrHJA8SBF2JibgnB0zlRjmDbLdv6YSsmGOoii
hb1WSK4J/PRe0q+2gLtsswDzTFMJfDEdIaKiS1TFvjflSje9vf2o8LLSDasu9imb6vMiT6OA15/v
p64Ka6XQFKrjLS7bAYbb/8LL9SIZOSwiXSeesRpneXk6mGoJbraoXLpuhEPEk/LkeymigK6ezJd1
CsVC8BmSXNC4RW8aJm09lNre22LYe/r01laooGhtQ5O1PYl+xuzCCiMhl/qmvqI4CpKVEkS9cGZy
vWG2+lDZXFZElqsVMZUT6hd4vN0xQx7sZt+Cjo6zVFggr3cTHEvhlFW6lnet03bLxUzqjD6Qvft+
htkxKvyBoCPTEZz+AwZxY5sE0d+82kmdx2xliSQtPTmjwWfG7wrvyOiysIzGemiNegb4eVJfFi8H
FpXlwpmb5jvL/vDG6yZTxVLjHwQft9FmBXRteWeEvJEQeGr7a2J+MFLGbWmjhUPw1JHei1/YJmQl
6t5wLDMDCFmKyNJ8UkRnqovJsWeLkVXznr68gAMX87hQE6qk0l9iSA1UI3uynUbelrx/RX15+14e
qq7O45OY2OS6XcxurMb82vJTnkQWgByebsJy5bx1ir+0p0YJ+AfK4cPWoZ3Xn5mTJnP7LYt9AZA0
/e9N8QfoChMaSY0K84Gn+nBgIH+GRLdi5HZJQpRw2UZ616LLcD+/CK+bgS4R9aIX87S+RGc6M9l7
0VBNc7KN/rrVPTUa/UVxP2uvxwbCxoz74i/uZHoCF2jjRqHgrsZGIOmhuEv7M0IAGB3UKciXF7IO
W+8poJkBUSCHESNCHStYlNkxlhGy/4sHUIj+aaF488a7JWFKINigeIAnG4RuTydckR7O12PC4/Pi
/AysrHgiqaLLo6oPETJHriFKti1nnaxjZgwh+mMEQ5/DWVRldSRX6DFqBpoT0NuLay2y2Q1Pg7dI
MIu/RTb7vSp2k0wxkxYMvn0M9i0IaEovltUcvLjaxm50bk3qFFpJjD9scdIzdrfnGJOy0NHiyEAa
nH+2Oer+TiZZrQjPHT3US87l1NjBtXP2I5r5UzC/eevWKp54GGzFiJhymnzGaLImrm0fJn+q2Nje
tSOMSzSpgJAQMnUIkAZoq+fyjemD7Psf/4D4QHwkI0LwKSNXd/4of4N5ltQZfgDxztTd/g4LOLFv
/vBDhor9srbYal4F0pKuPi5WrNTuSbaQyvajYKrnGWDzN6HHxoLZOU8PsLpaFezC7ttN8fLQydHU
F3+TTDhu5bfiC7dvJilw5lPBGk7GGcHCRlmlPXF1iBHwn/gGOiLrzi1NEnyVjl/8Mt3BiLU0psgG
CrXms212zQhiptSNNJVo4YR/kCoHB0jjjWjrUUyawAzZVc6mhuQMERxsCr30ytDoxEtX+UxctbNf
/0Y4qKO4taA4FmnokEwEFkJhc21FxFzvqbFJqXNloyjH3UugElEjEZT8ABiJy3geTmam/NFsNfjs
ns6A6PZpVxrYSU9NI5y47nD4AVZLfgjRmDdEbsKtIEV+aiHi2JG/SWMv8mvaAP7iAQ33uULrqcWz
bCrGY1niHhp0ZILvMY/cCr5jiogwVihkQ5q8LadLKLMXWPMTHrO1Eyi5Yc1pIbKarwwYTSNsgYQ7
c/vNX6oSnAR9B49f4nQofqWt7OUiRhQ5Aqdp7YOReR5rl99lGvmke07fy8x7S57VjQXwQQdMsLkN
FXthf+1HQqYEbKWx6sjA6fuJB3FZ8UWcrZm6lstWFTSNAw2VRhWHC/Q298asVlyaM1YqH3PKQgt+
1afVD2hHHoKd5r9QyoGUvVPVoY3D8DkVxtUYC1nOACDPAJCyfsokWSzCUwlzaQ6YmJrzspW4nuPb
A3e+ZFhuOqEPYhPXnsNNGS2D0fpfrlEyvy1btYmrq5zodkIJc4L0F0rZTaa9dfmtThn9bbtWkapk
djqBKnSVsCdAvf68oP3yp0NczE233gvqPLNSoGHxP1FyezIvpG/oGGB8sFPlGiarkocE3ckM2kvf
+tikk17daD9kR2KUWDAYEKQ2y1GlzJKiMqZqT8b55HaNeG1P2/gaOgoTIsoFTFBFi0+gGB5o6Ml2
VXcTsySsLtZIAcj4DebJef8WX+vM/rLp5zfli1LZlP+QAElfcIBUP/VwOnq1RjBd10iJTVqZ5hFM
39sOLfQ17ffmC3/rCoqqGbRWfVgqoc5JqDTCSZuOYJJyKpJjnQsqTfMzcpATCI4/Xzu0q9RRVMBC
7FeENOUg4jq6EnBAwpwIlbqfLjb6vy97ssEmK+9M4uCtoa6PGNgeh7tnRXF5LvCFAkxJrQMlHOgB
3kwakcVlP9zFJyH0JhI+3Iw6WNX7mmWdH/UczWbInttbbtape2n8XxEAZWSMEkiI3coBXON9Z6LF
yz8uyqLPIsqDi8bEbPGRzre8kGUd1lxPGJ5ihuCgcSr9nBary/YhpxG6plBB+Aqvy9lPS2vssTO6
/mDkQastpB7XkdIUZIqUWwdOH02ssMRSMtB70lSGt4ULk7GvZhZ7yWp+Jv35MgC42/fK2YLtoRSH
it/xcKrSUerWagtN29noZb7dTvcEc2pt8R0SGTTthOQax+OEhpZjcmLdtdjpRz0D2toJ8zdNfVeY
wCkl3zrp2FAm0TW6m1nME66p/JE/jvRG19lnrGzUT+IgwK4MPgoB37aVQQYJVEnGiJgeceTiwKJO
dnH4ARMdeLilwKZN2eAld+DmOtXqJCMmDP7rWBB53m97joqPH61aRJwCglN37zEatQeQg7mjkCrJ
ja85W1Hu5lADRC2adI7YncqhlXlwZPqObru+Ygf9uPdgTMPrPLLzDSZkUfE6/rypTCqJBjG7RIJd
GUNu7nyBhtAPD/b+RFwIDQ1wRkpCysXG8hB00Ngbv6I6/z2vhAJTrZ7BZr4dTHJyZCfNXJ/0+68Y
8vIImskfXnfMMS8oJIN7ADsG7JXw6ZJND/eNzR4x1t1n4Z1NbxTzi2ahNrPuJshMbv5JzYCFGcgS
HF6PrO0PiYwnt3fu+4IAitDy5F7aH3kjwA6xHSvUY1cNpTRSeNKvhlsDq5xNy5QrEe74YOkAe9fq
wp2I/ku87ma3424xMirmk4uIs+cINSteMK+g9bSkf4CjffTRTzdNL8KPpvGKMf3GstQ3lSs1/hiY
6/k9sfqtD76E/aHOwwpUJDzCIomw9IW20Jbgmomc6umkvZratIHDlvn7K4HOLW6tkIHaayPIShP9
aZ4kMevQD95KbENLSncbAP209qne1lObHPhSuV8Bsp5wsn9PYiVSwK7bHViH5PKrroF9pnWeWbFe
ZnfbeNmiN6yy7c848gUUs7UdH/CzQ+uzewSVpmWdHJ4+Mg3jeXMVTvTUx+299L6V3GBWGSuMg4Mk
Omwroko6cW41PHha9nD0PfpDGrCBSbox4tZsqUhcVd8/3VupdFPSM7anhBrxoqYapWWR9Vnky5Jx
BfKN8JT0yyenck6MACZNOIXYr05YDB5U7aN8t4Uqu4tZU20y3rONmBaem2K21vMobcvz0fxQUESk
OB7wlCe1iKCncrYA/kD2H8tjhrLUsknwq/eXDCIkUN2gqag66MIPhmV8jc4jVB4JR01zp0sURops
215gw6GYtzkpVne/d6jCCim5ZFGK28Rir9GNbRY40bj149TXtX+dQwjB7h8wGhBLkA4e8iMmi1vq
EBTcMeQE45DKeSpruX3WsF1eg5D7wx6anWI+LLnLlD4PQW49MWKCZwjvH/2fUGZxMVfRNG6mZTq6
wGvReSS4cX+Jv2rXp5wCl9ph3B/0JyRp0U83+V5Wed8Is2sJQ1xD51Cl0iP6mtA5nZuTMrHANfAi
iinSvXKB9TQiJI4DuY8KvJOubythIV9lZXl56GjncIvjO9FsCKWn23mfMOwPh1IkNCUeV4mbucrV
r70mBr9tk8HLvfu+Zgpca5m6ne2QdX/+SWShYG3MCqs2ko28wMRQ8TJz5jXYJy8u2iaN+IV7c4yC
1SEzZaJodXJCcvFDosbGwSvpzMr1JPzv8PAgRYXKyR/BJTY84JPgkJMzvGCGjohlKFiD6jsbTeYV
21qy0mhU52/njIB21SF5qa9+cxAL2mQsNb/J2EpckQ3D++Px4yualuL1AzApZmxTAtKqZgvodzeL
3sBwkqQJOnPOuiy4iUqiK9Y/XvLlfrQyGwNxhCa0PkJWdBuF5I1ATjCmv0LrAg97QYT2TBhNSIVo
xN2mch4JONQsqntqyUTsov6XF9b89Eq5QL3RwKd0REfDLb2t909Zvhi6dp6Fm71FMLycNOJgnInv
RtyoRhCqRE1BJ8KiD70H86wrXbzAq57UGq9l8XTG5aKkdnRv8aYk2jzW3LFXfoli3rhWKOMH+3AY
G/CiT7z2DxDZyuvFEl2d2mSc2KTsKonUGwkViOsf2DveoCgjyBTRCvxf+VB2zkqkClYsVtY3TYS0
AScdFH0OaggkGq/9egh+ej657ur2bHGrftVUFvEM0nbo4A2ydaMlhYFxQPMMvN6Db9hLtBqouyoY
hL0yElhVDFa3c8pGShBFPiMhng1b2EuS2jIihADph+lJ039MOSYQq0W3C8yzCNTPLwlCuqbEDxXp
pol0s3w4hCLs8AOQQ5XyQ9tnPtSBQYgL4fVbglk4Ay+Pe94nRlxDKmZsSXfgvJtrB8QaDRylejBH
ihkrWrhJwp1RrbG5NQulgUQw2NLDHuhEm41ZnoBRDkAr133EoFvMxBu2K104YyuI5MCtMpeBvUv7
SmsimkIy2X9aIoyuDSscaigUyBEMfotFf8ur1Z7wYIlmJ68DiAiWV/2r7eFu3/2oK81Nbw3WCtQp
GHTCXreEVFLucU9x9cFkAm89N0FBBr08Mj/uYMEWWtcE4zJrl8zh9eMS4OXT8MVvQGM3BwP2GreZ
TE1qzjSi/MXcCnCbW5EN5qkwOH9x3Qs3xwz59vEoaJQD/6NxMkA5GHefaXg/JzKvOLycLIfJNaR4
P5FFpRvE6HO5hHGptN8AQ7fZhea/d100SVjs5a0ALc7NeYi6BlMJZK447tnY1xb1JSKsgwNDEMd2
32bNHgySLJ2Xt6pcKTUrng/oHP2wTAR6RAYikDbO/ecVTfmI74apYEzDRv5N09t/uXPbRskXmx0E
IYXqE0fo16w5vOb5UM/XcuD3xpZpHJMTidDy/k+Era7DI+phLaeIlidypHb3fL/zIOV7SvlmCawD
+CKMDB2QykYJ+ZyFigTg76V8a7QZff+168I5JziYOYNLE6yTXD5M01dkMT/HVox335jLzHpQEgKj
EUbGLeA1x7e7QJmlmJMQiq7tbyrzGl0KEH7LhysvdKBFsgULJc6C8Oo3Rj6L5wc/gEBfUghuLgdr
iaVmoK4i7sDY08fGe12s5GgnqYxK2A5DGkbqXA1EYRIb4U5/IiSPvhxFXarv4Z1oXYI3Vz7kmmO+
7b8KC4zzd6k8CixRHd3vuLV3DVKha0cU0ctZYkPUAkyRkzWQRFWU0E8PL1MSliPpsZR6pCYuC3pz
CH3VZvpCgsCnXbdwY0S/HJXLWqmSlQ3plUodikrdD5Hnh1X1Ji5WF4Qxuu0guPiV+LBiTFhU3mA9
nVYl7FybBtBpryroB8Ins1z7qX6wOpF7O6FWXGzioTpzejEFrL2lbb9DN9GE99hpc25rKpPNCmtC
MwkLo5on7knucTj34QRrtLegCdgAKGwikXWie3s3gwQJahoRKteEylYQCvAM6RQDy6W7qaITTMgy
9+DiD/X5sQMpCFLOsiL+ee5bKJtCtm+LF53GLQh1Viywgn6cH2IzXB58IqCMzU+nWpTzAFZtLFzj
L8yPOWsjQc66ix5rbBjvHq0qqk1V8jGqKAgILM+qdeww8BGlNSKvKsZBH98oNdp4As3I1cWqoTgf
KFyuzqSdGQZPVbOOLIxEMginMXfn4593/O0nSZl1Hayu7ajtjnMJPbVScPfGegudtCSdHBSVOw/v
s6fKDYz2bIb6y2ro5eIsI27z9UJaZqM3gVdcMg10v/Lza5zc72Xq9p2KVY8adzaivm8V9JleGiaQ
sWTTqnuRWKBR9US28zPjbMZFDqHkGPhyoXFPbfwT8rsWde3Csxs7r+EL2Te6/n5oHmIQteTQfPvP
QWgAFujE8Lr1uK4FJbKn7xeLGPN/pG+1jNxOEqpof5B/ZZy87dV8/X2AZy/4Z4dOYKCx3jPVHCpE
sQqL4V0bHLo/Bltt4GG7YHyHJEfw7HWQ1zX1mJi3rczk23qFUau3GyIjqzNe+WjDgWuBA/EMWihP
o/KKJDzrZYSbWUL6BNgLWTS3gDsey1/suBRP8g98NubsotBEX8mjINnzQNimb+lMdbNSTwOBmU88
0EjeE6pbOFNt1VGq8amqbgBuSinAqZ6N7dtnwSF8yE4Ny7/zSCYuol/lyX2v3Q4HixBvycOYJosl
YIp7aHCAp94IcgBZFXux8YkFIr4sY8K3WUEihqInRN6tYaerVwOnYmOYUtpVsW1OL+DRs5oDpTE/
HaR3w6MG/gNmL28m6xf2d4ngWbw3yYYH/N2IjZifsM8SQuwIw4WzivHFIm98aU/Ge4ESYdsVXqfl
ljs7a26HjZYZQC3WXB8w9cfviNpmcBE22Waa8a5yGqtHWT5ohw+/TWFEisdYHSHQqZovU9CreppH
lMwnbkex1Z46IPAMIbUuyOHUuGSTxiAvJx9cbOOpicF/kGm/oHlcWDYZGUaEk4EioiOMgZ0isy3E
fWP5B2UFoYhDf2pq4xNlFgFAWNAnt9Mk/52DKt7hkmdGXzihkgHcQR6fIkYRZxSLNrGqXpLlNeIf
RRRsl9E2rve//6IX5z1wIyi8gFy8khwfRJhtRhUsJn8LxUUWDoUT25GqzdShwgG79aMnfbdDJZJf
KGH9zfyEu9P96XaC0ayqfaK82ACsBKcMd5GY0HgfNkR23D314GxPKBcS7mxnrSxpe4kDsUmy0D2L
nrLG+vRjPUCNj1WUCBV5+WWhF5XH9SXilAj2wlrC/B2kaAidSLJKtxDl0mWKmXHZYmFPfs660Wpt
5FX4w99AvHvpu+GCbQqABu1hBQis239OO4IPM3EfYPBh2PxrzDBDgzkeJmJRd84IBOjhEbgwuXsC
dXcYjP+OTNybJJYORLxBpU9XNMoP1qql7X4OnqQ07D0uGOpQtMlGy/82bBwoUkEpdFAEYlGjifAd
BsijXVqNunjqgbYhSsv+NmBHH06WwEAU7K7Yu5K75BHos5JIv3yzMa9NuJ04Nx61IdRRYKEaJuHA
FDMzIdokSk6WHlRSBfxBCntXkU9/IWot+/HjKVSf/m4c2W4FxFrsIGiXo2TNShVXPrDBSpeuShw5
3qADfjlmheNsjqk+jkGWDWhoy84hDxo9OCmbRnxDY5gATYrXOKJgo83u3HL2DsfrDEksWFkzJAas
Kw4weQS2B2RMG3CTvTUlEr7XTVdNplHoDDkp+Z+9jy3hXpgazLsXynBtqqk9SE+/BDfq4ledzbFX
HmtYLeWEzbijYXwabDQAU0GqcKs1lj6+bi/t2DCZvLc15jdq6+TSYKuMD+lYy5eyrPDWLaV50rwK
8934erqgDZhr6nSMrZHAIw0NPhm3PR4vqtGCiCVGoaUCTeNMfeU8m0Q6dUAYkyBjC+faX3rIr/1V
sbVEJ2a1Ps/aFFnVH6z5vThqK8G/BGtr8unwgP/kSOp9O/b6U8NWdKynxn4HlHrbYJL5AdI3v+WU
vYa8aDJQ0dDBt0gkOn1T4WSiy4EG0wIo4BWfnzlTiBQqQRVIKW9LlOfBnsvUJ9nLEu5R78noWNzH
QcHncfqTADV+CNnuh7VHDbl6d7rYr1s0U3oh56qlqlAF1w71SdirCT0WOrGCgoKjk/SZX55yR1CE
TZueOqLxTM/TkmjwRoD29Amv1gd5JMKk401txNZEaVlit4BNzl4u26M7nzcXMCH8lggZ6wwar0FM
TFKoCVIasSPzkSHEjscq6BH6/Y/XFDRjj3uGk7hCHML6oHgkqBPqZlKOeHD5/tP6vJsBDE0k4VbN
ZMgowK0AMEsm0hKEOIN7ZP7UJOq768FgXECiPfWmeCG3MecZmBeDPiPbVhSMCQXZvdzkvywh6WWy
HEhhmtdWB4Br5Fm74zf9PzKsfRc1k0TOT0s9U7udmygjl8GK6LysOzU7tSWiXh6UJZi6eeMyTBVm
Ywc1tfhGsCFJeDyXCvkh10tFHm0oFoS964sOQijBvHoQu0aNHiZhYqQUEaXpQEu6h4y0IoYvlDrD
C7BjZWvjnb+gUSnEpmTMyrwPuLVC0B0SV+HBeNBP7ykljkOkCczo+C2IdUjX9XEjmSt8KE+6UalL
J0++v9Bhlwkq1dpxfNak7jpZCpDTrjEXZJTeUbnYrFHQ5q8gp+Jxa+8s0s1wy4WAa0DJ1Gzrj00k
ZZWgFB0fjtAyK95rA0MharVJ3zA8lkyUft4xKogyVxP24lqmuWCAuVTqpFKCeYBpT8Qh+fSbnbMb
QKFWloJVtWRoX60qqcOGyrsdlXPfJ3rez6/S7wfFRyGRCfhZPUXfqX/T1pGCz1LBErtrKm9jyp1M
pcgOOUUTbHh6ffH4NGVFvNnpryDhfAU7Chyv0AIcf4+//Hx9fvMCV5pXHl9jC5pb+QXPnkarplgm
ZIaTyxLTf/XUN/rWwMrTR+B/GuIeuMAbiyoAaF8bubZjFE41HPKefo+Uqz0D+9n950HvGal25V2a
yT9WHrQMXh2H3hcw5RxNJVPbylP96yW0nZkr1pKFRLkqn6hm4212phofJXvPQP+C/LlDstuS+YE9
6Bu64ldkVA9tc6vYkgKXu1TyMiv9QXRQuToQoJstQc4sowIEzaXxUx0PE9u/79E+65sPaQ9H7aHG
W5LZ6IBOYbjb3+SRCxq3r+bsXC1vON3lzNLyqlrbcx09Lo6l6l6MVcRr7EjQJrDmzoFRhSdzryKc
ywNFDO1kNtDl8N81Pbhz0Ux8QWx/U85mBUogFrGQUm3UA+UA4Q5jgDOfkMOaB4+qcdQqTsO9+m2B
V6rBDcL6lOkTw5Cvjrp6+MYtwN1XFXvs5SuAaeiceKotqFhoMmjX3mPgb0nKTtaqMvFbCeb9P1Uw
wiGArvmeD1UN9ugPNJFP2XT/JerAEv1oOkPM+W2AFiCmXL8d4XNE6BVTfRb/xeDXMLktO8QVMDel
DfmVARC3dpVrTCeeXUYZj1ERuqtoIQDIkJM5Kw8ittaIb67cIYn8TNCkU787AnN5mruvtbPYK+8b
31CFAlJfykE26okul7gjpeRTPcnFF83X3P4BQLyG7JdXBQPAdpSmSCjCoVPOpUMO+6cV8paWtW3a
+fUvsMZ0DTFBmYhh3KMuKTUiB67sxW4C0ovkS5W9gTR9L/LtYdnB1CeFRtAXfgK4bNTRL3gk+Kpi
mSvzFro8podksyth9pUyhIs+ENeYdZDSb5Tx+iYaHmazay+1EFWmEQYIhPzYb7N58YcUlxgViduk
DZtW+vgLAejljkJzqluo5N3GLkP3+KbB0e3hR2kl4xhDONS+Ba3fku56/C5XKGHp820TLZMzD8QP
DzD5Li90na+XvOYQ/JZHrnHnk65hjtF1We3yPFwAyedMQQXT5W8lIYLgsXIenP3CT6Stb/b37tpi
NPHuLlkAiYU/p6gna9nFp6LIAbZMPXOzmcXh72I3Z9vhAKvUm6BJj1A37rR/em87VS9WXffE0vpf
X6bYFGxHZbGhvV07weOAZuoZS6U+GkFN0LFxdbCGWXuoSShY4RqMO1c/e8PDFLH6iOe+JlGO8VHX
TrblSoY0lB8e9+/XWHq84UU/mihwTLwM0R1LehWawMpgOIsVuFcTofylK/Kus8nwsSDdArhsCBgn
dqjd8hhoUI5jGanP6thaaidqc29OfxYZ8DqZmrLFzLRhlDRH2oaQIOc29lohuJagoIWVD++xj/FE
zUb3SV0xVMzvavt2tVVoMKVdfzmTfZq8Jum8gYgJr7LpY6Yndwq2hmciTTJK4meW4xbOD/aopyyp
nohBfd/0Wt4SUaA31pKuqXAcUeISPQJiRF6+GPci1CB+AQYYiujIjQN1C9GwIBPKlWdW4Pglpn27
TzTIEtlJm6KwE4N5QkSVKpHvZ+3efiiY5jK3AJkiX5jJmxCBL+ct4Q3KXc2ZC831+M/q+hSVRbL8
u+MYd5EtaCbJLsMT17mk/RiqGTBAxleBrDENOo6JzFfmtm9gYkbveS6u6S4hOXj0WYqRjDCpkE/9
8+vl0fhH3avr8SnDj+LCbYB82rKJcakSC1d4+CfgA8KfVPRQAfbITg0zUAFeHNEYbfYVBF4UgXp7
1moPvTWzA+X7x2KyDCq3PrKCciqc+uaqEWvtBzCO8pKkHsZMH11/Z266yCDzBTF0hjC2IXUCOfM9
DYtqgEiogUKrIC9c+SZVA64qTZXcodxkS4hbbW1FMOEOqwQiSnQxsraAIENhFnV6mXuHXM6y4m+O
waKka9ZLO+EesPcNxwAhh9b94o9NxZpRLS4tQUo19jMy83S2kLXtGvWx8NozvVVUS05d881tHhbc
Vh5mJjneI5IYCZ+nM2Nz1XCTRZW1ZDuGr+UAV7suAtwuK8OZsm1t54Muv3uLRAqSn0h5VU2MQfmg
1oN1lB9eqh2wPGi8R0/R2du0SFYZxbkyW5t+MrKPWus82drnKsHIJ7uizfq3ZP9AcdN2zN8IPjjd
cJgL5tuQe+3hW77zI5N3DgOAd+MTZzaBEndKOey2y8uiQP6pme1VR4GsOtOBoO4mr+0Kkq/PNXGU
cBS3YmqonI0nanR/slmsfyy6FYdcZyaQNuuoJMzhtCqPIfUClDIzlzWmyeyrgK7Zb+loJYlPmt05
vd7ImYyFtgLwpcgLhfkPcWOWpOx99EDwgCvSOQM3G3lAnHGZfhaOzSoh+wZ+sX/6J9us0rwu51NQ
Z2PCbQxOoW/VO1Y+wNNFzHpY3iASVSwkS851STTetiEVTozOS7NgImrbuWSN616VRdY2CETyno4e
lL3lSMDB2og4gkRTzinoLQgGN8So6D2mZSqzp9SBwOYkVvGdP8Qb/XoEAh8JzLVZnfXNhJgDHqk0
4RaVoVEho1XfbJl6OZaB+23nUfSK6qWa8OEpk+j9h4e8hOmuvoEHkH7AbaxTYHRLvFi9Jug4yR95
Lcu3q5dAAutW+qd8vpCfBT8oeChzfeQ76siBe0/kU2IMYBVzYLo9yGr08bemITsg5/SdmwGKv4Oh
tRWFSiobKIibEZnTvV5ZA8EPN2Uol109ABvVRU81IG9AIis2AO/URRuVFtUo5B7k5YDzb+KlpTge
p9z5Si7BPD0guLORwEwsV9zV/dpAEA/T6SqtOjxU8uQw4m2hUcvQTjUuW6+22eiwnMR9TssUSxZ8
MD1KadA7L8YMb+8rUdlRkMcApJGWyiLaBlxzwufp2/8pf1PP8AOFXFsT6hUQOZ827yisLRomkhx5
udyMi9j70sWAo2qXmqruDv9zDFxEtbO8SztXa774Sq1XtIzKo3fiN204HHpDnydFModywpJOmkhx
7I4U6HcJDYjzzKoa7r+gglyZ9v77MYzhLSbH9CTe65SqcB+1vFh2e4f24boV0WwIARMdXMlehKm4
NSveXRxmDg802QsCbDKSsAKLF2MX94vEfTlnLVxt+dBG0+2AhU0/bDwXy5jBz4/G3htgGbRRYzdJ
FRiPUGnN93HSfo4rxyHyCIaY3RAUTsrzXhFw6w/4hV0NMFYGoL56Fs2odHpdMf0fZ4R6UjCE45bN
SBgCdyf2bNutj46G39/TUdq5ZRRdPMY8YAPWMgs9VK/cCJU5JG9Zz2QrtsDj2sPf1MOoJUSSn74D
yXvnOK2HW0WNq8J5x3OKyyLEfb8/uEBhrR865oKNwOOlrtxB0YylpAOz3Gcm2w7V3jwE7HaaKvxE
bOpkh0IgUawHUsSoLzIDodhJf+h9L96ZTR1W1eCLRJhf8SIIl8ZjgtTcj8VF+bS7FmYREcafdyfY
55pUPEQzFYdfR+xc6TZweA97Vy4E1PRUgACSnZM1YwKMS/LRusSBHUtXSlwafM2MtKRdPogT4ZjP
81498kWM1Ai0U32uNw7JXc36zLM9KnGytq450qhcfkEXx6ZffMmz5Awm6Wq9ndNRv65YKLhk4pBZ
G2rvGwzkH8ZyvRpQ7o+h+wC4swjmEpQo4gLO5LF7lHzabjYrlTRggJOfEJNiLTO6t3iedW9Q3KT1
t1JFIR9273w38iWE6lWQ+EtNiAYyWgXRshvJ6sY11DC8RbVeErtCAkzH5F10dmqjNnjgHC3I/YSk
dIqvamr/VtFkVZXXY9wgmqvXnVqHgsziwfMmq0cSA/3a2Hd6YTqbddOOS3+LdS33P+CsOiuhwUjh
Gego5xuQy3gHsheVWOaYAEWbMyOV+texZaxt7aYONDklAfP2y/ZLMT6q9zqCo1QwTNo0HljFv1x3
euCUCfIC9/Q+Gq0nnQ0hXCRQngVH7cvJa6BWWddcDa4VOkRYzePK6E7EmZwiBr683VU6gpmVBw4S
ddsHGNU3+dHSPBk+p1y0488fuSmESUCVx0AvxIOiChoNsxFKAIZrsV5t80NTW+hhdIzj7n2wU4OE
BHrOKMZABJX9ZGepHXpt3to8GoTl9N2BlH5RWMEY007H3odZQbRKjVMqdx1aafu+e2CExJoK5rin
7IZzn1l9/z8JPYh81Gi7OOHJiLNAw1P60oVA2XHyYOM76Ix/TsOLl5Hf8NLCVrDNu4g+SuUfVpIS
tfy8M192+xsOFGyAXJbGqFJpTSlCPNAufuPLR7ZZBLji6eL5nzxOLyC8+GpWZQGRxxwrmHRVMrA+
XtrVD+VWSEL+nsbc04opTxGrc6hTQg7iYxLeplBzFD0y6j5K578IIxo/FW+/uD7RWDlJdGJ7f365
p5T4AupEy4ybouQ64VGGfykHbiMb64kEMBGCZl/MLVLt9G52EMeS91CXVgucEeKSAkwuVDSluKjb
E4S68WU8zHK8vzhLiZ0bCSzc8m1mTBopfRrW9r6DJwtGkeRJXyCku+Ssp8vaI2tID7XBADrifAlU
RiSyOte4dn+zbivdx9PoEDOzq2qbxUB9LKlh7CNcH+LwMwd6GVgra/9AAugSgrLgVmn2XreDjfDK
HRWZd5FjykRwEBFolOP89Hbvl6Xm7z54pX0ACQ8A6irBLdTp0T6ZRGZ8tIr8y+MOCC0INYOpcFDi
FevOsBrnW0XM/TYIsxpRQm/4817ZUGMMzb3hWd1FeqtVOBmEPSvW8Rb+iTSriZX5KptJmG84xPAu
qPRnNJCXjNb5Z/msIFBzIaqED5PXQr86KwlflbCo0EGgtR8meVzqv1+kDOGEVGZ0r6Jwhi4npa8i
jTPp9zu9l6hc+PvD/Qfrn7MpkpBRgZ4KAzjmcPqqDcwinn4QE+n7cBt0IiJNHHo7R2/C6z4LO80r
JguaNmCp/oE81WGQzbvVEqkyeCfcb1o5Vsa7U4TkyJIZN7CVhwIcfGuI8OFfxlZpMpKyTCqxQlPb
+Im6rRFTIDTHZ2BAXE53HB8Wr0DnnEmkpTsmf6wlnp26MPN1r0D1ig049n5/ld8MEE6eELe9JxYV
BScJqr2R80HDeeIYYT3Z8AUlrNvukkmwtSQYK6QeEsVG9NXj6e1wnK62v2q3LJ0gNkYVDNopWryi
gcJrm8Hqj0PKufHOfvKP7fS1SH3CNTPiFzXVs3gAp62YQDYCaJ3t8HiVAIByqAtdgEkquKLoSFBl
KCFar5v1jAQKefOuzGCnvO0ICRt6UIX8GI2GS1a5FtknQ8zbBr/+7mCTNaGHPY3KOMiw7RY8j4o+
DPz2OpI4hCtIh1X50y0ksBFb65jW3Y0qRFaJTTNU34hBDGXKhFznfmxALA2adLxCx5oThKHKn4Yo
RjRgS0zf0lWrdFq8aultqnzrGjnoYqCXVbsIXidjHFG6ZHdGGHe1kAHUVCaCvU3TZBSaAhEKT4qR
vGOP2vPRfIIXlFsbto2usRcXR8zNwKNj1XQDpmZfI6nzXREWWibnlp/IpxpeBQywwePPj1YRfrdL
swWY30Et0YjSRDFWPImYynYT34gRmHRUhrFmHjNjMmae95AeS8I3s6VuQEnS4sdzVBmFf4c7VP5f
7rYMKm4vGRkWxQ3ttFKyYeEPoFkxUpN2ZJOQHpTNX0GJ4DusJEWc8SNJWV+BvcTtu2hcAsaRWr2L
/U+21zg35s7sJXOP0YRBXI1q+fuJU/k6Bn/H7gLKiBpyyFIRKAY3GmvAXojXJf/Q8LlqQH0Ofg+T
JCU7mI7scs/wC0XOAGeW7jxyEAYfF89ez0MiC9fHf7TpRqYY32GOLI5LSLB/K10LOlDs8B3Kbs67
gNo+Z2OpGAos+EzIkxTQT06AQ4eAgMl2j0icIdZxMPCQgakLU7NgmqSmv+8VR1XICkNeCTtTGziZ
ADnbhRmiXkgQrHi640XDCdgkBwOHtzB362MYhZgdrMBZADlGtM/oiDf/MgP/PO9LNZjPIV4liU4U
9qqaUFSg/EyRzReXsPnZuIAdOj2FzYFrYXG1KretaC+ZkytBsNmKqOrIiOak0YdLj1n+QQg3jqSf
wKau3uF8LnTsy3CTbpQ8kRL25hsNC8mkjTDdUhfKVOuqfztfcfqStoqPgGJLa2uugUGX+Cz5ew9u
9I66nKDLqRtBLGYtbeUZK1jMGe9N7nLcMfxK3K5NLd8FvSDRQWI8uoxD1n0Z5gIW9QvsRvkww1eE
KjX30KyrLEz5a9nT+8tsDeS5gjvyNnaoYj/2anUkoWqzz7V1fiC4qUTspOVQq8RLNegduzxmTNcz
B1vZVKdN1KwGunp4cCUbMedTM5EgRFDZJsZMsgw1w7zinmiP9EGo01pueATZ7vUCq2X+z5tK7Vjv
Q2fd6uVg68+/reE2TD2KB+Exj7nH09KADgyV2gyyzNwYwh2LshSjhfC7y4Bjof9PtIINjd+SWxhV
hMeBxsBHxajSew2ANiEQuezvUDtwq1DwAAf48ySB5A9wL3iOK3FWqlMCLgR/gh4t8HAwCCmaUi5s
m20f5DIDoNAtFZSn4yBxTOJ8J6DxgCX69sYWKPkgvHNv+rWBP3VreVTIrEsuUE5PnrV/x3jjnCaD
jYfIFHahdue/nktba9dV8A/AAdCjKkUXPTTCcpuJIVmbH3jJNaayggAtngA8AqQXD4Mg/KeqcaQB
qTjAlcOS2KNPOBIvj8AlvtYE+5hUVBrpH/z6lB6uRqPdFokvTKun8wzGOjdNkLdgxYCVZf0wiWJ9
pPWnrt6hlpu7OhdF8/2q2YU0U226AWhsUxl0q8Fb02K1NC/W4AFcsAe/OW5qm17Y+qLqjtXuBm4r
0WAeGINjj/49QgnnrRqhd6kcB1u2qGylx4TYVmEvNAIJ+0m+WtcG4Bwbqk7+jMUY7/PPAPiAK2W6
MVU6CWfLXfYsERkVb5wqiQH4ZRn4YTkV0vGN3ZepRDVUjlmpLaHN2LWqwotRNh7cXwvZ+KiVK2n1
vlX1EK61/1YtFE0z2VLsNT1BjH18GQS3wlFQuEUhibKH4U2ez49/L+MUwTl3+6hnOlrfNk2PWm9p
IlWD3wCcDxDmzVeObh+qav5oZ2klJ1KFStjNom9jQtMNLNXu/VEjGiP/txsgQNwgW6vC0a4HHXwS
PDoBSXU3pYwhQ3rj2KjOl/8ZY8dRtQQBN9GTgmvdAhguvq31+EqfBaB0cY8ap7rPk6rWiIiPC0Cq
Rp3Hgz7HsaESn3MSrCG98W83OP+MIgpwXYAlWKtieqSRTy6jqBivP3CmYs2LQpu/e+5JBQjr+KEc
rJ6fO9vR/HymZ6hrSNuk5oQ96S5WLWXNd28jSsPyd9DeKWRee/ZUK5AYjruuZgupvlkrFYu8GRmq
qIUQZyCyW0FZK7CZl1ZCpH1fzdAHHD2oxoB/VFXYODiha21StDI1wwFXYjf+DXPiQF1SgJxFl304
M3puHhcHbNVHN5JZczDfGYa29gXeJz4ro74NbIF+4hJIYHrzNlVG7pc28Z+TmxonKN7/BSGwRz4M
DE+n9/cQWnNk+AjYZVW3sRgkzn6rw9op4uDymubZRCCIHpWwjWgHU/jrM/hE2ZoAPdJWHXVb236N
RwyFHg3JMvAnen8tnl1w7PEqgsZNAxrch32XMMlf3PMMzqHl1g/cLRb8kxxuw62+e3f8kS4thGsj
uPElOq9fVy+LOKPR6MKHFJyeMPMpiZmQzEmuGdKECux6rMrZ7L/VM+g35OkXSyK6gjEecRDdSDOx
mmV5li+EmnubHxYCjQUs6bXg3po8r1uGVODqqICiLX9Vf6d0wZf/ltDYyQwjBD5hhnpwb4omr65V
i1Mq5NScPgRDAejrn0ZDLidAtGiEV/wg/3tkMBL2pj3PKQLhGHCwYmBoEdQTfd//nMPTubNE0oc2
LbaSy2Rxk/DJBda8cI1NmUbRWgqF6jtXaZ6nNuFxEuO6nrSWIu43yplTSxDGT41OKD0fBMObrbRB
8nH++YJPnNJ84u9nY/zgdv4yxTfbIxLzSM3wehS/LlEfQZu+/ohzmD0xfjFrSMah1IaEG6gJ+WlU
0enzztVsLYMezdjbMmOtJdxoYv+Y99XPulj8TtFTUo0CAIBWu1pm6jo6rdVHVvKQPsa47RLRLO+A
RnFg0Fsj3M8IIF0k5pMshTjlKXd064+2ebHPrJWrMDUER+LEpfsf9ZNfpBdYQ9Yv8YUVCoDxmmGd
WMGeSC81rn8qnzrLe7mazgCddxSc6uiTB+2m8BJdb09U1P406roIz3Hlp4ZepZnrJalBFltvkP/j
n34q6e9zK7YRr3czbQZ/ZsRGr2rgayDCR5NuigHr4RZZY/GN8dGEh+yko/o3kF1k76tSdNUbpsX/
iHxUTpUIa107d0hOD6rXtjC4Nz9JRn8eI2apnT1SuBrGU34YFqxjXenXxwvf4/CcWPlQ+9vvpwXZ
fEN7XLYhjmGbj6nufVwkXIN5gpzYshcK8uay4qDsFtUG8URqaYTeqmv5yJbOPmQQFIF0s2FxyvHS
oP5JgRKONkCeobm0EbOCYBwJIzmhUUxhR+fXIhaROokpnNPtyNga9iiZDzoy4Jo2q1MNsl6U6zCK
8lYJphVrUB+HMGtNYU4IMZKC7j53fJQCmvy7zb7nqpGCbortbGm8aBDzkWZUW0jOddXp3fI96wYE
iKBbkuGJeVVSYmQsGliP2hLNZafzTf+VH74783IJ3TT8Sk6w7+t9oCw3gFAlcgDCZWyeoGVkTAKh
r2M7H79cn3S7uxxL2i7XqEmmooqbFn+6ubI9ZueMSEcTzPI8SpMbWpj35eCn2BUEiFuDeHzgqdwR
A4PKil2BfmVixU79O4fFtwnwZcvomvO1354tB8KZQZ6aZTiOTlqago7yTQG0YtkBwhJ21Ue1+W5p
y31o/kTQtR+88xclCq3eGVnvMBJYo5FMEzAkxWpzR5XNnpFejntQ7YILOYLjB14Wp6qNRqRUPa2a
DLajYeXJew3PJR0HWmR5UCJr4+Cc9WPC0PX0VgkHYNuQwgPNcK+zCXlX41j/pDjbHNxZhb9P+kJW
O4UFAnTDi0RW/6Q8mWxR/wCxddhF6V5+OIy1ELbaFVMSg7o/LGrnwwiNq2pM4oo6ulvM0u2Jou1f
aM5L3FE6iD+NtKM8ggh7FfrM7cHdbZ/JeKqi2cuH8lCo6o7KpbU5ivj5yL21ZGiAeKWBNezsCnaw
anMh1Rc3iH5C6durtbpgjdDrswhn8zse4KRi8HqyezPWYFXRCdusUlHfTy5s5niB+u20Wy61pSYx
pnLBwUaQGm62lc0STcO78QX8HwU8XOsf4BUAA5yZX/Jlm2th1vFPMkf9onjJKrv7lOt6y2U8CNbh
yIu0Q0fC8LKzr8GAEdesXkoK6a+RT9lTlMwU+o/jGnX42nbMtZ0OWJ2UDu846pPQlCdacpP2vlWR
/uyCmB9X9f+3VtKez9wP2aXe/+7Ql/fqTLD0Vn5IZCq8BqOR8KcIb/rHO1fn2BkdVczwXBRr6BdT
oDvCiMQwotx8AwChYIYdDzeY/ifSu+Tdy/magLMbJ/kG3R4/TdiKYBCSX1GChSCwHAjX+MQKP/2A
0DM0AjcIdXf7y45DSgb/mXGVbfNTyJq4rPf+mwDvZsUwpHfdgZv+OIOkAs7ilDy7Gof+sRTOrIdU
s2kI2r8ptGXMjGul+KDqpgig2Xukd/UyRiAzNeFVOmEi6I1hNPajEIvBzaOxxb3mbPnXF/d2/J/W
c4H4m0BEF+P5/GCc+MXb+RYW+db9xIx6j9IhlIpsP1lTv0WGslsc3N8m4Uudiy7dEA5lSWQ7X/DI
K1bBqQwzdXlH3oMDArOQJRfhzfZKQboOUQNfnEjZxRGvALSnFHDl5xBxtRY9GRK3+5wifeAXGwc1
fApQobFwpcVhpPZ8nbms5o1wZZPAfAnH/QF+MH4zUtqS9EOUgBGInzTsFRBKgZY/V4FwN9EUPTxT
QF8harSkL1Q5Ol8XKj92zWVmnlGmrpUuqERtKhxaubNT9UK6P06bAu2b4LYiRa/USJikCN0Z9oAO
bgGwmUjfnMUNKKHxu3twjgZVRbU6hhTnnHgneqXiJ5EiyrIk0vbqCGFN2lqnTW7CJeyPRsNw69d2
yGlGNt70hkndQXRfmoxj/tUl1l/Fyp/xCA9acH4490Xw27bqz5XO5A2WJGHPqSfsLGzyT9s66SP5
mNOYICCa0HMHd9HFIBZL3X7JSv957iJg8k6qOayEMFEkeD7NAN15cMJMm5Idylh5rx/gm7HN4U3/
NcUjpyl399kcygWq66bPxIQloyt6FdyXnrX/4WmKTCh+qDEOh4JGVWREmdK2hGb/sCgGVrJuvkuc
PtUFWVMnL9tUYwvZfGKMnTE2dpLRiFJ9JnwYsthV8hEY6sk3Dl8ZKLXaah4Cj9hWZQzLun14sYlX
lPt4U2Ui9qo1q8qKtPiE+0VcvjD2f4OguSD637ehK7JkBSzFqD+Wv/RF6w7Ynl8GEjbEL+hs2pbM
37nfKbtXVppvLQ+SCdXaZbLlN18uAV4/Cw3Oimpxj7tdS9cl/bCBcG3rlXMkLcKA6JcgzwQP6h4Z
o/5LbVs+elN/LBuaEHrFezNg3vmgLqQIm9Odo5w+18dpCuO1oK9DVJBhmv5aHReb1fkZFjqNamKE
2ZSjL8bx7qKO7+4+DWeq49Qzu64HWMaIo3cmpZQPb4Scx8u8lNGECIcKz6WEiY+8OXdBwnhhmjrF
5zPkiI43+ZWffiz14UFr8rL8jUTlFCPwQOM/s8NPY/FJtH67X0dvTTUMr8AmazPT29Z7bLa0W8rv
OTzCfDqs0g7XWpH7/96jbPCzQbP8fkXMpxgroynHxEBDRlWUAhHgpb2tUDg7e1enTtw1o9XXVrWC
9MccdunagknBZY8Gpys+iU+2b6lQxbdsbYnZfViSv+D1IpBn8tB1jD9JjFwd8a974q5PdMpTnIHR
a0rNIOLorpHpmMwhYFfnnFLIktoHfrwBNYp3kubsVZT8HulfSCKUUn27PR6mgmmcBUH4z0Kmdewu
I//lUclTSVl+xnLE0zOuHeA4/tOyxmi8yW9MyTjV0mL1Vg6ZrsX1hBmL498R1UjYnpC+urBXWD6H
vPHIEzcmqcpYXdJi4r3doJriO/MNKmKFQH1ujGEc+H4LwLYrykmmhy8Nv4ZTN5fKQuPEOLNmoHTp
sA7LX7JkjRoNGtjfhgAqFYwcUgauojj02jCdew/QWfFRY7b744o0XA35lPKLSH790inE7MRekwKZ
uJ/jRw94PpexOFKmQZV4wlHIembZtrV7ZMm0+MICSVLLBF5EAv2+bjFMRqZUp/aCjDt3FFJMqiFD
0Y2llBPGweqS7mjbvQuno20B5Z4bzLbFQvZRqIM+KjnhYYBHDvGhtadU+LOu08zgF1d8R3B2H77A
oHY0ijoq2s1bhP9XdnJCEHcbm1kScapU9tg5xvl0aTFaImxGEU9axjg0cnpKFJ1Xddy/qFBoDERY
q9yIyN38tBaq4fU22kmKMM7nn25E9VH7+wwYmXf1q+iQaUMMkzFM8zZIAWM7NlA88iTC2m5Bdb+C
5YmxZOSJKT7evXmBahqmPYfGTKUDOLLgkRAu+aC76OG/WOwBHUfJuiI2akcB+hGSL1V9hxyZJs/y
2REbehMS+gPdwO9xS8LVckN3cUYp59mPUOuoJS/zWHdue8b/ChQSUCiLWAqLinvFtMIpLCtTmHwI
Pqofai9x6kLgP41AbXvmSuxP/7s4UKNSkUBagqhe1/GX0efK+/NJaadKkPwnMga06GftXTz6P4k0
rikxUQG4FRV1ZMMwoAmh/6yajAeDkABjVflV3z7Xff661FhyeDUjEIEGdskqRAHUruBOZzEEXe+h
CoyfiMzaK4Bu/+7/M/RhZPadIORu9+9qQy+KbWhjBFAkeTII6e3r3YDXGE8QKOhLlttM0ctavi0n
Jx6VH7phTdcjs+6nvbHP1OSevR6SW7PvExxdMmqHDLXvAlymehAGcFxQfgSexyKcSLxniCBlNiEE
TXGqwKqRKxTBaCz+dhnls4ltLyeizGe++bwP2NpouKmVDOfYy2ZlmTL1Ah/nlQMlMQZ98Jaxx+K1
vWbPhWrC9YJccjnHTJbt7IuUHKdXqSg6rZcbbScGHdXuoHduygkQOHTPbYC4qtq0G38Qa6UdWCjF
Ro1kjpYN8bystnaAGy2yuvJFe0vve2T1DCel/ejXlBy/Ra/9hCEhmWsz2B7KjoZyycNUE+Fo7F8R
joOJX9EZrd2Uj8vAdsI8GgVSQHvLArsGoPMzGuzJs0CsnCcspqWkHMCMWz6GdDIEJ2zeRqnizMhQ
ClAH8XwZQw+SRVlDUK6E8z5T5sG4JuYvvR8hNCFJaGDAHo0k+NoVAD1kuKuykZsIXB+GFXnY7WPF
1MKQAZhnqLp8ZPPMDvWibOaru/H97ZXQn5qMLN5PcWVe6AXfUI0xpVtapAEEdjzJfsMb91T4IiRj
oXMYRgZsf3rbvKGKij0wgSSr1hEuGAbCSacaeFQ68jecbAE4+stJDF8we9GpHIsfol48gs2m04If
77ONcM0wnZuPktNw8/O+tVxuacn0iCCsxHU88BG6pOq2z/bIFr442+C9UJJGjIrzF+DdTgC57iqf
N3j+C1TuKF+D1NA3bM6vnM9M0qiHS1GX85Z8OdCSP73+X45NpEcrWmptNuYejVyFFaby2TZ+YgOy
UKKd7+K1h99YcX0oC7g/oGecEEWpUToP3KVl+XhUhLjUnPHH310ik9vrM4B2p7eaY6/WMP7aWAMh
xneix2kRoJWi0OWwFjauPutz7R5YmrcJkTzbELYSV2gfJC8Um3lDNCO096sxODrttVf+8P92XxIf
7DSpsNvcEOKkrVU70hgDUYkuXKI7SWk64LUagF7uLtG1xlQvzx4aOUKwMKl1pe2ABboQVzK8sUs5
5V+fTa2W7lAm0VBsV59ogmH37Awf4OpMuvCMM2D2h84joeOaxxxwKBLbizCysaQruualFlV007El
U7CN1Votj6G3HXCOlP1xDCU72WsFq3/ge9CVAMRQHzkuGcc+T0asrtaq0d6mmd4bfGFpLI8IX39C
0Zj5RNHDCkevM6Z9hW9rfPesjTMetg4VQ3IEpjMgSZyirhP/obqdxephT0vHSEVaqsX61Yw/Dj/L
69UvcxrNI4Dhg2bRAygRxlbDU0/qF2PR35igERQbbfO60Co0LUJ62IJEtS0FyqiaDgl80lu2fV3p
x1Gi/YN8oI52xCgjx98r3FY1sNtuZ+UgUwWIHB+ZMaFNaICE03wamLCoUxmO0EAdqLmOepFcjTJ6
S1LTzH4pVlh56ScCIl+yn/Mu01Kb3v8jLzk/PAW65AHBTIDXODPNecQdOd9mEvLLFyp1LWjh9TFd
xKKMKgSp+lb8Q4SYsJdM8f0mcvJAtgdZIo/ax5J85TDsoH5M7423KHGjw423vehRfQOvvzKboP3D
k6JO8ra2y9WfYA65VAnL3WNrIOOv5vO0GnfolIprR3RluuftgJBoNXvyzooA5qgIrbX1uanxZGLZ
FqROjhkmm4Z1+F9bRRdrJ4fzho2hrG+fmjLlB/IuCXT8/WrN1mTDlDKSTHmM/r/ASSWpE/lSrjA9
RC5rJLKLNZrbbpaQt1SIcLE/7M6nETAN5bFYtRbaGvFhne8ISRw9bX4dj+dOuLwOR9BOJdgZsI0f
dAVTUisudC85oppsebESt7cbsKWl/mR3/b7mD5VYmzLNfzJbkN8Dwbvpj5ed8lPLExEK9jh5IKHz
MXkTE06XJx6u7L74ZrmcDQePvldXmiy7uThOaBsTSuQ/ofbiII5QRAlvwxTFIJNYKpbJxogZs0f4
PzcezKM2aNS5qCwXHg2pCl5IzfuptFShiXSfJY+4DQ4uGz9e542EBd4I8cY0jVZsQy1HPi5YYmAO
xxIYnSMHTODWZPcRch1bK9wzxZBgzMpIJ4PpDu8XvvkbIT0qQZB6qTk8sqSOuDbFNDcCC9SNl2wI
sRE+c71UKK5iYojvdjmlYmPIYVvcPaSPuHtMjex4ySeTtQXMLcNIspW3eFZkgVoRtRM9KlULEeJW
zjdCnhQmAGJAwCzPxn0F6IWwNZplt6V/G3k8scMDyYdbfODT3rB+vKa8rZ2SIco3s6Qy1UmtbZtQ
FkpNAM/NDcVS1tOea550aquxSXW8Dnxp295yULLnr5ZJh84GWfvgzaJo+YJd4zdv4ltTRKdfJsp8
85DB8haJ9uwFMvV6cMi80NVS9TbOaJAh8MvqgVsUgn++2+xCEMB7Y7qHXaSytrqOSvRS3sQXfbyr
bIhu1oGhMMEPpHORshP/4hv28EmdnO8dgso+fNVGFC+hJlTzwQXarKB0JLnbQep0xkFirfFyZ7S4
CjOHau407SgRITd5c3qf22ndWMxyXDyVa6akdywnIi5oqVuqeFj9pc0JyG3Uu2SuiGpIZ9gGelDw
qMGqxb2ArJNttiyljQiQi7QJ+hA7n48XAcCOX0q4teAzf/2vouvVXWE4LH594fd7RDXkGvDCGyEu
ESin/F4y1XTDakeJnOdr2u39E/PTIzsbsFe8yJONoqlgPE2SjqIVOKXrX5wS5MnBhL9uwYxqfSwX
Ov9uSKSTfNNA+Y6P2k8rPntkhcTS7fh+4O5j6zUT9VlpHiNx2YzXRMd5y9QCLzeAzc4GnopQCQ/M
yC8HgC9ZDjmWrqAZ/A+V9qrf26v33cMc9mceAmdVsA91wanaxDHpsoor80FdKyZiKISYCksjzskP
peibf/Kbu50kdk8+WMhXnTI5hor10h/ylF8Yx465ghYRA9w+T8hFb5skHF3VqW6qSrbAt5eVVvdU
cWdUT1ypVBszXpLtHqMQWWuEtH4lwbJy1Qp0LFzVuFp6kmcdTmW5vp5aZqbJjyggdU+z0X7iv4g/
t7Ng6bpTW124eVup0kgWBpS3TNYe13BE9wx59Q70MLy2RoJD4IjI2E/WbBJrCL8WxPan2TkssHLL
oKimXHMuXelsFmWJpSvfhJ35U+l/pEixlzY2wcxWrxtGjKrUTk4NqrpdMBzzX+z1pAA51IlcZyl8
TY3oY1CXdJrlBC4rg0QkoSX/wvaeRtKnTlUCdZYPIid0ol6L4ljXgU2LUdK6LanT0Ju5kpG6UDW2
1eOycUu05d6OXxyb+nwO78scj/Eumvc+9aULw80iZFXFq8Q48XK2/ljTk+cqIiVr1wwhkx6w7YMu
+Z4ZRe/Oean/ey7GdXOkEw6HrHvN1ied3Qd+x1POUZp78X81KcfEVpZAZtVzzDBCvMcFzNPmOxKC
5Q9KIAZl+OIay41efVCcy91PIdlPB4wdjj6mgVIP2gMq5fha1uS4Hv4ufvDMwb+EadqR0vRTcE4Y
A+FU8od+fEKNxadzkGmMLzbjIkaVw/wJ2ivnRT7irmlCoMd+Un+lRtJKkOSnj/GcFo55ntR0D5IJ
Z3Sh9bQQotzU+VK3OZfW6E9WiL9UiEnlfzmTQa81+V8WNkBSskHouafVkCWEm0kmHtin3QHUS5Xj
MKef5XiUB7MZ6vC4bjjGo3YANNzRdFpN3EHYmPZ8Nw8jBcTcpxE7XrtHTaYf7y7v81/urDmzb5bU
z9obVxkqRc2qCEOuuOraaTJziyW8sGr0GLJfYWm7QYzpURncEB4m6sH3usd2MwywuhOLQzknShE5
wj9S6HB3QhTm2ZmyV+0L3IhrRsj/SW0hKcx39U2Szr0HW0jCdEdu7EKZjkg7O3e+Pg59T6WcRXud
OjDBWzI2BoaeCgPJ/aokaMlm94+XaXp2Z67ujclzp8ftF36uZdLS5k0dJQYXGKR4EXzmPs0Fgvop
FkOLG0rg+7VGK1k68sYQw/tO6vKkysn1OrbBpk7H33ORYQzILfyzcdso0TXhrZQi7Ri7oIhKlgy3
523JFc6zx2vYYbKecWpm7Lg5Jn0RBlEBbc+BaIbqNUXU6CAFMJqKmg/9uNEyIXdcWAjsT9GhqQYZ
Rmh3F5OW83gd66IQZ9SDbvvI6EOZTwvRglXRaWuBs9F6tKn5RunRx47aofSQF3/bxCMvG6YYRjPS
l06G4Ux/o4it5UKgN2oqQ016M1A3gU6AEWgylBKE2l5t84c2O+1t8aqBzuTWiCGlcPUxz+IEishU
6BTAWaU22LR2Ad4iEQ1cQhZvoeOiP6aV4nybuZNSA+OO0u/5UoJCxeRn3XcaStNNxRssqduGIlP7
y3fGWpVIT5aGV/Av9xwmRlzT26zimzk0Ss82YmP2U8q5SBeRj4PyiiAVVd1Jh3FOzfA+P2Bv3IT+
mXUrty/ELW5XmISRw71RezpIc9QQXaSF/Fp2Yx/IMD0k/WieROhqai7pjRQiIYKG3R7Mb54Dcj2i
c2T66Jo8rTuuE3utGby42X6pSsx07H2e0dKJAYimAjFIWCHWwk8b5oqK6nrVEmUcjwywbt9+juSa
Rgcu4lyyBJWeYPAv3oVTfgqzkWmxXjbkLDTT9Vwhx6WGfRZnK0DymGyddf5KSBpryLUHUb5rYauR
1ROAT0i5TF1HF75gukzgzdJQsKkwsmj0vxH67BcUI/u4oBP1Q8dr1QkMyA86O5Zo1n4RwnVPHfuv
kIZNDvb3ly8dAMQ1nGTiM85YxANDggjHJamSnkyvxZvylU1ggiW6JvuQUR/XVTw1iX+NHis8PBj2
4FHwe17Vqvz8LeIXW8f4qRdahvsetxi0Z+JtuRavvlRibqyJrLpNWJH7NwEz50pXtZ/07YiYanTE
TmO/9SYYnRIJ4QvXvQzZL4o9uvGTHnjl3CWOW+9AnkiY2X1wHGqyasBCzvv666G5+n3kc9GbvsKO
u4fDlERQKfz3ZKIjzWjt2UaKvp7LSHkVIw4odcXMDH0g6wK4/PVf/6nW8IBzjf4GWgTNSUmmhdIc
RXJl14qra9p8a+ypKi8eBFAUNCDLoV3iUGDz2aNNjq1MqXWThWKrlKb27OrE8518tznEnrOC+haI
rgP9V6KG0HBdHNoGpAQOxhesisZZG1uNXxS6AlDn+fT6+ST30xwfFVFTvY/CuIh93Tjxd7W4sqhw
zhF3y3lFeEEiR7oJJtNN9cgSDboy0caSdsQn0MREE5GtRnwHBChfI0qh94LFtlrbz9fd6deFqM/0
p3GglF7kchzvxFv08oOQOICzkGNJSnjPfvqasra6ii6d3gSzIZeJB8/+krC0yL+SPX5nPC3PZYFT
zLKjcFfjnt1ErkizcaIU8VSB4H/ZHU8SDetECwVhWlL5mKPRl7qTPZZ8w6I69LPEuzeIMnq/ECpG
PL+P4l+UHT5V9OTVtZvxvnFc/W3/xHTXxfFwKHjMdSWrRmUrl/OYG48F4Y5xLekT9Lyjn3MEpRX5
i9o3rKKgCWW43eHGxTyMbDTHbAo/XdqjkT+gQr3WugJ6oub6mVyGVWVskkF5En+9WKWYRRsgmsXc
z3oU9J0NK/90YK/dersI6d/oPtwHq8TxJX9epSKbMz2vnST12xFKp+BkJbfz0yUt4JyFKaqSK/yR
QA2gozwDM7zHhM99j82bi7QoVx9AsnyrFmT78Bi0uy5Ki9gUgjj/bJXkHj8JIgfxdgjPCoOVQ+6l
sgLvFTnIWv2dWHGwFSfn/mCo4eUNGp0MoyqRb/X77MSMpDYffV0kWRYItRuXGy/c+K7JH+37Qn9t
926n06TrFnI4BOhV9FQ9kwj6AXV2qZXNbpPdQBD4uAWUfAfC06cyDEDpj4W96XWRexoqepPz6xSd
90Ps/SZP7w9A2Dj1jwXNSe2hE94OpZJaJ5A+4iTDWPNF8KRvfD6fmbmNgiutawyNNtoxh3FMZcqY
k16gtMTa8oButa6LpgCYEI21/mcCdwDuOia8DQAW54d+UX8DmATFuFboobEfBAKbKw2Nj7HQT8s0
MyoCgx3DDKbymwClfWPVAZHAf/44LmXyP6frW0+DLZcxBxlScRluiUNqOC8tx9nJZ1ExXMn/KvQw
Twc/m5QyQemkD+PR7s51Pp9HcI8leGBP+13c1HVXPUYITeUe57JnJGY/COi8ZqIFvfb3M63IAhhx
LzAEFBCrx/Y1Y8pE06PfANo/3r8zSEjuWGwVk7jAHQSpPnejZ7BUCR0nNZGLl45BAvIfrlYPoPBJ
4pmw2aaO+3iI4+Ui+aofSLjTLxwMI816RkJBXvsaRdAwqp6MNFUStYrWSuzGb0VfLTdOOlHZ40Bs
g04v9tlJTK0B9CbWL0tai5CGpZCY/vm9A2jsxxn3+fig7XVc1tdHsCo4RBAap1bDehcrd12buiNk
tJKakIpQlbKA8aiXHwbWuvS4xwHglmSwR+gOfmawmWqf7jb0qqwuUXIlIjyxzQsDqczDOMPqX5sZ
33xvIUyIMdAFcVvwVbVg057erpguQJUMCducIu9AhEALF14mQZN9BqXN9ycKCQcu1G9ShrnLjvpA
FvNEF9mBj5HvV9IDAPgq8uwwOBnO1O7mN50TqJcfR0u8JSCwqzGbdomI1oBezAd9it68lSGx3AC2
rO89C1XnWuSH+51fxI6MSEliFLoZq1UGcBkESSWQWJkTQveIBsQi8l7RLZw5d93NqLmiCpUUOasd
2xcV9EO0k46ELSCbd2MAkvp72jBtio4ZQZll7W+gefrt05LR/O0f2wk6Vib5leP7HaoVR3pam4Zz
Xv8R8hHGZx28sjH5rnqaD/ZQq6vqa4iRDa+qe2hYT+l9HUr3bo+BFYrxT9KQfqW0SvIvHXvSyWjQ
C6WYT5uTuaUsNjADfLgbKf6BaTR37QesfsziJpyUKHAkgDEY/+fHAxbZkM5WOuwplCT6LSKzjVRA
FW/vXL8eYi7B5lRdNhceqngvhs0TccX5aMBPWIXgH1ydaatySvmLGainZNSGUx0FG9FKOEMK+uuu
1br8t1lnhCuErusJTlVMoCFzuW0fkoxb5PYKhEn2yzCxTJBGsd714lQDBgMaKlIhOXUQgOoKcNrA
mZLkMa+eDbh74xjbiTsTrhwHZNIML4cGghqlg+knfQ/FO3eGR7KkRvaGI5J1NANqLMbNgezQQKM+
mMylsfoN4TNcVqLcyHbmMj8n53ZnRkO2MBJfEs5lkTymtNv6qMMBmPAnj3C0INP/olGBePaMiGhl
LyJ7fZWuF9UPwzjPqe4TelauEf/tOcj9xdAOOjAryzjD13IabLdUrsTXdQLFIqNQ6z4s4GdPp/gT
ue26rMNowIk2vk3SmDe/hLzSqVIQO6DoXrZEI17Xmy62oVwimrd2YnLBYQmp4x95Iq+eyzS8B2uF
3PIk08EDz9n15fFITVrKwJCjK9RCERIdWmn9SJ0+T9Jz0Ts3GNMpBJcwVcRDfs6QRmrwQkK7REb7
kld0664OngpUxdJWyQ19wpPyIl9OjdQRyeIdqY10D4ITsx8DaF4YmC9l3It3T6ajJQwbmjh1v/Sp
j8iCL9t2QEs2v9Fe1CPlnQjawo5ZCynAFITf48ll0dhWIAfzN51hn/3pktYNEUw6Z+89hv2PTram
BRxFPmxLo4Q0akFAmB3lhhM2rfvuvVDDY57cErAF7OOgC5eLwRQwUXw+QYCmDfCNbJ11HXcXCzPr
4H67Bb9dItAa7hR3/H+qBnbcxoM0enMPg60GNduNVDccqylYhZ4geuxVBt28i3rJtqK9uFxNGppY
Rc4VFmSQ8sFZf6mR9XML/5QbFI6waGn1YrYF91bcdRpyzGpFb2smO2Iz9148K2hrPucgh/Xd9Jle
6bCAllZ0/WyjM3fvwdZSho9Bz4sKwOulsYNSF14R5n1dj63T2FU6cC6tQawNbsNlZtQLLVuGA+Ic
RnTRatVt4HPoAzDrL1Knjwo2cEpEOre4PaCjKzwdrN8DLyJCW3TMqBq0Db6tJghnMMgbi6MIeWhf
nbhAtKpWqNb1CpL9FAB9lbOU0JdBob+B6XfvXClk6hy503vTHAUjGK9noGzwzRvguVqEJKUMfJG0
GqwFFbTNI2Hxxfal8tRKhjCnLThttR0QvFv3zUai80Q4zt5okzWXutivsSodytWw7J/M2b8Gu9Hv
246dL3W/P1oUv3y8tC+j3voUr6sSZOu0jwVgu1fCevr2sVHylxhG4JeZy941xWzS8E1Two5h51M4
ACVF8/XElPAwF0T2UUsf/rrjwgGliLzW65yLSxDuwHldXQ73PaaWF5Qi00upNYJ6VxU13f8tiZdk
z3ORFMsUQaeX/+Gn+asM0Qg9nrppmo8Zdt2S8pL9ruFcuquKObE6y9LTJjWXaETYqI1WGpTOgzdr
HfsZYuVxfk503HigxcXo0quftEOZxg6U0xTZbWODKywkGBE9rVbkrYvgSfOWYxmYNWVGNKuQfrnQ
q9JIT6E+pcW19imN3TK9BkGYVFuCuMPZ6mJicJDgQxxNSdbsXbA/6oskWaSkC4NztVOYxBZWMayX
C4r9QaQL90oXlLKL9BD19dr5bqybvK6chF06909NY/Ks4zLKdVy3wiIJ1Q/wSVTIQJyqBT9HnNVd
MvmpO91tv2kgRBiDpCYJ19LE5JhpMK6Q0WGV/4igjt8qwUixXdvmGXx1N+uPqL5BB1KXU5H0kyIl
rm+JFE5P9q/WLRpDlbpJ6yvJ3LoZ+s8XuIY293AloBcQXGVDNgiy2aCDIDdGW68tHo3gXVTDedbv
RuU9c2Q0tiZUlYbT59Ja6C6c83hoUBnLNgzeoO4NnHkFivua5blisNfGSSwXBP8F5n13a5D574UH
8XbPZyRf8Vj+/+hpmp7ocYw6IhkLj9g7CCsq7fYMNINwN/01aFTMDEwTq/3jQbymbA5AoQkF9wyR
cmdWDajInbHwqzRkUcVsjLbZb3Ufuolzlga2vdnV8SSSnC0hApaIsJNRqgJ8M/23kB7aCgfZm4h/
zfYo7ThMjHl9vxZV4r4HgBBE8Q9DTVimqFWNmKQWAGg8hAqtZlJYFTEZstIe1KzLuySmby8RdKva
FNjHEyoYAo+4lIrPLRlOMn26zJ59cc63rGitvRtiN5cg2mwRNlTU1eznrdGVHCzDg18j9P4gpITo
Q2g4TGSNqJDqgCsOBE5xmhkzP9BRIdJk6NIypMQ1l8/CT1sx664XpMj6tCaj7vyDqyDra651eufZ
WMC0Ya66c6ZXmEG2fiUUfGDsFAn44n3A7hn/ppYIiyatim5Udi/T45KKLr4NimSVkYa3XdZmPO5h
mZKhXnU9wrFPx5E3Df0VWXj6v9CGZcOhB+mxsDB3ADvXGYh41s3vmkEUYSVV0b8EAj9p9ZGFCWA3
HoNxy83tak/hgp8SawDEOIUG+gbYWzBpEknAzZw0AFW0qjyp9QQJQPOsy8uRlrL1kwd0HT/w/qRx
1UUICxyZUyZ6seh7Q5/XRnkFcznLYx7izDYNcoP+/2HuNS5Y9AKqNlc5IPoQavwIXEmsLNaqf4zk
n5o1/BT7f64nHuQ5GU5zrCjFpRcfSA5gAKCExS5S2uHWbPEGbwtDJZ9MJ4JYCovxWEPKW+rVI9wI
NMdIBsfnkD25Yev+Gtne6zvtPqU2UKu9tlkKtCoQj1ZOtRKbymBbfYmNy9LrmJqUBVX7GkSv5DKg
PJHEw4wasyUQFyD/9Tf+eGIWDInjKCuRHk9GPTI9gtgqoRcFmJ4gwGuh6uf/vxSCZnQX66MjwS7d
3dPNzkli6cmeKRWXMR+R3sNdwXNgZ086+pz2gDldVFN9GcsSPy0bsPOVE/wJ85syCSk/Zn/5VACd
Jmh6xL2IixnKXMNlsKLp5bRKBfQpRF5S2GNhC7Vz3kPqTscBlm3+LUwnh92YSc7CQmT/IJXAfWJO
EqA9O65yG2rPCcr/+U05kFdopEdoGeMlB2phhXwJA4yjm1MPROlbZmm7mSWeI9543YK/z88zg8tg
1SBPT9r9pc8Twib5llrcHfe18A8Wia8wH5EUOfAhhhzxgLQeXe9v9UMnGWjd6HrHPyDDdlWlutwm
Z3axerXmBHayq5gKwtfUea+TH3eAGhApa4mU7u5MlLsggwTAXseZb5heoerbZSbDlBDxLJsf+TGz
ti+WKDOvSoTY59YdMaT+ggx7xy0xpwPghYzbdJHvyRnOF5GPtl8Zn9F2alVrgBtNrDj+4+VffaTD
02kWrYmlyoVo97Ij4reGhR6QIYi5UXlWFfu00qJ0+EvmfXVqy+OMoTFwoCdsotGoYv194nrmkWM8
HBsR7R3ixxxp5maWSMXZyM9gdqwTS7evZCurSlUok1dsXKRo5nxdlI+pNOgVcgFqD8RjlXa/O6bM
U6CXAACBVCHfPo8hbX9NZ1sq/Ldcf12/mC3iqdlx8O4rMs3qbNAARM/jtqihaEkA8Ogi24GpWzH7
X8RAgKGLBDClZ7kOpM7OxhzAg8zs27jsR7yrQqsiFCDKj7Kt7tC0kcLnlWncBoyQodsQQ2oY4VSS
VlIi8aCqi1vZPEMAP2Tvrj2MrrHJe9r6EWIDRFoyJB2kEQ0TpxN8rVUYiYU+CXMk+AsziPLpMmZi
31BupfRkNwpm6XeKOlW2ETNzJRhe8gPK02TA1S5BmLeFnQj5PuGDhOI9egPqRuORWCqB8TPzsGgz
j/rdwao7aXuJ7hZSxmmeORh6nMZtw3V/v7hKkn4TJe4YQmJbpAOL1KvO1cvz02VdQMPXAzKWXnuk
mceuOoGCYqhOCs2GiRBvZJcs0uirkvW66XO9keUrLXzeZvupe6yaXdFLQbPTIhIcKIDjsncChCIf
JUyrDwl63FVUFT31NQtEYlfZ/uP/52dylwqIJ6Faovo/YaeKLOZjORjg6UqdqIkwD6LFVVExQv+j
iuZ4Og+ClAKMphx6llWHUOOujn5/4T+sNElMxc64GalABPCQKDlA0BcQp88ZZWRHMBshm4XplfX5
vbnJCgfFJJ7Cc3AB2VgGMV9ZE14RghgPOvgteoiJZA8O/W8j85/JyoSRTU22ARWVdjncRt7S72z3
SbuzzzG9oqdpm3eOBUzt6D0Ph3p2Dthbct0QeQ+6yb1cDMF6RteutwtWzjEQkJqOmwrc7Mi6kMqn
zUyn49nzpNpBx43mrIuqx8oMz037cwkmKl3y0CCfO5JskblzDvbzK4W0yLozCz0Q2bdIPf7kLKuW
DzmnwQ6lzrzPyZlea5RfJlTw8s+jahKe6S0N6CHSq9/I0U7YFoHVqbTHvtRrXlqE4SjVhKYeT7uN
lzM80o88HmRUPBLLnDzCzxVQhmDEmQZn8/18Qb2aaz5OnrPFPmvmAyEfFVRXU5JfYYL0sg+PCiT6
7wUB9E8Uy6wtKQljHySAzZS2C68B+JMtYDHaPPyW7lE6d03fQtSgnDXkOuFaNuvuU3Oi91Y6u6LT
SE2nQUdx+xmvUOBTpNB5PBtvY9chzKxkOoItKZkvxtAfoL9ApqsHFsoEOaaetTTTOGt55M7kL3qj
Xi862YIOigR/yqCuPHZLL6fxBN7uWlN0a9cdoWIaPMGRGHf26hgrmInl6uyboLyd6Y+rMDb7NT+I
clcJsfCXJuruVSd+84oxQb3i34fODja8wSS4FAYwKzCw5MHXSuJ3wGjEMrSEhP8YWlWNdKHS2MTn
XO2k1B4CfmsanOJoRqhE8L6/tjNz/geMcBUxyafHotFZQZE+rDCTWx33BZzfFNWNmqwXLeU9K7Wz
RwOmEyPkX0B0V9FOo+jYN1ph9/m6zM/dxKYo0UARox7o2sui0m3Ub6u0XDMwgnK0xAVQMc+4ZjLl
hfqWUANnPJkRXIPHfzTjGbOtsXqMoX1EIp3ZM+SsJM74aKWSrvZhwf9q+qgPeHNO8I0+EIwNEGag
wLUutrtUffLCzbpFh4OZntmTitnjOJB/F6zGf/dDlm6pS5qL0JCXcv3PQdLfOZYnSUCAE+0NNgfJ
aSkuQ8wOwn4KrRZ04voAtODrYdept1mYySkO1v+PeSPYGTSBojmgcUgq9Jwrx7F13gcHd6tGz79x
Gbey+qpg4ggOejrr49Euf3gbuXU87OopoEpQvpt1ad49+woIhlznFud3NG6rmGrvCRqm4kIy4xAz
JD9q4yodB7+qRLgM1JGHLr1nkWS77rcd7ovuIixFn++IldF5Pz50Y3njd/NkkrtgkVmSR3bUtVLm
/+YJe5ugbvXzjXABnSn3rYOWvbdmBTLeHSjGQ1b1SHNC1A3rasx0lgq7b5wvFOqKBq8uqbvASBaj
nPpSETm1ZdLbo7kaJhH7A2jvMJeg/uM1DKODFaZf86PlT5u/iAw9XfdgPgq/guRVqQlGODVj08FP
TZ6g3NLUI5usXFYm7YuATpdTs4HFqY6VX64BOozrcuvGYnL0zvbYgRz5LbeJ6XKthYfTSHN7MWyo
y4k9m3kG/x+LzGm1GIP6oT9x9k6nKf8a1zh5rpxCdl2b0uA2ENnG8kTkrIszhdrzYpjTiR0vdpt8
mIbB3EhXjR0N5ajxnq/YPyNS8VoeQLW4sNJw9b4IgqLwX49y+0AHkDrJqECxbDIYVzQc4RArjopX
ETvu95lO8w85seqR7oTyswrvLu0MOEVviTsxKe33frY+by25pIb4Y43f7ILxi3reN8A/iu30Mv5z
MnWmB6vQZT7hoQa9++DWne00PflJluaG8nzC/81DDdM0ZqPTtgqI/QscR9iq1iuUOX8aEOcIpQad
JGxbEbz2L3C6D8JbixR8aQk8IvF6v0LlOrJF3SrPKgysreFETWX1nfyArRPPav6nnD/4+L0PSCOH
tUykrmGVkxFLbuO5FWGp8d3wnfVLWpUSuuTpQdyLI51ZCAu9LRDn2WbmSlyQsHazA81qUBFeUE/+
0SBN1/6L8G+t6ZAmWhnkWAelsmH9+gqYk8wsqSdRHKaRs23ul8oeHzqdqY0VGpo+4puOssYtlS9E
B0d+GgGBI5Mwt2K5jCzRblkyVfte7jYtFZU4bA5UTxUulakib15zq5tJE8B8T3KgxYBcLnuksSGa
iIM0NVJSaR/836YQdIzaGys2v8zL8wcjG2GsOqz9R7fD9Vp9X+qeA4nIzNciDW+0Vl+Bbkykgj5B
XFNaL3i6YsCc1rAwZzA1jiheTjewdgfDlRouD2XeMAz2uMW87zk9MCbHyfocL+9gsbibl4dpsWTy
k36KakRaE+6HN4WIEkjBfYBqO6xl4hnXW3iERS2/jUbA8/urKr7D55Wiq2ljmdUHlNyu1n64siIc
oAet7vZDO8roPjqEbzjlWURFNXHCsI1MCE7jbuzk8qfqWNlMre8x523CqbDeJdwdx8Q6QoubpVZx
X8jX3olnFx8VgAfjZLB4+b3aywab2iGWojtY0tQga7hT0myWPUFudlFuhMk9kHkuaKzB+YtVSqQD
L5KJ+38nKCRuWENaoAJ9FDBFQatZdM8+QwHTDn3LOESAg76AUf2JmWXN0q5jm7Qfig0u8NIzXUyV
EdlLw9rYHx3Q+YnVJ324PoE0RoAFV00uZjeAoj3fWg1FgIpl3TgstJO2HOWd9hZUedRGEZbX4ZsE
C6nzGEVOyl6nt5KBo28/cNB/s+jUhUb/+PtbF7vTJTg+kxerOvEJVhG4m+ZUyE8sSY1UqbdVbcDa
cleRME/HTd0z7IOnHZFz81SS8KuFt9tLSAup/ca5qYJljI3eGi67vZ4nOTQ2PqBLbKuwVPQB2/k3
GRCfplwlFEGWqUdxcBDot8XaAZ9v01XHrQAdxDh84FTYNnHpOv9Za7f5h/PPh226PP5T5sfaohFQ
sM11jMAiafMU317jTncAjYFCQS5ug6NwNPmBYGyaT1807Sd8+c2bM2O0iOdKTdAb46mxDHO2PdZQ
4tAIukSA1qI78d0AE2Zj3XLUA+fgRAEN/sB/+jwdNJsH381StNROvt+09sTNaiHcoi4Db9soCDKL
280R4Uyy6010yDoz0dIw2INA5KPmVnZEtiGjpIwyxR4a7gX6TBb4GVEqtqJtDkELLlp1QN3GzRBA
MsHhli64gz4kOgF+nNk/HFbptKtwlXACLL8hzLKhaSqJjVVJIyKAjOw5sPzn7MCRxU7FHSGTzY+e
o8ivtny1+F/ljdoNKnvfai86SWNBOTSMyoRlGHFtkIlzlqp+FyxbTDbF8amcXSM0rwek2vO24UOD
GEvS251YqnYweSgJfdhEv2Pnz85+F+h5MZQWTKocjQ1s7XKdtYpzl7jNxpuzHk3K6ndwIZEvuEGH
u1JRF8/TfOK90T3/TOnVvuIKD38hsbFegbFk5oicicZMzQbn4zlWxsMwe4duxJMRAokmAC9HZYFg
rAl6nzCd6FQgEmjA0WlnP4P0QmfdwoGVu/MhyJ5oIoYomVPnF90+xmStSV8Zli1r5ZiHIZBI07qk
lHz/DyMmGc9HAkptZDDCiL0fx5fmnFzMxRh/fRH0Zxh1azATDXzGiTHIF06IeYRm3XcKrYbDNH6d
6bY+wp8UKVZBvLXV3DG+NIkY6x1jFhr2lzmjFl56U4o7qqgUAihwoF/4RKlgFysLRbUauxVNZhvn
6hdEEnu78VBkaWgn7OHWnsrt6d0QV8adP7yncUTDgHMpzkd2LRWC0Dk0eKAdIFKxxnP08QmG46YU
+6DoY17/Vn67gPqQWWt2F/HG2baFRv9f2Nu4O5y2u8/9FMo8EXnE+u/aBBqzBf9gEcOI3ZZ7W1n6
xIKaczJrKvufO7PHuOpA7YyyPHsYQax3xJyO1FFRzFcpM16qxiXZkuJlCnve7cXQfxV+TSDFZvBm
S2dKZthuj3fLyCWW6orba/x/jElgf+HhbR6xc6U7GqLMrNYR1OoIPE5ObpV76F6a7rnGDFtz0Ajv
K740yVoyUB67CH71Ho6OIcOBKR43ggFJjDiE520OkkQWzsJsm1uH9dhZP009yc/z2/G9a3HyjREm
ogATlq0Gtwgjfv6Ct36FP1qC7DzgFH0lF9aFfRBDAhNDmPe2yd88VDKbZ4vqzasv5BXAksqIxB9f
9lLPyWOtWMZLn3M6kAtbYh0JnO8+PAxdkuClsmVBH52zPgettK2J3MtTi9AcJWKFDCVdYzbxEpBI
BwJbXctkJ7K7Wk9hVZh0vIL0fTEarxvMEYpQz8FLxmEfzfPBKNXwAKhjfUHRSz/0i+jzBptZIsu2
6mTfDDPPYK1vr6afnHQLkUKuOorUKwsxVx8hewcltJgQtlhvz1SDVT5z9d2tXivdJGm4AOhWTudt
G4pzxhvkjRexump2bLWMVDd/hVh4WmpjU7tZ+gEZ/ocqpEx+EmPcmQHf1HwWHYPieFEpj3Hpil4N
ZWmIRD8uJ2tOEAV0Y8O3duUo+QbI7RR6d89fE8dCsV2q7oryqzyUI9nYvlEMdEgXMz6eBUcC7+fR
eSOHsCtzb58IsmZ8W1DWMEMB04UEkX0f0n2cTKSXsUcqvI1d/zHtJ2GMDjJBlhfauaCtGkOLOFsy
hvgxCYyeaSUHaxREAw9LFIsxR9romVB942wPB8MIZlKHAa5AjSkN/3rf3fmpwqCgQj4dfuRpTtil
S2uUnhiX1cI00XUi1PkxxSygjgNDZ5qpCo14cIJSL4Gv+IIJDBtai3vA3bJd676yQ2OhG4r4CIhj
HrJUMTGXnS2833Q5lZ+/E4swux9o3l9xUmO7Zut5i58g/125mVDOxznxat8I0QKoYDf6JNXAmYYK
rq8FpMFxEpuk/x6kRozrv3Sjw42P4ZFh1FoGk2atc9MnutmGWJ2ieY//WwzJbs1IKX5wys//z+Jj
Pu+logdBU182kqvrMJd6EzM53c+Voeo85H344vtaPHqXQE7/RoFzvKPaJHSeM3nAfhBl/V6BJXM2
txJLyf55F2iWsF8JnLiPpWFholk55jcitsG7YbstV9GmczBKTKZx89uNwtsL5AS6geQS6yob2z0a
j+GFnSyZacqem/jKW/GHCA5ZpWLPgrGZCAtNKItAltNtXErHKLvda2d2VGpMKQLxx0SD+1kBF66z
nTG35M2WruF1RcjdA4ogO8oSyQdINlecxbg2mhy9lCmOw3mrNM/gf0JOPtSUUVeuFOiIyggZG+ZA
nWukZL8bE5t5BEE1zKggUdsHBqi1jXkrT6KCB1v36qQzCjBV7/5Rcn9MA70QHXAloHbRn1ShuvCw
YoZUw5Rj6dMwOrxJWDPQ/a+XV1n5cmxx+pKMlYoDHzxPFRqewmS7LLXxHYKKAUgf9bcpDkftYh3V
uUhHgqywO69sJAG6DtziUWZB+tXSywWX3sNWWi9P/NIgIo21do8bJUb7IXdhWIEv+GnCNmXHGx21
qrYt5BenTsblJ0ynF7n/X5D3CtNOCgUJP6zElpiWAmhGvwXJ/d8mVDU+YRGeoga+u3UZ4zNU0fy5
yp2QZrs0I/XsYBMg5ixrMgi+oVIr7Rbuu0mO/8e4SLXh0PlQT8Dx6r6EwoxGyXbDbKBVerv5vNtB
P/XcI0dfUQte125/euNxMNT10QxfEw0k0iU7XtkFM3cCkpTE2SPXRHO+eLCCZtA2n4rjpvnRoPim
E1xj6vNXrvHzP8GZnZZg0PaZK94zQ6fF0c/KPrM1sZM0//xvBFdC9UgBWPyRjEqR5D1aJEzhpET6
e/BwKvj1/FySTVVf4qVIG4kN8iFbaD2Y0K5YUOeCmyx8wv79hzlxJmRob2OnV/9IdlStJCb9YYWZ
ztWtu7KuO7L2n1wq9+UStkmadqbGaTwhtWfAy0XgvAtxOi6Oh+mAhvjkEVsLZMmmqyzIqlWtz1XM
aSSjC+H5Pv0sohJ3r2yJ19OJhG8Pb9SHCJrYWiIRuEu+NlbcoZrA0QSgXFgOhVTW79fN1H7YfKeb
eTUeO6rqj1IrrW6L8molmDrfM3bD1POAInP6kt9GtZlGUWatPI+yb5UYx0g3dGF4/H1jR/wDuIro
AWFVZe6Q2m4kWwpswJY6LBQYtQqCJjmmJJlr15r3dPQuSWjPMxP++wsqmt3IZsWP6HuEy0rotcym
3/Kr3rafQ9nmPaPUJBH2FgdYrlPDMx0WJVIvSEaRN9LH8vP0VkAhdZKn/f+Q4bpXrzD59qA5RS9t
3cwHNhT5kw+JG0iO5r+A9lvPCDGAZCtioO3rW1ddrKykVqGE/x9NUwg0pGxSEXEwWiG3P3gj4GlV
ueQSKZ3D6iaQAlAji2i9xPpg0oQ4VAjKM5xyseIaSBL3lSVQE9l91jGdhfnSXyrhEcpmfNKk0tdl
5oGUQYr9xtGnUMPpzA3nGnGbEEvmi+CpA6gslKXZ5OeYVcLflu33i32T9kXfQDHwx6AtOLuX/w6K
EDJTBukjh+Ru9aLl3hjEe1xqJUxsUjxJN6vU9ADQ/f4O8OAV5NbbWbFgP7ma+OawU+jDWErxRevT
GFTtWEh4Volsk0ovcy0Qh6VhiVcFgk+UbWNuRXaoyb41AG1avBJNhbL7YfeEos7SfFFAoJ43feR8
ECggEIzLMBPXEHq7QSjbkChFevoK/XmKeYCDbY3L4+BxZg7/uCC2sgSFFw8R8c4Ij4qbKZ/2CCO0
qXoFJIuwe6S7/p26jSBH13jA/t4HtyFOFOWFOeNJNry/JPU9c6SY/r0YBUE48Wsz31Qw8wUuiDrT
8qFg+5HBia8ST5S8BItpRCPQ7jbfrb9p7XPu627Rw6jAqC6LCqeQzRHnOVfXGdm7L2oicFSkSGmL
ib3y+FIHwQEyKPMkobw/+j/nG1bqxHsmQdmO0XXYK90WQXwuegiiWju8520OF3vYv0iwpWU5KST8
HMWU3/zdAOjlfDh7yE0US/pe/ix+2nhklrYvQIhQHujINgoL8lXRGwMo6Ku3eeKqGTX/N5tOtPTT
nTdHJf070MIzj1gU+JNVJ3bx7p/uPKUkeyr5fsZEG8FM9QAH6b3wJv6w9lunXQyh4/Xc1hBGfSJZ
PhuotI8UxTyOFDbTBxG+on5ZaZwMb76mjmnYnv2E9iN5UqjYCCfzsxLlmxskjm7x4/EQq/Lv92Ca
SxTSVlGQQI1nEvSmHk9f1S0JskOtV4OKj8E4YXbKEYN44nQi4ln4lUoyWezqbQVPPOGREn1pcneB
sa553FJD9Gawjr/5fig5VXsi7lWES2Cl3TUIGJYKNfy+0/xrJCCGUd5D50ZW5AOThicvTmaPKOeL
GhPps7gi3JfDH96tRlwKRi+y2DPB0SqviI4PZ8GgBWZxT/5ogPVhNpO2bOpNLaHDuzqlAQorMapJ
zLaANsE2YYYcv/HykDdCo9kiQ9xNWbg9Et8AjTh0/KH11LnJn9VHIfgt5yOhaymu/i8GokaLeIRr
5kvdTLYyQvCH0rjg07f2dW+MI90ij0jESDh4zRUm7+if672JkpNcatEDvokqyGkTlCbFzmBQb7eZ
5y7lfgMuShzitIHUqpmtuan+vE6ugMLHQf91cGe6tNF50R3tp1ornhAvUsalSIsVgvJcD604WOqV
6DtxJHCpzhIT84e4Fvje5XGgQsY483XCmR0A96TqcEYL4vCEq0k93J2RiWBGdlGZAZ1Nk4PBaQlw
SiVx89Nfi684pBvt5XPUiUub7/4Wwvphg3zT0TH79efcLne0Z00m1YfVLW/jCHzLmQbToGGq56Wv
gcKZUesPdB6wBRvy8geOK1tFIEy9oYBay6knKQyOK7eosp32zNY1W5abLXbDHJsccOTPDePmCwG8
BQPr03BMcIrWyGyOzYvDI8hm7+IrGf9d1BdYWxk+mmaYa7qp2Ou3CWBZCWIAYM0DIwN0t0J6JfvD
48M80IckIA+TfK3jGmAhglk5qpYB6nIf1zoCqeXzX0wcCrYR+I2EQu4pK7E/pwC06LyWgjqtNCGP
klsRHcyA21M4z9v4u7rvkSe5SFZNCZQCSPDpaxi228K5pLFqStQUK8yW49UJasP/a8Z/GWbh7+db
PknVYwe/XumxUT/9FdgsPERVF7CTofLG7hfaacXT/WdNe1FrqH5iGW8fCnU4oU4G3E69FqsMNtY6
apOl7Q3sK1iAcrlyblt+5oua+g97kC+ZhCug7NwINlOCQkUD0/qL5mhAahxurP5tWm8web0cEarM
JysmyZtcdXIv68JOA6gQFJF1aZSP2FFp8PNL//DkcLifKyINCS9hP3iSGb6F4mT6+5PMNZq8IOcX
yHgNrUGALZF9qzKJV7EkPR4nmewWlhcEtWa6rm+y4k8r3R1/7qyCKnmwcJuHWK1FmNati7Teo07A
xLUdsid3A6ToHqQqJevp28zhgzSCAP6AJ9rMcB9l15G9WqcP6mHYgncpSf8RFMuOstcPWyH8mh5V
sXpqlmn5IRCSdvQwFyw/OmlvsZ3t1n2Jo+G4axT3pmzSEkGgC4NRBaxjWXIQqYUIatiexPRm/AuB
T34Orjpy7zRIwuA5QPgcGzXI/+ht4+JVWPgQqHL/LZagVpPUdvaM6taWrlaT1WZflVO/6Nn6cBag
OPcfAa8QNoqFYGCBCz0AadADAynYoIr1Mb8RPrgD+B2fsp87NfJUMN53fG0K8yLECUHUz+Hy4uQP
2TR7KfweJ8SLORPIsutgMYwpeTGjoZeA5eLAvLzMUZfwFmG0b46w0EM3wTQOePZ6Wr+FmVWs/44V
aoWB9AtyWiZjZ7Mt6HrLkn3ahMZnyLHOuwKflqbptWxsNWT2I2MvIt8Hk2oPrB/1BbAy1Q5rh0Fx
YspyVwH3JbQ+s7zgb1b4yTrxzCP/eTv55/SA71WFJR92RSq0bJK9RcHWbxMjq9AwG74AYxoi8KLz
4K4oG4ZjrsiZtcuKZGIQdepy8V5nNEEOv7fgurxWaOEgvV4S9HvOYLcCjkfWLFUcY9403OGc5MOh
bb37tC4xNF1ZlgXPu1RWs7bgjCOSJYF23T5ofEaARFi9zQt2LtfTwZkcpjjxB6AuDhAv6QegheSr
QEgS0PpVtzkFu+ue3bCqB4dTsLxCQ9T5V+USJ2utlsD1ZFk95arVlIYpa8lG8QqAqscf0LIumh0+
zwr6dWfstDOfa0BVY8xZtj4tZXfQV8RK+EBA9xL8ok2pmuqRXLNI2Wz+K3ZUCJfM8nNz7Z1huzI5
h7O0/fLgYqpH0ju42o5SrE4n62+8/qDOXwYzBIKl0RcvW3Nf3iaWMb0xd84YgU6Rxn9zC+G/90xi
YURZX3PvTJonRb7hGOEPGF0Tgy95P0cN0dNHvz/F7fbgnX0i4KpdpWJVEiave2WXgcptba/jo5WS
O8/XRXEsfjLWxbyFrmXtPlLKeuhAzYoHZDYFdair/5ZfRYfRVB4+MvFSmCJ6SoBOz/hxtwKmDmjw
fwX7UaHEzGXswJUxZOn2M8fJ/pf1h4YS/XB0dXrImHV28xgx+Wk1cSrWlpsDuu6R+sWlPUM3bHwP
HXZjfZAmKhb55WlqkGItpK2ud6XzWWieFsFyqqZOpt8VU4Njs+9+6wDT/rhxZCJcoNkyfbiwTcZI
L0Ke3kxb4HZ/670jkAo5dfUoKcFMEswP6ac7eAEZ2kUZG8tfhRJ6w4BjiJkfz0ofoUlbbRpzC5Gx
FiSJsoenkwNgeGcM2CUw+Ljt4KpK7iGXC+znbR7TBIW4aIYmQZ5SfPpMr0ovJcfbDYT7ckOaJTMa
peC58quddKDuWn7FxeiMFlqT4Xti+V+XCk8wsfwOMz9DhGSaPZthPTtQ8f7efs+4uTy3B4wijmY5
tpkKup2QPF/asLeZEdUVSuTwcd1NqQa7gf+gIrU9su9Cpz4dZhPVEEb8kEHCBSeLqklwcSwaLg6I
trBiha19Qhka7jdep3iow54f1Pu0ane3Fyx2upGsKhJHNMKy62bCulWEq80oSCZDJryuR3d3EpBU
tweVPrXOjCaM50X7uP5FkXKELGD/TrcNYrhAmOFicYoMELE1PA4FZv8Bh+iqRwjOYKJVrNwrSZzr
NA5w/hgt44wYBeuOwCek+SQmIpgkZ69zo1luOzfXZNYWwaSXpzQXYcmEmGdN5eAGxxogBCGd/01k
i+s+htob4otEA0/yaVfr3DWzQTMjr/LDeJf9d6uaQ4qUIQx2VGMYpmWrvRabx/xsSbMglXs1LDsM
pb9gTz3smyUHPVi6vSIdWo81SLyEe8EYnavLhpe3V8w17d1HW+SceAPqIkJzdNBYXbKizMoibJ9s
caMVgc/RDDmyci1Mlg7+R3AvIcIqu7y+wFTYYh5Xe4rhwu6bjwlGSM8sNzb5vcAr0YCnrCL51vDt
PzntMKFID1epYUZEV65bHP/JX3NQmOJ+GJfmqiI+/R8WUv2CrnUMuDoSnTD5acXNzlb72MeDjefZ
cBAvB1uMpHrlESHcIPqLGd9LotRTRZGvNlNTSwH8KA2wUuyda50h0BNhAC+OnOHbrrB9pzy3iKus
FOn7J6jmftExQIxJub8araUAl20uMp0KjPgpp1mTS1ZMNW6/F3dVqyrzVKVgw7Tth2oltKmlE4Iq
BsudlmRh6a4TwK7k8/gsQU/s9u46AslRRVHWSeJi4/XtXAS94XEuJbueF/6I38udp+VmLH/eDYaU
IanpMO8PfQVtvtydwM5tjFowzrB/sHXyI6+KJXz/aZwujMtcTISrAK+ERVLhepx/t2i2BghP1jFb
9pvVVt2o3/NcI/n1fKtfR5ASU2Tbs3dqDzrYCOg1YZbwzZx9gq0yOIBCQYHLsllJVPvFkU0LLK5d
Id/ZkdwpExo0TSzMuFUGEXfLA3rdboOC60p3uP6ZwBr8LIwzgSQ93lCez8fON5jgnTqiDKx/8eFp
3EjbGbMrmXdgyX5Itu3UrDk9NyqRJsSb+hPEhVkF3XazJkx/1AOSgD54voaUlSwgrpZoH9BLSJZU
LVJbi2W4gYO5+Lz/2gTNGvTra/H/wIKf9K5F9fh388sP1AE3atI8akbIOadSJk9a9RjjmGrOV8PD
HwdO6JAwNjWv6/LkEwmI4EUSPpXetbqAygLHd5DmJfUH7FHmQU8wv+13nX6b1RPQOrB/NgafVE0x
w0MZojmZ9bH8ZJ4ZK1+oCiM4+qF3plQt2+s23sPmMWHvjwUM74K00hRUbIGBzgYxsyPkXLBaWpmC
qvcEtriIOJ2LfSfEhLCiE3PE5jm7zqQW4RYj0fIcmaV+rBaOeI4+rCbWRxl0lJeQCCezWWvCSrRh
zrIbnKR4bAE+CbukcErAOwC9PrVSIpMcEJymO02DuOWmbOBCsbt6O3Dc5UD3LrOFLMgybRTtmmlX
fkOSlV3tnexAZW6vx0lsIRXUuPdQy44pjsyze7zoWCd2OWZLbFLFfd8/TpN8JMfYgACv4AK6EagL
bl3am72h9+q2eXPysujTEEpCP3gzszd1byg98rWucXdckfBWzxO6EhVsNKocVKNXEWz7fDP7AVY4
BcuwzxLS4ieTa/CYPrs5ncD3Vjnajw4S8ZbN3wzsBIDhFlXS4z6yXHMkEchqxl39IkUeIoXS5RSy
mPywFvWMO9yvDHZnK19BUyl0iHSb4Ec5PY/PNd/HHo5XVax79s9W0eEoIvOWQFYl0DULAEmMh5Ee
6s71Y/FLDq24BvfVlx4tOs72/Khe/xKnC4MlAvxcjJLVJswvNviCemixfBEOERFUHD7R8an5oEXO
NdfuwAXvnKyuz5xTj5dTqNbJQ4EHXhD99KbmbJ9aGwtXtZ3qnIhitikXBxr5WbiRr8u0TDsXNRHC
ELvXv8j5PTk8F7yMbmJM74ykbBE8N2602Vugc4iq0JRKjw3a21y3g+TfN2D6xDMFWnBd0W/HUVDm
exeH0nyX3R7kSAZPs3jksfdBC3mos4iGvuYIcoQDZHEBUDFvEfdGpY5Tcs8iaOcGgDavPxBcncHA
2JvhQp/aNwTPnneaeqPXB7GaQOE8b9E61j7ldr3jNyvMjynQzUC7b2d69ORMKqljqncoPDat8ziW
Xf5SVi3EjT8IzgyNGVNFby2BlewHTYp2/qtptk+dn4aoNR1B7OWDyKjaf9gU/WG2hur1iMrr7ruJ
iAjfY3U0Vtel5GB+ghoSMTeDrEP2jk99fTDTikJXhYMaSYMLElaxclgrsxosjJy0L5JLd5oWcNYn
tI5IE3wY16kFIMQjxK7N3Hr7k3oSmR53W6KItOqDTrU/8CC0iV+IVQfTBYINtAdVIIJ1YcJ1Cfvs
kti8TCd+SSy3UmWus4ga6UPKLbJDZc6Crkvr9uQ6s7yElXJ0dGDVMcBfNWAydODbrqdeRC6LQF5O
bJyO3EedgYGQkuK9631RdwY88mexCTYPxqXLX78Rar6cFi/BeRdqoesumA2wv4LAaT9oClpzMQnQ
jDtoooTEBUFHBKKT41crGMmhVhCVFFasMQb8zFJNZ5ECSjCj2KrdOKGcbKRydv8QaXW3TAAj6Wgo
1Zvlb5Ym0KM5va8vkwlvQW8J80tWkWlue3hfZhmxdnwUGaiaF8ZIyxseuI2SMkp20BP7jhV5CTmH
8ITSn3M9W3CYlYLq5vuN4/sXejyrWrClLDVg8HUTec8FX9e2ducElsmdAgTNwneKqpdRgeEFuEGV
R5ftkhNbcd9qUiS3e3woO6Hb/Y8T+FHV+FRtHq5Dw37nW+zEPLRIT0k1ZeYkzI1iinRpemKXrJi0
177Ge27q9lSAmr1um4mangX33zmr9hhs2yWraODZ8Y8nvOyfJ4r350Dq4gKo4lGc3x06Q9x0rd+m
bWGsc795BopHLVQ4Nqry2Qv4P5cjgSahuB8T7+rKS4/rSOh3M359jNdQPJy67PV1aTbGOH7tZ3MM
FdmEkfdpmPrGmHr3MgVHkdOr72u2UiyoIDfNLVAYxnrDc5BhV/hA12CItbYNNwocTPRdMpFg8c62
sberAW8he20Th9PH4iRVXbwZhSzT7SqErIgGm5gl/nDwepJm5nwcNWBys0nPfjAJe+pXpDurkQbw
PLWs3qEC+VkAz15l/os3Dpw5aKdNNccNPOppzeDU12hVTwr0UIwEDsRbCLsHfdGtAyvwEYPVwGKi
ZF+1AHj2fj6mce00K3S7zrbSD/AlqZD2qxI1aTyqJjo2UnjtRr0BjN/L5pmdIe1iae4t6usuQj7c
59H0WIpPZRfjkO+hacv5x989qmEd7bpsXI1UzEwnFevvEx7DQlnC36b/pb60+9Fas/1PLp/ptypp
VCIijhZQUYVFNyfXsC1vla3ZmlyooBrj8k/cdy6VKQEuEALHJqlPL25DKxCpA73wj4rmrV7dqxO/
aZgNhogaPtAFuevxjT+7oi5TZXfr9BFMAwsgSiiUbdQyKRizbSgOZJGdksXnzxDoD3yVZodCahfH
aVtTXU/1UgNnDFvRlrWZTh6hlBx9z8cNdai2Lt+GW0HzkRhyJofy/GBCUfK293bpemsuMbO2tqZw
Y3J8e2DQlh8SVWcp8SQlq4FQt1CvRvKWgOMcT4a4ljxnaI2y8a1TZJik0cHM2YX62gdI060Ts9NV
0bKLC1VNQKAfJUW19xiMSjZ43AHTtIahG53CiwhJRemjrtP+oDZcE/1x7RVHSxkCthtFGxiM5ior
wn60ugySEuOzbd4iB6hg/wJlgDtMibq/KEQErwQq+shDp4cUMRfn6b3hvoUBbvgT6B1XjL7gR/Yv
HTen3QR5Kc8tR0wbd8HCuwezysinoSoK1IJDZLZI1bRLbcJKJ0tKmR5i1gJemDexjd4Z1NcsSab+
JWHCPBq5PqgJHtKG+qnMDvZC1h8qQxr14aqbQB4nU+ahnCZZ5xErb0QS6gGY4d6k+bN9Mg13q4qL
7jkq8CyGM6h3M7MrX3su9fHGAGSfxObjNqDGSm1vUz1f3m1fNxCbyPuFEnfP6Q6f+OWpTcanHZaK
O7SGn8A/PUPZpmE0XNXcI4HuLoPXEcwysjxbM91u6/c52DLgM4ojIy093Wc9iptpz/SBbIrn5CER
TUo5zKX+nvN26Zu21u84LY4NV6P6paeSKX+Qs+OhHtgP8Ddunk2VPkkTb2qog5rtZJnhmh0bKRFP
G7MsZ4f1VC1O17TvXLh+smzK0oqzqPX5bmTueKrF7Ar0rnIz3Z0Ot33CPGq2Pd8KiyEIDv1yo+Ma
3n7HoJ/pS49h+vNhIGtebh5h5y3j8RSgV6zjClqmJYzweY+o2o7FRltxn/y2T6MGRoN97Dwblwrm
pBiM/B0/jE9FQDKOhuU5/QnvZvW+xuXiq1Rql7GxyaErqham/vbA4iXQx9HWqhd86qMwrtQoK8lM
KeHac8xK0+GrqNkL9IVLcBGihvWaM1NWZm0i9VU3cxjEub3ErHTURipSKhJhicI3XFagQkU/Wee4
WySeilcjzk/U7DF7ZPnT6IjpiTUN698KOIuiMkSGBi3scuZJJhA4fyNuFT7djNtgYcuuYJ53v/TL
N9Km2ywx6Tr7LDsvUKfNqy6RCQ6LWo96maKk+3MJHCJOL3UxYJ2fPjBd4BOl3mFJBouHpAmvRbt/
fsEtMsGjrE0Nhh10aXtDQKxwrhn7F90la3JW+mwEAkn0I+A/gAy4YCW/jAcPbAklJzByGwS4xqgy
jeN7KVYj5xRFNH30djy9Gs5oekSqfeoMqEJZaJQpd4C+nOSV4LzYi8BZOu2SGX8e+FkMw1jN5lsS
H9agYbdd2NQUbtzLKWU0YRbjjLiGkmlve5CiZ2ek8SDO0O8W7vXXxiQNM5Pgxzw3JiyXb2Tmt/0P
E0nqTyzYWquaprk6bv5mluO3f0bJQ7NNd7akuCq6hO5xxD1VJP6cAjT23ZzEr3Pb2Umr9sDL2YVl
m00//WQePymqklJXBBg7QSt3L/Y1uUq/bvdKfS7hqLZgZz1GeYlUfcLgDTHl7fSv3G46UHqYJcgy
xnt/LKMGDLcemCIpJMXItS57VwA0YBMcBG3ta56H7D0HDNphaxFGP+VkvJ41lKfGoooCibIfzS1a
0VJV/gDb6UxztJYFm1M1aPrEPp2bfPdUNE/oOuQRIGdrJGkaZMscK1RL4K/gplVjziPk2X+Y4nLt
vtP8JfCZnrVDsbV+qqaNaMCugOFCFmwXjYBjxafl34a0IFKZvtWDNhX/ykfyGlybrwD8fnXkoS71
DeePUEKdUJp8KjJR+pBB62sM3UBEIDlLzx+duBtc9bACDqA7YbFvHyYPSMZZPQ8hCwvxvFgkyakt
mpnJ5+zUf2m1KJ9e8oKOxLYhJTQ8TnJ7gePgAzH/1bFcH6mHCiJTLPtiCDNO1Fb6byUxYnXwZrxr
WzsdsAfIL4RauEdGBck33ore3FKslBhfJmdGQNq8fMOdHIi8NbBAAcFOKVoz9tY/7wj7YE1R89NU
osNDqoluGgwum0umQXxIbvxMthss//xTTUTV6fKUIxkxb4mui5vpCsZUBs7/+Hwl7D5VybopTj+x
IJRa8m9J5O9czQWDiBun/yzwHDpgRFgEsNcAVzdRzg6n5FQbB8/SrDVhyEJIiqOsscobIHr7nKM5
l8BDjUq4kBnf2o/Y9kbEhk8f44chsdfdyS4MbD9X769RL0NdR9q/Q82IK62ift9DhasnYGuSNYEB
crRBDkMxcBaAnhnCvj5CC1jmU778Q6HCnsMbTtH2c4s2LM5XuLLtLqAn3VWj8nC21gQkkn/JMT1r
J5Tb6goL9wms+9IzCenSbh/FRARPptb4JnQc2Q9X1p3tEnkTKOCM2fQq4jq1HCKoeo6Ah0Ir7tG0
NKmYz5097D6qlKdssfLs30PWsBvFlRc7Ua2xtFfFdYqvlZMraDytwCru84vFSF6zm7r07JmiICFy
/iBcuBRsku4TirCX5LKbRQYVAWpa2G0kU9zsmBtZwCnB5FCnFQ+jCdO5g9LQxVOoHeF9m8LwmLbK
AWXmit1JG1F1i7KKb2r8xUvXcecg9e6P0eYbO0jIADFMCIyM6vNLE/XD4uC6r65OYAWHWUCrFV1s
g9a6kQN61CaYKyep/zMbOmcL5sj+WabIoRw+P9y3dro57iznzs8dGQSyEhDwzDtkQ/I3oME6uD0P
pH7EFrldk67feyhlx6pY6Gryb7Xf9Ls19hBYw+MyuSjslrY0HuVvdrGP/DFRH6UIEzlDWsq5ejaf
zwK9OgQQ9hKd5N9ByahcJoMj4iUM0dNqeR+ieCKlUUGoMeTJTM6WUlqLQi+NtC8vv4FoB3braOl2
guQrv/1dT+yTyuxSwyuXQID2KzvEeORKRufzWx6AqR6WrtpEe1cSjeIsZ8+VcdM8jBE10w5iEsws
AYsyu8su9EqTL1seWkHlU80VgrOIronS8vPLkOHmpTeQlSRo0bJQqqVq2cQSlcosnJ5ExFNJjQ6S
kYtM91hZXaa5QbWECt0tF0T8jdvSatXWTCULIujVgM+g0deVNLc51bN5xUEC5Ede/QfMBkZtVHUO
zTfwM0FJ3r2iUGuYEgqBG0Uw7SGz4Y+tSGhZCOWOHzXj6NKogsfdbMsA5pUOzbwUfjLSX/CP0Oc4
A+PWJqfdMJa8vN2ovAA2e6ywdjg0RvdlBZtoSh4BQjagcExKcH19ia29Rw3bvEHCvmN2lJpmWxE2
O36FmbHyNfK6izc++t6gNUxvN0eLOqViJG8OYoMj0Yd/Xzlrlo9phT1ntrpMzr3928X5jZkOyyCr
YAcdCQMe//kz8eyJXy54EnttM156yd+ETHo/ecQgDRlXmXbENGiHSv+eobzD6i6r1Z326rmkNRn8
/FppmNgeXnFWE7uPWjZXxqTMZ0fEBnrprOiseQYcee5KJo94+KbqMTgZOU9D9GFi187dAj3I6Ua0
mdY2y2Oygu9ZEf2T7G7bpyXOUdn8TYuj1vngdrjYW3S2RqoNrGk/cORB/cf7jzgpTuWf3Hcxw5EI
WlLe+6SYgn7zDogFfUW2mPG0/0blQfC8O9kOxbmdVq/sk9K4XcrWpBV4mKDwDbSo4gw2ckMelhEF
s1dvBWfLmx5sQy9VJpM3r4hV5nWI62lr3LZzC74xZCyBJPNYaSOy13sGu4p8UwqLVmFJwwhhec0T
OqDGvMOxnsPR2Jb8gV0vc2/otq/EPitr9Bmk3H1rnCbDW8FdU9CotRrbfjX9zVbII+VluMEGbdKk
QBYl4tCpS2+1EKYjHEzwLGYvvcxAOirkcuGCD1vymwpiQVnJ5Sy1j5Bz7q2t6twy7BX9EjgZCzui
IcQ79/7zXcqMa7/X9FmxJxENNGr186Fp3ysfsy6CKQ6nIz1zc7cFfog7d+hRAkUnEXtYOYwr+/Wh
aO/bKoiXsk+n6gV9ATKcUiY2U4FruabGB5imMO6jXNHAazUc3MP7/rhvL8rrwhKY5pd5N9RuKBBj
JOwbaTWkPm13h9ikVWCC3C3GX5ri33PaT627SbTZpx7qiaWs1+PfSXbCMIRBTLZJX6FDAxK3H84k
4yh5hT16+yeRDJhER5Idc6dSypeCrj0rFyLoT5CsTADJLhrqM4/OEFzz1D4Jk7USutaGMD3b0DpF
HvwnUOIEh99uY0bsXnYiHsdQH0GA208y2MWtVIS1Bn7SHHylq0EoKFk/pZ/JznuPELxrzFImFq4Y
PolbUdyQRjIfRNg+1WDINlTpbDfS/nQK1Vc6ZQLvmZUVeYnaOoj0ryDlHw/UE7lDwanwISxamOJC
7UcdGOS7hSnW5H6jHbs5udDQSVd+UCteEfxZjPqwwu4G3EhWB2ByFcs4+96TFGR8nLXvKdcktxGL
S6xk1+VacGo4QM0WgJo1Hoz8SdSulPk5MR+raOJrIFwDP+Cy0BURIe5Ca0LFTaV3V4FVeDoZfBfl
BVeO2mK+VOfn0TflFMy9+d1OUjBBSHTCaIP3bIAlSadEdedf/uZpjsqlgPD4Ejg4rSbkgDX2vCot
M4TgopoUVqXYomoeci2nE7aBC3VMqASXGXFYuNIjgTvDxi7YXTRq8JoqNVslkdTZxEMMDWGJZly7
NGHEEOmMTvG55yvVYpasy5cpSmhi2+W9XG7URfGKylUWGJDbPwWRFL+1q7KtYOvgW6LLr+RW6/2I
2WN8EJyZNDg4POZWX6IMHBK0XEgkPHla/rIXEb85SpbkDDdXG6MpcpNosvDZ9wc/Q5NBRERoGLuB
0rFvwq5PwUMdmph72sSlYQGP9SZ+VkK93vPKpUZoJesQ+q+wou0QxQAL7I/81B1uGP35fkTE8l+o
Bnl6bbOlRZxgxCuuXxzN5Y+ilVNz0AYaBXFcpBnI4gt/64C8Dg+CsRnW7gSUbGn/tat0SAslxwVD
jPDIkJsXN5/pbKRdoBkD7uEKvMT9tHRQxE7IByM/BQ5UaUdkL2HDZXuNRbsHVOlwiK//jj+apjZt
A/6XWmQllZAM1xrkZaqqgTm+c5U+Q632AJM2sl+SEJSlNYTSEKwbSsGL2geZCtvlsFan/10hz2G0
DXfA3Wa+D6TGZH6Wlt64xLxK9SIX0eyOzdizxcjPZepm3IvrLxPbWWCJ29neOhHD7jcZNkKeGKk0
dyJyrVkKdOmJIFA7h5JQUOgFoep/6ZoIaSLifuB0YKYRQMfQaxxmc83x+cWpHckhWMdZH9Uuz9Cz
jZ+OuXsmdISl37gwy0wZDBr+eEc2YbgynLkNruDp4KZrAUJnxsLtUoip8H/wiCAEnDBHRccswnIq
Tt0G9jRcYJNf4R89b6Su5+k4HfwP5APpyKXmUwEUNGGxOYinkn/H1J6GpIjjkuy/ZwJZ582scDVB
Otx1nOJBpjTee46BLGyQasKh3EkJLGc7vfJ52BjJu16j88VwqDq25fU108zZZlJXwkrXbRm/ABnH
iiK2jyzMy+fhurF25+Tb7OHeDjAhgMax0jiYBzPDy8IhdrQPbHl0z2YhjADGJ0En5iAC3/UZtY6U
AuMN6U8t0QrZQCicmt6aZEF7nCzk5UeFMB7o1fzt7z5hM1tqV76x0usd0pjrsplrNLsjrDt5o9bg
DbXdLjmcyUe+ZezTM5VQif0PwTx2iubCAxF6BFZ0pDe1IwiM1GFD2XtteScOSZnxyHcY1xWi1zUj
XDmXT7Z42dM9HI8LEkQsuHwVCjY3sjLWAyBCnKmEwJKQx6WkxvGZVZgt61wSUyGuCXqyMZDNJQiE
nd3uOAq7EgvlfrpSvb0fmhD+S19pvynIIcHxGiUD8RGBWk8LOi7bVReVCg90Mcpn26A8rXDxzj5b
60j/DIVVkpaqjRQxdYeGBa8LQ8ehf1ewpq92Cfa6o0dEBRUd+gkEa++suVMtySKIZB5pZIbDpLON
hdo6+ANG0DlgUK6sSkBES3s2TBTGkEJRvWe+0AlQdWW5MpSHIOZvhYuCQE1pHwrlUOu4tpCC+77G
HeOevmmvHxj+a1SNkyhL0SqeL+EA0Aqfs73rHyfWuCWrmFAYPUD4R4WvGiZG0FkjhZjs5SrkSDUu
lbeL9m1Dj6JlHy3gV1uDbEZOw9IhrcLpFGHwOvRTzGfPRO7u92JTlohpVkiaAM4l1NmUMEpPiCoD
0tuJldlNiW1DH6PU45hcXw8F5fHHxDtQALwETs7wTTeVtuLou7AEdKy6PdypuZ38ntdwX0/XBJlR
kQO7+FSVaz0Mfoo7Zw9/2MHXRux+ZqZi0d/ykwLECrOdQMPBjh2nDuXnq+JYUf5T92n5FLK/T5co
wHbfhY3znz8C6HUxkdLbxWJ0RjmQZStkIvVgPDlhx1s7/GLlnR1KA9UrWhXuqyVtVlFr87n1/2OS
6ZR4Lmq5T+iRMcqv4TwfzK2k+P9Rhifps3M9jhyrnjNe2Fq8H0ZN0jZnGWrBFMpVT4oV3FFJB4kX
0y3cQ5iAQu7/8fNasxkcyfixlEVtEKEShj7tM2U/W9vFh8URmHcDaP1k5trWUu3QJUeieB5ep4nw
YFEvoRPlw9XuVkcr3pQ6nZ4g2xLbZU0wCpO8bdJZMm2T7Si4hk8hW8LT9WWRmRHLJKU84ZbOOVEn
gKvfH+d5YWtiQXP7FPLV7SDnyzF/1+FpipTdujh1zakJuiC/Mvb+D0dU4kSAn112Vf674vGl6vJD
W6n+GID/ZvjmM6rfrWrH0snsGDsRHW737Qt7pXQBBbu+v4ArfAfV0AibdkDkDb+K6EJ0T/HXYmQY
gL9/DA/0x4OIeBFbyZvBzd+wUfrrqv8W28KmoK4GtQ/2FwMzgFW4gm+kPyWtovsd3U+IjxAIAevu
lVT6z0PDDhZBJ1LdCac28GrDTPpGa4jC+UEOVO8GC4Ks3pgZ7PvksnixxVla5sM8m+73YjzdFn7F
vr41l7BGevKZTXuTD3c7RMKXlDeQKhKBXhPyQd91AHvHnENZN+pxCm5+inDTY4bBxk4P/MPNtVFF
PELo0GDDEFnRfeJBmLO9bPb0UrHRtWNE32BPNo5dC4K6wkoFxkug6XXta6qk9C6iQx4gaLhvItK6
KW1bKDUxNas2k2cdVXcOeRCESwtgwnlDSdAt1QM/Uo6w5u2SGZQYUpxHnw+ObEgqtU9pvvhYvAum
ePvRn/oZt0wmzsNHnuES+Fggm/j7eP+dTQ0qGMjYecwlXB8S7mViQMu4Nl37RlLTvyjhWrWisHX1
l0xdKmB5bpIuiC3+9kPV6U5NeIfwDU6XMGGbAuaXXaSMKMY/kXahaihiDxgfc/8V8jo9Cyxa4aPH
bUhCjIA59SUO28F8u2ocmbCdRlp9PMFGQN2KilVI1Djjpi2H0qM6dvkm7IDoWiZdEM3JB9lMdoIH
pYPuM4QjoCqvnqlHAd+DwGOss6AwBmLLDKmolIR/gRhg+Uz8dnYgn5C2IoEiGEV7g0weX14eEo0a
SjcQOqoda+15DN5geJu1j5oip95lODun5OMpYrFNYf0vIpzdeF/iyqPqNiZofsZTZ5dbrhtGbU1f
wpRcOVgWw/ffLq48FTP9khKiq5pRbDuGCcfCe9MONqYLfl/+d3fLm5rffjPIHbzuYWGY3s/Z5Va5
5+DOGCIkXK4MY55bCwnGFKzN8kgb0qAxF4Jp55awLiwUQXnvE4qY8PTAMUUw3YzJYT7g6yKsDayG
m5KDK0QYqmYMVJMiSZOlI9dA90QwxY5PqePhPiRkFPX7/cGYZ5M9jNcbr1z2jjEgU5CiFPlrvc4Y
cY8yvLvzTYLpSbG1QXOQA6J4Gls59TXSuc8l+EoYOhp91afl/+VooPjS5Rb8/uryXpcq7trv9Yf5
Q2NsWn97uqc12+BUpcSxItLVLbdWAQgfMQX85vPJxw10t5rMjyxKSTIx7BSuv05d1R29sZis/r4F
4Pk5AsMwLk/m+NbEz62SwiqgpyNR9W1CdNP/ZXcqk2aWngVkSAIoQNeN2OK0yy4UIFix7hCyiui4
twxMloAfNaOYcGFyBc/tKHoumL7GR1yDLRf7eRRoqN6+E6xUR6Wa9fFvCzOLh0SwtEiCtrwX8L5c
fxoF3b3PD9dSUPi4UAd0wZ2zmaJrCFSPl1Ydp5Ph8rGUX6FGMGGfA6F0ioR/9wyjaUPLG4ihNc4Z
Oy+DykF6HGWGzsLw/LscImiOklC2eVG8OkKJkXCBuJSZ0MET/zzEVh9+rZ8SVQaVFSu+NU9fti6J
1LL3QB0hwAr+4jbYz+4B9ejROMl2B7zcolDzyH2OdMxPqAN7yqnQiw+uKPDv1qQNE7+03uFZm6SO
geqYGPz2HEot9dVobeNAfkMjnW/NiSKXczxtQtQY7XLxc2fyt8VNqU37aA2Yojlfo2C21oDKo+ho
GD9tMc1HuJC0opYPhMF8RDv7xV/hI5vI4X69Jj+VSZKW+V2fQ9xXhxtGDcH/GWMH24KB/0BnMrtB
DA82/GI1cfWqYNkwnIEIJsW3yzptOGm2DPftn/dI5NOtov46IC/zFOYPXbrXMay27BT+h8KegvPa
4X7R9+L15eFesGu/uCLypTcxOvIOYPDDIl8M5FJXyFCs0ruHWdek30RvzSssbO6s4IcuINnvAA8R
qAqsMPYhixOfMTWenEkg60hjSDeE1K7sTbaf484CRiXoaHABOxeKVdSLMG8OKw0uCW3dk0Fremro
0OAp3O4NxA+LHx24d55IWfB5pPU4l7039dcRnq4GWNM7mpP0fZhIec9FmswhIZgLqmbmACdyLj11
MmRb4QMoYfNMe96lGnh5FZBUpysjxe7wNiLDxijrBtBOQcwJmdyJn74V6Cb3y4SlIdg/HABv3grH
BYSGKEec8uL7zCwAa82CPka44nMTToiFO0tvsfY5kNdS82leRRSuXfwxsiDAmXebh4nKkJJSOqVX
7Owpgqptc+JPDv3gjWtipEsPz+HT54E2HLBBcg4knitkRifJgmZt0Lp5RG8AnAx5x1yrfOAt3pXV
FfN/AwDEtcarADEXZFrwgsWCegn/VS46N3p8wZDZVTcdf1Tz8qKPI5017mGAZSj1qdlJdRACSKCC
ThAz7lbHplpDXV4CTcHlyEKy7tPs4KTEvZnH6Xo6wTjIo1uVySG4oYokLetrGDg6trPMH8872/w1
LoBPGV/57ebTJ6z2rz2odrmWJFwjNwlDPA0Yc7ZYAvCeoc/wO9PVslUr7v4xaEi9bJvhCsMFj8Nz
1PD5kYDajNwD35eEhrMCn6OYzZhls9JExR9EG5dTPuAsLFztDNMDVHaV2Eo/qmixLyDUOnvU16ca
JDSx05hVW3O5Qv4t6taAtpkRU6fb2g2u2+A9RkvBMKj5N0wG/9qMX5fNy2NzPtorancNEoMNmsSj
RVyHKFVWM/bnH0suPtvzvxMX/aJxCtOMLlwppAraHYfYJxkJhFO1m4GXZio8YJbKd0hsguUf+m9o
Ui5R2TQfp2lP0AxTD1pwwasEgJ8Qrs4TjGoVs2q3s5r9qtVCsC4QqndOSbOYpVtRT8hfQceo0b7t
3IOkuevKpbN1gyhPlVsH+ije2qAPY/lks5CTeo4M3UU2rpu4SBFlCgvExC+4YKMxbdc1Rfjv30k9
MokdNcA//E9Cp15tFByWfYq6VFOj9TkdVmg6mZpRb5gDp9pYWPZNBb9Pt1YxNZNbT1XxPozLAjm4
W/Y26WyM/XG0F8sO4Xri/kHwvNHZFKA2WHBGzuntuOOLt1YiU6ks/01YZNCgFMeSMNirKamwNs4K
uS6XzFVKlilMymQ7wVPb08gAgXcc8c4bH65sBfSpFWzDeTCYDHWItY5pZqtZ97OP2deVKOzIVwYj
H3RRqdFjU2T7UE9w1mGKMANtyHte27Y9mxDD+N4GsMm3Xq2+TJdrmGWYAONgNHsK0UYdg6XEidHc
6Up97t8fy7kedg34gxusU/wV3gpeS90+2LYeUc8VlCOJCVEahLp/Y36DQkArVbUXIwJpkLjRZnWy
8Os8mtrqMDDtydEHc4a02CndkYYAR8CJPsHNBaYzQ8BN7WsOWvLDCQw4vchbkW0Bpfs/iWwQw+Cy
vdFCvjahIIn4NoLDPLHh2VoF1OSDOTa6KgVHFXq6122WLTmwHrYLvW4SYN/zcu8MM/hAJZYgzr4f
Xef0vO3dMNxOL6acBLas1Wb9XcHKoiZkpymUMm3pobIjKusVOYZ8Ci57FmjUrKdIel4GSzWot8Hx
lR79LUD1Cp8XsbgKlwc7k8JWFYHve9EUzOAtwo0pD5GTGGv1JcetjdCURmfvIrrX9jNzvrgz9PbK
PyinsZdBfonVEp3M7ZztckVNDWZKuKRvGh3Q9CeBdcqCbdKFz0EEO+invxkiM9cFgbumJ/TE/NOp
hCTfYYbLwyT7UUQ3qZe6wMEkcvGvdMiS6UTfcxHBpzx4fUXDj0A8Bf5IGIbwh+axNZ9g6f0evWQM
SxExRm+ftmuBDZALSG6SznF8P3dFwhKo1OnXYozAc6FtuFZ0gOVNHilNbWK51XnwbmDIPVC65LBC
KeW4tha8qTBgNhBiCUqQZPNtcjOGvNz4be9Jvx+6LWE0NSTUvJT2lARYoAP1u6Jio1mN08E51hLL
Bm7er7hINO5Q4iWfZTdYhGejPmm1NaPFCXrC0Qs5LnvlgoxznqVfqWD9ZMO3Gtz/CCXUX9WtLpS8
601k7u+3RDzV5ssBNtKlXC5mdguH0BTOizgIbSBHUu83t2ERMZd9Wl3JJ4EyzNI52aYNKVrdgryQ
LvwCs79YcrMC7mSe/DbaW2dc7zEKdJ3CeSoWxCKeBrwxagLcHb9Sn5BazQh+rmgh5LaKTAnTnVKo
pf/OOOJhPS4bbw8Y14jVjhwIDSAVysnWzCdmJxqzCwPlun77FfQfbBBF4tbsqB+X8+G68ZbmVVLJ
xdMEOxo+SgvVPMeIth4UiEDi0CO1CAlBuD4cERoxFlthHxZU4Uppw5CZKTehi+cOpOLWNwI3P/pf
tfNJh+FJWucWrdxXxqhmHrfkmAKy84+5UdqWMLkwixy39vVkVtLApsNempbjhXGEj/zh7wLKCT75
eKYw6mL2ZAXB/YhFXFdjiQRGm07czxjqKy+Af2upx94diwnThseQlO0E+CQFu9uWmTotElGHsxey
PraYcZaajB6YbMf5VPTGtcmm/8p4JOYG65IjDnt0MGAImNH8WIH8RvgpUNfnqGQRLK85P+BQNkP2
BEWr/cR1thzCiMzfXL42qWJhUWLcCewmTUBwdY7PI0F1gUCcR6Kr0iOi7Tn5VaDpfBlCEnTpwO7v
ThFqtjVnsKcLjRXFqUBKj47Dahz0TGx2WSQRyqpP96kA79hamBC3MatFUrvxtYwd2UcmrU52gJpo
LYReAGVef6CLF6Jitja2Mo0o0GAkBGGtGUlzZreOJbY+L4QWPzz7n1Xq8qrVPKyKG4Hi7stTF5Ol
53BBZjRevv+qLiZ2vVnwY/QIrPHjhJEzTFCoXkqr8HhvE6Un27BFa2t0uW+ZQfBrjBteBvcg7cWb
wNhcEK7FRUhxnbqBxATR3y5fbiVUGY6iMcMO8wlbeUSFUDtOenE2eCOnuHpRet0TpVdQx2RzmQ9G
V/l6O7yuqnT5p2zB2Q+xeRv/6aP82SsjcLssxUPv4cChUp1yZ3dtx2FS1JYY/fHzQclKHZd88G62
t9y2PSuVN1OKaXI9Jyoa70AQ/8vZIEyjWvkTC3z7l8UA8lJfYkH2xAVWpCVrd2lH4vj10UtGBYKp
9gU2iD2Z0O14MXbA+/EUrbSlvYoLEfmkm385+rET5ROI57n/Ak5dSZBq5t25qK9nHhIwZRZgLINJ
2K56E6YTOu0zMw7AppMZ59H6TjXY+nXl9fhMvLXWe/lMD5mxE0qvlacsA3HNf7NsBEvUlZ6EM09K
Jea38dVZGA+W89Y2GFsRqJqKI4NvqSdX/UXIlasrz/K9TPElI/2EJqmLckCkRxURwXeXm1b5roQo
+1Qe3D3mezvVW3NO5ltxl8by7P5S/3gCu9getwB2dJOrcX/96rMt4rFEoKElj+Tv5gIbaMCZbVoE
I10LdPMIpk9e2wjCKUWD9gFmtsGBjdd92hUmRbxUNU4BF588LY/ecAHKEN4F88T7M/+iMdZpqSNN
9IqwOf9P0XvdZv7D4eP+5rQKaWdLjqmUCA8Cez/RbnLVdy/j5xf2EZNsQCCA6ErvwX6Op61seo98
69484oB8ANuJrWm9hZU74abq/uooXKs+dZhvixcP+DRK5AhPrmdz7e6/3YvjgDWJM65OpVBIr8W1
y0hp9YZz3sYVjaOSbObtnDqidd2JMKYaxX6N8wXNWpDoEuKJZV84sMuZvif9V7CzeHTK9GUpYNDp
LiS9vUzSr9ah0/KXNb5xmvVGFUtEiRyph6Ap75FinlgH0nMwZPmC4V19FO3UtQcaoc7f5cmGEm2m
7wRTLtMXOgIWVJjOrPnkTFF6rk/461RJUOb3iO7G+RD8pubXJNrYcQPJE+BGQLWH0k7D4N/Cv+Gm
QXLYEGIlWdbD98qOcwEAu7ZOyFla0dctFmrYWIK7evf7I/qR6i55DB4ePNDSpLCO4htLmNTFK/6a
d0QtaQLbhNzvF2jMyZF7dOOdfz/n2AL/fAEaiyoWNpFcOQffmuCgjiDTsj/8x2LgueYmDhdukFTL
GG12SmRk6Y24DLhwTtx9XxHbQSTF4tmK3ZdxxPL1XfxhoYeZ5rU/9Ao187FwSdKObIQMBvTNiuJJ
yZtFiqVqkj5PZBdoJOm8iQMsbe7IXi3QwHvhsuedOzV6Sw/DeyoxvXlV31GztrgaesMp3w9SPahu
dVI5cu04Z5k9GJAW7fZsHKz7G4zCwju7tkpZftRI7DrlPsWOlFyBNNTLtlXVN9XSwkrVyHrVa3U/
uyV45nnyE1Q1G0THMELlGIeZvHEgCrMJE8DgDrK/8BWGwhZkzad47boM0ZTQD/rg8ThEX0XXmnOp
E27xx2mzRiy3YLttpXgCgOjguiz/c0Io6jRX4SDiR5oOZXCycNE35Y+FBZZy0CHdjeW7VK+7DO0h
EdGS36eNBZcV2kgX7Cl60BlN/5ftvQbJnov+N3JfBP8mRL6VUeew9MKwPWTMUj5ImMmgdKG3I6Hi
QuQgznbcpQH7gcHQxfg4iqwXIcwCwEFmxrBjBvKrXHLAxaJOG2Pfvd+DE0/5eJ29YJOlBCXr4ZjT
WZxDE7cO1cVz32C50+KT3SfrVTDbRh8xDMAsY5F4XHN/48zMqwNBPfH6b9CMj3k4k6jAhUuXlKLR
EWnKhuST4eWyvg9CPp1X3FA3Tu94HVMyugfUP6wPSUee2S+yPcv3yWxazyXYZOama303B5D+VFkQ
VKqMzM5hgDz1LKbefuoVccwqdCzRiB6ZKBy4CX2HccgLL1Fes90Y/MocPfOkqeZWklETP1PVf8Vw
5TkuIvWKhbxsdpjyarppz+fZzlHcXZCQRnkLpmoLWSr1UM0ZXzuEfs6AcSaSyC4MnwxWom6dBvJR
aUNKAdHoz43x0r83sS+oPJrB8eho47y4ST2cgQbieIIyvIo/WnN8rJpMvzZwneDdWAPh6Tl/TCAG
vZck+jarTe1QDaND78q9c6B3lPqbwd/IlMvAY7kvigRWdWl4DwkICXeDEg+3icsW7wvpV6XyQ1qX
Gygudx+23Wjx4JbnOxkwXkNKla0gQMROk5Jv+8QgjLBQ9OvyhzTFyJzVYrAWXfP91/HFRvdSLwV5
X6XY3CFuIrCp498YD+zzy5vNHyriI4Ryun8oy3ZqSR6IC/kZ62QYtoQaYpvqyJf6/2hUOWZUe4Rt
KgmUy2LjwmWlZBfVT9K/WyRukebbwDst/hD0B4N0J2UurUTIIEoF61l6edBObmU+K2nf6nseaN86
6M2VQ/f3GoK+MbpaAprh2ePe4ETLxTQuabG9vMrIrWbP5pAo9sGxYXfNK0HFMGDHpHfJ/927Vh/o
w+NspN8D7mCrIzL7W3ncAIr1LZvSPqz28AqkPVjUZb3Qp7zOMb0mRTlyC8U3F7KzVchuR87X0gCF
S6l0jOLB8zMXM44pVZOHK1fzegHrWfqiTQehlQ2OoYje6DMxk4j0pU9C4cJtEK2TTIp1/gDc2IO7
99TQBQ18yxC2x2qun8D8yfV2QArpTlCZNBap5HfMDcQCIBxyyS8CnGtIdVhli3+Junm9SKZFXjkw
XAkf+HS+z/YcWc/M7InLuZI/4UvZR1698s6/90jgTej3sXDg4kf7Q7AOzw8gJF49PfsN4w0c9SP/
/aIHQqY2H1znX4yLrT5b7mhRm4nWzXdy7tD9ZWQJNi9DmIvf2g/i//CYESwqW7STAF4eveHR91Sm
725Z2jjBz+Ji9VdluyyK8YK77r/TR90LP6oyPCj94X40IiazYpbr+o7QUHKKqqqSQ+BBiNcf9nDK
dTbi8xfC+b/fLBca1GQBEXE1D3Wmt3HMTpE1xDQ9VmDv0TSOTyVyeSrCZdAsD1lLkOVmmIUchA2I
h+W3Un0YfA0SF7PGUckl0RnT6u3NNELdTfow9xUUHe095VJxN5pE77FWStGQYJ5SkpIpyRh7woVR
1zOWkejiZD2X7zVpaB4D4cU8bkkg2kzSkCxd+bxMpDR2VA/i3FwUgwh5q3Cc5cLGmfpGDk8z54o4
yNJRY2B3rcWJx/m/OAKcVmhBON6+2p7rM3VAXgv3sH44hBUuruULDz3qjVDMfRfi84z2BMvZUm9S
2ANxRj17mv6RecFhTGGWIFe+wK5jcdwWhkqus48XzrJ2eaaCPPvA3rG7qJlClvsJw4EdVZt+unWL
1HhesutlWr6zIiwgOh+CpHX21Ilqada727TPxKRwbsJczGvf7+CrvzVKN1yPyn7yeTFEcURsyG7R
BxJ3z/ykvkXpa9QK7AEDh1clfnvOChKzbxSjW7Dn5RkuTV1DmY/Br9szmYCfiHdQp5cN9G1HPqKs
AewCvr2xb14dwD0XObx9g5GIBpbinixd6Fu15hc8BlP6/KhydqVECnmS+7xro0q+6hMenelxu13O
rXqzpJTJ9vL+dGlblqVa/FgeSKDUIXVgCEbNrKJQvzjTwbWOWyzF8RPoNq72ChYxDknDlyTElJjJ
/zImuaNPsyE8tRfRQd6uX4xwrjNxmEIjeH2BRnhvRre3jKbmn19iS1xtaxLUxAgkrR8K9Eicvvvl
J7shS1z/EqMT0+HKxOG3v8YCJJKvEgQcZ0LWqlnupsH88a9NU6U43bQCk4cfLDLmqAy25hDacgqZ
yoDGj7A5cOYNh32yTzdtprCDqAgIKYpgg2nn0pP4uo5CAUVDaizmwrCqLqZGH2LqrtyVLmheENoL
6l7tKgOi8jm7qmZ223JKeiG+uGN6SrVXYnitDS5A0z//AWvEREuWLVf4QorfWsNWJnptcvlI0Eoz
PDHzT0ZvKEpQmRWhKGNBRVug+hEV6bEt+0rRPSVBtUcJX+q9YWpuWlTJGsnHz79Dgo8Gb8KlrKgM
lNl4/IPiIMmuWBo6K454WBiHKHqGz01GZSovSzLTlzRQYZyPnrxxi2K+aj/DwX/wSvjC5HgjhVsb
s1V3seZs28pVucDQzZQeJtijLWaidR2ufzpXZU+1o1Chu3c5YdK1vQni2zX3+b0kf5GBbvykCB5J
CifTecKjh0yVi6o2dc0+7flOHKr0t6hG9u4GKGdu1vb702I69q9QBYvooL1HYrKBKzACm+mjZNx5
1ySPVGk7VUpO8IRFcHXi4OmDcDjj8A+FaIEiv7lR18QiFVxm7iS7PK8C8FyFZJhmo60CXuNRJyqO
Bptxn+6HRdouYwebs5meHj1VbDRAeI0FLBjy7+xe1gpAsWoDqfKzpFreXpnoXidWEHIJ2KpTv3Xd
slY6pVj1N4E1KMUABGVbN+lYGQpY0ltNP9OgTiDA9I2J3ejv0s5/9R1u2ckbtm+i1lURkYei8eQ3
8XN52xKTTkA+g84Tuvmvj4oEuePSVU4fMJk4yCxaJmU5JgleGaFNgun8Wd/KsMDCW1jqbRwfxiIp
EGLUT059GTmPg68VU0x/TJP5a0t1c0GLaKi8UJYs67Me7KEQVDtf14XbnC4ASCivuzTBrCr/59pq
o8CjwZIz3XGGZKW/KCLhuR+PuHMg8OQpyzaN7LlhSC7uJx8vDSP1CTY6E/Nj3uHeLZa31TAlDDIE
cYmoaAVxIysV8MgRSMOqLh958InIQr1zStctXRV/HSJuBJWKAGkSGHrj2rXSYW4ttnJzRs+SD53E
Rr/URJ9w6CVFJfHf5Sy1PIzc/ft3RFiX6EuNmPOFLuXdPq+DqdOkNshj5/P2IX8mmWc4KP+Vlrej
Xv13E771Qs7rQKrsSL7k5+QJnj1pTfwucypNE7vZN/Ljjtxln2cfPEHvlJfyqfACDXUKuuKl5/if
MBlQuNUCWhnjYrY3t8k3Iay/Q126/aVT0S35QLa8J+/iowoCwCeQqrgO1a+5jyWGDj1ncD3yHdjc
zp838tsMQBl0FpGYqGZ/TaZ49Dc3y+KvWIN35GQC0crLRQ3WIWNn+jVHQ57ZM+e4kR0HjqPVmMfT
qun76B6ph1BJo7VTk6y7JuA2uZtbTPSaT7kXTD0Ad4MP35l8RxJUnyzqHJywPakgxNMGloPqZzP2
kdkUJebdcCAGXMdy2qqQFM9VRxaZQlIPN4UxqauqBnHQEU2tAYpM4WgjsMeKrdOOA97DyWvZE0n+
jQTEaUHeLTTXBb55639lcrimdeWXl27Gt73l0/BFmBXtLRRbYdgkfkh4fqtISb0dQagTJkuVZirQ
VN2wZGZy/XJKrNtWmPrFCgO3Sl7xPBIXQkDAjd7IKSuytstGW/X4RhE4zhZsNFHnsiQ+hxGlBgn2
FztHWP+hHSpFiSBC5HH2RyfkVOIyXuCUPQ/hrItsYC6pHcRGzXqKnpCvNDBvUbFBNffPjDpzLWW3
Ki2V6iH7socayLS332saQfG1Y640jbx0VSNjUM1FSdfzzX6BQSxQx3RIa28ubpMpUW3P1uGGqDst
mp8nQ1rDCrE6Gk0wEjpzf4sP/bjVeCl/F3MDjBnrLXQVxj6yYvhCSsLtPRoVeZj27re6/NT1ffay
Jh8GJ2GdsI5A4xTL8NIqWGU5y0wGBS0drJoUVpda5nAZXyv9C2IB3vUKifpJyAGHh8j8+PT2poij
v7xQ6dA8QaQ+uOUJcNL0Pg1bcdvvyCHePlXRWl8Y6RKyYs8a1pnxH4qW+D45Y3DUVrPmHNbSj7TK
1uBviZ2XcrlaZhOEJTPYzkBaMW75t6AaUVrCZ676lDoN27UZ2D1hpkUq4s6A+2QC8sVPQlKCQaru
XV/XHKRG6G6p1xSSyGRcW4OXrn4kKAounezbQuaRibSFulHBwev3p9UrF6jW+9TSrooYaqtAh3Yc
dhUUSFIQfSnY84Mf1FGLh5ZmoU4apB1+eHkTxFhhOZTiFx7ZK/YrquJ7KsgJEBXMip3kRNrP2d4j
36dS+B+NLEE4SN0Yz3nBsolbXSD2d7KqYYOuAEWctInoB/nzU5uCGAJFgTMvmW/yLDJ5krmT+euF
3Br0MIHH/qiBdQ5x75O3mCn/VOcBLq6h4gkYh5H3W4hvzJWFCOAlKvSHHDCpL7WGOKG90DpxsbOB
a//oBpWHDxrYKtR+2wWNo7zkQti1qbPn2RNncduUyEoziwnOL6Nr+BE75oF8bb+o20tpr1rwDf6o
YXrBxGbXwU+MbR+P+3sX+5RSMAnWkRMQoN/MA899506RZHe+EeSs3GxbzEZLjqLhgULiCK3Jqwmx
+CnniQ9oUZmwF7ipTvITNE32YTanmPfrwyTdILUNU5iNdYuNTHtmDvoRA0PsIQYWw5gwj63jO3vu
/bOcv0d4kqvrfxMomSWkjbawYn31IKYhBKP1oLDQmzepraprQeXVwrAWsRJ8u8BZ9loOmsorIiei
vtoCo8MR7MKachnqp+W4IDsYNgizTfFN/75+8D27SKGpU1WhkTd94cxDMXpYYlSgKKwwLGi4esp/
PU6pzKtv1wYqZxt6lh4Ax7k3DLtDRMJzcHVPIqc0WZQRCQgiO34Lr8dAS3EI5bm7rfGMX7jLz2YI
h2tuPVDWXmb4Isz1X63VSBiSkF01q2SOr9UsuTCe2wIWgguB94aywwypuU4KInLJPkTISXlZLgdR
32/L4xt2zj/PC2pAW+/TPmJR6ZLXEAHfK8Vz/RnBPhqUyhLxXicwQHxdPrSFjv8WltsOLOaXBGpz
nk1tRZ+b3djTYYlsH1HR2e0KxmNGMKDc3Z15Xnz/+R2HOLVPGtjRkqMznYKu8CEBCh3pxxTvj1jx
TRXduta40joRk6h4x25llRtxbcnJE1Rnxzd1pWevsWHySxypEq4M07hrXnw0aUhkWkyYca93JHUe
dNQ8Cf8xa64bLVNYR6mI64XXVfSYYKOxfMfKmkivdwf7GPesBoHs8xTvnlWCMfvGpvXKdYj/em0Z
iN8MS/8DimllSmOd/jSoQFGfqjzAjkXaHXugGOVSTo5k2ZSmGrjOZLuaQ81PAscJAuxATVUWWcrR
Vz65Upwk0elj1xZ2vOCLIWA6uKbFhw6p5zCNE15stymoab1qtPRVuwAQgZRhjiwU/R5BeVC0BALo
6bNU3Y0QLzOKSWnsVpEm+OAJtK2/V7u5ztcYS0QYhkWpCWMWy1tcAHGBJHup6UfQAVBilyYP/9Zm
bvr9oIFmEDeYYF8mSMMmXrSC1sz2FNJpi5VXssx5gC1lVzl6YAv/X2aWhq6WTU+6aP6KdSPsNB10
S7QfLi06Byz3qxPKixzLOeOI99VLwKRoWKNVEUQYOWxyBefkjN9EkjUMqmwS1rkSq6XXbRlAwR1S
BhBFa5F2k1AdHUPULiiwlhlXHj1tV+sqpRdxmJo8dds3yKZpSofIglH5ef1/Zbs0TQPHMrxrvUfW
UxHFq09nukbB+WQwFW1qZRPzVls1/rsmXRmfdqc7ZFsc04xqM8rovF8Ud8Rn0CW0dR5vF0G5KLsn
BX6BXzBjMSajzA403/xu7omR1JO2pVq/Sur0QQVivW8nBs/gezObvFLMR99kcl+UgdV48lpYKARu
qZoqBzHSkRIFUnJDhg6flJz/pWE7Z9nLKrCLsDM/TSjng3ttBGaHMPPJx81LZdpe5kLCGGbxJiQJ
PRL+V9E1pYBKCPlBAgdBjvmnw46JgnRiagXDDiK49OTHj7md7OXk4aVfK55T6XPd4d7YkZNqL/Ga
tyh2rmHFTyyUj3ouwWE3hNYloqk5F3fGBU4M09+2duTG9m76gWnni2Av+wasay2qKmFZmxyvldwZ
OLNMdaA0th5jet1fZ4hgi/Kmh1zJGcv4GNmmcUO50wC/OAlPkt7DZxpYsd5iYDqtTy4sgTk1j7LN
3rDUS2zXKOGfpdNiis1HpBDBLwMO2SwEGKjZxODM5xGYgJjWrX/6jW/i1nVHCWxwEttAw9nzzsQZ
Eu5RHlpU4ljBpK7TlmxRaMwSqF+rDdtQmKc3aBnPhB9tGW4XYWAYMLv8WkPBP/Sj1dZdEhnQrjBN
H2Chx/QQyCUUOWvOSfEQsQeD6+7d6pm535jjGZTNZrPGEX2QP02sBA9Mo+6fW5aPExqktF6EqAtz
Km5xfP3pIiA8o/IXXPkIplxcStCRltwIrtDIIPTc951smB347Q52TbdX60yV7wKWrNRQ91HnHkwv
0NVtFQZ4vek2BMFA6IwenJucHk0enaGeVRX1YjFZXN3UF84E273mDZmpAKj01eJ5j6zWS0Bl735A
7DKfngtPlWJtdQa4cDI1n4Uf+Y/sKTFNfvM1Knz+1u3BktURbGSrKoEsvN0EhzznplT3LWxrIAFZ
+qSRMIwtLcO9sStOcQNyPlo5PNzBJYZVzwjYCCAddHChFw0+B3emzX2zdUj1nl9s27az24LGR2wX
JFtk6uBFw9gZvmgw3e8X4f8/10tw4VRCI1w7XQa7r2PFCzWasQ92Gv+cPyM6pcU6dnV4Qc62iJuL
Mn5HYfEduoEUTAiJ57dgMFgMIsAFBXgxVexB9If2lM6MQqLkG68xgaOv/xjnd345dS4wlPPNsxOu
g6mzWem4QoIjxS6utWc0sRtZdqdom5NngDP1S0q/m/zpSdWTHkK2fu1sYjELYcfLq0Fkb4dr6EaS
jmFD/IZbErQ7ICpoYFZPE8W91lQxCRR7zLjq0VlRt7p8qXQdIn0dOYGRHTuYithuUzrDWqLR/0KB
uu1iIR3CYR08HRKWWALoY9jWX9I8ccpVuMsc0QGLrhI+ep7d0p1fTs5t9hC32ay6j3X622Fb+8rx
jHouIZR1Lj1J7eTYwR7Qfc/+Lm+QBHf32x56TfMVALpuQX8wExqMixhrnTTNHXgZzQAkMxhMAC9X
mLwSI/EQBQGwJi/+a0jiH3y4cvcbjlYuQncOtbm6/f7cw8g2xP6c+6HMhY/L5ZidWje0TxsvdlD/
CwWaUEDBgP5qhcvIi6Pv4/inFglrhbH37BNbOMmXEVgrpKQtNs6YpBWEhfAVR5HYT0wWGSShIN/n
wm0ERu+tDvtjI6R9YlXRrJX3Qz8XPTtmAv7azpNrC43hvJOYAClN1CbWp9JOJnK3JqC0CV+qEqXh
IuAhgB4ThXhIorTY5wMHDe7+YwU7WjrAim4t5LXv1uOeZd3to372zvWFjzcteyCQd+5r7vaHsbI5
4WV08dCqSOGgyItiQoX+Rt092LkEmVZ0eKdVqLOK6KprWbjt3dQWik6ifCXsv7W/tiP4mAWFUk0N
kG+HqTdvr+HOFhJ8l5+egLNZ+Kw36qfNkzDEX3VfDGTSaKN91N5jKpcY1mzi9OUk5GtyYJNqTuT+
k/ZeRs4TXxaXfcdN5qPgI2hGN50J2rz2Fa+U+wJBL9OXsWhulo8Dw5Ftc09mDKdK+afIsDYBRl/T
6vQUNHXbAArSnTDN9tFW2YBs2ZoRUpPJl90kR46TmwZ6iBTr1xr1oMp8YZrkIUfUyK6vKRo8F04B
S6D0G8q8qKuHTem+0gQQCMH0glnddHtR3VPkuz2WGoyulmySPZLFJ9ILo+IzaNBoFr74PQeQ46TA
onfXRRryvuA4UQB0YlLsgFib3LDG0EbgphJW0YZUVxaVyAPy+NioSUn0TdQrnT/DSa/sD0IA/Q3u
WfXdJkBSX1b3jILIGcxkbq6RYZwKUg9AeHB1EEB5NRYrdOmi45HpqCnwfOdhdj2YEvccThgRddNR
WRMAD+pXbItUhbopx+3dY6KxlShr3GkxGMrkaDc7JVQze07Xz5RMz9CR87N1c+x8U35g6QNZe1U+
ZHp4pHrsFhtjeqViPkyILj2Yy9AB8arASRlqLOTVqELFGEB/0WUzP019GGG/AcNoV78F+d35Mafa
LqviMQnJsZ2q/nes4MWLE6+ErD8drmDpBB28ArnOshS/UywnhYbpCJXc5h3jG48W0kjvi98N2H3i
L6M3l5QvZ5lWlB/3yPNcQStLoWZ/HOojiQJYyWZLJVeF9h3aBPKYKpydZKQBfuoVcYkZlz+6TXUp
kNd9BKtgtdesljygFhX0Bp+0TXx3mdnWrGK9wIHdO4GGfatfxuzGXQdR2xq8Wpk1kkIgiX+wM2k7
sV6umUo1XCOA9eD/TphJcDs+5GVKdv3yKgvxOlwUFtm+cIlWCEbU6K7Uo3BrDcV6Qj8MXGrera5X
GauosZKbHtIRLMn+M3PB/lhVma4ESYKqRXkdqNxFGH9CThw68qSgCwEdeReB9EY0tfQOcRFGJmoj
c+LOZs2Q0h0jmVtgF2eDG4MsxTeNcioOpV6xQOa2P8F6veAJnNYLexN+3WAx9sNtmjuj+FT3GeHF
Hjj3ze8FGMlsNKzpqMs3+qvwAw8q0gCeIDq+BwYgvx5NZZiZ9IyV00rjeWA4WQ+n4nb7kgUk30RT
Ek6WeKHEvFruwSFMJ6Y7McFhlz0RRbzK90iJr1wYzRJjUv/jasI54s5m9PAfy0byEPxBwI8eeP08
jNn3qJECgDXh2zMR+Euo60FKFvhF/OCWbdsq1HS83UFg/Wm6RqypmypoLgH/pg7l7lRZwvNKJB/8
2jbTHnuKqZVuOgNUQHNvMI6iAlnZiYfZNkRzTiWo41ADbVhykPsSGz03eJLuzwwc7ajTF+XA1NvH
IwZoIdONuMfI88GfJjXGN3/UX9mXNcg5292GOE0xGY6HgFmWBpax4jy066qW7ipeGQVVNMle7QKO
Gn7hQ4RxcWyi7eYHDMZd+bL35j14or7T7kLrNM27sh2ZDIy9nfDsE9I/1sAvMW+r+mpQ5v8Vo9ZD
vC2u/1K9oxV7/0sM1ck4et0xhH4WvxMUnnP+b1pcr9BHrlueCDKokJqG7xWBQN0XP2FZoW26NIsE
qMW+iFLsLJbHAUDnWfsfam2ZBV99UNHWR25NofAXtV43AFWXVSuW+QTATOKSsZFduQ14b9zO5t0z
+aO17jm0WPrUzswtQc6qId5Xso+o0HUHs+Jy+vRduQzCOuVNDsYKN47PPahzgaftln7DKePWIMjL
7Bj9R15jqwp963zzCXcRILWNM2/soGyv5edT84eTwRDX1d/TwDnOXkFZmHDDANzp7W1Z4mexP54f
o46DJHVCTA7Z52gUJp8FLBYs9bTOJV/Ugp8ZjdyiZ3YOmHmzIpPbNzoXr+vzY/WWX//f6aX7rZGi
W9QyY3wW4pcd2bvofDaRIwUL01EPB5upVqLIchaJ3YRAPpaor8eAovEHNhZFU8OlzrtqHAHxQK3U
50RPkEFkWoh/pV6sCp8vl8TxqphDGv1ktnKH3k8d1jYcoAdmM6nKwxYLsVnrhftB+0o3xFKZ+5T3
yGF+Bh19HW/eEtzfA39QNyXFrFvYbAtr26z9YpuuNWATK5gCJAAx7433po28brYKgRCGu5UDShun
URITSPYi+ZWduor+U74KVqAWxI46t02nzEMGbrW7mrTT1VJw4CmZM2ix2B7TX09jSQnQmEe6w+Di
iuOPNIZjM8FmJ5BVyvAd85DsAK92XOJ8FyKAwP+Tvz3wr+bQF/L9lzMQiF8wZ90sk6SXGXucBOPn
Lq2RetNhnYvcTPpivCBi5vTSmrMUcRg79veapXQhLPJh2ZEhlDBFxlaMDkKNwyMndudu2lxbrVt+
AFHZRFcaPGadAQzYpi37LbFOxlmv7TU/tmitPVXrwAIo4b7rkDQvYSCAckKhESgIzxhjSwzvD1x/
+/hjcIcZ1W1hJNGPi+gSqiTCPmAoVmjakY9juWd89jrhwfrboGsfK49q/t9rffGMAEC9vb8mGWan
3oDernXNX3JsAZ4k3yua/u7TlPOuwes04r6yR2+bB04m5MgT8PVIrqVI9MV0586AkOq3v3586HOu
tj3eIXyZW2Y49Cbog6VBemUVF3NB9Ie8ydZvrebJCm4mZ6QsqmTAygkvUFoe8J2SOpMu06LhgoSx
TV/r4o8gIsnEw5k8qhlkUyeRWpZMCKm5J59Ri/g8EjkcKwT56f0noLJtoaUBb/y0GrOodMBmyVWd
7QMkeWPzjphGacOMjKKz7fJ8/ub78yhZ9iZ5t7kVhOLxlkBRz5lXKpU6XxnaeuXEyOP7huSCyPaU
ByRNuBpR/Ir7O1jfl/dMzJxjpC/feJf1rg8Cwwe8dqpJfWCQvx9304tSBfZkufiiL2/iLxRtfTdP
x2eVp7NK26EFrkuwHOzcy+kQctUC+I6L3ocAHS/GkUwJLdtxYPHSnrZBrGdfpCwOA+fMwH3C9ePa
ghmsYxeIMlbnGFss/h4DGm/Ye0h6sXjjzGYonrAwkcnwUoKO9LRsKZtGb4+EHibznLP8YcWpo2xO
IgxOUd3Rk2Fn5XDcSIteGb6LRgar0nDfn59XMrivcrs0EuNEH9/sRbYw0Puo6ht8jmZP76pyb5ne
0YTOVF1RBAAihdoTQl70rKt06l/MJbXrJMaD6d57lUYefjox4VdjQCQmVegnYHCRSsYgMm9SWbSG
qQsS1xzp1JnbgtrZkSWIuBQfQJ9R60WWS7LzgRVtAnaGcwa1k9pe8edkH7wm5zyt7skEFxV5d5Ba
ER5iXN7DGM+yPd6MjWcvMH1+mAEbj2DmV6Kmma9Jxq+KDU6X2fdj+Mc8rqYSGyQGDZpu+GWldfAV
T1DsvTq69otkaz85E4jKss0d/znz9YNmfp2om1zILkiv52nBhxovPkBzGRrXxaUeKuyafBz/63lJ
NNIaoek/Ste4wFLtuZPp6lelKcWTyBU628u6EqdX7dsx/mIbLUpXvpVl6Xetwo22i41kRtS6jxN/
B2vHCpkZXdt2KsrkHOK+QJgI2hg6VLfzhXM8lITLND9haeuy1Lu17ab8JH8Nb6YoO+/ZrEmhPkhC
5s2K+XzC0EhAs4x8B1TGJ3VJ7Zi1xRQdgApYcbq4lBwPDM9ikuR8Azlwz4rNAnPVTk4zxF/kezZm
DgFJMwYJOc9gd3zQNTqdibHj6lhlA2bwVuUvpv2w9odRqw4XaUmCn/anPkt7AnirWs1bgchdWOs4
aTnCkOxqmycAAUPP/CoRTBpaAdFEM/0YPfQNQegAe2WMOMTHVXvsVysP6jJBOpOfXtRak1tG/il8
C/6UEgLvZbNdABJlI4oiE1/c+QPkRZGU0L1Z0SGsXOo0WMpRjOQIGDBnpkTqZTvJSc4lSdntJp0k
ASelVMz53nar6QU2lQ3hjAYfPzMh1pa4aJgBQkmf1wv2LQv3Hh/aMKmJLWGH4H17JpDR/V273NHb
NnDckQZalnt+WdO1QORyW6leLpo1HvI6RXfMzCzkTgb9OvD6HocmKuZZbgz1o5yVtUVG1I+Mh9nI
bdF81PKbNki+P8p+jdIZn85QCHYHkL+ZPdNOKt1vzKJX7yoFGSswBlIyajmTu9yagJEB7XSTDjyR
nJCW83jSlOjFuzn6tL5/Od6CJGA53a2IhKB0yorSpBU6qERgLVJ/ZVH3nezUtUMdxMWSnIl3Ugdy
mKtcOPcyNRd5OtihRd59oVJTZG0trFbTyH0IpGSnB9GQPqAxO6IeYdMVMLLsvWVYAcsNaFl+Ckf8
ss6Ku+PCO3vt+thKJDx4E3HMyX3XMruRDXE6b57zgtLm07wcQ4BShxYcWnRgrD+rnxLzV5zf8vDL
QN2ImRZ3VbqoxzfTLu8kdIzO+Kw+qh7j+AnmN1gpNWjvBgFbXIjW3dTOaSQd8VH2rBi7mCGDPtwz
QZB+blXLHXT1ZZHAB5Nls05ns6BuMMnCycBWonrW0VFO88txgPnNRVblNED3HlnLlZx1qWo301ow
tiEtEX6+dmBffHW8hZtI8M+rqFajVUI+FjGQjZQ+uuhS+uznTSCANVzuPHFP4RsIhxTzvtrBzPNN
dDLyhO/haYKxclNtkMsKcWZHvUnGxQ2MxUCCtrp69QNTdQADbPfQ3UFAVB41GImz6YDCucpnAjoQ
AFchafclZtujlfQswrXL+HcMVYATu3TlVLsJhh4dE0+g0ZWnJKiiDKTV/faOLzBJGMtZKRk6bGDn
t/z7af9qvaZ17YUUOPrKdg6sqn7QFFhMBbGI5SlaJhRUsXmHW8ASc/HP5vEIt/8NiVfYy1090RNL
7u0FHAWShxeCjl6Gz1q2M89H3oDONU5dlarC3r3cxXRW7kHp9tgQVynlf5qwNr2i3xYHinin+CZh
l6hCHm66NDHVQ/Pwqur181Uvpii4Re9Io8SW6SU1YEh7ER4RzuWLrMNdLftSRFxu/oHTDu/C3vYa
U1BysfxxyyIogDKk71sXDEvTzHHWqeqp4yQGUKWItL8uOqkrHAtPNVPXygmRBJtZ3MyM+vO2M2gs
7UHoIUGWBP6tU5D8n4d6NWHjeB97HLiCW7yvfaJ/V/UysqGP60jBEAW08QZRBMA48WVzf2+qVy0T
YpM+3/AQXY1ThJeB3MbYIkvqmp1HvsTSiocjopZXkUtJx3GuxgggEE1EK/uSzHqWazzvy8FLx/1y
daJDCIdHhr2HrIdDiHzxgvBo+DpjXG1M0hNbc7gS/ThWBvwiBvrE7NpJB3vAYHSFe8WA43GcE30e
1RSs7lMpyF0NWhyN9QBZVQKkZBUzEgC4m+23a7qivUmLptMPKKbi5JZCq6dQ2Ao8uT5lSsUSUW/V
+8BytQlV5eUZF32TUSQ8BC17bidRXGNmoZXV03ZSafZHOxj4Rk0kv1lY2EdG+ooFFr0+YsLhkenY
XjP0ts3LMLzt/l9I0TA+HO+nHfets2EYLOB5xa1w2FwwDETr0MEGhgnWcM+riSxRdQhCJZy0BD84
8T18KQf6ugsIZcP0aWK17dA2gL12Q4ImaEuJo01aXrIn0KqRdodObMMkNooZYQoWsNlt0+Wn7Mzn
l4eS5/wws2+NuXrAVYtXgyPEIleQyMsxOj5gLQn0hsKK401Tmm0L+gjDRxOVmJVItXD9i3qGAomx
kiwzazzVbd04FQAefnIwvflS5AwkAdBpVVxMGqkRJD2ttGRicuCd9mmEbSCQKCrHGQ7+TimPAieS
LSru/ZLjU1AwNm939oAZ8jUtQJXBxsJP229HRbqFLP5PwoElTwFkj1oKrfmNcjIYse7o/mRpHljN
z1am4gnRVRws4FAJ2qvIlxfuV6SkssMwz6RVhF6Gcio6XWzXiQZMKPtLSTGu/fl5wSQyfzde1uYk
7TqmyvcrB265VzMH4cUrURgXNBEbYapmTgr6MAijjui8/TIwCwPuFYUI2VDLg4oiSvhxVdkjqbGn
+q25sMuhGOKlR7n9q33j9OiU5jTnPko7y5HFsUdaalw1qFvRMLXX9vVuJhPzMvkAfXxViFsRj3UY
l2Bb8UJaMNkN6UDfMKHSvpIC34UpnNWYYkr04NMkonZLFqPwN1JUO4eJwZviTmPUO2030/4Psf75
4NiegmWyVPLjuxgDR9mQTQADbhRLDI6H7RpiZUQOAFfW0w1cnkb4yxLvswoDu4HelSfoweivcRnB
e03kDXEOhc6iuBENLRjiLHOceAEnzgqN+1xyoCA1Av0a2ckFRwzmksB87s3JKHph4cofPdIZQUIX
+duReEK7d1uzb8ckNH+WXonD/R7rwwEyoEeNESaOjdXl6KOPM/sWPH7kJOQx3c00c5mGaeG2tFBf
uG5oCIEiqGfYdDJ8UApCBGxmph7xhdvYmNX4Ul+GpxKgOvMwh1YnORAUOCmWLfO1aDefgAPKSc5G
J2n9r/t5F05A4lTb/omKPW/gdWcK8/Ei0tq9atclDocVgNkO2hxil4b5uct5pUkpJH0FBP5pgBHh
junQeegB4Tr3tyUOmp70WHyOC7563PVzm+z0nxDOv5mzNo3HkA1anWzu5MpfTvNJs6RiQjwAXAof
81kjpCkE5K0UYbaYi/MeB6obJeqll1JrjVdx/XjQh2r5H1ABO+74risBeyX0qh7t1WvombKRJSDS
+JoGSoZbMq494TU7iNoLBG9qVKJgSct9iMbs/uKQjPXe5ZiiBfrG+211bKt2eYhp9pRoYxJy6I8S
Pg1aEuhIvEM3LbGuYMzxVTE9gI8xwWR5kp9wbWMO1SRAOIZp1lZaSXAwMV6NA3J/36GvrimF952U
8e2ybDQP/ktwQ9aPu6ap2iruJdXkD/GXMZnXlJws6zdiZWpMgmIHk7RHdqMtMBkyWqPm80Y1nmF5
HM70/H+Qb6uv2PryN2Oa4A+7c0tGxlWJQX6MVpvyw/zAcYmU89ShCYaAqiQAW13Z9YjveyAgfUc5
aWjouodDTw89sfo93h9OQZDjGxupkMPuX6E7fGDwYUqkxtlZiWfsGbU0pkOF25pMJjnuzoGMUBv/
iV2osUDJyPSnIIqMKlLRMj2lTHkGvkafkHbY4BSf+Q40Y83Waa9CueHriJqNxEVaAUa80SGfgA74
db/tm8E57PB9nCB6I5VVGH24G+fMmryyRj6LlPbnAjYnJDbdvuU20ROjkQZFe3qCxTWqdVM52Zat
rEG18B72TeVxSj6Z7m7jQexRY2tjGxfS62zAqebSWEwrxMALaKQPHhtwj0n4Viso2yoFbAmMY3ig
d2fm1lxpnjmziZRmF1C49LSMqCvn7WxUZ4LKxjbwU39bJunCQS98U5sObR4ir9RT9YvwYk1lzmzc
25hJ9rV1mL/sMqkZ1RrK4zqe9uoc43ofusyMeQjIfDmcOfwR/G1KKAyuOo7QFKaT32KwoCcjFuYV
rpiVzZIPL7SKIzrK4ZqB1KlD15SFXvOcDrey5JxciCp/06y1SARXSYS7yRcr7m2iV9fKPhwpybQ1
8ZKlUCUhjPYumw08/D/gAE89HiUzHpIYja6YpwFihzVjB8BkaF2RQ6yh/p8E6Tu2gQd+JfafwcW+
+0dYtYmklHoA1vvgF9Ez61CAy/Qhuy7OxKY7JuUmgEzpZHZ+kUVB55Pzd0TwhBCQDnL3LYh/DQZ+
POc33TL+1yA+1nS3RXaNO4K1D//5D6lzG9IYmgwofDfycEXz/aTqUWaECWhC1yTZM/Y40SYH3LkK
hMeL6mMtTDzYL9CmrKm8A9MeZ1V4WjhgNv3WD04YvWy+1xV8Vkh4VkuCmEr2WdrzqBemZpO2w/rz
nL6RZhOuo/nsMb5pesG3yRgQiIWMlj1t0fJSz5e3r2KwDTTmTy9MmMibDEDLm51mhFTdG40wKe1L
fnULWFW0pju87wNrV84jRFa4H946LIZYa+20aSD7kgoUUn3jl9cOPhduvutEUsvS8v6WxMpnC4Hd
2ZOiFE26Q/bFTLDf2h3GynxD5P/BkKp32398mxVDh8y/Ffy6wnsfUhUaR+0BWci9IIX6QDiwLzhx
KffdYMIUjZtCTbYDyPxp37x1qsuw/EfyFIBcbGXIWrphKRF+Qqz0/GgT8H2kIDkDL13NnrPK+m7Q
il8FDkebMdxZqz1eF2+4VwHQQICjN6cJ+ALDlOifuN08aJV4onmcIHINUpRYXLZNEtukA7FsSSko
EwMmnuYpo71+pQhjPSa8vVN3Awz/soNZedK3YYfJkTaR9I1/h0/cSf39owa2/KILnQ6AjODbiTUo
NBo4U376hLEcrKD7lvfPZHoLVMQbilZOgUrMDEjPt04KlZHwkK3FFLa0v4Z1EJq42wN+PK2dwnuD
mluyeAYj3KGFALCEKuPvowrfXgSZbB4oSfehS90BWL1t3wOfYfIxgN+jPPVH/u5ZB5YED0/90jwX
C54Sd17lY+az1EUjD9usX8q8UcNrNMPIiIZ4wPLh7dMo6v5FiaZCsuFPOQMXKMnBnxLgsNZWbOMB
NLEtrqD1jab99JRBwW+JXupKTL6RMX9sNVyRV1UEAkLxzjWU5MA21yMD/pSsaQfpl9m3yCsQ4H2q
m0c+QJf0CjAMoMiOrkEtX9z6m/iQrKr0lfp5t0zqMaQ7T2Nrs5bnSpjly0zVRmEKvU2ZrLh4E+MZ
Nn5Lp74LhlH/GSVDQmw3rIUCUQUGZ09AxLFGjGwXE26vAghoekCbmgyVy+KWYPJRiAHLc2Fqgp/X
q2ByZP/zQRfWYUo2Jq1raBeiKkMHrAZA0vp2qUaQ0NR7bPudZGYDEpjvH97pyw+0HgRjPE8g1zHm
420HEcFtqc0ZHhlKNq/VxZwbf5jYAn79jlOFxKpsSomMZkQS4DT54bPwPbQfdRydm4uU7FRPMaOb
kFaHLsZOuLhF2zy1P06j9wh/8c1KfS7jZ92MSOOAmRtUeFA1WbZlQPiTLP75VoQMwL/nL91kCHy7
wn0dJ7yhusqPANW8eLIYNtxCWl8tQvvWove9JE5NqdQdCoLc5Vew4CgpYQYvptcxFXn6of5Pf9FA
5slVooT2bxCtlQ7fEqtEHQDB69onu1Pzmf15jEl4VWpvdY5rdWhXOzRAoa7eZanF5/QlGJcODoJi
+cSqyUmaOl3t415nEe9g/jarPAObLiAP0P3MVo3Y1ID2H1vosI2sOxT4d19xQ9ddH4EShCitooQW
+5NA+7YjlV4NXE3nfTrPv+N9E3IJU+SH7vNX3rYtJlJFoJl52zdTLj+oQ6oNoHppEaosdpGHXPTJ
ndBPptb26fHnFFVbn4TsOE/hxvM9CviR/YqYLEHqStJg9UhBMd9xBjGF568otVaHQ6NIdHD9LCOe
olG5ulaUOztlYsuQehEpNy6pkm4EBA42hVLHJ1H/xEdj5V2kXdv5mHlR1jwcLTWliiUyGWxBp0Ib
p+YRx0CEsMFVcMIMDD5onabZTj0w/3uYhY360mZyxAFzkxDYwa4fbF2pxDtiwEDJxk508a1XYphU
W425cUpbF/y/bx3ROTUmyyv/w41OxCBjBApnPs6Fc3XcoB01+ZEWA2b4tzvzz7DKtGoKxhTKEuUD
a7ltsu7tJ5cWz4pMRTQOOj4tCPm9+9mpfiow8dPAPqt9URsW2xpqTA2X9dcAdJAt+pIFcPADhfis
dU1wsCpvvetg4w+JSoss0Zr0HTbibXN0YHf6MXU6OB2UtbZOuaQFl773iSnZ8AIkXdqZKOnUwcWa
CNAKLilU0kiuLnjaKgntkKKc0a5tEx63BEaXD/HsFFZo3OI4gfAhE9fY01tlEPrGq5jfe9TF5fzC
lnOCob0WV6+2Q2nkvLa2CE+GX7dYOfaJniBjSGZjANWL5KZ4bEllE61J1px1VyHPigGsmkEjxFpI
tfT3i8oWH/32w3fsfM/1KuseiDmB/3AZZOXyKCW5OuqAL4SZNI4nEdJ28d1gNV0GxpThAsq76Q1c
kXm0MCJhNKpN1ot+9+J+0ZY+ZgaoBqLL2q3eAUJ2ofNTBV3ZiO91Sv0G54ECVhmD/Mu2Ms8u/14a
U3bXWInZi/M3/XVF+aEac2Hyfsm7eXRPWYtuIMftxnAn0JkpufuoDQfjMSGfnyl9lrTLiPyOVYbo
yMRGoWNa9B5iJo7hAIO2J7Y35mdCmLE9NrdhGqQ7CW/AYEc1W1EkkailSuKA2XjmRE9Lq/u75q9D
9+SXO1uOylHQ69P+XdHGndepcj90osb1rI9H+nac6FGwOnUjf/bzfGP4d0GriErLJjYPWznuwqSU
JVp+jRoUB+Bg6Oj+CcWm1Y2bhvGpdylr0dQ9HKoMW42yZDv9AaqlhFQNoP0qxDJOuE6lINQ4pdJ4
IHUscImaRO/JCQpI0DJbr7LqreScYF+85wtdKgfpm7EBhAMEIwdgzqIAxxBAE1kqYRBRKw46ioLB
qUQuinU2sq2LmvHxa0U4FpsTbyDXXhZ5VVuJ3IeqdHXkizgpdVbdOUttO/nAV0u8hbQrQ4xd6oaj
HjGGaFRhLSVmTyxhIa+z9Gf0yAXru2UUNdLtBGHNq9oPPyJiPqMPM8V26mkhRbE3pkxzjJxJUPdR
GkSg/4YVkIGjj52Ea+6UfaQhvQBqaS1ifMmPWsZ+2boZslMauzRllTa2yH/4ULaWCgbhvYsVxmX+
IV/WtCcrHwJ0/lNb5A6ESgWhiQu+h92OYyxqho6YkIPQFtXGAFAGNYB63vtR9uhmjFDLoqX86Sn0
GNNGTMTvwyIkFY7HBceeNEO5TIw6EDvTAXfpQ3CzoaRpQKJVHPWqHMXiMq15MqoxHspPZQKb+7sl
rUgTxjVafETKRbQl6O9eMruSsS83vE2Aglo/5rJeX9k+CDoxGM6lDWXFlxCoF/o2fidYdWBvdmyC
TvETpTEuaOJ6JtRs52BHL8ygPxiDy1HKB5jEv0DP/QzwIZp0jSK43Jz9O7Dg/vjCpBCqm6zNNncO
W+CX3nmeBeZjk879XmCLVpXM8y7kD6QKggiN8INK3RS1eOPFjcwC51JSJQ/1dd/ALy41Ve6L+gZO
xJ8s6WnYy79FAQfE60hqF14f5hG2tGNnb/OM4B90j6Qk+QdqeAVWS0kTstHBkcdjOxc5O5Yt469N
fIj2w02Tx2PttkfYqKIFaYcCON/T+srG0C7nEASzmx4R00+tnVc4BuaTvJ2DwG1WQmFlwkMzIZ36
Xvc3fM+ajAgFW8tifCpG62V2lrFuIkUXhVmQcjT5GlEIKzS40iNh3eqyOA20mozFkQgXZxZ9aC64
abCeWhEyDB9ZBznHwYuAYMGv6w7tBurJ2F6O8Sr55fu9TPwJdjYIRsK3mY27RlbazPh08tsMtIvI
NE4CXzslEqS5S1kxpKgUmfDR/Feh8b1lnRI3QaeNhBqQurK2aoaMLzfblxRaYaw7cxOnsDqN55UO
6yw61tRMt8HWFTQRoUS45UKPGRaacBsYbuPsIMUsx+6qHpgpaVlskNeYjNzM3Cmg5971hvGYkX/w
usGzHD9lPhivkJMhOahNrAxBR5LTQ9UJyIgMNipYeyndlCs/c4ArHnZoLzdBYcfGJUypNkRbOGdY
9d2Ed4LXnIjSK1Gc3fNnF9fsX+Ux0xVdsFM/BjPBNOpkIIDexe4PwyamvZeUAn9QmGr6idD/bpEq
DoRwve+NouMS2rGNP7yQmJAfPIr0ELz6B3Mm7PYjuqWml7JY/FYaK0OXNqTkddoAy8KyEexirpQJ
b3+qrWAAlfq9MiRLS/XQsIumRTCfBtFG/Z5PISx95TFZNmEZeKYbh9hxatLO6gNHwZ4Qh60zfrKc
hzdmGhX4dmQzyeIHNFKgz+4CwzJ6wRLxiDO0nCqv5m7Ow+tp+lu6XI9xkzqgNdkEQVFfAHtzTl3j
b8u31sG0f0nojXyDdazkCal9+4Y2yvaon7nFgaM1d0c5CFf6CXmp0w4CRA3j5m/UOW/i5xZkw+tJ
jpjHc5NY2WYCDLBxle4tRfhs3P4G5CmzJjMa1wzpybZBna188zVETRBjtQIid4nyVMKneDLXBNit
7OpVJvrB2B/A+4+s5PrFYOLgABzZfcn5s/WtkS5hHLOd1pII1UwmJnCYAg2XDJH8buT5L4zfkpEe
LFz98u/72LNM2q+kHN1Fo5wpWCjUcI0aXu3sPqoEvv5gW879uQkgjr9mCSZP5nLI5IT9cob/020j
CqF+OKuzBZTQjvb9V2If1qKX2DIqfsD6l/8nCnmgszkIGWASkQke1WOsNTKCH+3uc40/pva64z8z
W/FihiylCfqa1WJksM/hE2pwRjrmNo0rKLLO3f1UKzrDLdROtf2QfX2YHdyRt4ZaVWZ0VJl98ufz
Pa/hswOlAPtwFX6+jWpKsMFssA5/4PObJbs0Wfsa7InmZ1ODqWFR+aOH5rflu8sViixfz2U2i+je
2Dz+gGK8MkwpTgEr4+X3K0so9RV0EiqamVtlu7DRzq4/Aut3yPPeJvlAbVtgutAp7Y2OkkfwboQK
7k8G6ghQjrEVi3j82xeo0TaJAZ2hsy/gsD6CZxZMzjPHT0jBia0Dyg76+cZXaqGS4XUQ1Q0XCuxZ
x3d5pAju6ePPKz2nCPGQJWckF32zlunWxYa7oVF3frQkIWMnSTB/lBf5BjOTiVTPodFEHWtPY+w3
7jRVy9Wtk5+nIjPvok9BeEVNVZBrca0zuVCdGS96657gioUuwHRRWq2p3mSMyVaukhigMcSE/xHF
Kf7r3hwk/WMqoeEYLu8d5s7i42OlMcABcrlIwm56dT4kwRPvDkGEpxnpjgz4D5ZEta4c45S+uXg4
vPHbKeN/di9vg/PhGRdSms5kn60JnwmAi2HF8hhGV+zSVK6MeCC9Y7+qMCG+eUNXuTHLCoDLosvL
wp+wdPusFTraE4NhaxrVifSvWJRUKEy7vufmOlkbHUo3ugBO011H4kdvzP3JyBtqzr0/k13ZG0eL
nIn873mUeM3/nICfUtGmnP0lpwjRSwT8m3wC5Z9R/bDfpOFrQiw7VjvWY96tuIe3v1+54QWKhISr
XXswjf07JlOYAPp80aDrf4nNLJVlbiS5AWP1n2XvVbv0WED2DN4EJbksDO2/JNAus3ZFdwB+TZ5Z
ZUvzDmn4FaNaPezKx3hPt+DzFffk5tXJh+JwwnRowNSWTul6pWWFCQT3d/MPlOrBJVB4gbcNqI5e
dNW64IXpweBwa3LeS6++WhwACjaWeMvQWvJfktG8t/56QT0O+ht6njo0pp7uWAX/ckWYZUHdJHkZ
ly9VV3rNiEob40rN+xb+ioIwOXcZ3UsrddLnLWTFRaPZs9spcjTBZTapeKoDGW1wMPn06AiFDc4w
t7zxY8BxJ1p5OsCqE4vAJDYbpbu0qaRCLQVP/rEcHOMCfwBjJKZwGOr2idX+XWOPMxMAoQHVerb7
hRXGekSnkSxPonPVBRW3ixX7W9ZEbxeX3Q2538IJ4tRGUY8ElNAkU3wvIdnm72Ig02suHxnertko
sTbU7q16Z4S45QXfUfbN4YDBKcI6Ioz3iMmEK70Nvfh7LjaxNDgY4xhDLT4IUTEjPHudmuOZDON1
EWJFfQRPdCnhJ7QLen/rouSwkPjlDWox9uyz1ZCrw2YxggIBTc1Yy4M67NgNj4va1U61qUX3R8mz
B/54iQIZMJI5jWVIO7iOsJW5mWrkixatn+bborJzsSqS2d+gHOFMs5eW2xxQY1FHJcbmt8GdqQH3
SEgITgL4/sMt24mS4lRPuYCueOSLDEfiAZifoYqPuLGLqibZPv/j7lgu8Cvvtxe5jH8BBTsmlDoc
LIR9SRe903ZCd8gyDj2vmeciRqSLmteZfD7gwYNxXAtqnjcwqhmkGgMJrxQR3v6x+1yugLBrKh3h
LB3hD1R464sWi427nKUQQXTaFeGqv2S2TyOhBlAy4NIFl1swGX0XTJz7R823FYLasdRcNKmN4GY0
jwzYT78YezRDWDBtkCMxFUZHI4tfSb0kC5qcIGcE2GoCeSqeiVB1TUgMbWiF5E65d9uupVjYmI41
Jlg6ESZU606RHWs6FGuNBVpo0/ifmhPkk+Jw4bCQHACimJ16JiSt2yZUfKa7K+pDN8FL1uBhNLfo
mvD7u+G2jJHsKtCDb5CgyoBJrHLMa57PbYC8wqTO3HGCSFJS7/iCrWztG3b/in8ay8lV4IUjmkxB
hOb6ksPWoruUyEhkTbNz/Y8IoqebX1l23IwoSPuXuEsh48PrI+SCDsLh2xbtKwUY05LAtWrSOv8U
W/6yMzSLEXZCDEPQ3QDxz1PUSyOMfQ0l6wbZsc0x/l4/quXn74OD8dOUje9jWKbuXVtc6A/LyUPY
KvqERKV4tw+szKDpXxV6NzH57r3B3Bf5aNWLqd6/iVlRzPV6Bk1OROz/+7zR8Ee4WDGgNYZ3fXdH
kiAUsDXk0UrjX61132Oq6JqcKE8byiLodS1vHVtiwOWNa1eK2kTiXf8LmHV4svEV0FT2ORM0ZGBV
Dok8akp88rAfevfl78cQ7lqAUmRe6KhPwNSvuQf85ctKs6ygFljUBZc7tJBZtvrIMIXImGWiKHgB
omHpL7iUzoD4m2RL/PoUD5Ka4/XG5D5Xcpu72GKjfcBEI5pXlVa02hMiBRAqgStU72muZdo/tQbb
yAfYVKrQQ73D5e4yhCDipOvilCjmFaFCyJ4S7/co4iEgooGmDzWYLe07E/aB5sARLByBu2Py1DD1
52Lc7I/2bgeIjGdNdBYDui31R+FYC0NGLjI+df6epjDe1IHxUVp4RZ1MpuOMY998Gfcu/J1wkDKt
Ksz8wPdXIq0Sqv9CSeXtTwLxEXggDHkJShSij3rZT3yiORGnAL1aps1Xrydn2Ez/SEeRMthM4oSa
3gel362iZdqRMvvYJYiU6OaPjQptrddIRrBuITRftd5/yZbxyIigoxpkLOHmAE4k7HOyf1TVMLE1
AqRQOGxw2StlOgRLlOj/7GnjlAodEyZw+8yRNj8jbz3C/X2Ap86xa42l2CoNpW/OC6oSgR/OgzCf
oIktmHF2LBu8M+4LEFSl7SJMbvamCs6JgG5WI/6UNLafZXotxemeWV5SFM1N3XLgNtz1ho9E8QON
49K2RQyA3VEMJAL/RO7FciAGMwkKkLbaFWoZePwZ6mqF4+0U/tBrEUPh04wEk1J/BDii8ga24niL
3fgxDUNtW1zmCtEy0rRauSIkEjeTZAekJpkUYdonP2tMpvktHgJ2kWwacFQtxrLLPb9MaVH1JoL5
A44krot70FwymgdvTI+/zGHWdxRI8HtC3f9t1TsuptG5U5zqSxE36w4koqKTTQY2T48U2Q1iwNiF
ackb9LbiUbsWwzIRVemTxTue0AJ5+Ln6+GlhK2xehyUGfWlrFLOI/44Xcua66c8AYNkGFvyVLW6w
w2pjKxNJVJL29uWaBhhoUbput/u1J2O6pj3YVVKljD49XnAxW1tXxLrFpO7945M9JXfeL6ZRtGR7
oyN2iIdov0k59ksC27ARE4GStI/Rs6FV0XuXBOiWz0cH/xjhoHJHiUuSJPahxLPHjPVTX6xJXJR3
xVDfymSPYOtuJOEyDg/3XE4hiuCzsBGhkrqAXx3bS5T9y4mz0QLkUYN42e6xO5+hUJ3zsbMDc6Kb
TR3dEhfOK231NRWZOPsxBDIZnTs0y5XRG+PAaE6i/0U2BFME6frSXsqyB1CylETNgRuhGaOdCvAo
YfHyu/PvmXY5qxsoq8k9ROgwMCQg9x7l/oq+yUlCsgkVniXCBlKGi6aCriLYkA+98abDr9oUPzrn
ZTh23w3+C84P5ULn44qgloNISAvwSgyHnBhbv4qlwQgRI07ju3e1qLnyRFJUpsEWkrWVDmemyjeg
rso8EwEEPaYJdoDSprwYubLAUSa3oAcKlojjvH7dXQzV4ifXVzjweq1iaTkdXLAsita8L7N0KAtI
JzTxiHTIMeYZcL2p3tREe7jQwATSABabeQxYt2fwzFaSxBtHSe2TLlBAvfBX16IWqtiwK8HO3RQx
vbLL9IOzGSCNt0gOCX0NpJp4hlQDkcGlaBLl/crIvCkIlieF1pPEkoCpWME6N/kzbZf87MPBCG/N
77D2Oj/co40fFX2+XduC8O5ELUNPPPIXIEh9OOg92V8zWL6QcrW/IxKr6+SlPkceh3oQD8N7FEKt
D9kLtq/Z4YLGG3iZnyZ/geTM5Nj1iYSfadDnsJFBFhCWo4VpsvHtzqiWhVQtTvivqLsmsyo7aYXn
T987evJHxv4aljy3bed2X5M741lzvNJMloZ3qLSmVcKzqlD71QW9zqrOGJjepg7J2ZBM0hdShKUb
MSFtYYcDLLJTrnSGsikJx12sUIulkE/54grcxRFRaRTrEvjyDoLgzlcNMOHti3pZm+PC3cuDq8y3
LUV4OHg7krz/VEGzYspaUsKTjH/AG6tg4a1yL36Jk6HggRT8CqO07Vt+tkoHR7tnr2b8KzNcdNND
HiSoNGLao9sx5IE4KXwe8UgpQggmDIT1bi5eOEIIjxkcVDixS2K06JZGbAhoffrPXP+mvN3lOTkK
h8a3AWj5SfJlbO+DfnDnCVaXUytZphTP997PGX5J2es5QlS0Zd2f1fdcuYwGIwKLfWv5TZHkfc7R
Pv6P0TH7z/xsEP5f943iyANKv/YQsUb3F/+aMWrl4b96sb7GJp5sK7CyMbjXesg2KZ7Y9o36u8rD
JBrXk1SsKTIqvvD59bx1i2xVd4cq0lJK+raIuNR0I7/j0hdXjhWkSxr9m+rN1SLPvKonra2rVONZ
Byd6xdrdJiODqGCnDji1EqxWpQy5CBSmzZLGUIpPnDFPe9+gks5832SdeLLTIpteJDtOuLspLR4P
v6noqjS2yIGvLub/6dQeKxEBU7ilZ1h+JEZNNrUgOQ9gdSEOvZgolnYZLOUGVxLy9uiymLLjwGuJ
eqBpUfePl/dTwLmRtjApU/68s+UCJcgen/5SUItsr1rBKC79s2/1pOpCCrtgJ/209MiJVOjivcY3
tpG/MMjuynHRCdTWAYDjpg1VW0vY6/v0un/JaXz454LIRz+yomGFEJ7PSte1ROrya57HbjJgpfWG
xbem9A/TB8dVmjk7qanhDsCBc6XYIB0Y9nflOfnKPCXZkFMtOtcAcB5l/8my9Lzz87dkzyfxU+wJ
AEgjIF4jYyXv560CzqTEP4usddzaAq1wwGICai+D3LybSeiEG5CQqJLb45/7E06ilxO5S0odY+s9
7bDPLOu8dejZAWh63emTBFjkYK+PRXE7tCqxiI5DT5jb5IYKbzE07/QgzPEPy9M2NbeM3Lja8lLv
baVxM2MOSsgCq8/E1XZzdpYLQWHWDeX67I638rerDSnBV5D6zzE6VUpgn3FnESqv7bzltxq/TkFA
Mue6ABnhhbe2kbnqzXiqYQyKzeeGRGAUCBkqs+6IvV6EgD8OGUZgJ1ksFS2Rg++zOf8m2aybYDyU
Tq2aJNxvKieUxC0gXryEw9V77FPJdd8Sex56cWvLdUW+rYVxM/vQbKxdxIkE3wizQvMwDzRx4vtC
rIcSOmFjxr2DOGuvxsLqdpZKYfyXq+HbFVoR2mnr+NEAejnlU04LJYGoeXYzjTAN5lFRlcYDWH2g
A7HeHZ6KOFtTS/UMo1sutPR3gTfeHqLTquT7U4SuL4cYtrgltNpKsZtqdlAyNW00OPMneA5wjywV
urpVgjf2Brs8GsNCARmmT3p2WZj0giVY4JuBfiX2g6FMwaSGt0uRQTCe3SBFwJgqGMYlFMQanuNi
WR4zAutCyCsPzWz6ykjy2E/cjqTRty9vbfyhggjG7LQdR3ROnazQ6f+ycPBKpf5bC71xBjvv8sUH
kZZViTWKPdWJs5d0iT0oVkUh3dsu0tuw41XGgIipHj/17K+cJiDoMNlQn74Bvk1w4Go//Mtb+76l
fpBJ85VGYRyOyLgNHDN0vruw6HcQvpsov/fB3ZMZmDKcLy2UllMouyADMn1lLeLXRECu2NGzywF8
da1cfU/xIjoNj3U5jrsLoTAVq24Bfz0jGq6OGMklcHf9KdV10TdYy8wLMawN5WWDAwhxvtg/DgdO
qEjfOx+EVTdE7I4B/F+g1/ET4KMJOADIKIF/K9q5guLqNzJ2sogf0wk/ay5yExb54DUes2qm/UnA
12l3cYhpg90fqGDUX4QMeGn97HcZEf8/7W8h3btZpsqC54aFwE8A016cFEAjKhugCj1zLgXb899K
RbeAcBhASxrw+Ineb+/qPGtafeO/8Fpj6RegJWWeQzQiJEJEqgCF43EGFqRQf8m8gcD4kGKUi3rF
Xm3/ghioeP2FPavorvJC/9saPG0ATSy+A6h1QhtqWPOJJCIvBRm9Ql5uiY8sLG6L+hihyDsrY839
ZLAZu2vBsOmNP7U59rkbm8fAdEG/EU58LIlfPZdnCwEjNinol+naitIcujSh83tZY65m6WIz0usl
W38tioHu/8Gp1AvZXF0A8m7cCbslKu5CyyYRnjUTM+nQwhovlviwW9ABL3QWtuiVv/7AXqlev5Jo
zu7do1iIW5NWxGNkF25yTrvkdpxGrwVJxRqOavOyvNNOIUvCt92o7bSshokTJCLq5rKrAUNu+4ch
6m6wL59UAC6rrzjduiGsFUmSnFfGR34R1lAA8pUjtQ8JOhcHkT+L/pvYHsnx8MaPwyV165IXJtey
casVud79DXJMKmjiVuEIxty9GWj1uctHz0fNQqlc/xeuZ/7mhCTs3iM9idPjYe9M1o1H/wOmNL+Z
8F2mxik151ROIwoLFEbgNpDx73qRXNWcYpBQtRs4KXs9/oBreSHwSaYJoOyTbJJaLKY8g967WrIr
8v4vWsYfZzVPGTWNCslYiPcbKmhqM1MPx9JTRwsv4B1Hu8kQAybg1HMPQtU57auwoI8Qhws03sFM
MiMUkYMCkfzcKAZnbF9dgMM1MEWdMD8sL0ViiB57lta0HmrQFwPOzzI7CiWxDMU9xxQwh7d7yNh5
5dROxj/GGWOCQkkt4XhsZReiefXUtSdVOSJAOcYChzo0WSi3Hf2roh8sxaz5u6KbAO1wJlHXHkVH
2SP2JOeKjZsBtv14YN5G/MUBeN2u4FSgnMjCYBhkgIzxfPSb9SzKNRnJSD67asO+CHw+KMtkghku
KCU6DffIVY9QN3Z4FYz2hch9Bpy4SuSRTi7q3NOi3h/apY/FhGxOfaB1rm1gcjUhJQ/Nj/GpkAg0
ec31Di4GH1OGkVQI9DSsEWml5HgJgQg+Obv03QeXT/+lI8FCcu3SbMKezDE6XnPRUyuc556JMRTl
+/HVgCVjhV6xRUMjMiFGuW5sCLlMSVDjUAD3A6ukqZTppW0GqVX7qbw/VnIG+2nwVsfs0rSbX7U/
GI980oWGNDvj1CYi5DZwqMROerCFlxpanpSg+eMwuVzwDaJuUnlhRgBapp+Ok0CJy6sZ3slbfIeW
1vQsiXyyLUvpM30ufik/Mm4y6TVOd6c2sKBGJhf2k8S6RgXA0pehktbDbhuHahRLEqdQRu2amu95
8xBiSmfVAP0KbXuT80NLhawl6mqQ8pr2W+a+33MaIdaOz7J8RYwvJVVATgEHF8vfk3UGo2MVtajX
8dZz6GqyUM5/ICttrFKlG8qqBQ17NFhO74IKzq339SfWwBqGVQDc0AjQ6tRDUsIwvKen3toxBSOO
pKsXbHOGzJbDzI0w49VAxrAAewilUePjKBJSVQuiC/glnOWb6qzuN8CFbsdAecF7snw/2mdnAgA8
K4nAhMDTr/4k+p/yVgvos3hUb2TuqMbeGJSbo/M/2u24lhEqtcu+nazzGde+JGH3X9ct8Jz0A9a/
74C+qfJYwy865idAcioVeUv6BkP7VAMrG+btKW1IHwiUHTJoTCQeykCRJBaujUekvhKGkrhDjJbO
8+KHdE8N1w56RfMqSpOZkQQZmPvrqK5vTj66f+BabKimkOfthAc3zxr8pKOjLAUUDlD3CctqWpMn
l43njoA3gWzv5muHDHw0/HI2/w9YGwbNvafOs6IygGegs/YZURk5dOPe2wkeWu+zyT3LXeCzbchG
kBUzBjASR76Gc+wVH2OZ/QVHFHbnG9gYBS4yD+JBRqYWPNbihIPOFVtuhmDu5To5xPOTu3qD8ePL
Wh/LfzC5+yIAwfmkBmJPpxnOT19fv2dblUJk1luMaVdzEpIzvuwzANYYbh2fJjcjvafR3uzPF738
iQ3onsSc8DrptxPKhtaZzchnG7LAn27yvc1PrQtbywLhnst5cJ15Df/uCIAzMSh/IfkEI/CjMlHI
95UXVUtOFsbWTqPoGYrPH1c/neG30+zB+jEWDIOhm9FNfHQwvRE9YElk7FjEeszhTpsng/6ZOBdW
T/8goDJRv0vSmOvgzW++j7ZPXCVLZtpL7LDAkyr1YMskUTXfmWl163bY5dKh/Pucoh3FaBUCmhVj
SSajeYBsDdXCdva0Uv0M3JWVFXOFse2lPREjjByVVUXUP/1/WH1sU1pQzV36b3hRFfttXA5klC6w
krva6kNlYBQc32GsvKBOcnkAxIi8/ZG6Nca6+wQjdgBIpjxQpk+atfzKsbR4lkzXmV55uTgEtECg
wppvUUUJiAwvnAtzNOCHoH7JmUXenERUevgCIeMqjmqJU6/NpOuUJf/pG707hMAlbwNoLTUgO7Iv
RUCFkrD5n9MIHYZBUTnC9NEM45NzWPNlKYKaeEBfhKxO6+w4AGGT3C9/huU7A7PBm7/C2i3+hSzH
HV9poySfBGkGb+Al4n8A6BdzAKAuIBOyNlZI/Hlv2UCXwh45unFVkgWatC9jQXJ2s5jYK4Skkoes
hh8LPBgU50wuyjsn0OJT6snmwCmGuZC97p5AvnyqcXX04tSeiWYy4qlHR//oT6+5S8OYjKflcpFq
YucCo8+rqLwAps0/Xc87NcbVG1EaOIJC7Vfw19MwLzPkVxC53rGeODanks7Zc/OD/CySrep+PKFt
SS0JCc1AP+YGT87cPOCWXInEr0rPfLl64JYe+yxxj50scCtuQpsYiKeyVTx8p6f/70p0kXetL0Nd
YLd6H7owY8KUqB+r3OaTS+61JI1bTyPxuFEImU/A2D0DqtSBZ8n2qmC9U9qzPUE/7ZgLVja+miAa
65nas3d+3oIZunKBWYJ5sVnxbiz0vpiRjcHQHfqJE6hn9TSWPFY2HgMh9JW6l1uqwRpbVwXNl7dY
YEQfTfzUmTL1nGsaTOawbn0ygMkTr2VlYG2f1vqRbK18Ud3pNoO5t2jGdRQ0V75PJ/14jPoNZA4c
u5eMSIGIHioA/kX8dXjWce8h9dRMMDKtmGx8C5bEZEMBPpet3tBc2ehjkP4HvpykccnhPFVVGKPJ
do5Jdf0At2cesLtn6Byd727Ua0eU1GVk2lMiqUQFQLVUjb5N9UtNHknOKrNDwAHD04LOnf7JTb22
J+S0WF0OkdaP/WGqu/CGh+OAME9V/vQOUJsriLSacLNt1bIEFI84B9bzFGGLJlbRk9tswuymDU/1
tw8aSMp9tT6KXAipUIeG31S7FZhOu9rwkdSn0dSqzBdx6qn62VzjZ6w3zL524DL/BPJezA1gEr5v
/tomxItgnCkyKirRReON6gmqil4f3bUvuPMnYKx2ffJbHy9RIzMFNrnL3W7pC6Y7LCGHnIB1TkWJ
Q9c6peY3i5h3g3vQTvb3UrcS2dba0aVazl7ByXq4mZu24zNOxCxDPZu9CI9PXkdlUesCbeYtK1FT
vz9jXGl2YIcwgfoE07CJgbQG46fR1cgN4Nz2WfRwl0mxTEs2T6O3kuP1lnWZJ31LtFKvlgF9NKeG
vMdvWrDf3rIlt5S78k5IZMK8UzE28RL960hJ9dQMX5sKFCOJrqjjQBRWYeEr3ERxzpNuSJcvC/xW
KVCwFTM4S8W/uD2X+iQyUsK7cS3SQ8oUPXfEhgpLIzkw+UC0DI20wsNqp6foUyeee39XWlPvO26a
Mh92Q2wjaA1DUXfY70dF/u1m2RJxhCRh6U/wZn/kz8ey/LleJhs3hBRBq61lAAYc1CSCb8pzAyD4
yf851xRi5eDorjqWjLyhih5Vx5ImQJzZBqOC9+b2wE3rhpfB/rVMn4D8kbD1p2KjLkltc4BOIrQ5
W1MiwaR3P+vAj9HTeLwzrYlVlyHq+BuD0MiXT23ebVKpg/jpQMUSNtF7uPQJ2Bm7sol/T5XiUw1V
lI85sGg2PuHLRTqmIrOwXChL1XPO7COdtdL06Sndu4cQPBnyoXJV9sXe84hioy1WI+X7Ccwui248
AOYl61flTBefp49II5Kh5qh/XHBeFRTJUGDo+0m3puO8c1AeLhNPYKLlW/gL/CX8zfYyYFeUbOtZ
mYa1+M6ZH3K7ARzMvMEVwtYKzNRcm9zG9PzXb8jczFg219yv4X9JzpGvroKr9eZYy/l1wyB/Ukga
B1vK5y+SBlUN1IEBdCaVr0sOID7T7WrMRWkneJJPbpYjxkE3jrjjiKWVz/HKbvMOB69nudCC92cH
wO9W/xZhSud/wEsP0rR9YXnNkCAFVmw6w+j5M7WgT0JcZhkDjk33nWIn77hKKSChig1vZfLJ6mQb
uyt3AsOjCl7N0mSr2mUNsN9SbrmsmzIwSD/r0BsJxP6qSBF4GzICzP8aGJvwjMTpA0rlzLVcr4E+
nQDRiYbsbqxQHliXWm3ztbGcKn/cH2Blh4HA5Y5Kt9BiTqHGbvwvm3rLca6tPtSNIXwbxz3DD4O9
h8bnfU9c0qoMHnupsF/IzScx+2YJgaRDgkCFm5OIc5MUhX+pNNPlEm2CwEFU17K/mOqo9XMnIv8m
dI5dgRuSqMgF9IyCGMxJzXL3vTPSW3M5OHkfVt+6YhzD7vz+wGN5ABhdfuoDH1I5er68pH1aL+eS
l4DjCThwgQ9Tg44zgmJRcjhhclbRzVYmkCbRrvI1185fEHm0cw21rpbGQYYlRtqW5kyOJC9Tfza5
fjovZhZYRUbKuBka4dD1q1smxLCqp+mPhi7bLrJMmw2z6AajewcodCEuwaFZOW4fBmTjIj+RpbyB
Fh6qHvj9fcpEYG963XJ3wDwvvdB7stJE65o+GY8dgPCJk1lPUVj7/TctGZfyjCc2bOFUoc1peg0G
Z6/iu4SKxwFtwpjaf8+0/LhoApJ+lklH2SExulcfA/kWFxiApZLQJ/KQc05tNVC7Fsye1tFJmseC
y+Fke3EOnEpaQrBD+jt7JetVVW3CULWWtzZIPakIeFGTcut7+02CIEpZG+vKGjlyW+UdZEevgcWy
e66s6usBFAIjnV1u+/vSJmhEVzZqZT7MkMH1VNhLWCiGsplLNeD2yeS3S4ju9Zj3kmR+MUd8rfXg
t0ssPCSEF2HFC6zSEvVKQEAqvWr341TF/idb1rCo5Eq2zq9SOHC612TA0GoQNP+hOyCDMQUKOW3m
dG4jnpEMUKRWOr906F1Vm4dF8eszPPljWM/Gp9CNFADMy4nznQd++JnYiVqviBJ/8thHX+5ka7jX
qE7H0mwIoIe7c2QWJjEcW0/94glYjNQ8G6Nvw6+U5VnsbmpR5cU5PG1FshE4wgd/+ThcKf5NHfTy
WBfvEVixww9AlrzdhnY8jCcblNpRCdJmpsZe5p6vwKF8fmqYkgvUaHM3jWoN9peFzKyYsK/zkYzY
Zrggo6h/IABwsinwAUPX5CMGVFPTrOh7EJPKFudWXY7hSgh85nPnOcxls3gTASGMKOo7kN8a6oQ0
i7VXBQExp9pSLljVA2IbwQRjTpIolGn9vkzpwSo7u6VzgF6pKLBcmBv1h/YTQA81jVEWur24vKlB
fFK5lij+Ns5DGfFbbcjDT7tgFUjdueNfH0M3EnZn5SFuRNxla23RliHRmXzWVqFjmy/Bu5A/4vXr
brEXS0IU0lpiYM5uXrZ+6lrsX5RE9Xa+a4nGzqQEXIRaIhQaWIqpZNaqritN04tB+BFcwjq9Urre
mQ881FWVQwd/Whhg07FUuWgpVizn91CzD/86pAItSK/DV86tEd8ZCUGko4dQC9/FFXDt74CXsILS
hSMJtJfxkzeC9U3Tsdo4hI+xBxdESHY8hnhlkxcgbU/qih+u2NTUwEfB0vRUD5kx6hTeDOI8gsNA
ZsurzwzAyiPL55vSkNLHCEB6FYXtaP+TU9+AYaEO3iIWRsjLMrLj8Cv/fOARtu5m4H3/bCtmGjpq
k+H7a/h51v7bhMjBgccOkQPm0gk2yWH0TAI7umSO86xQEOgLFDYx0HMdld5IEdvDOfK98ZzZXL9O
BYk19AU5oJwfFXHhlXfZKME9/t+eLxU/bgHIrl8/0eKxovyI8pn1tsyPSpZD+wMFnL6zd4VG/EFA
+IsnLJPaerbxQKpqywz0nespAlMsCMC7UsoMcjL1IMPXKwVKAC8y0j0xPaMGoNUgzGABHDb24Ik1
i2BtgJicy+bfYcnjDy/FWY5kXeih90wfys0ujJPhOjVnSkXqSRQdjdKC6AgKxHcNJJOCBzYPT9ST
xz6V9d5lW/dIbp/whQO8jRS+1KXd6k1mVr8Xu/M3ifSfmurO6uUNTaywUy46vf1cS0888ZXTfxaC
Yl4Jb1nDGFoH21cjPGeDv0fLbjp+itJ3u1v8tak/dfv8ujx+r8zfWle9Sn3BXSOEIKQz6C1Es3kS
c5wkIPt0GutHXejZgorQ7HZ484eBuMt/W/A6GWatE0xLgiVS3oOqkWQbX/FrzEvRcDQ1RhAY2QxL
E2MdAaIA8arf/dxfbb6r8TS36kMi1GccgncOGzOypBDBHCnuTAfkUQkG7fjaQRvj5vo0YorD8Yx9
Ysi5nE6OFDAt60e71m0r3+ruTsfk1hUf806gycbqx1wEjN5eMhIE7B+I/DHmeljYptHdYQNbYVWe
nPx1EsDQz3NVITG7LLAZgaJ9UZnsg8M/M7jv3a+T4eReFZ9gENqcUqlYCD9fGk8rV/SZHv2kTGwM
yYgUbYwJ8MzPkWy/lotYKLa5VacsHLaAlQQv7kqDEmiWS7JWN9Me5XQhAmsNFhLvI2J8gJILpmYw
DDccQphsDL2+He65trEzq50a0M0/Nm5Ho3ka6Im6gonU2vGx4l5+GKW44TBTVy0CE6GtkqnSpsAB
Rj0NAz5RCv//piwjPJzJrHPYPBLPXtTmgRJ8q85BvuFssJKM/lwjnYVGQRcztbWUfnQznWIeJ5/Z
TlV4NE2FUdCd0+hcc8orYuQGoPoSU+azq/2BJNQXxr/QZ043D6G1IqcCawOu9df+hsZbjjdhepL3
zr6S7mF7+/h6tKaO9/MgBGtN2hqT2sikVYKIcOMZAWEea3PGA3goOsYa/8TbT9luN54Nffi+BEa8
8T+D/BOoO86l+H9L3iBfES6KlhibtfUkAZwp7yeKKcCbwnwALYOUioTaYqbf61VHDnlTSz3K2+XR
wjk8T5IVBJNruM0xoKY8EcijYLRvpV5w+whAnprQBIzRmyOLQp2WpjrZP7higlhTpuh9oTcA8hy+
D1C95z5cSqT5tPl855HcJn9BkhXXQZ8QEY1CnK7bIIVPKPRHjHXaPfC3lbQx//uco+kcVjx9d2Br
CYQCypFE/oj7jYkpjfzw+VTwgfaZZx8dx+Bl8onO/Wl8rANWIvngXXT2jibptMjQVxp/HakggvWz
/JUdE0Mi7jPIDEgOKIiat5MArwooMlF30LgKkpXezyih+kNkCTMpSG5g1hrrL6XlKVuik03bWVni
8uiJ/DpLs+WYU9PkgtplizPoHzbZrTejfIwaJVBYs1hQ/vWP4qfYKztHLNHVSKYfvDOqlRboEv1q
rUhOxUxiXvl2MqObpimzwyEzqo6VEXqlAEprAL9jPpoRgn8ppAjbMCrdbyRhI2G8rRrqPt9Xep47
FMOwRXFM7obCo/3qH5nJ8S3JBvBlMOYQlsXb/k+cLeqjqqhpqExdGqriiI35E5GfhdBHkWjMVLy/
8/8RSBR72y/yyw9r/pe8kxNEHxHH3Gm458RCuTWU6dtVroDAipP2uJ/miT24lbaSXr3b4gjBxmlw
4Hn7oRseRjxH4zrNf9asF+rZhkqLngFM7GEcHK70rPDJp1CpSvsD1SUZjZw+hKhQWIKi7Low8Eku
//HWC7zvZd6uBpStschvLqHwFWg2lHQOA3Q9H9bhRuHVpvrSkEVauPEWAgvPfrt/ZE+1Lg1YzOd5
X/jUvYjJzQB5/dfUvUhLwdlUoLphbrrbECj0mb3DlYo/8G+HI1VekTIgqXR61z5sBYfb0TLlq7G4
xBkIIjAs8FaC4i4tibD+MjlpHrHfB3YY0f8FroJa4xtOgOHf32lDPUlR6Y+1pBpy/qYpblgbWUmS
3WmQHl2Y3TpBl+WsxPGttERRG24BkCxVf3fS6WpWSLXWOQnyEdFTxOMvZUkh742x/hPA+psoJdWT
RUklOCQI0oqR2c3DsP+udCWVqN3z+JoQCUanV3cXf0/tYOMLNs/914C7/kSTji//K0jk9phz8cBy
d5Vum9QC4UMxaMOx61Id80EZfaeTmB00AKa3GquuljCfm4tf1/gVnfhLcFvrzVKN6LB6A5zEc2vY
6VopvPvw3whFkRHwLYQny0g+A1vunMTIrwnZJAvoYo5QQu7SPl+A4t/7/nnzQMb/9cSP0rREGJm6
dog7Y5i+AyuLvPKMi3SxHW3aWzJ6qxksc/nm2jxowPNze+0pnWRoGtgSTe/BTMIMhhn9whlA+yje
bsXJ3yXEdgZ/PNb6YZkwu9ARXEjaZsqdu2q+5IJbfvlr5fFH8znon0jEeMHpNbhkhv6BHpj+uUMT
G7Ft+u8eGcT9OqJkeoBFFFCj63V1VsmlxxArHNKnclZbUsJOCQ7T+NG8+vlogoTxZwAcuA5Iv7nK
EURUARlQVXP12WsJbE5pnRou9L4JeXNzIuvyWxdAINlTbcMNMO0dlDrhx8P/9HaelPL3A7wIBzYL
2h3n3zcZR2Xx0bi9B1XG+1WgIJeovg9b05V5K10k2xE2WSCgS84VoUYclPFQjAufsqP7ykIYWuM9
J96LoAWmAJQ6/1p4xddwYLztww6UG6E2bICdyRz0hJJMS+P5w8ZsBIRGjfrGthZYtdl3nHYRxCIP
Hx8nTHKp0Gerw2mS+Hh7o5cM3kTzLGbBjIar9Ducwn7Ltf19+AlTACSArG0PcOpop0VpaiJDt5hs
5yUXaGIF7UV+F5WW5hsMtuPnPEuylibemWznDnb6PBovVsrKb4i3sdOJShG20hhtM/nx2qaGfCSQ
YzlxxwMOSVeNax1BBb6pMPxH0+0D19qWp5uCGzA9m8NHDPF7KQ1xKfOMWYqhbuVyl8CmqrMR01u2
JUUOVoUDOfEBtqbkpRj1z2hg8AQ6paD9dsuo1QtylsfR0x+uPbR5ub3wvzjR2hzYTGO0ruKF8x1K
i03k6YbGipPdqE+R7gU2Z03F42I25A3Mq8iJWmaZ/cyGn3XkmcLoGyQ6ucq4+Js+lPX7I5EimVlM
WA6/Iw8XJiLzlMZg0BlTYV6aLrMx5jaWD/sVLXrzEFSJyO574KxQCOmnLFCsG7KnM/NyGI2O+YLL
a0YpZzPnQpPFzDHU+IoBR8QwX9C24bsPftfMJ550q9scQU5hWOIBTcp/N8L4LdtStXLbYcsQPEHz
wNWxkUc9qdIxA8FGHHoLzrh9BvWIsnAWzDYG7xgwGA4vOuvAb3K9dZflAzAA85mzsDlCkWCRDkrG
SbqIbtrAC7wuCNEv2DI/Ym5koyJQh2kUhZCl80rYadK0scpyHQhevoEAUAbQaDzhjWXFW3ySHDCT
+HMBI4zxqNlHKM2DM1LJroOTGgBGlNM63SJDlDqHDqJqgujw68EfQARvKX4x6fmSyRFCrkpPb8/g
lFFu6HJnK1PY88aoa5txnuNZLtW/UO8dJpg0XflJPzxHly7RL36h0d6KGntoalkKdCzUUjvZhGzj
Mm4iDrhbflf3fe444hQnLDY3TL4E782mzH/TvhpflNSDaaADizq4yvVsaVKPBcwXhR7oJHcTMoqb
tq1doK676HLf5s1e10UvPlO5J/pE3vVEysS1vZd99IxioFtaXdQtZHpXE2nViGK8FUSFlrZk4T+P
4d7UGO38GLctJbQxRw6cBQx6v4rzQNc9JnFTgiRjLtgs7dA9ipe4OMwgI2/feJqOBYXeIgsBOJT1
yDUyZt9hI4GmB6ivyVbwTIskuXCadxz8AxCYQhv0XQnPqRG2/2Sd02A44X/RiOgPYGpzZv/3RGB+
AEzi1wb7xvqJ6U0rSwHthR/lndZ88HEgIRCa2jM4d2unEDLQVbE80qWJSnnGCrZsAFwpdFlxq1c5
feamy624VG8Ow+jmsAyNnOv9l53DftGNKDOo8zKRhwoV7ojlV+NiJlTObbh8Sp9vPfUvHoP9ZiEN
dPfaG+aHc2FrePvVBLlpL/7PpmLO7DXFg0xc8uIalGy6RfEJXCZofyFRklQ0u6UYNoQ7lEjmhJZb
MziI5PKHAgQ1ZpXh2WXk3NZhH7KDyGWMGOCfsIhy0qYEnM/oNrhmgJNi05nvoCCtO4pKhX3BwRYD
icSLIrYMHAn/e/6WkXitS0xTcz2MmHBJQeM/mKVvc+a1CM3Fl8t+9MM1liR2kPLizoa3LJD/YtzM
Pj1Pr/V/S2jFIbh8QYP1Tp0DXG5IHZSikEq5NYoX9ssHba5wDuzpk2jAvDMJ8wuYdtE6VijUDYc4
SsYaltzxkUlsFgbhAcvUMpArbZenRS4KQ43lsWggHXE/eSqMVh1mTb0doZw5IKUD8CIRdkYCpg8C
1HHltspZvtPKQhJUR8Ia+cK7RfUfMPtnUSlRTu2F1eKC8HHa4OGrV1t/WmvGS1GB5LtfORLyjKwB
eyH+qjO9nQidmYDRNB0s6dBk3JbBpdFQaaoS//GgdHjO4Kr7AZgFnpj4vjJec+J4SSNDs6Uu6k+E
13Y+21HZDIb2jNse32bIFj7o6nzqe+GV8S6K6gGRs1rJM0lsr9Nfl2jtk+A0kkGj4FSaQLI2rdj9
UQKnUpqXIF7lz9Ry5xyQgX8SA24zt8VI7rtsPqsWwWdFb8ANjzfEHDUfnYnMj5jS26KjtoKx/U85
wQ+KwCZV2R+kIpj16xYMjCG8SzbYK7IagFSyHp+WrPtCQt/6zYy1CW6eVAPUVOgcfN2DyX2e+WWF
M9R0SPISURnRAHRwArGkkqh4oFwxNMH0GtXr5tJ/qJUpJL8TFL7Eq7FSDBby8MPZUyiDa4EhEuou
7Y+lTLo2/MQjsPKiRY53qD9RPBKqbVd4Q7D4o4ZmvJuWZ0TCzytmPmpOsZG+si5BLrmw+APvb4lM
b/T/bbcCdbo5KGV2YJUQfaa3kWAXtmOIUfQo/XH6uNcn+7Pwz0LxpFBldRxM83YsVv8qO/4uftZD
oa6o0CskGmHTkOHsPETlS/zfGuhyxK5CoGzgyCYbepmNFv9yADTkvgHNQ15dMBkwQP+AuNMXCWaR
hsNZLPVCXWMIoTfqMnK/Ouy23gN/xaW8vn9FQzGp8HmyzSOlTeFImk261f2TzCo2GrLuu0Hnp3jS
xM+IXmlLbUTDEKRoHLOZMYYj2p2UZQkNywoshuOXZfLpF4p02Gvc+KYJEgPStxRyzFswfLhrzQHZ
aMagSbWTPGNiBQ4IkAT2hJtDfcKkfr+ibyFv+GEi4TTJYxIKxsb4VJbTJbXj9kObe7NPivBWQBwy
Js014nAmCfb4/79ehUrJZw776VxzvT+XkIAr5+bbhDwWqpwhKPw5V9+yclla1l9ynSzTTWZxvPsi
/RbRKPtdEMIJuHimmHP0mnyjHgshuUfOVvNTvDfCpj6UVeOJqCBs6K93rdvDLxLwqsSfDGK55Xqr
hnv7IDdE6mEpyxtZBTcExHoE90Gz9R+sDU/itwJhOXSQvB9xsIu7jFf8GcEd2Qa8A4u133c6Dhuo
6g325PHB8Z8PlYhGldgkOwBZ/0kceqCzFxDJSKwqYW8fMVjmseTTEWvR8M6ckgNrbMfC5hbrtp/t
LsOT1DlHG3eVj2XmWtQbXk1Z+ktDVxAAU+g8y/O24iFjF7po9L/yshc/TLZVQaksgoQDXuzBmIdP
K28o1BTUaxHr80ldBm1/RKh8kBp5zuWL42PD5h0/a1hPx4DE0+WOKsaH/SYoox5SxxV2lRHd8mpK
e8yxnZUxkLfU7QAKBtTVtXreWkC3xXDEieRcWjYPLAqOs9EzBOvp0Mo79gnV19hcumxDr3JXYk77
EiwFbf4vhIS5O+L8RHQPP6xIwOSFLwNzBZZCtxGh+6RCIx8JVrSunEhES1jUQ6yILRW3lsCAi8YJ
goauHpuiyrBckMRLrdmBOPoVD4UweiB1KYoCH16lfyNfSQCTi1FZP4fEThTR4CkfU6yS+Lec4yep
TUd7g5kTa9dNolhk1+VZXTzLVZyn0momUtGncT9BleUIqAh6aJ4rbQHQ/FvouxShgK5S2TB0z60z
qNMaNAGRwHbYcg1xzMVkJFUeRe6KI3F2vp9S/tDUA19W1wQY7KrQPw3YkP+PSdWn6Fhrqyitn/A1
jlT4gsRyzZW66pDAu2C8qasZrIzv6NtIWt69eqOxV5LDVs7VUJb0OKGvhFRJiJXRW4F7+8D1eG1i
Y9JUtiLB74j4/2kt8jPCXYK1boilgqeTHOg1FfEyxNXKRm9DIymTH4jNetsjBBvKEJlsFj2Y3cGY
mTBeMqObCZVqPCTVqzggQkUK9z92eqnPi/Ro443SHtMpsAgS4QSIBqIlipcfeCT71fBqat9h7La3
hZ3/+EbtwjhtGkMizrwEhRNbqAJdEfqNyHzHDslF8mRV9l8JFYcuFobR7KQ8OqjHzlQGXp0kS/mW
JJId07Ab3cKscZHA4Qb/VRDJ0hqbVy8bplrKZOh9vyhGmpkIEjkqipvivFxNJg4MSZLOt2GgpP2I
7OSJgTvXq6axJzy0xTk7/QjWCxGv5OuT5J/TQve3m4MTGBHd61JXpnG87zCGDpWN5PO9kL39oyvM
tGyd1ig2RJgfvCthnYZywBD76KwmFSwbjmfUioi6x4qlAXkP8/0uIGz3x0X8SLC1+9NBhP6rFw2h
VM1HgyZ9/jjSYNGKXUMOXAlMuKBlVArl+cys5GJin+3CDn9M5n83wq5dXbEceRuy7qgbil2Gf0De
4G7K2DB9gHX1kpSyB5MEMuf7gGZ1up3S5p/+o1/E8ogWqjOSd7GwxFNsX6FbuU8TzOiRni+8VLnf
t7tCOI3f6Bl8RPboC4oMV+13sLT1QmoLZxVR4gIAUlgbVTXW0GMjhpMMNmJtb1RZVBCfSUhFoYEa
9I7scUaJWfxa79I3eIK2ped/LDrIvi8nNQq9y14vnHNKIjGDZnJnRPU958SoV5b2AN5onTuiz9oF
cphipdKBCmgGTJqO3GNDWJcG1+vMxSH37kd+QlF8cn5baD7m/N6Kpcwyp2b+5C/3tARGRS+GwSmY
YpKE4CWEB+moQdVAHZ7qoaJr0exGlNLhKxGVHrC7WktSMvOj36QbYGNgFDxG3ySzhuFahTSojnBy
iyQBOQYYFFK+btuBcgKpDSxBppoWJOvGVBNYmtl4d2VdGzFGHNIwRC6o3OuWvVWnJX9RD1iD3MxC
SoBzycMBpfIQcSGXpKo2jJq849UY/kMu83SXzRg2prdJwZcQjBYfMX+38FTLtfeiXusIZCUVJSoa
V7kmAhAY2NhYgIjhTzjzwu71g4ybni9DqfrHPYlgBm0q5vwn5jEnbiAGBGrEkgRUQKuiIBLMG1oa
itF69R4roDK3xoyWaS7mlhYOPM61SyaSnPjEM7vlvaMS1eIFQ2cq1QXPBPZDgfzbti2rNCap6q0+
iF6URIeChY6nrEfE4xjwmgV4dQmPy6ofuuHJasSLP8pByZRp/pqNh44YzwZApsJMmYYf7//7JzWi
QKkCBd18faKtTQRU2niHj18pA8HIHzalIPsODwTcRNbdf1eAueD/nXaVIzOPYG+W95yDqvSZboTz
UHMCrkeP8aB2O9WmcQa96yh2fNKV1noXwqDyxR9geA4WDzEXnE8vXkVEVev48t0e34/G3MUstemY
nLvbdp7fsgtOoIvo+ZigzvKs1TGRk7UUxgTlCLal9MuQ6H5CRzcdTN20rP2MDZl56pRbxLmPWSBX
NBKUX1veWOQ3Dw9Ejrp7UNzSlJchWWDAJDkBMZ3yfyyHACadCK94Dglx82BYatjpmGwtB25MRYSx
Ug2MFiaXmwBPeBXM7/gSLQbe2HG540J1CgwDxoyaE7AbV4lac29jLy6Amu11MhffF9VjxN9WpOr/
wNsr4/jZJX2TUQBqsOaMX89RrF9VZHU/l/KF7moABcykMCDJoE8x47FKY0x0Ws7lDmQOq0xUz98A
EPmbFh9d6eHad1zLkHcGgj6gfAeqZx79/rtEaBR4bC/Cq1XebWC/+aEeaK0ulau2fi1+Jsm3bUBV
ZqAXjf+wWlPaSoEYD7RqtVOVG+v/Ln8qWBt7kJPSwTuyCJP2oA8dNKpbhQ09LqGfAazGbPBP2PFj
ptRHE5pXR2S78FKzxq89Y82ny1aTrspUlYCXMgLhwhv2BPeVxRig54RGG1OxvlA9P5/ugIm8grdO
3XV7DT9cOxoPMZ0AFliDy88vi9pGZK0YIyK3/ZOXp6ZbjUgIlBK6WaAtLUhsEShWWmDsSd9fXlot
/kRk+WYU7CbOzW2Mqq7FhXfslqSfs2Kc2/YrbxIX7ndTLUR5ODJ2K6sFi6daIIukPDPxA70HauPM
j1Q9ehdyr/fF+kE5hF0urmdGKNG8gasK+CTZzXU5azxDuyXH12ZmR7pgg4XiLM9aBMHMzkbEB/0P
fwsxEnMytEyAvOsk4H7jN2HG4XtbijcJnO1sUUcO6En/ku/r+UdZINPpdNGABf48xiJ6fyoLFa1a
Q7Wfp+4DNPXjl73czXlFCw1qSeA6wK6JDuMwAwN3kYfYifx8VXPNQMjLaT62TE409LLz9KAv0aCk
MjIISdplZaeMZwMWCgUIddU0sekg+qBcm/XnwG7trvzRDMUHhZy++BmC529gD2UeGbA1FHVubp9M
EVT01KToWUt72hFuOQ4eAZf3mv4nGrvv79PQB8KRPrxmSl4D36Pt6aPCjyWh2njyHMouZG3a7xIC
sSjemfH2uY3TPdjCKcS5Kw2gz65p6gtAaSwww6tyWQxdWxRAfBoJRSIQy2zdROmlwQeHxGGMYrg9
h3tFU99Dw18IdGWrl7IszRNHBWAaAdh4q+n1UWBncSYh5jEB9mU4eai9SFgkaB0mI7+R/n3wg4Jo
yaBxR//6tzIAcnhucZnZRFXPkPYE0l20ry8Q6eNJiXEjFyS6U6cCK6BtyM13Ns8QXuER2yDe9Sxx
DroEtdxUKNaY5UX31XHYFBcRftO9e0fQChf28BV3x0ofq8lDJ7hjfCvtj7UFUGsP9QIr8+VUYy4t
JMPvKNWQE8jpCZmltY2aJWVrrmQdoXtvxo9pqWXL+Lpr/73R0RuQLct0Z/dBz+BgeB7o5e/WlYnE
XV7GPIe+vlocwEF0JkThgGANcBuSzSE+zI7IINePs8fEM8iJsPDIw4P5x36wS0JtYHpbTv6aHqZT
KfNaa9Q5r33ObEyaQpvpziuiwZiJLjeNrcFhw6HtFLBKQkwDQFFJqogJsOcMMaYL0xDhuEJs0hpc
W5Xc18jZM0mMNxXis/OeaJDzHIu+5qim0EDB6zEMjFyAzxZoPbL2rUfQ5Ws0f1I2+wWDjtu4U7JN
NTvuQpXbARSyWgQUToNjve5oYydKZQlzxsW3aeslCXF+722y7BDH+UmXTCs4NuwDjUPKwIrQUdbS
uxc1JV1eTf2KlFaIngej7XGNRQoEcjPAEJZqPNvaLumVhaxILLniDdyRXIQ/iY5jOBu3W/R9+9j2
h3JZojI0aSC9LcZatNVQJuk5Jwj7xlpFg0JuHHNqgFCSZyZleA8nYfiluRmy95bWgCtFSMkCZCZI
F2sMMLxPjeAR0K1GFKGHICG/CkaNN1Yx+CNFlumRlgCx/k+XK3ZSh28xqSV8x0kRs1z8cGu4oMBb
QXeV+N4DluBbDR0382gmhvoaL1MKDSKDV4JBFLohUukgna8eQV4pMperSpIJ1D/b0XGYS69b+jmv
P5KiUqKLraTcTEkMMEg7rtG1jig/9UGBkQmHpW4pike6qQcdBhoNCbMJl7c7MGnQnyCP2iHT3Agz
h/n/s+091/Blsr6Mc3b/QL/sNDSHIHX1a21g4k8Oy9ToHj19uAGh1DOO3+YFwNgsE0eYlDl6vLW7
AUSaRjjFklUe7XA4Vs7auuWd2coD+zH+i5jOTgcVN8qIpK80dv5iJjeyc1jhZHE5VOKtXnmR/rAB
uKfEIG51S1XouX7Oy6+QclIJMVQZMh/8Vm6mE/I+okdQDqGll6vTZwYU+5q36v78aVgN6JywZ323
f6QG9yZi2Syy52n/72cgmTtJU6/Y5w1bhMcSnaEuSMn+IhvcTb+uX6Eim9UNhnjOMf7dTeeL4TE1
NITHokCUThZ4/ZnyDH/Kdqg/8j0x74AObaQ7cOR3fdGhQKwEY4IEesgiMp2UG6TARqQI0SJBad7z
+CZNBaZyswWsEA/mCStPxPsBPJPY/JzSHlLQMSjcm94bPooC2VPJmpxI32aU7HXRz96yd8FLiguO
dXJmXTXrP/BpXyOh+6BhwG+o+LYoTmYSS12OptAhlsQwcy3dwt2xai8GePMpt06HEiywk0DOi+Qq
6B6y7uVIjZ8jM+MRiPQqbb/g9igqMIYsBIhzmE8aZQN9uViNTzEG6p6qz+WZwbgKJu+n4hwylLvF
uDDmJYhtIKa6OM95P1Pcy7UJNTY6EvHAj87Bv39a2R9JfNtHGrzmfdHcV4vddvi4ACdQM32AeetB
iq+ipFP4U2PcVKlcm8keXSlvRGR1J+cO3cIAHhkVuzYuqEpFsjgxaDq4p6kZ601vZRNs/w5zP/Dt
nRcv6qHO9PxlsjpZqKu1JnMLEyq+uB3mB12MLtv03qzoFSBWHzUBC28MeyV/a+mXxXJb/gKwryII
N4CDfEQHVv4PC273UDjnaCVYJReHq0VGeozNqPTRDYjiq2cSmSUMzhC8boh4+IyqgzICejkUfIWp
2N2EuuLKgVcoaV2MqnaYX+z2t9JwECQgV0Sg6escWEGW5xS9KiK44SytxKM0vOpTMdb52VHHwaOI
A0fcsKOKy+Gr9lmCCTDJ9xbSnWDXHO1AoW8n8PICugQp1p1jsH9a5/CrFDAjvpmQ0nKV4sbEzKei
55wvlE4uV2144/5DZ/SOyZewjBxmyclVUUdfPL7KmO51tNwuJug7XfMuw3I7rwSqPUI+23ulL0ZS
RFIiyGCam/EGo2wfO7BSpyQzw6U+eXUWGsFa967p+R+HdiXT24vP0llwj9B19sOW3hphkM5rzYgH
l613r1kWKX0nCc6Ab+jMVEjiN30oe8/znf0XzJqNdKLCYksv8ENKsH/vCqsbJa1J97rbHzLKFPaY
xomHdD1jkHuPs0SjKpCN8RCsMpRKRdrQMf44Wg9xN1mx348AhEiKYJXDwVjkApZaE2pfN2zOvM4d
SG73QnGfMuzntnqlYxxPU79/iuMhzMAdYTuB0hc9vvuuos7AiRdg44Xaj+5Ursz3ps8MbO/T5ybB
ZFQ/V9H35F3V2iGS/fBlbjXBVh2xnQE0Wpxm8p93zP+S2Zr7kyNnK1XzD7M48po/BL9C1hI2Zb25
WMa32XyzVrv41Yltqs2VATU1cwK0hwyhtDXNgH2C4JmbKSbUo4GkO12bSCgzeOvRG9Zb0J9lYbQ4
ckQ41AyqQ9wkMmqgFQ13JOA5egZQMMxV0xa4NRgus+Kfu9zpy523K3+Y34aY06fBt9yaKjyFs1As
rTxhlE8mZ3v9nHCjko6XhRFPP6u4eycrXMTZXwPgOHq5kYEV4UKDg0AX4SfGRjZZ+7/qaNxEOtrR
WNF4eBJk8DH1Shx+q/Cr4+m8sRMSz8ThTn0w2bqr6FHfbrtFBkPK+n/W0k2S/LfDwE8Cm/vMxsD5
o0xppjzcRHllEXL4vKi1VE0FFqKgyXxRt5wLRaGaFQ+RNVU0WSHujvAv9hNovikgXsLDctz5qzos
FEZebsf0xYyRO+RYxa83aZGAlVLrErHe43c8t1IYyyo/soVM4MEG5cVkxGOZkds+Vxm9u+hwSS1p
8lZCFymoQ/rRy6nllB6qYz4yhHJzZPIiis1mI/k8OmBZOqbfP8BJ2TKMwDeiAmUX7X4jKt1Y+TW6
BxSWhouLGU2Rlmbt+u7HLeHUKB//ULEjRpZP9TAWqwQ0xFztgxHMPnexg/q3/83isMrtu7plPZ/2
eTkuDbCyHPuXpPWZy/9STx2PYQzXvahx2ohEkZZvDAUDf6+N1gqGBI5NWGZuQS3Yyl/RRChdgd62
c5SXFs1F87cKaqebKSxZMK+0vX3dnyb/AsrdUf8DshyYTDVEGgQXD3oMWpciKClfqSOB36k8EjeU
VfZBcuKc2FJd3FvPRc6TD+9Ha7I5Qfw/bbQi1v+VkHi9B3Rbpw5Q2wqUmBOGi5gia7R4JCl4B2gF
71ewvUm6M0MwefijbPhcDXmmR+/EGij3mL9x/NlehoVd6OGCpX5mXJNX1UR/tHo3qmwpcOwsmHwr
tsaq86T9fw5kS/vT8vgL0shxLNWQbhxm6T/SMA+qM7BEDydp1a/kdYfgUMlg79PSW5TCqdZKfFc/
RI02G1MUI94yzL00qkWEaf0odQeNaSOEQcyWrI3zv4gxrto1wcw/Hj7CqYDT9mzGXCXFmuXpVMJ9
q9aOMnxQ7ZIHqQB3Qx+Fs13C+gsdOztG5oRMT96465DV4sOU8xnTe4Xf+CMzkqOYhlO584zu01Oa
2J310V9BcBtqHQrXu2YMHgS6hy6eHw9PDPTvcciZbj6GkEbjebCwWa1ZviCf24dvt9aMRDqGZr9Z
NSsRYvsu1WZhIWXv/bcFx+jVy2E9UVJ13rk9s8WcDrdy00YeNuPUrj8KrpBtCUMCtuf9XV1ly/42
0f6e8bkkIpp0DmcFb2jvn3I37rUknuhhcMmNxV35d1lWntbZvqHvA/ADVyIXLimtkQ+s/3Wl55dE
E9D8UOsoxjNsK5pfdQeSalQa4yeZXr1ZoaW8m4atKJkRf4kp3LzSjYQzEIIep67oaAaB5riJ07LA
bvTZzwha56qYCOnOTRoRWeOYdUbojIH1z7dEU0R6R8hRGG5hvmaPX0WZxz7zaXyyjSzk4BWBd1xX
y65ZR50KCutJpq2rwV19EP8pqem+O/8qnrezCeIRUFCTCWhyPro4P2vMMggmSyyADqQTvQ086wUP
ljnTwXyHSfcajVm7+tQrJcnkZ3y0T6bc4hNuZ3BniCC3h1ldsgdECUpRYjXGxfljli7/MAzRM63C
O4h6vHHvZOo7K18Uag85Rz5QDZNqm5sH4fqS6aMn7kYAEcXOFD0pXEK51BHCF731nTPcQ1VMMC2G
nxVo4Hl7/jz/jNUDzV61sQdgkxJc9N8Oa6edjXJdy0/cx7JxQq3oTigQX1K1rVIW58iuR9gKI70C
+wpbj0vdII5SpL/7k79QgRfH/t2fcNNNHg+mne6O7ARElTyDqf+QI8IZERe3HCAOKJEkL8cBj1Bn
XJPfBInJkLW2Bwl2xFZIp+SjviKQ2QPhfzqoR/bGvOtmlIZujlbWVi3B6c0q7Ig6TyewhgYORsbC
i3a229fGHujqwdJdtdQv7v+mngyLUsY+d/A+/YnKsJBW6pz9OTVQC4tB7csf+T/jANGH4nvBEmSE
SD6hiupPQes3PkGnZpKUat6mhxMU7nDdWLvDndkcLIqPFPJOeu+lC0EJUCpxe3guuHkW6NVZs7rp
U/Wa+XCBChPGbmZTsaejtZMbTxZQcSqPLph/SnUtgpoKobsPaGj13B3Dca0V/kea9+eZKMSvdGO3
o3M9gMVpTR4i/wnakWwro8tJUNK4JZNpG7U56uDJURlwWpE/gjfJA6AUtoNEePooLHUerbTWntGK
4lzKo8d16719tGfAnEuM/19lwCwltpXfTSxa2uhTcXnBY9A+JcInKS2YUuDmSG5ktu/bKSWniib2
H5x9jmm9yd/Ic65wY2vXXgXgQv6NBnYPtWUG2L6kqjJ9MM3cak3VGul94YhU6mq8OIxYYPncALDr
LQMDirKFZhLHCyiYl6x4ciPgwpXW5Z69QCYgl9N38xdB5Mk+Z2vzIdSdaw3CiX3P/zl/pgrPv+9j
edFdBxxiLJMB3g3MA6cVc3/NWhNPt6ABsulVJ49d0MW3Tn6KYf3RK0O6bCm0O0+H/kU2Ljxo+7g6
8p+xHTzT1Xn8B5kJdBQ++vY5WIBrosH3MkC1wMGsZ/cMi+zBNnT5dViV4KqvGgwraq5JiAvwD5yM
Vqqt78R59zjlsHdVkuXArV7SzqT4nctLxDGWIzcvZhoHCY8shJ1c7iGoXqjokMFIpyAtg62NB4dt
XzjPorRX+uuPZpwkMyfJxhOFPT9ONoz0TkcJX88ysW3ISlvZ4HT4VXR9eOpFGpD8MGCRWiGF2rl1
TxsFWCFgEmJy+ha0WC20UgNWr3BplNOue7IAiMh0OUjtVgbLZO++ZZRAIjgIqSjL+Tu3O+GVm5St
joZWXQtJFkE4zbyg1ZzxESYk6C0MJ+QQeuBMIHbbk9lBo0j9vCPbwUvgaPaKu8iZaRJzai/gBT9h
jdrLNXDntk+26ms3iXaojDpq6XqQ6i0LYJtqstINZ9DhTVgdxWiWAuIiVIt8M7kMprCjcWukmNHC
DsCT8I+ZzR0swIFTeNv5dWCTJKf2QTdFRj/GByhzpbHSz8Vs8kVJRmRloG+j+PArjacrO7cYL7Xg
UG+czRL9WMCOa4BL9NuOsoGeH3CF2NvhvProH9QGJ9vEjDT3bIjL43pT99OUBylmTHdjvcx0MBj8
87sM0PXnvMkiDuGANJk1JqCDAXTkmUh2k6HIFbhWCRF4eqwXnC03cxhLzDfquslkRcKyQ7/4W8CX
QFb3rBCcAHifaqzWbI0dhs37hff50JhR3GaSOGcFA3Ccdi5Gq8xuwUhqd5iw5exeeUV9UJN+Yzkc
uFAsoAUhqYdmrky2AOEI1LP/Yzj5WgBUTicfGUrNFauU+6+K80YvD9zZhfqaLukNnLrvKfQ+4HrR
1wRuSB4lM9T9muzPZ3VuMlDnqIMFIk7NMG+3iw8xE+daJpQibsi3rB9T5Lu5Ue2HE/dI6sk/e4rm
IRAOEW6fuBvxYJUhIslDH914MwcnoSigh5jorHB96/uacqHGPWmnvzW8Ti2PgWfsSD62ASy5Cvey
ugi44IDC/mfwLUTBapaQhQSZarbehMKbWAaGxiKRfR6R0oxjBVHylZ/zFhTzGFglYvtBTReUq4J9
88TizzOzxPRU7nRb8dL5r292nxKvXzDDfI9OZPSH7+9IHC4GaJXsaU/wIAeSIAJM6bAN0Hps2rk4
K+yIlf5bSfX4yi3wxil1+bwrotfribif6VLg/N8jmWr0OFwRiayx8MDjfeT+SOpWXCIpLvV8EqFF
y0T2tQA7kcCr9LPnKnfM113U1uQ1MZLAKIv+Wk6DJaQ44rH+iyyiK2pLnufj+nvWncMD2XVOKXHC
ldhMfc6EFr5s8EMT8WcE/37cwtEltSj1fW+sR8WLX3zfM+Mur66nQ6qS9yeloVgf1xYfMEnUauJD
nW3C1aMMpv0DxxN+Kk17h/jkzMUpCzkhcAi0EE4mjLn3D7zao45tDUD2ixjxCz7JDRDeVtHXTDQI
EvsU4eeEcoAUlcLbR7k8cbr5RLEiZqr4LPmCABrsuWA1fVvMNw3mvpJwKHBWbS0gQfMPZQpSZH3G
3+w6ts8CaVoAKxrGvbpm646bjdyZLQIuZk8zJHrF8N3RQsfRhPfPHE9rFtOeu891yhfcigYxpN7V
lnPwRcfiRpb033WXu+rId/v5VLbAEyNqKK5u+OFvezAbxQUwF2dFqtJofIbwW95tEcRy3PbSq04i
Y+idkdnW25AUH9jkbrW1Qsnx6wf4gteGWsk8q/Aeve/WyaaIHIVzHf8dgSHBMWvwvFNI+tOmmNwZ
L4msMmgpn6DFf/of3m9ZSBhqPYeYwGpXe2XECbM+XgtlHarmPVmgcWKc10GF8LQFT+h8Jy1IRqtc
sB09KBFK/JyRLKvEMY/u/2n2qVQ03270aPBrwjTYdiWOcDUxKF2n3totRaMJCegQFtpf/RshrH6v
z3w4LeZ+eXrtTua+ku2hEiKut7iYSfbt5qQhyi31FcrwVfyoJ/fWtgKkd/lPYUPl1akQiXdKl9Ui
EhVx/r9md4ogF5j/CZbKpFpuB9QXv/kV4cf/cn6IGeHVdQjazBfPiz1kobEMT5vf+u2miI4kqTzT
VTr9OJRfoYp8F+lwpDH1MkTf59TxQHJzAVYS4j93+HdN1dL3LGjaRj7qgmZPXqAVkDdPUDka5hGI
GCJv/RpESWpgQWf2vIH9RRVLrpLjS/S1avYV/DVwZ5aDib2vmUQQUMzpy0vN/9CF3nSCaBsm257V
/KN4AvJB4EHdZXJM7bu6TjaJNFZfiRMKcqyl9GnJJ+oaGABhkipGhfPVSt4+iqV+jDJC76Yuj3rg
xPl1j8vI9eZ/38JJfGNhHzU8zzrkXT5ZiGXsUkRmU8uQSZoNjnArTbcfueEULUeBy4lQwTfNx2W9
slGCoOEzmAKV/6zqrZpstcXkNXctI/5E3OlHvJpq128SqZlfvjntBtuVXYyeir3f3oBF3Sb5vrRj
Olppp+DvwYLdlzx9zQLVoFcuaZJS/+VCx0jKW5b74sWe0I803PmmTY2k7kFaX4uLnJgcGdnK5Gdx
aJauaFcS+TVNWj4pe3IMoK50cvnYr05PlFACix+/dRzMadTYRmHatHgxagFIyh7vkZjG9qTbsHls
1COOgNsLjfhGHByMO9Vc9XJevSSgv0xsHPx06REuHbHa6OxdGrVOYag5391x+LG1UZzbe8O7mLtx
sukgwXdnwJuvWpr2JczZJQOHwIHdnWSuXZF6gB99Jyeb7a57CVvInMNBaVxwDJFRqWkZ1tEHBCYI
IpRl/cFAO0yovp36HI77FQ7Wu0rXClUWB60qyH94CEEZ+jZcdgEXVtQrdzfTBzfLJ6+0r49eQbBJ
8u5nSWF9xsBigMu7x+TuG0xb6dfBvzNyuRc5N4h4pa7jyaK3tD3L4wE25SeflSGpEgpOmPXNjPWA
AHokYg2iNnkUqpUnsPwwgvZu4ACSW2QEyVIAmbI4qy0gySEBGhnytsSjweii2wq/ovWOdxzoytvl
sc6zrFD+Ym/zU6I4aFePP+opFO2myMsJ7Lp+0nVco7jRS/H9CqYzZg45/9/dmjZ/UKN9ANujMio8
6CP//g2QUQ3lQdTHEkQjO27+DmSy0KoH/yMPHUErv4x4UKp0P4o1SsEVnJ6lHYyOEE2K2yLt7Wls
Le0cB3ISqdeu5FR/gYuwVnYjniXmZqQPojCu/XgjK/l3k/1g2kAQnVO54MstnHrKnX5GXBzMRHV+
mzp6Lyw2LlPKCot+JSobnhaFz1lPTsPkF6gX+RDQpGH0HduQy1x7pE2jU41d83K/xNW13MmnJj30
chE0QLIflk69+CJJzehm4LJ0VPykn2XlaotdMdiQTTQkbkEXqLAbydfBvLDPvdjo4zg/G42kiuSK
7IVoCgbxTJ02rehClmRyAb5J9J7KKjVJaPQPVzR7yf7/Pt6VM70ENAMrLWScIULzowV+C4/agjFh
Z9ahjo9TD21v7qOBQBLCVfFqEVEXPDQx5eDxOxPNgxb+2KN9Zp9glsPISred4N8Sbca1gnvrdIJ9
2xnVxiq2xncuZ103Aipk9+1Dvhw7cKFiM7y0zg49l2d2PsysvX8oD9VNAFpmSm/NaJqf+MdwYC9h
dVlXxTZU5RvD7F73a1u7oMI0VjSTEGNXpigD0NaqSDc1uQ43uS9ib89Cb4vSMUR8mthYjwaw49Ia
rgtvfQfmiTZkeVDxnAz9DNoutMxt5Z/4lXfsGlQHbNGwkUttZtKWPjlf374b7O6g9zTTMVK+nF4Y
iFswfbS/yFdA6Vqe1ss8jGfx8cUKZlIROLA1hF958ODd6Z04m0AYj+3fX2aGmrJgfjxdDNBy7VNt
dgKI+066n2utJyO8Us5SMeWDn/DM+nHMp3n41d9eTMFG0n1i+3/ee+CFqboNT5x0DmnX8GfxbR/I
ExJM43IBR1MK93Eyqb+fLRrcrH8v1sQoI5qKB7CQNINF5xtYxfOWpyzbuykCcAWDxFXTpXZY8b2h
9vwS/PKBgJR2sSSazyCr+en/gRurlxnHxLmhf8Raa9+ZGNxziU8c66H/wfHh/4hA61/UadHX95jn
z5Hwps6VahWsVg7KDcBjuK7yD0AkOZln10pnBeuiXdjEw5F6jxXjbVvX8BOfFfMsfhZzROI0fiDK
5elZmQ2aAQ9pGHhwaEldoO3FZnLFO0asbVMnbJVvww6yCoL68R32Ak0Y6InkJlCL90BP39ard75n
RfDUMXhJCB5OMBBNxA0/ITVr60sF6Mj7bUOH7xeuy3GEhmLEY3ey7sOVczXktR/cDRVu+J2zgByN
Zblu0R9zAZbb/gL5oTGPNn1Lo4mlbGr8sabKM+TdP2uZ4Cl+SGqgbNBvTS3woRbw/CbcV/EPzaUw
w5TUJnLcsVWEb1wQQI4IizSGKcawlTKcOPjsejd4egwTdyMTJGHs06dQY0AzPjpbUt4nRJV2g2dV
vpu2eQ7MPeeS3etnZ3ApRGPRKsFGgLGRAgMUe29Q6ZuLuh86ugHDDg5ljFXIRirLGGZyYRUtNwTt
oJdoeBzWnC2WlxzTkgo5LpcIuKoTX3URvxyIq59H+67rcuLTMXtiTE7x9oKFc1zGpgGy1FU1xLyH
OEJjCHDPBMgMhafFn8WEAeWK8tDViJ+TuuT8dc8FNYC+KaldAccuqR0sw/HTE5OwGRWG1GCZJbp+
onyUBddPZZhWHh90LFQyJYb0gm38U/HQwVOZ1bcOo8h3O3uSmGJ6C8fIwKUUqk+fK8x6EtTVMPtw
TnosWVrDsvPEUuS1C3Rqklnr3N68bm9xRkS5Rkir20gbvwNDO6qDyFPt3oM+z86nYmObpa+Otaw1
tEb2rIh9JYg8deeBmFviNrGe8srCzgWPdGqeeu1SYCS9/0tm5buy96nKMEbkH+FqsEeAfWuNhn11
sAQuBzQi52szNhBnFF0aaeED1t4oT4Y7FTjAMMyq8nc7hdCxy5CNEYR9eL1NNkajUAkBCeMQe9+s
VKi7EyWFD92biZ3mwEn9f0EexHDhb2Zj3EzXrXo53pDOUE7b95LUfmyubQOoeKsvZTKHBAeov2oT
FvrOeQLfDUVMmKQuWKxSiMmAiiEvCA+XsCeukJtb/BEv4pamYG5+rjbapEAnmF6laspgkxlIAIKo
Phsnm82HX8xaiyvwU1aK1CUr3TsM0bHQS7QsjAtaj1sanoDhNdrlG38cXRMTRqH3qM1rFh8XU5wa
CVF4W6Df4YpaChb4RCb5IdpXcXwPwzyNuI6kcofyzHlkjjSinSSFRDaLaYHPJxqe4gWGh9zVXcvb
sm+zqGERVpInFmgcSx8cZ3BUNNEg0k08CAw/CQ/eEmPIj0fADqfmtzJvSZzu3Zhy0JSQoWSxaMdV
a1Si7qhMd47hemfpTidboDiBiTW2pAJTPUwx3ciDkDZjNRpiDL4yKilP6Q1+wLMltFPfk63ZXZ0o
2rbTSgZ4Qaqzuglwf+Ue3N4nlLH+YSLX1p1yKVC4jw3NtVrcKqDID3ZGM3DDTtcsVhMh4Q64hqAF
+/nJiSqXCbquia8mPDJ+mfwU0QIk2+so7aDw6c2veqfWw/x5JIlqMSoTA0fkGXCfb8nRoGzU2XZg
9hHy7e3bq70RLzpLf1tZ3GenUMRJIiWnLZ7wIhOZVHtgcoM5a8smLOiA8/R63H4EdteqH/dVInhs
dylc0H3HfJA5Xf+6VuBcXMuJ/yqrchkCNFZNSo0Fy4c0iIlK1blFKhRn2rO7OEDaN+CEzg+Zi3aH
8GMjLBiVhNPmntmhn3K0kJ2HnoiB9ttnuB5FeKZa8+56KlW6/fj8vYH1JxOKQNLORvFgOGvcQcnc
cz3iE4JocBgMfhE9iKuARguh/FFA5XSiyzsx4nHkVL/jVcNWAEuekVijUyNInL0dGnemAriRYC6k
BFCPuCLUx9yrklPeFphHnTmnoPqgUOA7+whhKBzyqXPBfTAkExrAUzP2kmMKXQRAho3wftqIYLEd
gVRh2eHQlmt/Q7wV/dJccYUJ61MXLI6oY1Ea9Gs0oC6rbG6kpjr4BXq8yqewTyRaIWJwpgwswEEd
OrqKXflKfvdA3mZtq5dPJ9l3+w3uVOSLkl1IknmhkwWzI0/syDCveTMYbfs1ruMD7sTGKmCBQphh
vK5MqMq2zQZjWn3w85xf5WUzlZJ/4MyjHzuFrou6ZDGBLxxAQiQqRyl8Qygo7v52kdMVuTgsxu+E
fICNLj9e2kAfSJ6JKUX0Vkfl/1UlL5NTa7AuuQVekQ/2RAt3wR3DVmxrhUYwIB2oe1zqqbxbQltc
/j2zsH1V4j2LDsw58tPSW3jkW5BzZKOcKo6lYU7a1OqnVEF+BcZpjegqGQtvSbRgMbRxwaX4lM7e
csjVq/zWj04r0DKRFJi935MIHEXyXGz7UMQFJfBaGri3ugUlMnNl+lqsE3i0Pi1WiRw9QNdRd583
0OVTq7g8FAjqQwtZZMIlUPMZxW9cNdG9dQvbOvf1X6Ce3XzqNmNDoALnsWKIgh0QvifrnWDKdz94
MCqDPCo45xAAV1aSytl74KnIRVu6a4CD2T7DyE/SRubLCdWkZhTy5nOMtMzRmtNhy0ZXxkDXFngb
lVzxmi4SetD8oqss5UN/HFVVG3tggr/UORx9rjlAesBDIWcL0Fi+9c80RIBGxcT+cBLDc0aAiEmm
aJFnxKJF4Gf9a24qBfx/Hcncn4OamVy58w4d+8Fy+2QN1tZl2uIhrP7OOXkygXBD3IZVj8nSBjgr
I6d8X/oOEOnoZ/cWm6C5usSfiA8bKItPYL4x6JI1W6Nux6XGyVx/vBMAZOtYjdr73xLEXLvKkX2n
fzvHPQGUiA4WLJy0qPapzEcLZK+mvoRxsbgeacmHFvNQ2sCVXBTzQXkkUHj3OU1pfTUx1pVDRr9d
yY9zgcxYEIarD3YK43/sXGsG8qWOoTi6/qpBgH0QE3ATQH3Tt4d0vDRp8x/BNH6ibHjvFovx1/tc
bk+iDEzlvvL55i0Fwpu3kzoI40NNnmcDDL5LSMPRjWv87YQNE/yXkQNkal8iMw2mLQfouW6UOkgT
uT5ymBzgmYgjJqaxFt+/ETwpa0BSczygWspZd5OFwLBx39ElRDT0bmVe4/nV0dZjkVigrdTjL1fN
oEQgKQjzLUaHx7qJ5nF7Jm2UAUiVTk76NLwa3LfV7VkpxzmM7Vjtm8ngFPVDe94StOJEShEsYXOu
BkcY5yOrF6h7yDeodAQzBK9bCwvbrRKXbEeOuxu99pvo2HdVAYFFb5OhMogSWmhsdSBi5TQP6he2
g5//nirzfvDV+cx4GFo+0D1/GPseu6WLwapHzlmQXUQhK/eyYdatAyzatsU/2d3N3/5Ucr4X+EC4
qUcLn70iQcBw8WMtuqlIVM+hq+Eel2bYjZJ1nD/jGJ5n7eDwsZyjEaRh3BfRfkcnnwH6soUYkNjm
Z1UqDlaqRiEHHuQvYjStiXcWcnvF6CE8ynMX85GKXuClI3DYxzZvZM1SPifqBZUWdDeehQLJUrcN
yPEWuxb3AUgzHXQu7L0FN79Jy05LscF7h/lwj519BgU4Mgk508cGJK7bNd82x6iQ0iimM0ordomW
3OEqVl8InLFT81xJE8h7nFHOAYVTsXqmybv3pLxetxxoAwAK0hG2I5ll6NuUS7V884GkG278VleF
1yediFe7ULw067kvcFer304izlJa9kG3FGva7jPmvFRKSO0ToaRchKQoW+pN0VUmvkLLl8D26e9X
Z9IJRNe0pqBoV3bbxET1c4SYC3l7U0IJRQlkQQ3QzLkFuJkNp0ZLbHqWegc0ODMosga9C03H1FjY
Hd3ccY6yL81ZK43m4tWHimIxgwFH7tBH8aVfxhUDTRz2w6T6LYO2ZWR85pMuaKq+Ih9HR4FdsoFK
B6znJfvlfG3bG0Z9UV06aiA5Mk2+qztQ57U68d5Y0tOWq+6ZlajONOXfh9Y9jeHbYpSGU3GIVy7M
hlYYyNxoucIsPf+7LcaQR90DWJIaXU3DggmvdopHbmbkBRgeMgtLBJxUiLxg0cqO3gfgquFqFtSh
dgeAw4aH0ohYXa5gNAGdHLnxKvHgGA3TJRFM0oI7EFvRLqJmwXHq7+/EuvBInb3OtMoTgqDaexY+
xqr9H7ROBgDP5r+ermpb6L+hn/pYS8CF2QrtyAe17SWukIZTpTr+RjSazvrUTixfKPzNSwNNZrLC
Mfxkst+PmDTy/qHWjw8MuEChAmlrgpNzCak6/+ZL2lxyURtM3p1gvN0raTrbymvzeBnDvj0RDahp
w/7CNF11Mozyb+6EDzU7sdboGHPYJ9yIkKl1zZ9UooDx3rG3VQ692c6S8OOILyguPn4Uqt8r/wfX
b/ih95xJgVbDwrC2OUQjpjt1VJdkn77ONhrwNbyGKnW9gC3slh1WlLd+ws1KQZCiABLfcTq+iaAN
1k3Mv357ycreLsY0I2WBPYXwGhikNO9N/1RXsVTWINpyWhRpxs4sGcSuJ6HzoHqrQlcl81KaR+g1
afTVSfeBgsX9PMQ727qUGEPZw4MDnbt/gK8C3S8YuQvLA1M7rV/o8kYFi0xBQ5re/BFiGTUbt7mO
v/rChx+/6MSBivBVUPcBak7jMuIbXwdXnghNYJo+s5yBR2eDsjdnfO6ZmMhQ0Rxn3uNGO+dt7a+/
tGDeZf0sYQr4IoBGZUC3WkkaeDg9b+cZf5MYIsVldPfiJw1aP1gert6MiBeB9mw7sGedx4369pgn
/sha0iwL2NCk4frMlTfBsZXFj9efg1PZThkUoGknnKWxeCHUpB7mSErgxEz8auyxy74iZRX0SpUG
yA8zbMflmh2wdYgg/raWgrxbxmqB6ynUP8VBH41tgpnasKz2A2vfQ+ZUQhowY5j3zAjCBrr0NsWB
KGyPr0U0IJEgWIXU8ArW50O1M1EUfGGNAhuvuE8Rx4VcaKZJ4wVA641iDPypwKwcVWQzOIEIaD8b
x2ZJeQD/+nikk8oW3h17WJTU50FgRZMKx2jtf3MMV3RN1KuwEBVXEnXOvI7WGqY8kmrHkkq+DFvH
oNct/WFEiEtAcefisxN9AhVAch1kLU0sOOS0vNXoCD2FejqUSq/s4CoFmpKmaDtB2+PL97CMfoc0
LwUMofhPz0ilz2awUkblnyV4dD7pFVzSgO2wQ+0kYjdB6wv9wpY0aqxQCitVKdZrISxFWKR9Va4H
Ee+CpPYNidZHkoFQiuREjFpzJ8yz+Flx+xDvWGiLigNCgYAlxUxllhsL14lbRHtWofQ3B1KZQZo1
5/Gs7P4dHkpT+jZjlhXcqT53JMgkn+MdDn0XdEvaVwCXLDlo/PRo56GswBnK/2Ktl/wsg/89h/BS
UFgYNwgDZrYZzHVmJoQlxtziuEBWE+JQM+cenTUCQSJY08TWuScGdbvMQBRptP0b6hPi7QP72ox4
YG3AMczMmdnjiaisIVxf1l/q4Sgo5jI4Ge+tXU6T3chkD2DZAl3wiGnRrlhnDlT/8Qp1tOfRYvut
Ju7PUIhNSqTzrkUuEAn0ToDlw6eq9vsH7k6WxqNKX7v1Fi3imu64TlpwIsS+ARaadL+pUOQKorY5
EFB7LlXckz2T+1egQDdwsduOxfx+tQP+epogKIpi9Rg0MWcX3S2OYM/8qjndQRKHP5awMg6hO8c1
yL2i6UN1HoG5DO8Rycd0SHOmHVZyDunNzxFOUBb25g1qxiaQCgVpq5B64VGgniUaOCo2wD7Vbg1L
X8/v9V+pMGwCq01/t7Jn0LIi5JxGpwOuk8nUDj68YCRUTcsAiYhEY/Ldm9XkGGOgiUyi5uQIsJcs
rP248O2e2CGyU5whd31QlMu5OksastRl2cyXCubKsq7X7r0nrPv1KfSGeUy79dZl9yAio2Z7sTwQ
e8m94Tfobkv+QgkMWOqWAjCrIKPPVMJCXh0d4cEBBJoy4L9Nbktar9feKxSnqFVrbfr0Mnv68tWM
6miwHCj5FNgW6WDG+oRkLWQmgeKmE+Q4UM0DUJFYmP2VX0vFOD3CQkcZJ9TWS8bAg7AiMlp+us8C
gg1dB30q2l/+95MOvlaAU1vzyzPeqGhssdImKYKk4A7wgfMrFXpOBgvVRP1vPHaA32uD2LbuCxXx
CgydJKih5wDcPPAMmyV0KuXazNS+ouT6A3fHHjXULi5lZpKgz52tXSbhAANoMh54qO3PK7WfSOA1
ZPje8QMOPDsBCdwdoTHLP8qAS73tOp9QxEk2fSsFlTKhWKI3TiEcJfuyO/vqZLC9Mo+CCwxsNAfK
CbEmjQ30JqaMyEzSgxC73BG+JjZSELap/joe738tI4IxhCkxMRbdUo1nia7e38uUfYumSjoI53W4
vK4ksOALWBDk4VzE3dvBpdWW6Jd7aGVstQT+9wXaPA4Xo1+3lxEJHKMlj9Gn2ufw86NCofsL7Nir
7Ge36N8hsd95TDMAhZ4suP/bU/5v4SOwOpcypsifSAZ5/du2YPUSbPjynNvgUYRmtGJk3HJI1JwO
lXsuDo6oEJBbofRiUM5hkwydVItQHZDwCJ0FwG2UMAXdaMX9xUZjZG0DWG4x5y/yrbommxMHoZy2
7v6ev/tNBUuySSkFThPiXWD0I8Kjfw0lTwdpA/fmKK+VOptzNudiQeIv3Yv0+YUrJQg6Ww1HE4Vk
s1O9T8B2Ab9HU1NEACbrG389YCJqm5BqXmtabPSoReQF5stulaDEkxw79qFvvG7yd08E9ohbZ5ih
dvRoO5gu+19hPYhsw7jCi2qMRL5AaMDuMHqakPRSzy5Y0lnklZXC+l9huBDS+GBNd4s/Ea3wFmOx
j/lyO25O55qHSticxu9JtF+qVediq6WKb5Qm36MX/7BetqPv66LoKu+ScGYpw/uhsUP+QFIswxIx
7nc3tWDXzCNvhbNRXgBsbrhioMwufDjeTVHDK+Eym0hmdueNkiNw8GnLjntKLr3ZKAhiwzzXpiaq
ppileoUEXxMJTmJc1Yoz3lRXDrFQ5q7APtk5enVQ1YObl4Rz4Wr8ankvFuCK8lBduNDjalQF7kWw
5rmoD4UmUJ2+i/GJ9ZThb6jBtFOGAdDvrMtWFbwC6HsWy95uGe3iTOkWnfrleC+9KOCx/tYCu3B7
CSd2j6Rstf28F1evxxEvKnEmhbFYs/DVk7GwH0JPbxJf/GwNllrMUpOrfxME6GKN0WQgoaNRHgJc
1eT33GAC3SyeVNFumhtYpdtv9Jq+RoS7YUZTPWXRiwyjWyU5cExK+LR2EwA/9eEDOiu85aiUucOT
uGd+Rl9KGYIGhnnSfXRVY5r4fyz7d9ESKlHLj1H5yTqur3o0Cf7tAPvhoszCOIvCJWq5ynXkqhsj
3kTVtc04exLa8cGzEnaQ+iSAJZEWvhD3Zfb/THEhsAqaRu8z79DXrMJXFCgM4XznKaTVtcQeC4IK
Bu7DcoFfVPzbRnsF8DJWBrE5lDsU/ZkJGbbOcXVmBbfeHOwbPNjXlDx9ybzEflETCxS2lMowSHQs
/5AQqV+OQXltHDcxOegWuGkAPY+7Px96Zb6+i5eRvPQXWncZo5cQadZEAZ8fB2DxcJfDtCSx9x1P
L2h4azlNgJgxle9zbZxHbBJ6BjfbcxXINzmZ8+6Q7Km0a8/emEnyI4dQgomXXR6VHs56T6G63fja
M2xdcXx4oeKL1WViL/fyqpN6IjBvVKHqGNuSVbQmntq5gOZhMk5+22qxGEiP35F9UGFHKl8fYJEa
cmdGnFj8m8l6kvpzxvcoQGSqRZ9Ru/RJjSTvAEKSdUUm426Fia5CNHOS0KOqepgkR4P7Tqx7PTuM
hyMCq6AXkLVnXZ7spLybwJjnMqPbR20WLetATPo/YhZe89JHgW/LDosOR27Uv32/rsqPRIuShKMk
SQuao4+dZTxpJ3UoVh9sueziWfjrmRBX4pkwY+Mghf48U8YaCgmATsjqfzs/Qe2DgjKS2pUYRV+F
wMRlqLEkVNFMefqzyrzM+vV8Hav2lPlllwXgLrY9P9Ed5a4uokwFMVG2547MVU6/mDT5HVBl39Al
Yb8mUO1VBmr1CuEc13u9J8+XITk9yAdvZVvnKXk8rgk+uEZrbsg3TSuSfIii0osBivZ2sYcsSjSo
apjHyVs0iSGO7ajXbSbHo2fSfzHLteR4cPAriJUbfW4GmnNWRTDn12VxIAjxcEtCzspdxdpDFqJQ
L8ARS1Zq9UCKwUzZwjedShGE1uxgUaQ/w9e+TWXiywVNM0OKoDHIr/mnEetiWojto7beKGpqTAVv
yT/Dv4f3NhqYd0ZbQNa1hgdqD8k4QAZQNS8ufsi/jV7UOr3dG8BudWQ0Ij0L7zqn1qJgBQuqdl5H
n+pk2tR7AQ7CprcrAVJ0zoUwLFjhMGDmTZx3eEuMANof1AOOgTC2SNUsgVUI0fbk6EDB0xIF+DSv
faXcfzIca7/JMLbjh82lKS5jg55fGOiKpzrr/wSzLC1nlapf4phh4nmfcZNFZThdCWWxlYldXOxc
EgWJcTDcZVTYwfm2zE8qexDN7BedvgR7viS4KlX/qgf/O72SJec4XL+qTZCwhNKpeGlO111E/1Gw
Kz69ZO+6wqaBeIoYq5YpnaHSAsJ7D34ZzV7oxlm/i7m9EXeBAYL9+h3f/epbjZC4JWKYtmMtLuTL
/XX4oQxS2IAkK5Hn/GIZ8dRU2tafCKGe1NW/j11l8/UxCPlRoSwKqKJpPqEZLJIo0rEbtr24GNMd
jC8SY3nqY2o/2LI//YCbThOJIVmK/izTxCF9og9rB+f+nx2pAGCMIeLnZwUf0DVn/MS03OWyetEc
bjGlXwIrT9eX+Thtkb4qVU8mv7t9D/0AqqL4APMMoAxAHbfY5XAClDbOC+uj5nYIzAWIu7kIzHoE
6BIQVwFuYimYNVK0dKXa+wLY7y4RGNXIPv+2yxfP+NGFkB6UF1exuz/rKE5sK/VBnq3tmdqSKbzN
1tg2a/j4JATdZlJ8jaci1w3aweR/Sik4tC7MDce4Ms9sO0o0sx5+NRRsn9zy/5vszp+zfKD6lX/a
HYGnkcALghyVNi8bnNuxLDWcFoKToZ0935YEKKe2OUEd5AS+YuMvBk0TpUSjcwNqAaMT0GgQeJtV
bCDsimTE2sc4Af1EtTn0KP2Z3++vDhWpaPuVlJbdMW07dhfjISqb4pa6iF0kT3m1sBlIEAQvd0to
Vly/AJCSI1yDFeUsW3EvWjlEEValUYvlQlK1qUj0oZcCn49+h+KnG36SHPBoKzSxo0ntiguX6y5q
8jIF3Rv05vW7wMgARYbnvBQj6LNgn7Ue3IPWTcU5tKyIOfi1BB4b5uEM8eojIJffi2vxnkQd5G3A
XvzBAn1by4uECuMDQjVV8svTA2pz55KGwxJOfwdVKjrEZ4fuDnNt66rP0RgbOGNwOzHOynAR2Wga
kS9A0oeBt6i01+hYbK241WmZsFV3zYZ8UKKl6Q8ZBmKQYYyjCF0nfFWJa+42zvY51wuH/kR/nwHy
FKjyfF7pH+JVXu+1Nt3wDSxzAGWCnQm4FTAJ8HSUmucFDYQzQHQI7fnGRZw1IJpYWB/mn0qXAR4T
ENjPe4uOeCGkBw5WD6qYRnuukLfxEQQqzZARNYi8EBc+AG96gIdx0trOr5S20tglWIpzmKb47ILo
PHN+U86jy0+BD/gvF9KGTMRhQVR9eVGjP10zF5qy7inR2VkzzkmcT0WgWRizRET7MDWv0Xshvxy5
NW1zU3Q1bRP9ynE5pTOtbEjhWUfuGtosU7bAGNRF6qfBGMOhULyMvKjJMGUUYh7OMK6rEu4f4H8w
bFufNjuemleD4WmJHTlsVTeY4jhFCr4E0zeow9g3+zOROF8KBC/JLiCdsfIyuMNrMUMwqBgaNiJF
B7RkiBfx0QauL813XpvSMNBU6OCEMuQpkJZZ7DJcrmcvCGVfSCc7MwPU9z6fR0+ElXzFv9x/OLQl
IoESFRUHDZY8aGtAxUPscR9MOVPBNONEWuwyBrfgUJTub+o0+k2Weu/Oz6x/kbuQIsgpa0q9n8Gf
XQ02pOcVzbSbTQzum/0CjHJqTrhNBc5QYpNK+dXkol4epiFQTa1NYudXn9zQOxWNqAbi9xRVQtn/
Vq5W2l3Y5Z4IdXHUCGMWa3k5VXdGZO+/dFv7UDd0u2Zj1Iqhl2NENlWTGlYpD1AVwgFbK5A6h7+c
NpyRC3Wva8lQKGbE4tvj1xarP5H7aHT8PwoodWtXAk8GE4UFI8Gs4hgvjLaPVAkppaDdlHYgMxn2
kv57axfRqrVHKbBUmdIcgl+hjoAu50PHNYJn0qvMclFD7wy5jEqDVCGjkcIs/cUlb6VOghOx1hmS
4H75F0Uk5zN4S32rqqEfqzWiZF6cDJZ/o8YAPftuEcPOpWy8wSNZUtvD7Insw3Y3T0iVwmWd6bE9
G/jcMj0mIJ97elz/B7XCbAT7BjgbyWOiaQItJMg5SGzLsRTHhTE3cCZUj3u3R/d6ObpU98+j4EFD
XB2wIJ6+fGfVk9rqNLv4RPdPYBjDs4DgrxQKe1YuwHCMNpJOmheiynKO4vjSzgkPbUW/b+24I1k8
3ZBBzcgWUNvEaWpsvdQuegyp5yirEa+sve28kJ0jwjV2U08TgPX0Trsp8cdNrCwCN4E6tF+c4VpK
zBa7uBxkQhsD8UYSmv/efvBjjyJnn0+2JvV6zmB38Dh8yqZftfdEKCCgyNOrzVrWUgLPbQJ+9G70
veGbnWSPlPlSLy1vezJPfR0ihXliTC5dUB0vqmVdl2eOqrYBMnkE2beow+pr7XGmdZugScpXpDCp
vJCEiKQHNBVIo/mTOKyebHV+UGiQ6lQjmcj6coTLuvAAnI+LyxXstgt9XNtuElkqAY5ugsgzInmK
KsG2d8YdnSj1WaxbRMthLdgy3VCjM7Qfnn+EuDb1Ro2FomSoLxKPwbrokpEFZkqsbw1gf7Em3ocQ
hmTtL6u6N4hfJ9OkhGIfLtXdom2dIPjgGeCE6KmCEG/oZd7oI3HQ55AE+72iZdSkfxTxFxCElB+b
9BwYodEqPpdQ+1y9N7JWqcKeuBW9c+m38cxtD3sca9F8Uxp6tmqG1fZLl/zXdtG4nAUHC92ut7u1
v29YND9vNDaytHZA1UuZ++82W3K/G14cRungmhAgnR9Vui12qlkKNE35kTWsdjEU83F29O6zKYfl
fpg03DHf8NDh6Cdf2iyfvhN2zf+0U1wm1mxNpxapOgefIREGghR6hz8haRauwZ9IUbi1jN+tSMhh
zQ1CXzd2+tXm3WGQpujPKVeBWt0l5NVYG8gR4WaV/mbdPBchb6WmWxxxn5qTZpo4QiEO1oBbuq8R
PCpRuZcGo+UMrkOuGsb3wrFw56fOruFEF3/f6W6YbMHHJGmKj72mmGHb5bamSR6ePPEVDHSDaYBy
pGy2eaURS/dlrMRSaGV9C0ePsbyL9/i/LMU7WlAnSGjJ4uDczTOVvaHTCRybxcQvXW3MXxmU7LYd
YtL85AKGd4x8GLTLFP2D6McEtBM3jawRJ4ae3JuXIJ0ouO1yBC/GSbhc+8RmOu6OcEYy2MqBsha9
HOahFqeWXl6Si0BdNDJjWkpbVGhiP1eazdc6rzHXjSeLM+JKxz8S6PQ7kAXuhBXNnKGYBe0UTVMS
fAYUZbWrynZiQB04WT1l5taaWOiMCsQj7srF3X+Eb8Vn6IEPMEoGlFeHHTxGrQECSvWquWpTBhjN
Nb1JrcEbYZLsbEc/ehruO5azTJQDe6SwjD9+axaidsJOdRZFNtnfPngVtMppErKiq5NcnRRm2cZE
Qove2BWTIgDGOawQ46bjl+qSZStP7QLHaqdnyrk8W3H2PZuWvGvhprDtcVieJTtzlhiWNZhARgYm
BlQFYn4Inq37d9+cIs4rjYVI8GDdc0IscKvrf7G/fdPme4aQwIhCq0xHLElxWzD1iPG0hR2sIQKt
ugwajgNIdFn/JNodGfKMzqw3BhlzfNK56raHpfnjlqv97G6k9Q48bamTLbrjyKUM8gjwrLPY5Zu2
jLTEtQoUYwApCfTVyk80lk44eiJUM4eYMY96oEWB4gKzuszsRjRmtXUZryXYRt69Pu1ycAcUb4We
QSI+P+N4C7ySTS3cr/Dzlavt6HdLQfgQq7FVmVS/DbIBCjTayVW/Jn9h4b4JqkHdgt3Xpf/OS51S
RSGpxWhClYJY3E2adIzYZBSqJRGJMVtt5k4LQXb1QvstbeTwzXIJvhB3FbTcG3RPpaa9wTjQa3ag
8pXlpLC2t+bAC7L2EKVjUMjO5WYndlwqQ7YrV+LatZfsF6VrcyKl0XIPkWpw19GJsBbPLhyAsenw
OVH/O0kcHxEITNIsEVs+l51NBJKafJgNlCmY8NKwstsDoaPVvO9VrBnz6fkZ4BFI5Kbrz8Wp//Re
AQkRYN4X4lyNu33oYkfpxUUZWf2RYl1Dl5b3jlxEFcORx7FrxINBeGn5T67pL+zf1r7PxkvsOuVw
Rgl4VizNzyLP2r2j05Lb5JrDuey0an491P/2DH0mFHhrlnmY5wh/d+BAgNrs//sUUJRm6DzgTFZZ
J8vN2Xd1xgq3T89M2kbPuW6ai5KrivGaMdyEmxPie9hMskbIDf4zgZcZxZ4WDQ3V9uwEZaJuhWp+
o+fh0k4e+cPxHzjy838rEovwEIVwLJobZmdVaDAcDJEyK6rzM7LTmg98+gvUx4VQlRsqKRRgtEz9
jFQAQ/vlg/ijOay1F/O36L+fTCevBKVzVRp6or2zQSIfoW8a+08FtJx1+7s78bpxyUO7po0PxBRx
QElhpprJ8qM31B45nJNEwMju8jccH3kK+EFLDPSjeggBmCL4ICxw5KI6dbCeHDDk/1UHmG5URCEe
yineL7wfaNi5YQchWqKZDj4lKsR1GCdgfK0bLPi2sfqVvhiIOfpmLDXIqrdBUSoCHRSmWl50twSp
oU1WgSoG3NMOktcsMSqsPBzciS1dsa9r6K0F5/kWcYW/YNTi2v3FlQP8uDxpa+vsSujm+Sm240PK
yS8xGSPdwJ0nc2+UWb4W38lSxipaTaCMFxgowc4fhjbk6MupD/FWwcTEZUGx0MCDHSvMEvKqMmaS
4YanoZp1ZGGlVrskfM9fwkL5thPQbXTFYKBMuq1fpSebE6GBNKypReAJhJQf9CkTh7xiCpxScNBc
AfuiOXjasOB5mbpjLT5+DO20m75xizw+9jXRdPHl+dAeKHAULcgzVVfQr5PC2hxGYxaKB9FAtHOY
Xfiqoj/yn3BQjbDCkpjJXRY/1sFjdd0kQmhkM7neUE7g1syJ+qx1refItZAfBW+PJ86ZjeWgOQWu
jmPr5S0wZtYHf4BHklYLsB127foxDh/ARuRIrIJXYoIzMbubR2OGbBoBrfUh+DkaLYo5ht61G3D/
6UjqITZIkdURgu2WJoIDvUQFjlAnZR9o0bFaCRuw6SDD1i+7TFD44/hjiJTdMHgYj5v3gFH3fQjW
N9j4v1ZJOxgqQei2xSPdDhVvHcfKm6QkvPQxH+4yh4ocM8xT3BGb/W25dvg0nETmNpVFo8ij/Qmd
kK3ZlD41vTWG8f0Qv+zjuzR9d/PUtmJ0Oak0Lhmg0rGi7MI6byCfHScxdKFoKx+ryJIlL/hxSHfh
iFJEgCJlWr9LXLMA6ei3UMkLrrjmoT2433dzgA1rKB9/Ivra6XlQazXGKUa8B48apaOlhkE4SgId
ZxmgvsI9bq2kLXbtcd8rK8bM0B6H1kUa5aqrM4mQOgJeGw4fRV652zOXPimsu7yRBag+6VSVMDhb
TekCfx0qroI1d9kpRMjoBXsInYFJJvX3Zq/mVsV7bUp9L8plJKkLwuzraAFC+wT96z6Ub/+1fhT+
n1Q0vwRBNi0HhT07xQjJaNHt7TILVx1a3w4SjlUSNwNjwo4hcOBs7TOG9UeN2Sq5tTAA6dhbLmuW
K0C9MASw/yfrjxIbRilLsv3jYXXsz0bLoVoPdkX9SeB+qOXzKfik0kq/rIIgTMPCJ6nFD9jlyDfc
tyBgjRvLggP6mlZo33w/ScjgUnG5jZHNn4p0dnfMlD1WzOJBkehyLPOsK8/qj/ha5mULkTI8g3Sc
ezitUA5m4cM9134bWQRN1PaMKEnjyOJTO70IuEybt80f1kB8cxKzrqoOsID8ZuZP5lDws0LEI8Kp
1y/yFOQAwY+iywnKyWg/3HWZyVXWkDREqvE4q0337qbf259UsuMMd7NDcEkjgYYh0mfrwKha08LU
Yb6g9D56iRvcgfgA4mE0b/8/+35HAomWSy7rKPhW5851OWzY/f90+5qbntjozBLYqOmjMxXw2Qav
93JpF0m0jlZNebu8nnePIcHd74aomaMHzBu9/cetuBqPPp364S1r/fFlrTee+dXT8C+m5oG67CXm
rml8fx4Y75o4K65iRov4N8af1bF+b0wQV3wsI1iWaFalO9Bt7872Nat52bl3AcUHUV768oKwT2m/
FSn3qHQKfqpO7/T6AZaKrDj9cT8OO+qzb5owwJ+jKlxOAbtIPynB79lAESP7TgPPB/C1ZttK8ZX5
2Lp2eaBqyMFUJ0af/Tdz2YdqX/0lWouZOeReAj6PpFe2yDiSl7tbAm7vmYihDAcRt0NFCMZRlhRU
wjoxUnQfRQqKWn/P5TjUEkmw4YaFax0UQFvihiWosW5+9zVy6gVmZctErxA6Jke+CYRu0SfNvFia
kOXeMpe2wWWrZvWjFv3p88hjPgvK+1zeDnnB1vYlWr+PpOWiVevfokOfivYc5JRm3Tr4vlbFuKst
NrVYX9Zo+TkfzHRkhDdfxaEFR3RoHcxvl0ElzONW/gB1iE/eoCbHF82UTkpYWGNVqv7RO41Jivry
Dgj1JDC2+gKZIU3D9gz5e4jrzYwTIXsxl5FbToTDZeCvsd9FQKLX9KcswPIWOH+Hh08RAVK6P8cI
rfGZmShC2XOKclSSGJSzru/PeOyUneFcQFlQpWjBvqsdVChfvkQ8VXkuVjyZvK8cFuSX9ey1imRM
SZNOooviX9oPP+ZtYA/57Ctcj8/07fL9d2ag3zkiynrGoWlBnxPbM2I+A8hwX/IDstFSOBdI0N6s
NeoDd0JE897D6vNMoVms948EXol/wKCYYuamrFeX66yy6/7JWMxuiBy8Iy6nnjO26mou5r2L94WP
mUZxhBZdis2XGej71sV28OUKi2x2Pj6Fx7hsyZbOLOPiCLKcNZAkl/XGn5iieIS2N4iCD/Opo0uH
ePkiBpOUVwAvembMFbmSuhgiX8GInSsDVf97e8wJCa8DbtjOWzxwgByMb/nemkxMaG/Thix8dnmM
S7BgzGxfumwK2QKq1S5MTIjNoGjoTuaikzSD789A/N7iIeE2v/FQ0fX4Vahekc/vCkFhsJ7wnByf
IKZ2WL+nt8vMQ/Zxt5VoAxsB1zE2XTJL20KrzRkvXdUuEtdqlsv46BYuJioepgqF9DhGHcPIUloa
+CtGpUNATCeubrZdUAG0vbBvkyK3BNZTBl6PibfH5QWIfi3Jy33U857+DoqK6kpFh0snkQbdK2H+
zLmHEq6wmGXO0PFVwk9fNdx+JGX7W9Y6/6pHqV3aqcXsV57cHlKAOVfUIwJHMCBLSmS/xqRhj9Ev
2F053X2M7wE16nvn6g4/7y1h1GeLMasEyXRKjfE0kBtbJl4NIB1N6rDTUai3dYNYSkfIATGRa7xY
XI+0MqHCsdar/mLxQCFmEehSJ/atohr0iqscGftk+qAz0LaeJURlPWCGzrNnCEM1oE/JXWa8lTc+
knmhlaofNU2KdOgQdslql3dvm1AjGqtD8MEB8PHmvxVaG+BrX9d6Qm6CQU9IR3wZiCV44rLelHkJ
YAN5e+kPDS+PdsEWa8QVyI+Vdn3alwcge/wfgnN5tPweTzTHgb2XL6w3HX8oO/HsQ9okRAQqB+Vz
apNRaDAbSIIUunGg6sYtkdslRoiBH7xwWhCNwoPV9SEbhId0AMs8Y9HsLsGswpQBXBe0Rf/7J9J3
LxdoouaxkR3+fG+ruApGt4ORT2ge6P/JIZ6gkNWlGQrg4mNJkMFPZz9Pz83md3fY0Mgh/dkpZMg6
JxW9ghVTjvtMalxnCIuB9D/FgFk1YQzLA5I4uppKVS9pBXZDXBH0Yqgs7Kw39YzhvDo+AtKMb2hX
3ZU6eFuzRs0zyPBqgbiWOA/ni0d/ZX4Bu/8qh2edkZgqona2NASmN5nhwIC+V4VBQ0PExcYWTssL
3uUikULcfvRHhD+Fdvf3tA6LukBDG4BIgaQnJteeyeySpGKQlgXC4FGMHll3xy4OBIOqRRtZDND4
q7vbLpxH0NKuTpErqFzjJdVZMoWwrYrwNO0RPvxAZW1oQggN+Gw47WKl5FmTvGjyjQ7P0cd5egHf
Xj2+AFNWZw1B6y6e8Jel+QSUe6ACissv5CW5fq/UjTIz5uTwIjJYht9RIbOKCRH3xYk9FnvKoDeX
HBlTdvaOh4pWnMr7KGLg0wINO6mfnlpSIYpK7gMw1B1pniqDgUT/VWLxKnTFj7kOb7nEwtKruchQ
qdS/PAIZoR/0MNxrxYGR2KOjDkr52TAQtxlYYRUfKCj6SxIRKevd0HiolZOTtFzh7DbVVSlyHa4Y
QrhVPhv0/UyCxIu8ik0Xe374RIYY7i4YIA5bwFmWWh2M7P7krt6m7UmRx5YLUz4RDXglM1vvseNY
z+T+p+i761ccSKHH4vga5plvFUKGa5Tl9qf6hJLUxHEEvvPgIB6P1ndiy1iaF6pNphCtTSv+Kfgs
eO1TyC1Hb5dduiUkWOpDIYT1FCeoCmTQEKrubiQo6fRQdarKl/Xpq3pQaGSmKW7kyKDUAnUd5mR4
k4MsJWANaCal9ABaavxZbN1juIZ/+nXGsgGLn1I2G2SPe9fVCkvA91XnGnLK2YwmPfF8CN5laA/K
mclDuu6Hzy8gtRrWZ87vZevuEBiTPUh+MQ8dG3lBwW3PURA0636X6tMcibWtU+hHelAmRqjABtzw
/1j4C5HmDSaw2CB1zxFfI/HLkPSNby/sHrFjeLC+cmtYNYg2sV5k9rwEf6YB94HMDYznD3Loea4c
VlYiv4gxGecQTbQLa8kNxoL/ooxmvxDuqDQ+hioG+4MBE5j4RO/taWIFvvxDJm+U+/rfs6yHuIQb
qEo2IdJNraePEedQuC22kq4/TKFupuVBK/8Z0fBPFZyezd13dEYAtIvjqnY10jY2PRd5dJATUvUy
Or6d5yfD903auNXRLCGGs9p8hfnh1ijX50DEjdReWf7Q6tBOiovFmVJNO5mab2TkueRuCw2XUle/
4dWS0xSAzB2J3YQ0I1vrmSpp8xZUVvhsLLUlM6khYoKehP5e2u3cM4VJa2Osl5VS085dHI5qp8m4
iPvF9B+zQzoJN1yqSw6vwtt2YMpcxXauM32ybtLonUE+i9iep4vYdGubbEH/J39oYqcJOoyHI7Vh
sZqh0qGMmiR/Njs9jBU6dNGOC7N6wjQTNdRW4fUVIDY5rueZWb5WVxJMKSW0cWAdtk4JRce8YoNi
I5RBAkGJJWqTsERhgWjzTzxkofVejJWsFaAObWr2hdVgOHE4JdMxq6iZ9uTXsbt/BsRWh1Lu9fX1
EFEOHTIWIVpirZWyDgTMeJSLRyV375EJ35rJBpUF2EZpscLcfvj5Or9bHd8O1KMO+diqU9m2LY+U
7CNygm+fpVtxzr8ebhX5s+oXDcmT1S2q4oycMrmeEa3c0YlM09rXuc4DVtfGIQHytgnwmmcf1nmj
HDVPC90qL2EBp02yXcNkvOJTuXUm1VtkV6huuTqAPByu8ANvyPAsxpkqrpi0HGoZkg+DZsufrqSY
31MDwEuexlcTP1g88eEk9RJGZhFkOD6ms7FHfK3OOhya32Ah9oy/HaQyEbzJPVevLPaiUlXMo9wc
giWGpK7Ukglu+wwh18PnJtMkGgwNWx2X9Q6Eoi+QBqlvLdidprPWxQDyPg2qxPVF9Px39tK3/tr4
WyWb2Uqduph5Ypjdt34U0Vlj4lNNEnhq76DgqqoWipPzBaTtFh6cy+FqQbtaU3pC6RtOiOLiYp/S
pB+Y4yWBdd7TThIBV2YEZRJsfGknViLOoD2xCh/G7Qb9GHZ4VPaERVhHd8omCa5nmRTRETsYmoej
sxKo5B2vLvWTfFm/VqvckFqKiwdSI69UUA3n2Df25cYS7Y9zrG80yLG89l/pgk2nLhslkp8ztf80
YS5xpTo8UuBvjkFuoNK5GL1lGBiIdMoMMRTJd77YCOLi9CF0RH0SAQ22MRhyJKBZ4VDsq/ra9+nL
A+lIrFwcI2sDO/KYDXRJhz3kMZTZdnjZvmq5ub80MeWVaVbdBP/Ng4t9tGlcQUKJ5wZqgmygolHI
IITWUF0biB8cHEL3lEyY5xE+S1mKK3God2cHfRpydlbqqusV0AZRjKs8lPO3JNhg3rDPey7s/uCU
DF/MIqhitWROZoKAeD/dXRdFlV2In/rsWa6cs8rM/FJpWGxxW8XiffZaWqjWx294lEIpLhKmSoG9
a033s5WdzlcgbUvVerZFvWk5nTUIztRZMjB57ar9MUiUM/bp9PKuZ66EV9mjAVs57/ZDBy5vSeiZ
sznh4xDmL/88zajlHIykRGMVfA+Szjh6V3NKLs9GGCgOz2BFvTWztivXD9pOlScdKRdmJSXWnzce
mQhnNky4uS7a0S4znwJ9tOr5UbKewW2Z0DeGwn87iT3rhinl1eYayQjZpTkhZIsNVQc7ZpmUmRdS
kc+BhL/aUgdcufnEk94e8/JwiJri22+KoTix4TacGna1ukXcPGjk69i8+Oy2OH+PDJgtCSuXTnIC
Vsn0dEf1pM5KcJcYFiTTZyja0v/DQACF14X6kXdLHXismUJgKLaSkGwG4JcdFgrZX/LSeilcvx0l
ogWi8lVFQ5ZaIXzu1e2Yzl5EsF+1zbRF+oGGoK21dX8IgRgivFFR2KxlYRKKOwAvteXnFDlcMQKj
b2hTk0JoE3QtyB0/RDcn3CquZ9MqG0FPwrXF4A58dSwaj1S03XL4uKh97zvtJVqgQFnsF9ktJZzS
xDIDU47n89bfFz9Zdqo2qffO4/PxK+Dhfn2f55tgi6kj/U9n+VKfTXjaWe2nstrOnlZ3/ceEoCDY
iGapfYtzBoHu+LXbx7rScsVicxYUgeR9cgb2JQzP64o8UC0MtzHhyDc5oDPltmbPxWfVHj7YJUyW
eJkk4NV+3/kZ0Euxlc+xqkt+JFVgzThW+5kkoSaoRqyR/GDLYmnpXdH4zCQ49kGpjxippc1JSeEM
Pr6TzQzmzBjRiN6iykojhNyCNsV27AVg2F8gwsrCmAAvETFjRFGhv5reYbVC1+DqLpJZOxP9gSPc
PObsPONzGLMMvRqiu+NCnP11eaAYabvcQ6bKcsnLOxW/Z3C/RKCx3Xp5RzKGvCrxhSeX3SgERtTT
4HEyeSnnXnhfZzXjg7gDJ+gtoMulyCJcOuETT4C+kaB0eIBBYe8QTBKME/jEskMnZ7+eoGvPkMkt
fixlzTyS391Nj00njHFmsFEXj/SE2UjlJQ/ctLRWtTcXR2bLEkwTb5R/P+0CziF5Kxd9QNhAYYsw
kqMRCtqmWk9QdXGNwRWlYW2S1/YAsL2v7sI3Ug7K4Fb5C0m961REnQzgryUNXMS0Fmp+qaoiJ7X3
7FBmeh4A9Lk9B2+0ORcfQmRRRNxLpEdl4gIT1QJcQi/oXoaKX1NS3VCNlG54f6qJ3UdQleycwejs
7A+V4/vBb2DD7RmMwumKj9o2wQgLos7eUvN5JU7B/XIeSVPMVahZiULw8BG2ILvLOa0Sv2p5bTLj
hauSBsQ+hK2atT2WvfiIQQpbSTRTjnMt9f4zZLTjjFZuwzNF9L2dpLAN2DKFFTPZy/dTAVUKa1iR
GAEyYitclCPyD4Qb731xoKzbibUlFgP/9tWSugWKfbIWyq3cPCUQ/s0hpRVBQM9WZtGYPFwsDbo5
nvgNHyycZoDaBuKweNV65JAtdpJMP0S20+MkYX/EWvT/eiQclQpv0kLnM+tDBgC5I1uUNJs12/KI
YuGx75C724yfCS0Q36zwcATQnM8kjzRHA5C8FLUGn4Q4kY00unKOp1FPpjNnkUC/P68I6Bmm4tQn
JTOLI16WJsm044F0+3t8mxreXXB2/cUm9Z9rOy/CVJ+2JPXu8V0rzVtClVu2n1wO6Q+3AKoZ9SmX
kPHDAmbLsuMPPTC10Yjq3E3xaBsNVU6nFIJTp0PRvrScTiKUYCR3nClS8S5OMxi3gHu/lC/1JL2P
42RopAGErUcZ6Ev5ZTODE5s9fuwie/79gGfZojNnZRkFmvzk6kYTEP5rxrudR0auRGmTep2ejA2W
1MJyZQWPvialykkSSAr6C3K9tllVTdnhzZ6q/N1dkedw5eJD18Doc/IF+ZLHsVc2tcTFHfOddD3Z
q4g2Qkb1iNerZ5NxEd+KFVN4iQeOZfdDq+fGsTHSOxu1celejUKcUV79HE47lfT3E7TJ/yQqVrw/
W5Xd4J7xuLSLyW44fjgAPToWYF2PGdmkE2bnb14uEitmWpDoEnaPXLbZPlmL5z8IAEtw44lMVI7S
8ymyBMgB4ymaejZo4e5NEPA+nAie4N8ignNY6VrhvVABvAALMpy52/NFMyKE9t9W04Kkwd+/ZpIU
5okAz7rqE2KrhNuJn3V93uyZAxdu+ZKX2zb+VAn0JHsbf8S2kOyIHTUIgcfsYHent6hpB7lt+Uh0
PjZDSSqa/rvvhzJvDeczF8EYdbY4eBR2CdoP+eIEjGbEqbUJ4+eNKAyKaegm0Q9rOukQOpX5yrxj
weuyc7hYueLSYG67t90ucW5vFErH9WAmS5T4eEExqxxzRBspuqcl41Oop9FFJFxKFb7v3u9BbsJI
AJILdWf7YkS4ET58b5uKikk3tHQU4Rb/qSotNE7NCqhemM0j0DItWVntcaD4F4sXZ00nUV4V7LZG
NVyFTLGOGM6EVQNEn4PO2SJWFIaaZohz+QxMe+YIrlNSGNrAbXn3E0YUv0eaHZ0buh+ppu92isPQ
nM1CGYuDLjPHcWQNda5eZyKfsjuRAaaJWhmh1zbLBBRIqbBIEGGHCO2e2mIN12TwlnvGbOBJFtZB
WQcth5Pir3vu2y8ihQYtoYEBrQdnDmMvO0dNI+Z7cewYfpizy6RBJC+Ju8avg0modbj+eBNL3leJ
pFKIV8GhNfNNBPJ6iZwXaOUOHL4UfgCQdSa4vK00/7Xb38llUvJ83W2bQwWLNG6Ri4IPbNT3Cn1A
+5wCEYDVeKmPkYyR5yJSq79IvXndAK3BKrc8unMQy8Kj4hH/WNKbVAxYCj+5eEHUFbpPmC6HBvYy
fFnD9JMr6S5BTuaR/qZ7Rfjnd1GaE+Llemz1RAG7GWPeN6b5Ns0mAQxK5KQ6YKoyoGvHTMDiK1KC
u/xvM3BgwLgn8Srx0T485hhfcDAXQfeoFChuGK/PzaRTQknoJwoyFZmPrexCk5oZ9eoGTyLgJcxg
J/vtlNvsxuK/WwvwK00JsGPWBbCIJm3s+WRH5ivHnK57i3/XR0D5VaeYzfevMc2c5OsVjkzURQwh
Fi3St6ugMKXtykLxUUqs061y/qdPlk3uZB7ZZ5gHhouyyckU9XmQiddj3Y+orPnOFFYmTYYiGL+F
A5pDt1DEOr99LGCi+ON9r9WjE2Rx+C1jNk3oTXsH+DBQ0a5UDJOaUeEDWOjrEFOOUWn9HtcOoPWv
KT1snyR2E+7e8aM9gts8+CcxHcLGtrvOCyCZbgkwwTBdZo88Co1MtD4ZEmHSCdTTN4n5m6ot7kCG
vA8+IYO6emPZyFeIced51YeC5zgSqbVGXEdA1lIuKuou6SVJt4bxUqPgANWQA+AQTSamKuc7IUzn
0UwkH/KoEk0bkFEYHSYcP3/Oj+7Ct+/wSUU4qj4mgThaR0qwQjN1t3lo3UnlxYQJKlN/KeoWKLVB
+BRJ7aEQN7Qu1H0RmEvIiHwKHZvemIkFTDn3Vl3gP3OzfpPKOZbieJX+TNHUo56h/YpPUxFAs5Se
XUsqfFuCGwcjB4OWWE9yYK8yIBZFMmWS9zg9zt4PdTGwqzXUA7Rc7fdnAYaIgBdW1hCUpyC0vmrf
qj4V2KH59OOMe9BTYE0oHi+vvbMe70OI/flc71z1C9t0QNcWcIUXJcIo72YLJePr9+qlfme6PuDv
2onFMYbmjb9ju/skjJ7HhjztuzAxsHfwJktk/doixGIi4s9fal0X59mnusGPVYQl7XF97rlzUWng
dsxc48JOtQ1mdL4ze3dnP4j2vOPggSIeb8OH5iBPF7gZQbPReHF3o13Owkud+u2EYYsAgACLFr4U
/j/WR55fmaTSyihATUZVx9+N7c5O7L9mmZEniQP24SGquWjE21dDcVfz2JZLL8I3qig5xu8u2A22
WPpwyNC1pDLAs5KtaQT5NxoWTyPHz7ouZmq6j3Qbb7b+z2fyo1qF8HzAi2ABbo8VddzBpV097Hco
u5J9jUzxIZ43x6ediqJzR9tubwNPw49Re9R8erT/VuWTZ/8cXKr39cfpdEDu09v9j0H6sCc2lEDI
JS4fhOEuiS2nrKPGZBLE/OFi2mYN1UN78Va6aE0wkZdybmbZnlUqk9df6kA9fzo43Z+BZE2y0/CX
wFVjcQHO0gbal/PH1lQQ05CDpO+psyyIbMyjAv+Uq85k3j4YSsM3/oPFWewHX7epbdzjoCU994Nm
AoaWKasc4a+fsCjDxCPdJLJOHLkuSLySjFgmR/IFwTYCVa0bJzXebDLbmRd594UcYJOFweG5LU1D
3u43R7t0jun0VxBBu6FcEKnKjQMeA8s3Xb6TJdUFjrFVw6B8053+ksohUEh+gbDiE4PlU0tut+FP
0L3h1sir0LkDClUyrGXvy3At0BZtxlfbXYhMJQQX6VxNrZs2MaudUeonm0j4qNkWbTy3Dw98d1sV
iEIbTwxrJWfHp7QiU6P+j3DA19jT7WmRHULvD71kxWWTvGp5eumScx3EPp/DPhjFbKvPbxmsQwKX
vjPWPq3zST4yEwSRvLjrwmXi9aql4ine6r85uVeGSKIAWN9xfgzgPWARjz7ifG2vCuKRNI0RC+Vd
gGzZoQUiIcglS/ZzXJUksZWA3QnM97dH3YXna2vLd075q0U0jWI/F08WHOMiaOvk2XQ31LkvyxHC
T9v5iSRD/GksNdoS5Yje9ybq8WWnvU9CTDAp3yZI45tfC4z7lPOhy/ZFDIcsLcKip0cxOi5P5VA5
M+CX9sKi+71HiEGF9puRNcvF2v8StUCy7jsahKiDzZmh8Ob+kKQ9d2r1wKjP7guxR8E9qPrxPC91
EhqObm4B5nx0weiOiwL7dT0bW9q9pM/s73dE6m/rBNquEO4xcHc6FLW+sojNzHKdNVP31vCq3VKT
ksE7wIpYujo+VWeGYtydPeUCpxaHiRa14VyHC1G06A9b4uD98ssiCheEwUBn3iVjbgwuRM8X96vC
8qAATkeYLreFe+rDoS19vRRcjmNawvjCt7jpZ8Ird1EaA62elKzzxWPryAN7CkwBbvUNHMFYxztw
lhyHNxGuLVcRBNHnlWfPVdsQST214oFGhgJajVNWLcGf/AWPythA8gHkRw7V9o6QTfKrIQ1vcGXw
ZX1olyN8LQgTlcyYp8785NN8qGp0H6BEKGMhrOwZ49a6GJrM3xdtqErL52JK4z2vA9AZ/BhRYbHr
n/3ey4zit/3t5zZypUYtGRTbH6JaOQ9KSkxz8+/MugblECpoAPeUxX1M9k3OzHLi7HUNvmvmFk/c
`protect end_protected

