

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XpL1TFj1Z4ZooJGB3dSP6Pc8XBohs9jsfkhCnRPv/E0eBWI+lHNIXEa4u+PJkwlVZvWcONLhadzL
udIJCZSJZw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YotU/iVRJw4SZslAhIDvcJ/D97KMnOVr3qgyDEyjv8wq6q2fLHhj3+4ICqb6ugcylGrOPKTM6GCu
GySdwK4bI3nrS9w0oaYDzVELEOvqIm4XJLCRGucgroBYyoA8PVkBaBN/hy1UZ2eFbtpqDZTDDmUW
gnhHXGIQXAKgWs/2+Vs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FTBaXnVGlPEYCL5pjYNf/Hfv9XxLlTrcGa+WNNYupZxR3vhtfNpZc42MK/1NS/s40uJdFgxDtyJC
45US5Se8hJI4b4aDwCX364idcRnwiaGry68POf9K8M/hGFpyZ9lO5vMRxcwi4PxsPQ8qmw8HByT4
OYHJzj5VZVht/NK8xDiyoIlP036O3ULaNwMwFHKTcQi5PfIjaD1Kf2hlmMtRmABdZgxWPM2aDyjd
/VJT/RN4hCqzU/34S/Xah5tV1LyNxh8bcoQcleD/8qoNOksi1KJWJ4VINA38up8YMtfghuRTGnUb
+GbLphUSgnxkE/cYRoPFpMRVyCe+M8TQljtPag==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RVJj7ij2TGFxBIQZaIX4ashUMEnPhUxpISxR5SCF5aX5jiCNzK4ERRG6UskPCAjcM/jCqieLq27C
qmTGaTpcaUcgUesfno54IOnoTxDkZMAiDUFH/1LlefExhF1XPDvaM/vElL+mKPOPIlno9IJyNJc1
zEpJkhiPrTqkzb8KZEd0vDlGi51GzyO61dXEmY563+nDtGW0yt3UDR/7Kr4HrnSZOXgBfBllkyU/
Ltqsv1GP2HVOiHJjq73GH4jn9otgCggzWxZ2YJvkIgp/91ApwOMvBeAC4XN6dZXeU1ne9oj2vr/m
9sZH5pmnU4B5jLXGlgcB+gkSLnMODUbub08jEw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gyVZLPzK5/qGBvghd1xSzWzNxT9MZeYl7bwDM36gyqd97MSrHl5ctqmZZjV8VXmrvWlQtD5Wtf8M
Q1uYUw9jLLjLTNHK/wG1CxJ5o4twhIAQ/1VqquXRCqFkv0p3PNpB/uB9I7bTd4AWiaBbdAI7BtBw
pQG6NzdwiBg+PwPRZDs=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SLIEG44Bv4xTjB9v4fqBf1KZQbqfKca2IxfLjY4k9zESKdmwVnCmXrKEYqpYUxLJzCTdHsKD3S2n
FjbnjBB5Ipr6GLgGv0C2J70oz1d+i2v/Ude3vg89VTUFxsSxGevMvUSBnGTKAssdquUhBgmjAF7G
f249bTuKJj0kavAU86FhcUh+zwvj7mCkzuDzhzVkGMLizUdnLkDi41++Sbn49x7qC0fk9Eb9+cn5
hntm5QZ0vfbj9kz0xoreeY4r84nY12XBhaXYwSygISZfop41dAR5XcGn5qNOr/rSd8SiiAMMrDYj
bn5CvJHdPgE/d51yQsqPbl5UBX2PADtDQGjZTg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K6R6rom5y54yZsKd4jIAhbeBfM4n9MARJNMDeVGkxY2OqJ/8cW2x8wLAR43wEYFAHz2eQ8HK+Uod
wOl5zhtkBj8ASe0JmnE1aOBYUwHdGul8g2DXnoYOtrrNWJdyzb7UzcWutvF06RUuFZXUHTkTFySq
9cG/9L0pTjR1ZeNkI41RWJuoD/CLI9HUdBkfyNVMA7/98+qUdXLxPkH7NF1T17LIxenn+sQWe2Ht
xjAMgqFsM8iYLzuIO/iXG6rJy5W4SvrCeYbsRdCFERnoVKysadAJf87JmeuX7FYBbt3po4UMrumQ
UvSHKd09FRolFIgQRylhFGvGUu0A0do/Y1ezAQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ME17zFeYzdk7MyEYnQGDKeQBSCGppuWnQkdAdKigBsEhKvLNi54UcdCP533j6otidO3IOFIfZOvT
pMFZW8OTE9YcCi7t3SN3ESV4Ir5aC4TZZkHyt48WD7/CafAtx/FEQHYa2kknyjnkA9Pg5WKfZURm
dGfLQsQcFoVj/oZXtY2eqoP2S5YVXk/CrUH/dVkRBHNQEYPtWd4nn7wUI/CUNRtb+97SEHOSdvcx
q9+zdms5mWPPOj+o+NXjDwoX4ddjh04v7um6NEfjSx2nU8tdrSXSvP9FqYpHJNdEnzErIlKilsxO
5e52iv+pPKSqAPqzyQPKlRxZnf89sPbtqNrwYw==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Dl0p6TZc598ihI8QgsRd5Cxs37R2VCYY9gICl2cvqRWv2H8CrH9NUPD3aLwfUZTl+Yd8yrntWj9T
coqvorP8U4zO0oRGRPYsej4lA9y1iDlXyNcNumO9c1K3A4EiAXv5UZQEYGbDHFL1Nu2rAC+tKJEm
pe6NMC8VX4bchoEVOV1jra1Bz1ePqQ8kxNwemoTx78T1M1R5j2lBlNrk53FJuqo3P1RXoeJaZG7U
rPLzQ1j9mPvF0/mzJqfIZtE1a97g5PKv7TF/fI23MKSg3GyNJh3xu9dc97DLqEqPwYvKUgS7HKFa
oGwejJ0EI6BiVfHRcdFq6ZTSJAybKN5mf6PLjQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214096)
`protect data_block
ABWlIQAAAABspapjsX8AAPbTY0Fv54I0Zc3I1sGq9lx5qQZQndPgvFHKTCgNWaQFEOtxdQiLzMH0
NTDDTgsxOcAswFeD9Yztn6ntscfwmOrHaDXnaJZyWNqhrRt3iD8f5G0lNsMADqr+eI/BgmSvmv5d
8OVqdJeJ0khZ6Pa760go1zDz9DWP9Q6zCbSqi7EyxOdaWGfbZWCF0xzA4Rsp0M5JHHsYzknDNhHP
+I2ltLOHabIFGFMAQY7ox5A3PC+avyMRUHSt0a/CVeG91z8ELKPTftwbl3ucquimqNqsHSlgBid1
D05R/llMXuqnTBv8zFuyfZ/TNiCpQBwxktz32ytini/X8GGChE3sHrZ9cZ7qO0obK2hf/nH0Umxl
BihXBgVqF+JvUP/+5nqYaThqs8XMkBm7kTXtewNF+1aeTQqg0GNBE0syahOsPByUd+9+X7qPzNmt
vbE2GULRu/Qw+CR9+JXmSiPnIkXCylSOyzs73ssZrdJq3/DPlrKbyWlI88BV9arsf85EV5bCCIhU
ozHM1qZZl0jX/QZpWA/5VDBGW/60STW0iyzn+trZVcaZmB5KfN+Gj8loOT8OXAS805jwWCTZ54D+
Fes/GiF+8pYPzp+M3b6NvADP1WXPyYVFtAs44CxyrP5GT11pvAwg5QiLVs2h/iQXq5JXaTCFDxtM
Bk5cc4+yx0cH66+d1wGsrIXdceHlfYSBAmuG3vpSPM1kKJcS1Vmn1SbgFRKfKKgISFltSVISiOdq
QDPBpmFSoX22LZcZ72RYPo7Zg+zr7CRsrp20/ZEXU/uPs4EO0SeiV2V4OGfcQtPviDxT8RyzriGa
zNGNXbCSNEpGgzAZ3FaBtEjZhw6JP9txIK3ZGirajnb9J+UBE4es5VvArGaQG85Y+2BNHotiBAya
zPKKbnvhbKu1DeYZJCo9q40xG4M0G8d1EDLJUveXTZJ4xwx1s+temhjIGAYFj2ENPM2TmRJLHe60
a6zny7A2SAEyhfQDS2nrpnckvAQ+ASqJS6afhCGZy4wh7F/zC9xVEZRFuC9jyX8GZMJNx3wRFIlc
O8Kgz+W9hetCv12OXaivgjDu6TpR/NTl8p/FcTZB+FmFZplaWFwTchZq3zE0rMIk66w/H2+SZfq8
p5UzTXlo/Ll3jWxTXv919Llkw22t1Djpanwg1M4Cd9PEP53LztDQXZYbHMkp6/OmTjiWq0FQ6PZI
I+jbSwUs/MfECSBLXdoqX5qtZWAYEI4sIiTiebSZP1BMnKzA5fUd8PwCyX6upOr/2V99QghVpcwZ
13BSWi+58Q8fPNsYgcRsUugrBmr7zCzJIgJnoJMj7QY6BhznT9lVC2UvGQacokoWwAHeY7Bk9YoR
mMhKi8iIymS7iWechdHSijFbXLTNFaJ5RK6FSsgrwNxNaOyMjVEGHAsexco6n/D6a/zN8UNYCzSd
fV/OKxqibyhfcOT6sYj5zq9ANjSrlWSRaRNvNtPjEThOPR7CjHiMjuKmLBdn4KB3+SPYCqA8NNtf
qOWQ9d04fZw4BSEN6zRIG3irHO1LNy5/dLWn5gHu8Q5n8esgBDdmxAXJfRTgwW9T2HnC8oJgeh6u
VVpfQsQyTEDRQYJbA0tikr+/Fx1WOdp6QAhufC+2ZH6ejU2BldggOQDlZPbt4gVQ2g1pHwu9Sy8G
tJOJdID+dn4G+eS4hjf1Ah7JOgsa6elvkbAx+tk0y45MAn4Tq5+eFNnXN63g9B4u/xNAyKZdPlil
tlpxDfqXNpv6ba9Gztb6Mrxd0OL+DqJf0PCQ0zdZnM60mwKY0W2tOYSnicN4OW8TI3OhkJ0hqSzs
GQSytJv6oCr1n5N/PFcyqT7oNAlI3tX6iBX5IhzoO4dqe6nY+iip3M2kaiIHgzhGMfIWAjKemLOY
TSCsZUX4/w79A28yfwD2p0qRu898gBb8GA+MEfqVzITrq1zH6UhgVA4sTQZ3ze+71b+cTtOaBsHu
hmX1Sx1wFR0JBzDNF9r6ORoJl0ToPsZYTP2SdCQjmpem6uc3YK07uvwBUmg8LSg1S5olN6FvyzXh
DY/IgZnxGWnVwQTB4B7dYR6d45FhJEKcnM2P8TzuWb0DsRT4LuPZCy+NPUtrZiRWX8+vMhXNoVCy
hpeKAzGzo4J3gB5dCdCvMX5eMNy+WAoRj4XIGKFaJ8JHvmE8j9GDTxRpbkP+0xIL83vfMFdlTYhm
wC6yLjDxb5Tc0C++BQir5t9OtZ/RdBnk3jMY6Rpbna6kjNomU+Rjw5ShKInCRyGOwCq06k4dYsj+
gsO1vRWttt+iph9G65Iu+0nlFsnb2lsQYzooBrEm1WUpA2cK3lNI19pdJ1JYArzEFSfapMw9L1na
bxdUHrB0JaiEjVd1MO7o8Ad/BCP9wMLPkWr+cfa7piLV+8l0wChQfrrXOH2lsiHJW1iG6z/lD9qq
u8gCa9T5oPVvt+wnnVZou90tCybfZbLJHr9XpRybE4GfE0ZyBUNZBjkMUHq1h2zP3UOzjUC/+kD7
sOb8PSlAk3AFiHCZReMa4S0ihHjc6J9CEtlM0o514Y7xmesfc6Mj/f0LSczerRHGvPWMhMWw8llN
u+Nj5oqOIDtBxUIILTIoYkQvKrP/kcBk5qPbP3H0jmtlG7HPJWu7LDgSMKjz8frEz/BXW1P3/bqp
YZsiahXsHJdVpuyS+VuppIklz+pB7SnHbRpc8lWrcROZck7aHgEP6jzzpEhIsXfWy5Csov469W8w
CVDV4oTCy6ZnpVxLGgNjnAHTJOATxV9ANe15F8Q3mGnGT9s0mKzLTXjj4yVxu9PdikrYMJSTZySV
U4DG5cvG2nqzHIg7HdvsoVfIdzkv2v6yAsgP3WAaJ0XlPcHD3MmG9rBx5OEZ/w3zMjTMFGWA0Vs9
MEG1GWt392McqyDl8Qjq4m535jXUA/+Sq+sgxXiOTS0ssfhI8kLebu5XGwSHm8yT92Jj2J/d5N91
SQxfMJkaaupn6L3JRutXd+zRQYJfd3ij5bD8nyw2pRUicbD27AwRhgXh9cxEx/3YGlzZdzeoiZbF
chtrAI3GKl14YC3WHbSV9LxMIVPK/7hi49NE80Ia4rDme3vqGw/1/VG/q4eLNzCb8JjOwD7GZWKK
Pak2SZ2XkS90Bg826J/LiVcB/ziso42HE35zVp0etnSvZcLFGNRH4u9xPl0XzErtIwVOirY+Ov/i
DPdZAVRj0vVQQ3gJTuqdpVnZlVKqBdNs37Zvp3WivfpAom8Y52THtiHDmhu2AE//u0VrLzM8WRWR
uN1yR3zNg8BfT8mSPtJmO7qNJk6ZgXyIwDkYzl+KpFxbGtZR9d6W+L0rVH40I1c3OTBd0plnAyfv
grQa7vxEzBVIRfeobhx6pSx3oCDippFv9KqLNTQH4IP83hi9Clz/XeXH6KM+ioZLIaFSuH1msoqj
DPb1YHrLxyYJdQTY7hiSICEOGw2jZpaR3P10DIvaS6H2kqlxQNiujDoVzMthyN6ktnjupn6rrjzs
iAMBUa/ie89Byz6SmDKb5mXKQxx32W9cSSNVX2tzdHvoG2dl/SbOi/oGEv2Hyag7lDOnQdylAkIZ
TcohNbx3oKgntZe2wZtkSgwarvgWql7Qwpcws70KK8d7EVLe2MHLhaV2PAZ/UqVO3PoufZio4aUW
RFxmzTr1J0xliUoG8IOTvS/AcLZTGdeOOZRokBpSMF3yRny6YkUrAaYbQAYxLaqXDcppbxch5a6L
zZV/zIHXrbyGIT4wbFnroTwEvrh5BZFp4+8Q8iv6IYxgD+BH8IKsWqsXW//AhRFip9+9qYZu7SMw
IBOlXzAaKl8o7cMuE4StA2uAb3QlioMDxvm1N6wss4wVhv2p/L2tQ99wVXhjr0f4+Ix7XjHxe+7W
OlEWr83wyupLve/1eTVeoML5VaxW5GTEdM6SSMDRoKi1ZAhtQRFiUm8q/dbzyP2w/L3enM27qAk6
9tWXBAmbmMIl3r15vkKi/gkv/MRMH+QreCer5zJ3S0jRRnYCpXcbHzmn9Ckm+5QuehCbi35fIiPq
zQxTbhZQmhttPbMOnqLCO5QxXvQIuZdvB8c88CCK4qPHcscLLXtHr/ex3N8DYrCXhp6KaqGAShKu
zxYVD9NR2izCiH55DG7Jd0zCwfKEnQ71GVw9quXXQRxYu3JqitLYujj7Se/9g4TqPED/qVMwUcd8
darPF4lNQ7Mzou2tGn95m3FdpO0coZOhiwiR9GRSbCrsAXNEsFLi8hCqaMCziPPQw/WHE+cHWlwT
95Tx7BmUUjY+eBV1eTKONURqJvNd5vZmVnvU49zwACMENpgZ+oqrb23PKVRt1b5k8a8wCPeZ4ndM
+nEsb4NQb9IA8pOZBiu69ZvjLG/yIEOy1KnIV+ik9Pdc316nDI8ODClx9VwVLzFQEYk0Ec4buh0Y
cPd1QxMAtAHvafbVnco0fLkouY1GoDyrz7bvW30l4pbW7WWl7biYWmHgxwCW/gDmq4Banwhcdlfd
/mBIFSV/vAxQlCn14r6PfOSgZVQPA8pyjtQZyVkb8u258e/iTJTAv+1xW0ckaKjROWor1wuXq5qT
YA5/PpfziCuZ6sK/fVjw6yIMqkLjQvoECNmq6J9F96VAd2ywlSYmxaWo6b8SPtbAPyhACzvONRAQ
tlc8ZfO8u21bGlHkkrhUKfnayMPJuRwf55hG/53cCxoAcxwM3JM3OQEFxQMHmcJL+PiRy4TH8DHr
QNVS7ZzAPB0M4kQArA+vVNSNtxW7nCcLn0EzBJXn/SmNjCRZnqe9vLckCQHbUHd16aUSHQGIV0sm
/Bl2ousKiZgbK03CjrJl70LUoRRsEJXb7Tq6X1UdgSSKFlBTQguCdIJWkRnISAPGJ7TgBQczGEBo
5dZFIp2NC6JsnYXu5oLerszl1YcHKpYokwPsa0zv1iTHSUFq4xEhggj+fG8A1QaoicAR6fSGw13a
8DBvx+avKcIBJG/JuJFBHtONzhpWhXPBHOqbYWbWC7OIa4/uHkUojEFjwPOHLJZ5vbThfMvV70xG
GfFyKPlsiUtC8gRynF/p2Oz7vn4rqfq0mBTsfH3ZRo025oJriUT65umNFxqRXIy620tsjbRe9wCp
WLzMgiNgFhl9RndNVDzaLS6+dUuT+oAvimyOZynihFXDX6/6rWYP8R8dbEfoKgvYwSxeBaXEKAub
WxZq79hhiMPX5fiyt9r/gOTadUy7If4eBkCxADjESbnLr3fDGmb5wa7gwI2WkUpOjSAMcKUHrbwX
qqvYQ8HM+4eRFILSU3yCajm9gUDjHDzrtxGgTBe64Jl9tGaznAnwLITvBNV8/vnwfqCkykwNmeky
QWJ/Gcz5svi6Hk2vLfSUA1L4OSYgADqslp4ysSndotAnsyLy1bhlwjLvfY6f9qG+7MU/APJPzYCR
T1HwK7U2j2iAKOW7a4eOXrWBn3Y3ylNYC8SJYvHLItZGJKBFHPvT2EzvhhMUVQc8xaDaEYjfXrk/
DGk0f3oz906CpILJOsC516IWCov6abYYflA9qdQPPHeRC8pCdsx+FVIwLN35RrJ/+GeOqYkALJY9
7lxlmg8h9zELhV/rf8BRGFNiwJ1iElF6FdgtPvFf0UzcMXAiW3xNZXaidxMfGgRx4kiagAmBMerH
wH18SCyrvz7kZ2BxTdRHKckuO7rdpFYTngCCCjUULsezgc8ytEc+fP2tmEZ/6lnHK0csbidI2p65
4q62JbOLyhWQZxeNtQS/dckCzdHZD/EasfY38z0C9bBDGnLlyXm1js3XWsXzPVh0lm1bx5gri8Yk
k0vz+nS2i7k8BB0qHptdwjAdq0zuBG44fhlyDMl9TZbU2qJrTKIf/t27sZxK0Ktx6i0Lzx6sgHr2
k3QaAcFi/k2Xt64lDevsXQ/72tQ5Spfrybb9Q2dJLR9S3e92AZirs8Atbj6lgElTHeLj4P9yC6ha
WjAWdp9LXCwcwz4Qe1FwakN5Z098F2jbauUHUmRWgB4VSE29gVOV4Q6hOwFAi274B04gHSN5xO9x
3BAJyGaujOvsSzt1HoN7sPTRQkE414c+xZvuBV41j8YgB8Lm8AuHeUpCJ05+NloDdoyOiD0yloWJ
WuroR08p3VKAJ3tqHbd9pN9iyn9wVe75fxl2qXqjoMc7HX69ttG0XSy1o3Iki8wOEAsrS3NdybLp
JGerPntcH0fZx70YL4bkzveH1wMN1Akb5jhfLJ1CVzKT1lzkcTDo54nMg1aFCLBuDTIABpwQAmEV
iBme0a98QPNKoEV28Fq1z5S5+HVc7Nginc13md1Hvoe+331jr3sRJIlDp+ugxcwVwcgbbTNURbYM
Bo11ekxMnXAMCTuCgor/Y6ojCl8AAPBtKyc8ZXg7BXWdZ7L1fUtiVHYv8+3tgE7OVEASIRlOBu6H
NsWumaPcMfUAZMcsidQdludvytZOS7EGW86PpuLJ8EmkY/OLDexKFJyp3fXI0QcuAfBy897phgTR
kBPWo4CPxKV93HhH+9OqD+olrmO8YIu/JQBVDIjequig7NbiayXFfTDGHZfX8jrh6M+b2eMnvTYr
u8TdzrER/fRQaeCdkjLXWkklkCWjqPPNbaFIy6DtuauNFKTeTQ975P3WLeDP3E1c5k3/3RYz/R8/
pMTKj3ZMzypSRCEuQE2FxbPtp4+jk0+hk8vBwOoF5A2Tu9PR6CMKLJjZcjGkYoW7lh6PY2zELW+h
cHwmV/9ZStCJPp4XhLk5uZRzAp0x3WUn4SSer39mfEifgZ9SzMbsWnOf+Q7zZmZYC2wtNSsx59B5
0ktOuf9wJ1XWAEia9rkitXfrahQU2SuL3K9/o9Msyxu+c+/R/EfMhxgwWpKQ5aHpRLg6sTSURSZ2
h/FVUDUqaxCnfxtOZqT57ExQzbb1OGwbLyIkgw7eFf9wLCCAfyqCYmkrTN0WQVwUHZqOr3K1P4mv
brpOiLjI/gO92qOw28v8un31UEpVsMFAtGjg6Vu64icFl4GwPZgURK2+ZgWd5B073nc+9xihBEkl
o0ifeUAL270ZwSURlD9ZzrbqYr7UnnqrDz6xkYmKhuoFe+dTLP3fHb2cCg5EjxgZyt9CTtI7J1oH
//5Ff/usmc+Ll8eDzhOdOSv/cmkANjI/J3e9OyOZ1WEuS2xS0jDnXxZZtMoeNk8yU4d4HAIZzYmp
Ye64R15fJPJ/d5MtkAFJtELtq4ZLPWGoiRWXF25LXyqLugfuOJL2PerjARy7m92JMtDSZ+vir34F
KTjBAbR7J2IakScsPSvvP9SxBRtCshCQiX85F5mmRucK8Ow1jObevhFMT4x+9GfABt+NqffQSrTe
1CEpI+eKZ4bv7uTnxdcRFrvhs4faHWbzaURAWaRWV34Ym/mK+z9QqKWpdlQMIp2/lsaY9+x0ekky
aVpu4IHXi2zB9BWr+J9FOohuCscc1G41scjIpLzPyZttzQEAdmbzW/koCFmg5BptVFD/eMadlCLm
hgpFDD6KmfQpymjI4m9Js4Xr1edqsgVc6jXzVocTo+D2SmBROtWDB6DOpH6D2J7rQUdHulQvVjA7
dTY4RuVyqqaGUoy72lXDA8oOYoU8bmAxf0MrqK0ruU+ELOty8C/+vBI+nOM7Ro+C1DZQ9MNfMo+x
wXxtJVZ2fPDclNqNBS0tXxPO3t4gTlkd6jMCb0ckQ2lx/bmwmQu8PhYCM1GUTW+ugcLZ+HXN438i
p0WGHnR42NjmfySWHoAY260F6ZcK13mDSUlgtdT2VDvYDc2ED9hB5/0We8xi15ZDmLhqwW2j/aJm
YMUpMeTRgE/82FP0K5f1cA8ZQUZpbUB27kao4InbZ7tpE5i0h1zAv+j3s3a/pC1CKpPPqlkA/YXQ
FPWkit3pyQwBt6m2T8twreVdMHKp7ANExNjFXoXb4MmkU3OPogqmIPoTXsZiBlLtD5BAzACCOOGr
MBlN1OgLx+Yj7vMqLfnhy4xEu+kxBzaIxVgVVnB1jZ5qOnd4Jkr/u+2UsLQPRKShprdUagCPV42N
R8trNM+q3tEu+xZmoYmry2xeyFkWxMZrylb7gjyd5Q648hb1HmLpPr6Hwez17ExViGchfOqowcGk
dT1SUCTu3zGhAsbnwZJRO+8b46dlx4SvrN4AnfOpYqlSHOPVWSEIT1KvuvZy4iqB89uRAuii3DnC
KdaQTmivBcshxtTP8NprImA4Mr0od9MoRRSCPuHkxLqLqNtSMVHoaxBv3h/F2VCej+AVZ0ARDZNl
NiyWPAJ4d8gEuBlmtGTPOcT/x/J/B3UDLUeEhOU837hxcdRrRjUktTP697LgYz+JZQvcqRTuYgs1
wYbZpwM0k/jzD2XLKy1D3MijWUvKZR3H1v2Lgpxvzbvmx5ELWwRRjOErRcc0lO5cWkPq2v1bfgQL
svbdWsJlaIpDwrRkNVRmLP/quMTauOm0+lvscdu4j52C3kMmh9E1uR1hncnURN0kuOefsNwMVm97
brleUXWQKORvrL+YGSD5AdXMOLq6E5yrLubDH9YGpOaJUzEl5yppGiKiO2sDW+lBClXTuLtcUet5
w+QZ3mI45//+PJA+MxvHawZKlvlUkgYEZbie0elWgGR7LsXmpfGkomLCX2/voiuHyK8zMVLm1Kgm
to9AlASAUN0IpzvVEBif9KXJZ7/BzhCL0NEcrtCuwBcQMCbT1yZKT6RGzo79+qLjMBCz2XI3HmVa
66ofBNXB+Ovrvat9cM72LMbPEz8xAugXmG2LUuR3n74H3TjCn5wXfZAyaklAAEQkoPC093vUW7N2
G66t+l7HfdcHpNr6zyXTPuX00zTUzlINrg1J7IotxojgLWoAWxDPzKYyu0Sx22/S2nHPgdREiZ5H
Crq3C/gnHtj85zUbeJnLAkJLegKkstAljh0Ms0+p+v373FXM6nwRBlVAPQ+XeOOpv2QXCadhR1el
cm0VrcxieN+L1Uq1nzLd6ayzcyPMzKi9kenZ3iXj05h3w3xx/4Ixl4bVG+WrySus1s4VznNF/yWZ
8GsCNEM4yhcojInpVz9vBCbk5VImvHJi282DpAwrqL07jye/jHdTuxqApOIdToCcD5BqQW4LQaEX
m/SK0+AVgR1xU2+20GmUfvdzDCWdyGpG7SPI6xeZdAICS+7OIZ3YoCBx+S4HwnFG1nB7GnQXTuEM
9oDWn4/dQrIMELn+uorCVJ5zHooYKVD0LVNjP4SF4ELvGMSNu+iuHQm9DHqEttJFLONHhorDuLdf
vCYUgnGEDF1dC2AbfmhWkvWInQpn/TrhMa6KG885+Lc6qqdufGEF2don4nFe87YgZMM2N/mgX7et
d0LOhtAoeFAxcWtIv5gbIOV4wyp9F4V++3NIQW8hhfdEYKGqAFbt26wT8rk0xvbGblydsy5byuXV
qOZnIfQCP/nVxHwlK+Ne8WQ2t0TxBCa2FTqPIqaXHZ/kwZomI0oajGPBM0b0Qd0a2y+ZZjoCPz/Y
/YlekEk5Rn0dZgHLi5QSOX9bEXAPU3/yyOxBvJoRNVQ0jqP25JxNlmyznCPdd2jfUr8T/bZeskVs
s9CHJx69tdmLQk6amtHmm2nfOvbyZ9eaZrSzH9ULNus2xfKGRB0gmJoHKaYvgJAqW1OKoUh/X89x
9RciIkNIvb5CLtx2bYqNbr52Yk3aXMBUvSh4a64pnE2EdXTYHmPLS0trYaS15KLw4ZTG0rkvkAS1
MuUivVH+zJySMOkY0YuymEXCtrI19kC9gvK/Xton0b+rlpK9prT8Dy+xH9iuQy/KaVM5MFPC+Qnp
yH2WF5XibDOWYD3Hkxrj97Xa4Z7ZC6NF68PzKdZR21SEJsOXwFD5U46d/oWXm9ruWpsSigTs4PP7
WJBCvsXRMUYe76tlUick0UF0edHsaEYPVCuuuc4wJauiFIe1FiPlQNa+sLx9X3N1THBgs7O9i8Pl
Hm6wBj1G7KAdJddqStpWOJLp1HGgPDFgQkyd/rbds2/ACy7AUvuDlXZp2Lg7MKFaIvCx47ePFYSU
TxpgXBr4gVXij+bQK3/WaUT9uZs9V3trWuGwdU0lpawb1ol4h4PBM3aDJV42AY0Y2wKT1GQhggIa
WC0Yi1saxI3UyWjEFXMNzOwUH1xSDDeQP1Bk5dlYjKQTV5b8nPVCc+BUswhOlTrosS4Y25U9pP2W
8LNmCWjz2+pvnfWHJxQKpsSh9xqEU5TrhRops0DxLWBpG4tRu1DBLKer3952J90NoKVNkpByI1nd
zMH8mEEoqWNXLLwOATgHCW08O6y2EBlTrx7irLXpGajAjvh98fC5nJFkZnca8WnpNA9FAFomsDA3
6gold1QQYIfZpm+fDxYbFd9y1/wufcMbcpteK3Zf816Umra36Nl8vm7GZE+7U7f6572bFvzBjSEb
iX70fKkTeBWBvgT3AYh/n15cj8VTp62Kp0C5IhxzO+PQgkeO+75TW5cZMDb7HmJfZrpqJCjuWLg0
vir5XaL6eYQlX3V0DPsqRqsMv9Iy/yOUPJ9pYo6M6l8ivrpF1N1mbbhMGcN5JyW6aO7JOFx1gDMT
3L8LwURsK2l79ZGN94deYm+3hTCH/NMW1AFPe/MQHDyc6u5uZF38xv2Gc0MJ88J3aRmYp2B74G1v
uJR2GbbF4Ixc87RQ0mBauw1goHydrGSYusIUvXIrPUMA7BpAdFaVCAgZCacq4n0P7mZlZUgEyiNU
CjWSixvtW7sZJEbauRkiEyMSobRS0BD63WdRmFWi07OYXVicYZMAwkiVi8/Cm7GSbFRGI0vK6jEE
6fDxJ/Aqr0SedAC3TUbTnqXg4Id1BSsOlW1HPNd46iAAyz4min+X7hwvzYt15FKNeVV+0S9D719A
tS9bDCMMi0FlyTLydZZNSoALE2uu5KIXn7PtQRVumF7mc41dn47QxHHA9dtBNcl0CoMOG1LItogf
EQTQST06wubZopt1JcWV9Up2thPyX5j2epq1Z0VO8yUJoLyVeUjMiu3uu49sdr9/A0cvzgGAiAjg
NOWDAoJJhNoH9eQkDY8hwxk+2GPp39l23PW1eCvYQ3/+ZDWA1lsCu4bRwuy/C4VLx3kqbTMu2keC
nzPkDjL6Hqbb4SdwL9J26Ux+N1pyEy9dHfV2DVkHXbhRSQ08nA12DT6AMUsOl/kk5gn8KoNKkQTm
B47lm+h5i1hw1mkU+75SxRrO2ws4W354TmjVhVbox2B55iNaWKorrMkUm9gH6xvV/Y70e749kCNZ
jo3SqNKlFtu3VrAwGZSdz9MzUaEGceNeLA2y3ZxC1ehjAeW6aPN+gi8dhvI5PqrLzR6BQm0eLj7B
srCq5MTumE/zGvd4HSmkY7K7nKiOfM9xTQSDweR2Pc1mChV8SotjIITq3Mh1fOU5Zd1x3sVDeKQM
4FEhlRep8Lf+0wqP2OgC/LoJ97bOwUGpSYa6h8dXn5SssNm3s7JnSCxqOJ1jxuL1Dm33DdAuna/S
nye0ULE9nDDlpOGrjGc3wBbmVkxgzVZaIuBDh1P+msPpMcMNQNZiqy1tm3D3OaahQ514HH8zLhqE
RF3qN1hL6Hh0KIuVnvE6ni68aj0JDQnNgV5hSCSmN0renhAHtsxSQy5xqYQec198lHV6lDTMzfEq
KbJFTavGiEFCkFou3yIZWRN6luokAc7jjsxm6sYGF3Ov34LdaD2oPSbreMIuJjmgl7MaFqHp7kTu
cBoWNKgEggyi5lONJ3J6W0BOeZJNYXNoA+eU8XcT+ZiUWZDC4/AkvvsSRFsznJJXnVjLQVG5M55C
V7XBqcJEqrrbDz+8cyPJV5/N6PePvIlYV2AzZfQiJzmUJLHMBXuctHRfuIWVtjpLvH9xZ8CG9M4K
Ibi+RfRPZi0eTHq/23xi9lwlV8sjLitcFXudh4SbVHOeO5Ow0/31iSQXC+3C5EQpaohoHctMKVUr
+q5Xg94u1XKzUZ3ACPqnOC8eL86MX1A8dAd0EFTTKlZE/mqhRozGykqiEJJvvwgeK9dNsBpNtGBT
V6u2/9N20i2+wHc6Xvt86MRHaWo/p2Wpt7jXNa9xVzgmkTFZ+y/iwUFIWujMY9iuCezwO2w8Put0
DuxciEougynX1Rv4uvAoo7qfFIhZ3GZkGMeh+iUW3kDsS+yOsDk2QoVDP6FUKd+gkUPyT7BFUisL
h7jSBPRaZDqfKGSCFrQOKLFiEs51AdsSSpzfk5ilax+Y8PQCMmHdB2+hEVEB0T436BsDHWzwX6a1
QQvL3njOuopICi1ugiFF9ZO8TxbC4IDXSQTfmO8hlr+aVXAGvVN0Nyps0ER52gPM1aiuxZCOl3bD
vqz/mPFaAREMW8heN+In/CTvdSugfA4VJFXoAgfkKMtfScrMl3cGRd3SrrcmYWJmz48rp0y5TIVI
RlVNnANctll4J0Gmi2cCcVcvpaDFHqPiQhlOhU8nfYFF+uRxxYP8Vb9Jmp3Z1S+KZP/cJVhAXSCE
A8AjdzovC+ZYASoS1muk4ucMatd5rbXn9CaWGrLF/+cH7Fk2apt+CJcb30JQRf7bo2M3oeAuUF4u
AOIcBvEKSCtbRjz6AWArTsk/+T+gjhsutclWErH5VPJd1gxVa1rRDU7NeGuRbvak8X85iqBpwISF
fdccZnUKGkt6LVqPSrWRX/lsDZhmEG1+gUy3ozbpoMN36W6s8URSTX1GEBQIUBeqo/Nxfj5Eg/Gh
bUUkEejzNzbdd5s1+Z9HzoOlug2UGAEBeX+aagQQ3Yqsc3/BzXh33I01Ft87ZV8hy3uhvspSp49h
sEiiUSjN7vObq4ge7XknTJq5S2xMHrgZ59BrM0uxo/zdW20kkG/1d8p5Z5VS9tcuFdZBu9lsuJD/
rYXJgr80uTC8ptGaPv+HLTqbm/rG+g4ALQF+wJJzNZqM1P7NT25+UfPy5NL6mE7fWsOIgCJ/U6Ah
6BoSNQg48CA/9f2tuTOgamAZWESsM0zbpqALMgj8VBsGB3sx2xgCpXsU9M7OucJuY9C4EoJk56To
BlDfeG8s2udfKh9vpgXlvV8QcLSWmYPeiFjkgH4bGGIFZ6J6Snu3B+fYPxhSMPLucKRNpEVVmPFB
n0imXI0DO0+YS+fHMPg0FWCbXwn0QHwTrslphZirxahEFcXaggr4P6hQevdLt4KbjkGsWbFoug/K
RjBgopgj5SmCX3a71ULEuggofLm04Fyycl6gvnJ/o+uxf20yKwcJX0dp4btZcZJ+JU/jZJBdpoaH
v+uM2wTlJvesn1u9kHMWTto9lfELWh/jdZfCDJuIlsYvYe8EGpEYMR+c1012idAoyYM1DjRqli5H
xFgBV5hrS9wiaKlK7J7NBYd/1iR4Gtcho1qHnIkQsk5GsephP4oXxDNMAwEwMCtFYCBXxEg1Lr8g
XunQS2hLhiSy6b0B1nvMJnKlBDGZNxJG5p86HtT9d1AEwNf6n/FBiR0Q8k403nh08zBFvsvxLToA
z4eJ24SDzhwxP8YPDk6NXkTeo3DCD2BgzmbnJjkTBa9liAGkTnbzTs+5CvUrbe0y1ni/QO5Cw+0w
ZoAOba48DCTubDzKp0Af/Cu2u9akUh+erz85kDjq+i6JAQkjpWJnKRpNSyRjFHAtDNhCRBlDWwT6
/1xjFOu5NHEmcbra6eydJTbnknosc2dkLQCnUS4jxNyo2eYtrsYsIM1sB6RaVxaLap0daj1aFx4Q
Gh999EiCgW94QawkBG+3e5Th8x6XE2z7T2OyfgG04PldVWVFXgIwUxtIFYjWgdF8muxWxJkNamUH
S9CVfBfGGwVnK+8dTexVW1UYnGb6okD4PEDHg+H4sq9Yu1W4L0/cZgFXvMeN9rI4g6hrGkw6jRYf
h3YM9t04Qsq7AiXYqlfk0Nwvi9dn3AZz9nKfLyO6ihL0u5aq4iEx/wZ5TUcdlq/Czf5dQoG5O1D/
aeZ3Wr/SJgASevx9VTYTgl+mMAroH9+uBm0sjmkAslyqfuA0IgI5JNUBU7hCdUmdeny8terAXaab
x2CQk7AJM++twmy/mSMs6rs7HjtA31X+KB7/fYPtbAl0QEIFSm2kk5ftbkmpWM2EtOzox2IzTUB9
FIRmQv9rnwVPnwy3YAlGF5c9hY3HqO4w35onPBe5gekOFb07OTH5GAG2qyKz0vPRzRcdTL3LkJw1
liwFm6RdhoVUlsshhsC9U1TYHk6nnLSzmDSjRaZzRt2u9t4Kl0DwEjqmbF94nb3yQn4pylIdx+sv
vvogVFVXqoY3rLN776sIat1GalBWih8wdE+vkBDYGR2KUynd8eU4sOfAr8eB1TirWo9Bi82kbx1g
PY7UTzhGLfWcgTAONhFNBzvRlAYOZ2RzBVFLYUGDmqVwyr22eUgWEOYO+ItE0oLaJg+ljW6vn7RI
pSmyENMrHU0yPFV3G3EiqQcrQZA6hzbDavzx/sRHFKozc+wNohS6Q4UWLucnadxCjV5GytOMyoMm
42AdYyw6IQ8j2TxeV1UNGdXMZLSM9Gpi80Pva0ywD065FEROLLCKEHGjPqzHkPn/EcPTg9fn18PI
AZvlMmPOdw5xvoH+AHY+1+WovwvIwZ+t/MYhnuI4X1QszBTyWa0B9KNAPRoVzCcex2urkth0hMo8
28HzmkdbHnUFm4vnL/Vzv9Rs9R3oYg7DeO17V4U5lsNGTRWGrQE/fswm9ZNOxaRx8maB34/Gr5hW
efg83RrFeg0bdTt1JmRGxsxsSrbQsPoWDMHnFUZqHGZvnu64ZCq2iRfXjqyOKyfxW7Au0irKGwDo
HOHhvyi7y7G7nfyeIEWYhqgWoEuBhaDdC3qyFxrnxd3AFo5bWTodA0a1CSdUvnzdfmnv845wN6GI
2/ptGVkNY1xR5RwghMrZhgjR7WKlpo8c4yVBjYwuQqQKXwM7QpppWaiPJGZASLdzrsg4J8toD+1N
X5G/XFXPRiWTuDKYg1yxdm+qYoIrbxXGJ/sMPCSiru5blh6HMG4toVIoCZw0D74poK9DzbT1RW8A
Y+Zx+baM3LdzpCY3nkTpukGwmqbmym3b0OnyrJLAVfe3elu4G4JwI3h7U30aL31fy/SyNM+d34Z0
VvANdocRElYJm37oRlbPAMDfV3xwdy0LAJ1B8nH52wIvlJ/OncdczKKzh+oOlihO/PCguioh+duS
Fhruf0HGry2pzMIvljXshS7aptWQ3g+Y0w782gxINDr6X8ewOHs6bKir/D70PhCE3FHvrtojR/fi
d123EXKiPnbdJ45jV1/bTJYhcKG3h0EThkssPq1XLI1wsPZm7ZDHOL4YfUhv3tBkDsFiKFqFOhUJ
uvyjGavBOyaXrikwWTZzCXkC522Ex65K/U4Olk2bFdVy24/wjLy/u/3U+pk3toNoKu2YEK4Jntqz
bKMEmeNy3vY8sdN2htiyQo8Ozx1xjnH9s+AWXdOtXq9e60XhBVjWKTxcS1Gtfpfnmq1nmUspc0oc
ewtOduSqEWruzp0IG7njhuGfr3grdEp1vvyM7yiZ9hDk6VNgUodby0OroL14bh7D9ROKVWasIjCh
8vtV51uNX6OyrY03CtPZnfLsKQNDUoT6Uw6L8wJmCKr0pRxPycQ4kvc9KhQ1PkwncgMQfU0e9cs+
aNQ1Jy6Iu2Sc5ok1HoqCFp3pEr3xYAHMoe9dFlXR/ucz03bXMeL6slV6Fv1Q9ztd4EK1f1oyo3fU
TYwyAhOKqeFYa6dR4YDNUsE7PrVMSc4ka9mCXH5GTxHFpf+logX9smOAHBtkgnm+r6Hu6C2ECKrg
RUGvFLMOJacBzN2zRn6e57wQvpnnpr3e/90g4G5CyD+lrHDzs1tBhPSZdHFhI1JZlSV1Ut9rTC1C
Y7/WxgCbSwTg2fFjTa+NQdvaiXTaqFY9IxbwTWfJJsBBp1hxGtmHlYGv7NhtjbamQYbrKUoNsyYZ
3W4gzAhlL3ES5Y48va4iUhSSz6trjdijPBBJMAJfE83Ng15EPfYvZP3Ttm8WEuQOz8csBoB8N+S9
959hAw7sbbuPtYxrfFjjkGqyCVt3/3aZvqr4pr4lNbRQoo1JQp6Z7MCXnfcOjgb0t8H1yfL014Kw
ilI4Fvt1Dy7GYTM6zE1yUEB26aSgyn0c5ijDVEX54k72R5fFR9ee08ZowxpYPEU8cBLA94UrE6h1
zwXQe2GTfz2mi+/vwxBk7Vw4bdxm3FNpen1LdeCZ8ake+DtaHrZpILlexTFQ2BjDWRPSVDf7ipP1
3WSWFx00AYTmb+hpKmSmnhbJbNCglNH3OooUx3ryjlNFmfTl9Jb9tLN3D9NLW5SPFGGY+CQJsJg+
jJMCtNXshBXyqQ1IwEobpoaq6kaIsXfuK/6Vl0aCHgkgmTMl5istm4+jzTCS7JGbD/mR95MlQZMT
1pIVBVsl1Ilp0/J8wdt0wbZl0VlOG0heRVKLMK/CvMB2FmggbL66VnWbmmGYKfpF4QzQqPt8fnIJ
wAAFyiXRxoG+0L0/O6RA5gLvPKA00NSh7ABDnDGsX5W8iLFymdb02oB43gFucns4eor9M8ZFk2CC
SiSu/2CKEmUwiJ007qxeyfNz0dGg1s1Ogq1rAcf/hJYAat5aLScNvWuPCd4sNdZsPfuS4x1vzFWu
mlNcoELXEq3PXombyHTze1oUxhEP+v50o20gZmOOGUwegFZd9NWdrIV62NYtJAtqdptzw6vqfmu2
x1VrikYxLUq1OBrGej3Mi0eii3pMpEtIN9v2Sz6RH7GetdtRnbS/IEcEniKvdxnGJGdo8Aux/FeS
Xi044oz4MHbFD0YpdSpQuVMKp9VcBji7VerP2x20cFiZyAJUCBf3RkQ9olDtaveHQ65D/k1x0pwP
UzcmUwa4cRUfh+t9UnvPt0wfi4Qc6VBf0rqNJwJs3C3iPhDLLXg4O3vfjfO1jHtxDngVhCpkSjsJ
T1uztkVbWflZLJQ8jzgZwdzzjMkiSOGRgnlPL5HwFSjCQYlZfz0G1RCOLwLuRS8eGga+cBLolYtl
NFRej7ECxONURG1/3YJ6rjbDqfG7ffGwHKYaYfQabIta2eakYN42NtDKiX3kBP+gLjQ7zQiiNACl
qLG8GloHlhdskCu662ocSRINYUDCUx29jsxbDeIgLL3FIroCfttNqSH99P44aVDLcPii0xMlXWNl
RpaBIpC2XzahcXhun+lr6tTYD8VxH5YJyADAiW3lR8i/cXQGfWjca5mPUr+XnuES7uWfiSzHDHfz
4wnK8ugWshR8njokLwaOFVeak5yP6pzdVHPwEcgsQQN9KsebLVX8Bsts/pGu6NS9D/aaq9XvIr9+
JoG7G6mxEZcJXziFJ1ZqubGeOxxBRvHSrMPSVLGf9YyaTwVPPueDwYIiVGd4C1SOUjX8ntpdFFVx
WHBNp2+w82B39I6153tkpVMFsGhnXJhuWBU5hhXlAcRo2wQyMo3mwipLCZ080i9ktZQIdqRQQ331
D6BtBYO8zF79SyhX6zuTPewuWkdG/0Iida0J/trd9xAcJCDsCKz1jW+uJBm47JmHkgRqJVMMK96Q
DYtAip2KqH1kkfy1eSbhj8C2ZEHfgtXAZebkVUEvowwdSwfnpD3z28Z9Evcmi5wHX/LOvZusjsZP
K7Vkr5EYF2A3T3ULkOmNdQzoeizso1iD9yyOzL1fXU3KjBZVM49SzLlTiDpaK/Pdjjy9WV5eraz1
4sNl5PJV9pvujyTZRVUZyvS//VXKIFzmUgW+MJIrLz8matXE5Ol8spgruWVrzlYFyg81sDbzelc9
Ze6oQ+tgjcuQ5lL7UTEeZ1NyKcpybZ5v3hPQFNXPBQLWB7gAxixRs4hQBCkxFr6dha/gjgYb7rEE
p2DhXxQRfVA6BkzFUUduGcV1g4fY+OhUvjvrjJ94tMANzW0tyAKebW75QVn6wI1RxE3HT/q+SL3j
cJ0HW9lwwgkupm2K3232gqCK9vaoKzcqwmqQY2NKQ3gpyjNGobBiALI77LZiaMJwoYFtOOEbaSlQ
shVk1sQuQzsVWs75ViOIqXlBaVRVK+zVniaGfcJ5U5O1Q3yLf9qQGyknSlf6gJIDDEiNDFs+R0Uc
5WrwiB6QQlkWgGaITYMbaq42NYzruGJ0L9JW+tyX9QrYkHOOySgtsxDkjfydYlSRVMyu7U6cIaNy
FCCYe2PcOzut6h8O6XznuNBC3EBRfT3IPfVTAaWLKYF+yyXRlVhqmv4vsHiE3laKqlxZhx7tnuiw
YSuwaNMSGEs8fW/TdyTcAZnBLN4jQ++EXMfpwHmFE6Rom3DHSePoKOezD47JhcKxVcNumaEUap0S
NltjKL596nXPFkHaHIb4nTfWZ7NMa50AuBwPE0OpwjwfgRR1+P+VX7BaK7W9uzXX7NsKf9YG0XBZ
gyVg8HOXQ3jFmECPuH7z+YmUyyHzf/CHwQoH0mqsIbiXVOB3U+66U6EnfHpKTf4Y+6/jzKyuKXSF
mTqEwLyxuJMeZVhCmm4RszXyXakmA/LF5Y5Kev+rrDzXboWy/9FmhRbFSRQtyLSCUCwiGdTa+Dmh
rptmU0vysOsMk+KGzpUNELiVGzHanfKTifi4wJs2ffiIqtV9AKIEjEyiR7D0Nd0xmkxWZlyi+NI9
ix2AqjLfOwiXMf95Ws/hafp3bI2q9FQaB+M0x8cgrv3Dzf3HZuk8o/qDCYXp0uoXXpbjOgIwpN8O
cpvSgdb5qK9GJ2M/bemm0cNnYO5K+p0fPe0MW1jdvzWpg8Z2nLyxGoUK1lz7Al1zk62ClTwvDBeM
GuqwNJUCabBhPBm/dOU4JnAY5knAINLiODP/cw+rFHOWPRFxtqi9cnkbiaBS+ut8CNCImt/Lbsmy
QEwA1VWvNMnHkZddNMuVj//OkSqtk65E7uUqAITWprIKV4kS4+OLE6AHaqcvVdlY1vc/7O9LRM1S
YlSNTSj00HOHVGArlqvDOSB+COD6MSXsFKmPDkUQ3Z9Xe8xcWheEiODAxZvEPxCA+tXRgCZMeiM1
MK9BBtedrEZwkNaTs/GJU3uNcT0aKAl/XuP5ze6lmALUxDdcVEialP0DnlUKQn64tbuyqvdi3ReR
I/24PLAOUK/tLaia0x2sjXfgSEOGTxrcnPd0++gEnOhoa1XohJZBGxowbC444JhX9pPUFIvMQK+I
jPLH20UT3MDpxfkr8/6wllqczBTYNxEXV3T3Lgb7ovcmWVkZMb35uJkR9b7jQ8D7b314Sqyc8IvF
OlW1ZXtxFKpHYht8Jc7X0BWOu+VZD3XIx2mk3t1WEKXL48iGvBV0ov4QfHGBO98cRu28mtO5mMQS
rTzyitnzcGIvvwIoMb6ZZtco3WwswBHkeLtYZ/RVcvo+TCfLk1lmvV9gIXAxaS4RwiQ/RTEE7DFp
JI/UqkpVPyZVvF6GjEisnKowwDdpkVJFvL8eBi9zQjZlTuMZr6alZMPLZ1i4Dj0DCOnVCgaDgiAw
/Ad0dg6DHSS/Rllfiiz4iF/+W1ZfcTkoBnJ/q9J7ILnQevYGPLwNx3kAlsxpHPPzz2xJXsQwIqoL
UWChum2UZdTUX4171nayBeRU5LqmTBLYc1wPpt6PDPVJHyj10SZ+r2XxBpoOCFnvcupv39uWQBcs
yBFAZ9ZLq/6Y5Gtj9h5DQklZuxgZ8jfwDnDtnxS890QmNyZDVN6l/2YE6z6ORljkTMDyt6l7ef3v
GIz5u67FbrJkg3Z89nS8j/f3K+WZn+g7Uu4a8KOAJeh04IGmOoO3Qw/uZX3yiRtKyi3IIdNSpfDK
SaKbX8eSZcg1sIb7btARlJFElfQae0TJdtX0bti47tpALVUv3jUS/P4FMLlfjY1ZroLJptjXX+s1
LqejtubZCnwMSJuPGJOPEWxKqHeqG7clUO/k+gSeTOf2UTf0wVUQJPWoFFASpm8IUo6bbL3P5bdl
xZxbhx8bx9tv0/Dc88x3ellc7/xNIFKMgs+ITYRpWA/EhPN6UZqODDEX18gnrEwP6cXzi4QP4cNs
i7SBsvnmphzeg2D8e4vNbpCraKFULlOJkfUFjCVE1HsF15rQiuN+/9r4g1Voucxk9VWUFSeEPQzG
x95mNlJStLzAmqdMUXiAHFZvGGwx70BFQcF8zTyt3Uuqe+6pGqq31pjHN2bLPVjCflPq2fMyR3iQ
GEA5sYKIrgrypku3PW9t6oapkeL+YgQsPdzNhAH8MpSrwO67w5VHWv8mWryzLo2Y9fTHkLaMpntP
I4mz+oVpXblVT7Q8qPivFJdGphSFpIeuJ4cTbMy1gnGoLtcuRX4EqBeRVSd9gPwplrSQkamLq4PG
22o+HQ94pfL4SRFes0ADdgIWoCx5Jsxt/wRoUH1KNdK8TWchriTM1qYvYwV/oE2fS3L2ifGx+1G/
600Iny/p94gbrrvwDLc8SezgU7e2hNRK1vJNGFz+ZQ3GNh+MEo2xgt9h5J++x1O5g/O6UYGo1BFc
tevwbDNrdUbfA9FWqeKCyGvzniedzPkBKqYnr4u8eWKLNB4/p+vxfzMWnsf4DdN6ugX58+313ZKd
wX4OcimuCLW46RiR07ar0/+hySnMNUitR+xo5T65ZQGiZvIaRMmGiy433OERRGBen+PR8K94IO6g
msxTJzR7rMCjqRHEjHwNNZtKq2v9x9yFPjwTq0nflPUYqarwzbGLoIhPr620DegbcpXUggeAjucR
ElnVb2s2PKFsa6rHq6xpNARtcbnD/0kFqTSOhrMYFxFZXL8VnWU7x/xPzkciJyFSHVfwHJQJUGfE
pH6KH3DG2klzULKQo3uHv1pFC/G5pItqH7nMwXzqE1aF/s3rb/LMWUPYOQgXfEhXCTORIor+WTIn
4eLqbq85y+PKvknOxXPcO+qQzql/QPo30xvf5cmMxqx/3zFx+/N8fgvLPJNWi/bLYjiYwCv4wF2A
EN4WKmI2ggbOr5NBYN/A4bg4gZiK+NbKS27UQMXpET8HpLroY+ilheWwuWDAZ+JFw072SGQ1OWvM
29bqm63HbnPaylfTlJIo51Q4IJ+9TM8obs/7E/DktZvLz9x0lpUGfmuEGGKsbGd9JFnoUJyVweo9
IhBpbDHcE2axEwLB/mLiFyhsGCW0Xe8j4PMkCz2TvU58FunCimPS8Cud5OaMjk0X3tNJo6Nviyiw
pdY5u+rLZ7+sfpXXOybJeIiGbfPh8BADK8/it7/avZWub1pg0dGxqJLzWMzde+n6Lw8fUmZxPsyD
Z6CpGI+Z0rB38LPehI+efhlQ5mWjaXjtkHY5XQmRC4oLxiSNN+PZcdBfz5IAuHT///9HSVz7ZCnn
DbRBATsAT8GRFm6gmvh48Box7RbgOVpS1RcdsW3wGEj+7wet7mHvTl6FRerfCaU7l/a3Km/muF0e
7hF6GMRCwEMc+/tfS8r61SBEAeG7pjLOtXGlAKgWJNK4A5iMaUbgbzXNQBnxe2kGNVFE0kD7jXuz
ps5cF/FJPbhUV7QHTSYZLMeFXvMLgILjrksWP+dkZ6Fh/tt15OYQliRTfI3gL9p53q6ZRpnR04+K
CQIjyKrFIIiwuWHT3eltS6rfttI8RULPaBjHcpWnJ3EtS3nF3MiotJo/ZYKnsM2iZRFtw8t5Zovd
kqWrM1M68Fpwsds7OeWYct8ASWCfBi8QLnexT7jlm3g+bvDbeGHHKxYFVv2It/dW+pYv+z36m8za
W7YNTMXXYxjKxnKeyoH2AZNxh0MzAS8eH+n4Hcz0xqDP5unY9jpIkGkbUetf+KUOlPy5xiPZDflj
DeIih79ISEPY/v1UMDha+fplbI05tYRW0rQMZUaCo30rC44uWzqqi8MwEdlaV7+Y70LcqfU8Boq3
xINRhvjHo9e88M0iZBw0Edxb/TdVOsdSdYTw4PClXHjS4gu1eWZTiq4hmPGFfAYTej46+kSEa1+q
VSj67vySoQeA0r7eQtNgYYLGerRn04CUHQ7WWx0eUH/PnLxqULQ0o/kQLilJMKsjyBFBisl32xqJ
9wvye+c9nvrr0QI8SPiUk4LJLZi+1gR8VjS90O3KykJLQbQ+4et/NLH2LwNsS4XyjzZ+u8ZQJE7u
sAwCqG8lQkoxwmsRg8N6wtqTMvRWWtwPgBkkVlyuXyOUGJVay5SBILU2Q6ywJ/taZ86UwW7PkntY
bqQFQUVWALMUCVa523yjdQR8WeahJIVdTTECWefV0lFtG15EStsc7nkQG1LoBkkWgglXGLVfSXJb
rtKoXx4U8r9FuqqFJplPVsfdctiovLkMlF7xr8AgTvSs3CDVbm8CW73/hjn5VKllbi9zznkAIG7U
mnME7NMrd61gnifS9OSYottImbrs3Px/IIS78P0BkEJ9Kg9USI4ABv1f15pNS4eCDdWAlwNnkmmy
+Ea0sPFilgMn7yIR25rQX7KQCXMRYtsdX1CMYHjHi5zbcA4NkYIDu1rPKBFC49vR09uWN0vhxBux
GXk2WCh/XKFnie5EPGj9oVRn3fi4BwHPdkPa0IUWRCeXuXwPJpXAWxqSRq0WJjG78OBkjPuQfPZO
M62XnWI0PtqX8NI3K2vCBS0HLtbtl5xPOUU6lG+G88pryxMbFZHn42FZ1NtC7W5KZfgpZUJnHLow
AfiZhSBK+Wsw+/YB25vaVYBXNGPeNsQbLYpN+DCleSLUbB6/CyWnoVd+v1KNCtMrlLKDotNr68oq
LfCUEo2SnwcI4DtjJ4pae74HrM59Gg+ij0NJmdslfKouajSL4RObwseC7J/uqOuoF5ACpsH8kY57
mxZCGXM1QtOzEwTIFekV+eM4b7R++ge+351WRnW5B/BKbYf09jonBzROZsNiEg640GUepNLf3r2t
YXgKPCxlku/7Pzp729rIIVBwFGrYA7yVB5JTURdzRCjGrYbrwJplJKU/FhzDASkCC6wdHLZWTxvJ
Q4L9czLUQxEm1Q+zVaweFxFiJZUYHeXnkwJVMIzXmUjnAUwvl1iA3Lprlz1C7Fpf5NLAfFQrikp5
jIxuS3Nh3Vve4D4gaJ+1WU6qGa/b8iJpSx6YdSPnbnTw+vTIG5fXU5tlIZbUhqkKR4j3tWo+b8dJ
6uyZQj5KW0khA7AmIrQIfPmmaNeifEtZKdkoUiFcmb7NKSRjhrOdBAMI5wEXvvf9MxZglv1Y6Rbe
vl11q9NFc5cJAUF1I3I7b/Hj1gg7zdqpi2O+vCpAJRvaSwVS7b73syo42NtezynYLgy/wd8pPSlr
7eMRuUjsZiA6Su2hQCyEbGoEXVdCweM9nd0kGEApfpGXuQ4rXDiTnFFvPTZ62/d4BAqu6DDujPmD
xUUmipm/0BO5xpiFzUT/lzNSGb5rDbvN2Cs6BFcd4clGwIcWwPEkDxeWVuSVfclr7yMglPCq/2lS
VHTW6QF62zXaEfZIfSxqZlalDSq2ZzDEG7grUni084p0tgMi3kATJoqcm5Nzk+0V1/6Z29DfuZBS
r6ZBNAYKq+651yOgcmlY4uvXSqXHcBHZ+I6gfnB5c2nuYoT65M7Is71aVFpKHTD5Rutl6KXCNfEI
6DjAYBsrO2iEQKB3QniVuJzra35munsMCkWx6jB40PTWkEzzHtHkn8DoI7CZ7Zj9AydSP6x+cIpj
OjbIiVRRMFT6unWUyl+zfHHnTlyeiTzNAC97rao9oPUYxjLMVFKuzk1zhBl/b/ormjWg8NGarVZt
a7zogkLz1b1EYqHjJINfAm8UzTtcB4RWuKdZCjaoz9WWld0v2NJRgeJ05Vbp40iY2A958BDHy65g
aQkFXaV3qCLfCwsuu6YdlZgAvW2xjh8CDxgRVVQCGUBnOTWBxle4Khoy3fuFU/qWJsJ9M8uwwKvU
06NYxAwQkGh4HHLAnbsDKsOwEifvgTXVj8sx6u6JmRxRNKC5xOmD6sSUeawlID2Ds1G8isV8lEiH
LcuXGvKsbcuJpYm0UHL6U9iXRd0FfHNTnVKD44Dt1Wj8moL5LzN/xWJt9g5wwl6NNEGptZYST+a5
LFSTjhEtMn2ZirmqtztRhR1bv9sKjx0cIymfGslwQUr6dAc4ijjtwyYiZawvFRZaP+EhKTcQV5hi
7MIHAy0531sgxic240/LbfQkO/d5XqR/MLIZJsNSYJqMKlBA75sClEQ1gdMlaM3umymKNM3+/gMO
2qNPgmWbfqfbOfpTwGEi0/ZC0NVhHppBgf+l8KfPG7HUFaucZg1zbVI0YEXufkUd2WOPr4HLegHQ
g/pETvC6pIYeCCi//yj0MlqitN9YoYYhqfU2lqW/f3mmQivLcylhDADtrZjsffzqqob+D14nl1s+
dfyXqgEmPVHBOxx0HZNEYC/Zfif0esYPd/heI6dlFhZpOjJY149NexcksVm2IZ5YDAoacj/LL54w
EeUUdWNos26pPgSUNtsuIvPlK5t0Joxyl/0Poqw4qfhaZyn69ml+VlxC22R04vmj4KdlQ5jf5Esh
hK5dxaRYHen8xo5kvI/nG9eUJOO8iZqhNMYyZBOqflGawW+HBCkfXxEMuUnq4T+IIqbR1vr42cXy
hNronDO0MvDG62G0wYX/rsTYQ8XHWWKh3IDKMLQzJWkBAAAD2cN8ucwXioegnzpXApHU5lUFwFig
ZK985MdCC/Gx8YiM9vylQUSmygwFDGNsXYOffJfaUWRHX1014WTPaocuiQR5zhGPhzEZLi1waPJF
zS0HIY7duv80BC3WfbrtbwPBBJGWByK6gYgVd85GbGEQ1hW4rCmUI4kjJun2G1T7LmaoBbXlAIyi
hmiBM4OCJ5MntrB0WzfXfehAQB9OAn3lyv726y913W6AnEOsXy2D0E6zkS5xGtspv/jZfSJGXvTk
VotxUYYfay5rI3p8pCOJYcr+gNrSRslCO+kFtWkvkcrpXksaQ5UnXcVXVatwL2qJhudcLieYBpjs
1S69Yi0N5BfRMzcm6Sog7fiH3LuyMLNRWVSvX3lkRoV93yGnTCOH6OwgQKoP73iBIZaOQ0qVlFJq
c2lZYjb0jcv+AUruJ/7RG80fKoncMJDBKCAHOlO0viuShF5SUooKZuNmIil2YMPdFnCzLz7j61gT
9hP5CXaFg250lSWT8+QnTZokoV7Zi3rmYQN6zuJpn2wU88ZXY9oI9hLX/w0hWNyJjtqxQiJVDdIR
ziX3bdCHqM0Nve27ty4qiXg8tEodjFmpDYj+gBc4cs+IJkA1CbxfxXsYVfm6eV+abLhnaXfzGlgk
eac0Mzu7CoyqrOBpB+ne6hZdbeqrtOK1nYEvI+/qsj/wlR70dNNfei7o6eQoiMlqP1R2Pgh3A0yK
mraYFGKQKZkkPHivQQK+gIe2p1mz10mh80ah3cauP8z181jumsXWVeJAUnJfMXe4l9qrXlYNVk9/
XtRSBEj6uhanPTAQ1elazGgm54HZU1giLh6+6U9wtc34yJzyondldl67LmveXDsaYgLHHZmaDH9P
aO4nzRqzM8nCco9gSZshQ9pTAmClMcuAuPBVfV+K+t/lZBiEVUyaXu8kcOlA892EWml+ssizeSBU
5r4FpUm7OPTKYaBgmRl4wrxVMIC6cvXnG4OKpTJxaiuSwa2xqkBSKgaq6h53HXT7li6U20Z/OcR9
TWhGj/2D9OXsZ0UvcUU7GlQ0XqTXL0WAFfyoypiiX374Xw5jQaylrZtKMf9PV9DZ8ZmnhnIECLsj
dhmXfNr7pi4xCWKFjWS5QqhkEGPC91cB5lloZEaPJ1t4rpxtB1WgnsEjGAYGFuvwZyVpH8Dud5sb
amj9wD1EU7IHw2FKff8BxrYnoHT18RORi+5mG0y261IZCf3FC2D+qp9P+kC08Oa84UBFewVgiscX
neM5RBwZqJgr5PwqCIT53kdh3KC2h5a3xSNVneZE8T7GuHq2CLFtvUFWV4/Xyt0raKOyS27kP1VV
FW5oxWWL6ZOl94pplo2UzSUAtLfPFKb0KBy9bod7fyAESYwgZgbUf1+l+44Hth6IfCjW3//0NXMw
++DglqOqiNRQ16091vqy+kroobPaIinP/WaIq4Cau/T7XV7eNrshk7x0DMD0MpzJS6ltG/BIPp3l
QGCxc9jN2nIXumnnedFC5C668LCfyJlmWv9DHeunjyb/NX+aTo7pFubT6WSO0EpSVMcfMCdnw07O
e5Aab4t8CdVdW8eaLs6feJxZldai1DcHNmeb+gq9ok9PkK/sqDGLBWUyJPFu7BaH3YySSFcUAsyS
APWcitsQnGm403UD37KLnHRWbEXRfMy1EcPrxww7bdhiTbppNuqieDkJA98Vt0hq8j1xjN2VcyZ/
04oh8NtqDBl5GYxjiPADsyyPDZmdL7Sxci2ZJzKxQvs3+swBst1p6QHfqPjY4IsDQAl1r47tgXMV
8MNJWz8Y7U1zDgc1aWkHWYoN17VmOX/PkUyEK8Dz6RDPprXNj0f+dB/JcyvGqmGC+vS02KsYMr5K
0wi8Hf79dbRAp8aH9MFfZ4W/a5oi48Oedt+v+/Hf3hQ5a9AQTyJJIpsMqO25J+ZDqxnpW2AEjoRD
43PHHzQUGXvqVWKP6BZi5SaRTCSejlah/ix3UuLroQxGJAbDumJJV1hqTkfYr11udxr26ae58G+S
N3+XgbC9Ie7E8oWtq6fL0GW4HPSDnM0gNcgWJ5WQRk1K2YEK08ggTuLNwaGpAeObwLauKod0hcJa
Wf5rVb90WcF5TxCjUbSTHtsovNg2HVM05+EbSSEC5/PDg2H7bemIDR0bVjNgWYQEZXvlDU7jeSob
FlknqjOdvprQ4UdcEfg6zupMgmcQu5tOqAYOSG4Ek/8P3rV6289yQ3qJxZ8PsAXFGuWQT8th44Gl
kT+BEBBc/iSde2X5SCCPduvbh0SkuRKrKOEPr2K5al+CRO6AiQshqpGwn5ga0hEMSDxwJtLfKY5D
7XzPkOETwe3vwLAYYXK8cpRkgtiRk8inta5r1tQHZq0FNK7/dIpQW0jTgjYPRanZY4+h2FvNkIiN
yKzDEvVMeucrn5BAv8ldxMwDM87xkHUAMvfyn7fwm6XJ0kPZEPRgtQZFRX6iAW3eEPhyLqpELTih
W5GQDP8SlmzQDGe9sylWHR5mOMUY9b9eC66QIE2w/d2gZMl0hU1BAvE8kMXT0hrIotYdxIE38Qqx
BdUET3f6BKc5BblOqXwBV0nz/Lz3lQJXgdS10DIerbcRPGF9eyUP7ZtkloZuv6Hlmv7kJChD0UxJ
/Y3PfKUU+0ENvo9TTAY9K2nP+D8pJU4ALYihJf6oOskvt5FPuttAZ3VSOHHIMlrP9ziQ4h2JWuyM
ukem9JliZ50QevvqXXxYBeV/PxwDy9sswL52hZZI7kDbPqg0Nse4eOof8A4Vgl2SJRQLY/DZO+3z
gWgsrW0cJ+YbVGKbrPkIKvtiX9jQb8S2mmI2x3LCcdlg6/3j6wGM8KtlORund6ZJMYq+xNmNGY4N
PX2+Tpn+7NZK1M6fNUwU0QzrJryxkzSUb+Ffzm7BKgm44c7WDi9pseoxbyHhjJC7v/mj3Dye1qOi
wzBt8C6en4cGaXfEDdoAKFBWEAalZ86F5neoIWcHjdvTlJ85PZHPKM/aA9W9ayAB5QGe4MYm9mxY
AmBR3bSP22SxSPFpcT0lYv09w57/tNzbC2lGIuWkvUoZCwgleuRMHBIWKX/VVAw9tDx017dI9egD
Gn6YVJW008Ch5rmylH5jw8RR+b93QaL2kPFxv4AWxovQjvA0nAlyAJMabRCg+XASo3AEieJwFT/W
L9tjzuRZ124BWKkFognmh+KakKhccYYENSIipWs0yWowMbq0akiaWMY6GoSaqxpQEJNGc6hn/8U5
5foT7cTbWKtTlU0YtWxhKOZj65Ifr3aWYvQLvAl4MJLT0HKqifeT79mPg10riD3xbHJZ2GEhj2s7
Y4m+PKGRtMOEvm/lfzKsPlHCRnBQORUuJoQ3RjNas+PMoyF8KYaX/PQC26tqJeun651NAdeAtQt3
JHCaDnEg3uYjVJG4rGQYiF6DCHjUK/5Ol7u8iTFGahokSuPBdFLi7MfDhlQBFCGi0H3Bhz1sk/H6
Ypize746zx05HEarJTaiKXRJ9SrMgkFEu4lEF5wwEGtbMNPB/GrZstVGTTly8SXwVSd3qGy0Spwy
0bH1lN3QKswN4ei5s0HGp1DjDk1XVpZ8A4vl8QPJi5b8a+AhD37PE6hxQ5bincP48nHfyFDdBN6V
/CkIWmYPthl/i+Gm1pWiJyW9vWsUlwkXzVLrNS4JLC7NcWfdjuxTWrekDbzOfL/2tRSvTMWSZkiV
n0gjbU5xG9psjFStSykrjQA/vxTWd2ctXdqViHm/CwDOHXTqCsrEpsi59f48Hh60keN3oWGBdF5J
kWBiG49reqqqwuiZy0Ai6QuEmsNZrtuMXalu5JjAoFOP3Wun3Q6x5bAcB2tCSvJ9NEMN5USOnjid
BaEtHoA8zm0lBO087GhzYhPbE7ds4pJ8FG7VoLy++EM6NfwDCWinbRj+5+I+VJGGqyRSvOS/xmcC
e6zwv0OLHCDuksu8ZJ4bdNnY79uR4S8rNot5DN/FOlOd3THwaaVVq8Z6IdxMjuB0fYDm5PEKJ2TN
JpeIN2Psecm9vCwXrnUw+YHUBOYdebDIbn0uTOOhKzx+0BHs2eznoKbxUaPFrYirBgb4J7u8nkJF
BRMwYQWfK/tnE0jRsr39kgWIWjgP3b8RT/LBAqi2T7CkOdjcTKkcqCnXqWFU8T8cvtx8XZaI8Efg
hU2kus1XSs0bAn19lC0Naspz0ImD9YPG0wVWHooDlJFjYCHrPADrmnT3nFKo+PtdSOJBYr2NagOO
s/mz1Kwjh1meMsC8iJe2DC4hp8p3tN0HYXoUZ8GpCMTlvr4lONZn5cQk45SeJX62xB7vTI1MqIyY
X+EcXIxaYg9jFeYYl42hrcJbRtSl3t6xsXVc1sY2b/X93su9uQ4ZBJJ+8zyWt8X7Tes5x7zVG0ZF
Vig/GwfhBnAw/xoLU4cq5h9Kq+NgdWh/avPMbrXQ5oMXiPVXvtcbiecyzHb0DObnfAh6pDBaxf1N
9GEpp+uflttPkUYtgAyjvxxlPXmeQZA8BDbVHP8p6vRnSw1+xrmZ7Sn0A/L5piut9taxDOqEdoL7
VRC3aTizTKXUemoZ8Pw16h1G6g6UY0+1wnBWSNCzB6C3+DjW2WeGM5SNIPPZcUl6cp5P3cepxu5c
7BJR6MHk37vtibyO0UEm10jM7Ftih3hvaZzpcZhaiZ7FrOYa/scFd28/s5opVp2mp5f3WUARVlsV
9kwX/4nSU5IazlIU32fAU7cZzQzBpQMwulGEuV92cso5n6iVbSoXwNXdY2pctDdOvH2byW60uLUc
eLyX3LtiKmzFw43A0qTGMPqWRgnwribuJ77dwJcmDlxePQBJoMCOEArYrdQEGlX/4zIFWF5eCafa
Th+0MsBv5GqY9myJPNEnQWhjfQW3nr3xQjKS1P9ZFoGF5uQJHN+Ae3OfNUgGCKlyg9QKqt4eK66p
zXSOF36/gGTIPadOlDuWA4djHaEk8Y13BX5cA2kSi5VVm0PndASPtB8n+AFTngfTbX1Mn9+6GZt5
AC7YNLeq9lS3Jpneu1OmVvNDMZaTWF/n2+sp+LETnVkCp/Jt2vR6TYoj4KQP0tAJfCTtibAi+xFc
9eOpXRVXx3Ha1C3q0jYEIMrFv419REDA8SuL3XZyOxEIuR3Pxi20ok8Ttys/ktSePL9H+9Lud9p7
8mJegFJwNG8tO9FS6jWRCjzSqpeQjbguv7rHw2ebsrXXPeXBH2AW7F5E3VQ+tL+BeV90FEHp8ghG
pGax1WVQWnzkls629Eqvg7N3Hcc8kFpPZlvbXBep/yqnGXLOQ/2005bEfH6t4CHYrzhbT7ZIo58A
6h3SxxYI5bjL67S8QNJhatj7pVMPlApPWxuV63ofwicBOcMWsKHV8oFPICk/FA0IoWJ+ZJj+PyUk
+Ay0s/KxUUdtrYVxS0lcQx2yTYgr5o4pLQv8v0twrAA3/7uo7hHRm1foLlliEX98k8P7r4rIIJrs
Znh6OhIPh2bwDBobPpb+ZPyqLzvh+2APz3oeQA1dJAZvCiMssYHgMzuQ97x3JUjMR2SsYW9MpmsJ
unpwce49Yx0dLIQWeTmW7jCOqDv0uUeFu85cLwesVtG46LUzYHbbKQ7ksaS9QXZ3qXUlwDG5Ycsd
PDK2nxyuIvX/BnPdvw30k8Hhbgdk7vdMTQbAJJv/tlY95RWnBOa+WwMZdQgGtX+g49fi63mwBScL
hOfd3Sj1oaJpK+/s0c5e6l4Efox4v1GgQePJ9Bm+gl0si/OFCNsoAxY37fX/oVR2TixtcyQPkiKL
jvPAyNsxmdA9A+SX4CabQl/IW9B/f8bZEkxaAwoCAMv+IdjRHKyYTxgqHGp+OTtYbEkv+Zmqfs8P
GBtnFzlw+PDFh2PMSeO2lWZMmOpjxP3akp2Ytuh4+1C5+Vmg6UswOsCyuGTTIZ/YZua18voyzk2N
CxhkV52lQ0PFoRSRTCqEQKW4j2KRrPtHYEvR+ylnJX//NYtbouowoHMJ2jSCgNii2U04ziMKkqHr
ZdgNF6TOTdpUd1c+tglM363etcOYdCIr/JUW547u5cv4/zMv9yIPOZ1zp9kU+EOt9uPe1UhFSpqx
Gdu20RyG14nMO5R5E8mpiP0pYK3bdjsDbddOcagA5YZPJ/aj5gttoo54QHsBA+AqMZEWu5Ap+xsA
HystV8sjT7l6dVfxn8qJtI2FmvC0jsT3Vy3ejGQgDuV2cqupI3Zgn8d4dGhE/vIAU5LtTILXFgZR
AN5uN1SkNMuT2E9rpa/2NKtAWo+rxkpvbGOZ8S2UUMQbeWo1JmtHMwhFIqbdkrGFpgIzlAA7tDQ9
o04ukgl6QykhYnFHTGWSgQGp5HqbhGbTp3Jb9fykyH7RjIdvAW3SwAx/FNocUMpeeFMsHJ1U6//h
77gJ9DSAxppV0NllvuK9TCrugFFO3NnZWGMRZEuXasb16PL5gRBn68Hla9rIttsUcsEErdFBjrnW
LaFuQTWg7tK7Dg37gOXPLNaKrSYalLXNr/LBKAR1oAwA5Q18w+yrUjKGLYemLh+Vdr8JcurjUMDF
IaTr1uVbIMg1XvM8FG3jGUAJT4BTaEn4+bF2YO2uQ7D7jLAgEoGioYTYlAbYIWhf4zk6VldLK/3H
yFD/DABgVJwsKFSGtUXQEEFpDYuefnMAPg38edJEVeD+e6Ra7/dJRVM2v/hO/L7JuUQfcRPf7CD5
U5Vi5lcWmN5y0wHwVRfASEUp/1kkGI8lxgnZSDJC/ntx3mUr9/FZWjjjTPZgH25oDWhOTsXt7zUQ
T3yLGvAyrbDtTfZgy9EGNFS7UlUfRhN6tJY+ZfgvTTyxoZFvfv2VTJowhZuDvtiZDQP6aWRaHxjF
2zb9t47WJm3Gl7BPCi6yZniLp7JnsdDoiaX5ZrAdzAgGGNEUw2sEiFzYd3ajKZGJhMk3xQnNzz1H
O9CJw45toKUxU/83xJz6odVNZUBAFX9TaCgOgpEHpaGu508HE/WOf7W1yfBcTXbirN/WpqDl93oQ
iabYAMsGXShRwaWVuDFNRDF44MSeK2oDO4Qb50yeuS9xd6Hzm4T0wuruxbVFjBIzDalU3R7XC2g+
wQmRWasvKWUc2JMa/lv/r2yipElm3NvE4tMpLqXH415ewLluYLZnMCmPEKbru6ffxLHpnuK6KvMA
WvOKPsinJcJx051FANKGan77+CPhzM8JyjtEnkSkp+Ax8A/D0hQ2Gq+aW0qADlyqxgtmhHwpQMqq
/Q02SXUnEiq2RqLTLoHeRRrXGcVo9JfDhPeBrLZn/6WQinYFTWKx5ESUB3SLSVO6AmdKjcvSCnvH
VG0AaBTEz2L2vwsDl/ySDDNxKN3do936ZcXOy7aotdWhAIIzZSikhj9reSpg4cN+8HjpgUafHhm7
YR/vtqv1WDpDJESJqVdoUu0mONw+xGeVtCBJPMQxUP9APw7oZKVS+8O0eKvkKm/06nXM2lXUT9Q+
4JRMvWCnVWGLkGTJrdU9ufw0/1+FruiClAZvuvEKWafqmTyje9WAZ0TrpoQ5s7JvWNRWUu4eQnlo
+UV/4vnXxCIXWeEyq1vx4nktR1zCYlziV+DzC4U1QhkeT/qbZR4xwSMCFymZ8dwjqBOYdm2d6gIl
98iUI2B6BZ/eCibdwtBFG8UtEic0wlOI8wQtazoqYrGGC7NtVIJGFXtQ2j6h45+7sLtsTAwbyd2O
llc05K7uBaw9MMvFg7AfhLnmRMD0nfiO4ugBg2v04yg+P2rnvx7PXRb/G59qX33hgUXvUP4NqQD7
m9+UNFqMfBGd4W8IrNQqSyGAtdUKr/0ha4BHMbhTjLZJuO9tY225rVe8Y2nvmZEpIExW6RPi4b4w
wBTjtKHWrtsl0KcHj5GbZpPXBWjsRKjox/GTQPiLLHB9GQS6JtaP/yDUJbO/7MRqKN8R3ENeUpod
w+hzv9ZVXqxLYtHeMZOaN9ztC6tzW9HKJ0T7yYwQUd6LbSe4C4/GhT1x06UsGmurJJzVtEr2CxLf
9Zw7Yj7WhCArrSG1Fgjk5/yBVXw2B9+Q25L4Hayh/FgUSgv/aCW59oZcVgshy4fg8p7Laz73tc47
Oyslk6DgMXJwqq3U0lTNCHKvRB6NieF+bs2hJZtmaeuQCEIF+AP6djOLG7Netylo2t4W7pYAtnDp
dFPrM0IZdbGEvzm8jWPZOLUX8h3ZMZIVWgdJZye3lJrls0arLk0P2md+1xHdra9xHOYJXbrVhSRB
0NlDy4bxOWagIbQqvAWxZLuEzh5THCU0XjFFLTsfYfSNPZENRtaEYL3psMOtO2EJKSRpl2JYVklf
eWmbpl9ExDakQwh82mnziina1JyoetOh788qMkSM2U1Ign71vVoK02vcB3BATn08LBPfO3yMoAfz
fN42qFmUwhg8vlskpQcJoFCf3TZougbYBEd9fIYDJtIXfr09PkUmwDOMxj2nYP7hkwXuiFo33DiW
/gKVnF4EZD+ItipHw1BQZeoIQ5wKiWxUli/LTIV4TqGexrHijC74UMN2BAv4VJaRcuTZ/c5Zlhxy
OPBf4unn0QI5/qGLrnoUWcXIEoh3ygjg5beDYMXj9w3j0nPY0KTCe4ltrX+KHFcEd1ZMh81lRcSf
JIX9akDE81zlqbZuURDobe6CqC0ZCsgX8KstRTMqx38f1OrEB8iLXdyso4taMZ4AWnbnZjH1irZr
kTl9rIqOc9lIGASyCq9P8mGcOe2AuLaiMi9MWOD1SLpKDFV8i1ZWV3b56yv0cwXCHKbRabWEXiqE
hXpF2gwjS27AUK97xFfZOaU6imjU2Oq6kEdat2bnJ/dp/t6QNLtwjmw1+v5GP7bnZGqHrUeH5Uzi
j8FS6bB/qieTsF1F5pTWjHiXYIVSvCuxI4CMQ4e5Xs0g4LwTC/YEZaqfXD+fl02d8ERcaJSVvAgw
RuRwArzetn6hn186J/0eJ13QfFBUvSb+njP7h2JiRmEY6gCmY3K7PtO5bi/3koEhezEufYU5EqTl
gsS3cFLbLtyacnFgKAY6Ykt8ZjR7qjDPxwGP/CA6bN/K5UAIRLGKIs0hnxBc+Ln6f7FJxFT4yhNL
eI0FQLQQym91iKTBjeSpFTBn4w6E1L/l42YtfUUKjdqZkMoqJo/s7Knl9IQxHBxuuBsPyqf/FPuj
5nQWfktLMGOelCwpcPs5pbpnhMaPmovI17bgD+8sJcw/C+zgm+FuiJ/E7XiSIQl6frSoFJWhkeMo
Dnj2eIHnOudI15kyWrGL6v6lHtmSl2Zlz6W3XYVtLxLIEbArH/9yWjlWymZXklIsKC5OsocNy5Lh
ALBG9GTK/Idi3gTdbr4kILUjF0xn5+vYIpUeGVPI7hZOWf9LDK2XG0mRDC2buvx5FxShq/qTskqW
IgSTs9u9P21/QBGeRDd//KGcT4vLH9hHj2Y+ueX+R2wr90o4TsfD3mCBHvLWqqj3U0bly9T+aBGt
R2EeeDfmcF4GYXnPp++9OJ+2gj8j4I/94EqrxIYms1tF3epPRIsdC98AnkEI6S5FC+ovWUq4RkVj
kKOBVINJfxUzJfKwHr/kxmIMIR2fgFsEVnuEVyt09+tRAeYG6ThW22admeAPBME4gY5sdYr7uh7V
4FjclmngbaQnoAGkyqD7ddYtLOGPI+K4dtaHRyKRwO5N+awuS0HuVyioKKi8/G+Mq2mY26cwlDtJ
tlzm+0eGU3h+B0JohmlEHtgFd/La4X11pySWQHQszs9GWYjwdHs8lqaenxEWHpkje5BvFqwwkvB5
kD56qJ2OZhtIshyoa8On7pz46wW/duTIDip7JIDIoXhvoT9dSOpKbVADHvIfc1mOcmkwP8Lyfcom
yc+xQMQAEGjLIg8xI3bmETX72wLX0nQN9EnQk/r/u8RRLXOe+zwG8YQeTsi1fYO+oT+wwxXfX7Z1
/apFYZkKAumBdwSD4R3Ng2LI/TSalTAvzRPTeQxbJ5DtDcY9cHgAcUWz2Flp0FENX1arZ3TTmb6B
RgKTA+kWcZcTbEG5O0gv6xcXVhV49DSQbCEUQHHoErXI8tdtyGkMv210qagvF17D6BZK0bA9sAnE
7isYHqVxwK0NweJhbHxqb/KoldV7oDlLV/hVVZuQk8megRuhUvsoD0RTaHbhGPJrJWd99msdF5N8
sKsqVmwnrxejn71pxLSlU4udaE6gvCcEXgQ6uAcrVt+Zg6Lc+vvH2laacQiRTtm1FXl2QaWU00O+
8hTHiwvE5m8jChNUxLoprKL3ZN6skuhskM46ePh/ZNKg8JsjcA/2WIcU9+D5mSkMxWLSREbe5fAC
rLvEMHG/jCEeGvk3suUCg7RZE8DtI2UmJHdnj+/4a90kmARZa430YfL6sOOoCg4Y2AIhS8k+BA/N
21BYH279gSDiyAU1DkJEkVegLe3ZZlZxoAAVd6UG+ZdoVOKlnvyWs15WCStOqjjKcwtTsCIsBsvs
pOuGHDqX9To04WAGC79CaBAsDT6lQ8hQLZkV3ZVyfoOEgLroroPjJOrrL2fH+cuiWjcBo707kFhQ
UrOFLcgHmoP0XDbsRAbFll37UUB9AFjbsf2N2WNuGmGuwIVNQ6BGF9Wctd0PhdqjKXm5PtfSLZzf
Qgskolzv4Tfxbh9uv2I0gyXdZQCQ8HxqcV3lu8lxYpMFk2fuK5KHm7sdhtSX949jkdmFJ1rxe1fE
i3aI/fl5pm+IZXZMZjtbfddz8g0AzDLwsePD8r68JVEaJmK287bfvRQGUOC3WDl/wl6phzC+AolY
MoaHbIBqmuz/fgWkUggYe7GmXPnL5gjzOTPl51eUIBa4LURYgVvZeG8JIH2on1vo4uDCySB1GI1M
ThN/6LijrxCXjDN00yKj9KRFs1wAiRaYys+7m5SSHt+ftNHePBM/3DndVk85CDHkahGIr6kG58ac
Nd8gMqAspbA3ftMHp5N4XdWYhK4YI0YEGqEqQk+0ywR164B/DTbnBzSr/ltDK6y7ixCNcufQJUDV
LSjR0heP/+QRe9nC0S0QqxvgrEsehHdkLgO3BTW3jK1JNzRTzgGYTmgrm0tsT2TVW1p2XiPlSvxL
z779RAkD5MA7zbzMtaHDTlloxZavYL5kAfOIu4R7AA5eaiyrOqGDzrdpmRIqsv5Mi2njfP8IQFc5
amhm+43aFKv5r0BBS9FLI0jEfZ0gFuXnxc7Btkn0Wu8G/jt4Dz9JEEFQPU0ix7cTwPzrpMCPw/jT
L7id0bIsVC5zY/rAP5DvoRSk8XxwvuWxLQzGpCMPzT3fdxAHbxQhMA/2TOOx+NdNeS27RwjmRLix
cyCMHr8BXBFVepsYb9ltWRBN9c8dfCubxuCdpzKVs+/mXEgYF4vLLlm1hL5+K9Cv+Dih1pZPq48f
nAK7P/U8glhJmjbvlVv2Z5xF68JwFr27Uel1KXaVCkipLPZ/WsXjzJYpMEzJNiVFMbLgmwh1ojmI
r+LK1DXo7hgLzVNT37bx0LqDfl8t5N17NbNqAZ85hfWMoK7t2e7q69LvH6nqTWr3z+1gMKE43MqP
hqJ9RFrKRI6lCUUyGGD307YVrkcweoQbsAau/oKIMagQz9uBr4rQ0RpXCKSzjm/aKKvFx5zwWaW1
632GDXw3aMuB3sS+UC91NKlehUELdnmItL0V2slOvnTXTqVbap1byI5Twg1I99r2SIDy6h9iVxdW
fzSsTRzQq8y4kEEhf5StWNJ2uYuoucRm8DbQP67094b2X9CzpC8SVu8w8EN0BSBfLBxigaSDqJ5u
foX4M3imZhEd/aoQK07ZMcQqEMpJVzPtAlNlY+470Yo5i+pl5Pfo1TZgE/yjv7xfHIAsREUl7fpN
kbBCcP4cr5O5E7TD8ZuXQtilbFJ4PHTYJ9qGKNwBVugK2oCgXQLx5l1uHMw7MvQsn7wCg2Bjn1CY
TWWfV1fzxT2Alt6a1RQ9zvB9CYfVBAVAUmlPuswR/Aalmd3wsC9jK5EvQ5aynxrgwULJIw1xF1o3
VPxc8YjhvM2/h0Sri8bZETF3yrF855l8hHK11arONZi0PakG7BH1v1gA+UD8nnTHPehHUoP/Vj9H
qSSoPtuawFC6XWb/13wB493At1g6QwqPFPg3bAGReqCRdZBY9b5XfzuWL83OV0savlCYSRI+f41M
lonzjlas+hNaGafzpwNVhknm7OWZA3xNt1tS51OyWaecTanGTtHqnZge2lhMbKc31fnxcPwTstfT
a1QBYbTI4/p7cgKaB4ni/Ba36Tc/VF420XC2u8xWcRf+eFOfpvV914UWnKGddJn/lrNwYrOX1V0d
WtSyRJ4lo5z/VUWaFbU5M96DWJXNYbCMk8SEtftK0CUXgtwt8AGrbPBHK95Lamw+pdbwxgVcr4Nd
ZNUdUSsmTGWHVHWtsu07YxsRzE9J7GCEAd17EX1+Sc2gJdBK+285nosR14j5nfR8Y+++fTaJj+qb
z0iyZ6Q/7eQWwpt7BDy5s9a1fOuaK23ni06MaaYPzbWXvVitQGlvBdn2Y2joBSjpnZBwg2h5HpZt
WIXec9+Sd4oKGSKHyGSdovu53r4STjC/fMUV2awkYgdlQXtechL4+Eqh6BSX04462M8OMR9STSpW
48pYxP/IvumG0rL/amN2plGP+AAmMb1/EgIysrg2GF3YQ68I6Cs8apuumehL6YYvJfSyEUtRdRUb
t5VIxfa7t4Wk6vIArVNdQ3U/TPwxW/4nfIiSoM4EblQc2gyvFxC+NdKBZXHBgqvjKOAO1OSgnREt
HA5SeKmXlCBZenylhIZV10LcjKdNuY6E0cLiH1OhvGMGXnB9utx8JkdQydrnhDiLpFrZY0Qcx6gI
kqoYCgmOZP2dX/HGGtrZtkw7NwZDApo0vOh61gDnk5N1TVN5WdGWDaj7OsJEyIbII2t1eX5MVoVJ
WzxeNyu2RKkwrNoWBQuUOoLJVCZq7Rz6sOmHQGL51qyHFKN0om9p8vgW6R3cloOhNyzK79OI1Pb/
LhfBrwT6x3EMV/WakwqgTnE3tEUr0QhDNVWNB+S4DPG3hCD4INKl0teyVMO66/ptB9bjslZHNzCU
Sdpj+Oo79LfSjCbHMP4qE6uc91Cll83mFNGkCQVz9uCvUE9XK2oKo4jMAjxkoVhfY5u8FZ0BvEfb
FziynsM0m06vd+fc5GnJQkaFl1PS5mk7iQ3J1LsksA+vcqsCPuPXtvm7iH1lU3jc7jKKrDUqJEz/
/GFEhrYXLiUTgVrnklHPaY3dijW8bpGK5K+ZBeHM/qNym9pggjgkLAdzIvBoCgjdhuLxJY7Itt8W
VgfrrM0zFpT0clMK1hmNzO8ZjIVxb5OTreB8gXTQjSzrZ1THGf/zzbI6cxssIvhVPfOF0rYM88Ip
9mGiHrSCnrzS1NhxBTtQ3iGZXu4uJ16uiDiSSS9YFLYWwgReQdhK+dccwBsKk2tBgBTt+4+8qypV
BuzDIxyRtLhqKc8giAweLkV/xRpDvFoVo1SPAus7nt7G++np6s9obY8BC/VaI8CIpCuv73xtAxKj
ScNOTpbghPoV8dxT/7gyyLn93VxrVjWm6Wyl1Ik4RWrR6PnDpQNEtUy9jU0opdNDmygu8wBrDTU1
+ndphmE5BfiCxhyCC4yo3J/+aQK11/ChiOR4KpPHOJmVdlyw8Ur3Z1mrfEq+tAxQd7C0CPEggQTz
ZkzhPyNAuh4fd/0YPFp9efwfbL6tHGYWgclRZgw+JIWv6uLVPZLbglViRsHgzdtk/vS2M3mvPHiE
aRXsapmxxYGeWYTIQwvniq49fYYPeO67MkJC4xE1SxC2+6g05QrNUUeoIKCpa6RqcmFfKLmGfpwl
ndZq376fSLsGcun0xtnb59pyBiGOfCoWyh+xgemIwFO7rHSri/d6N3VetOeOkjTZcuqq37uAyw9I
Zoca4qH55i4MEMA2lfF62hkN86CjoLn5A8o1oaAyg3ScasnHWqkYP6tjnZhY+veI+rfkKVItnCdU
p42/bP0Vey6de3fczCOXNXMG7spTgf6MHQH6ZtwYGTGRE0cioFAGgfOux/VS2Pgnx3bsUJ455ipy
v4QfzGJtYA5JnD4M7nwLophDkIDBX/KhIdJqOyDI3ha84p6niQalIMxmLXF+h94+J96sOaFnILZY
KEmbzk9QM2oVrEgrichaxYsZVy6NC8YBpqCLrilRWKfWnMsG8qCVhPhijAoDotCVW/AVeUiynu8x
JEG07DZzmNkOII3YcHiU5sQEn7+nZHjdO0SWESidDV11cR86nkilKoHvLuLBpMCsOcZH8sWLwdoq
puFtO9c+iGgDINoN7jhLcJ7zQh3gqLdksNcADaqzywnBvY9wwXSJ1MX42dgvVW8Yvey23yKzZqiV
Ut79W9CxVBk6OrBqkD7kfXz6UnMMiCT2VxCjTzbhYVuzfNT0GuoC+1uqtVMn7ssH0r3L60bXNRgx
WEvplcQq6O9faWRSGq0GV9+NcD4eBc+AbnMd+SyIsjjgNDOkZlfRGKzVTs+Me8SySVNn3HLIzWeV
5s45e4tZtAOwbQSTyxbLgYxflKwKiM/hfKIRdR9IJEfIK0R8Oa8d5csvBoN1+Mw893LBK8iL+xEC
o5U0IPrUcZI3PFc2LStj17ibejTKhgTvabgWONbYkct4ar7ZiKUp7P9M56BEtvTF01lvR3LtPRvw
lT6gT++by0wR4JWO4cBYHhg7Q6Hj9f/cp+TVQFiG/ymP8GlaI07xmTtqZ1VFQQF0bmxn+3dtqYtx
tjD9RzLky3j5c3hxWBSwjVu/D/uPEjfyN6l73cxoVRkN3OdZ8O5DSG5HuZAVNKLRsB2bzCGXUHbm
Lja98ni951VNu6uLRvsP2KyBgBtYS6UqypgRQNKiuh/bX0yMgb+Qx1NtNtuKuJ5tRUKMrFuT0FtV
T814GXLJbjeUk93uDI1YK1UioC0++DYk1tUM6lQzuxRErTlS5OhiB6IWB1tTC6XqNVOIUJKyjElm
KVOA3o4DbX8WNtq+81XrHO0XbijRY8YwhBka3cPpafdWj0s9d10ylYphmVv74jJu6AB/P7W76KFq
hTL9HFNWiFZPUTlyDATZ6Kp8i9WpYQt/uu6YhKBdFva4SJrvhslBHuBJbHQ1RiscKD53wTJ4CYFf
uIxwB2O6wFwWEZ8ZpdBXzjb6ZpXS8ZYd7MPnmugTI1pnpJdvWtfTMKH5gxYB+PVVBt33ekZ1EpOR
8hzULkkNS+XiOlkfN30rvoEDRFhm+0hiVxBLyXC85+lVgYVcEUnChnjrD95gq9sXO11aBntWy+Ul
4iCh/ZPXRz22+9eOPEe3eTcROw3/zUsDZ60254gpOwjCH7i0Zr2mpkhkTT0OdhTo/eGQ9N75j2LF
9AwkVAs4aP9JmIulES2M9viSyJPH12VpUVRKGxQDms6+FudgBoAe5LKRDJL1haCORYbWEKEGZXuo
b2JA5gQAKSSJPu3NjQyEu3szsLgNtoQaUoKMg+oS/hvD1BhtQJQjrV/0OIKL7rpJ3pjL8RclKyfm
bRLGn2O6B8o0LjsCrcMfRbwKbB4yiiyHlaiCDO7PnpjB6vMoXRF0T/CMWlkfts2ZUL8a6b22RkRR
/aeI1IebhigFWHbkzbhqE0Ejv41NzWAVqekrliBLK5SBPadsWPzLqx9TMtmyWhEcULY+D77mXZXj
oCbkq/iQILnjPTv2kyJNhm0bUAiqK0DQ2l/wsfD7o7PVneLlt3AR4jUjODh65rhd2zQE6r0pj6TP
OI/UTCDwd72fiykXEoT678ggjBCm3xmsEObOku6gPNnX4CjAdgJAE1jEQ8xjX56a+FM+6ekX2XqB
oDiyPwH1QK9UU0TCMl/rxBjnOiEeUH867SL658CjjbWcpDJxYGT5P97jDfMPJr1wKqYY/aFB75K9
cSq54N1TRPGqtR2K/JsTY+mgE1uSHWble1Za59YHItaxx8LKTc4hDMsD7JA6TvYUKoIeCqFdiHmj
RQhSitoB/etObBW19/0JmI7lZLdcrnpXmXwLlvsyg6He0jOvrFzbLBV0maBKcLwfG7LvJlYIZAAf
4moQXPjejGyzjVKtsjK9CPZO7Y3Ew7MbzNNSWiYX5uDtJBcF4QurDZ+ASP5ZXu0/Zx0S/X+Sdq6r
Sns8qR9G5I2uRA64/8lsQt0wkxPRlwAvWIvkK0YoNn8DCwPGddQlEe6z9LulqPA0Ypa5Tch0zoxf
vpH8S4JluIhci0pq4EkUb0blimFna8I5ML/RsY0SvFbFOG/ThHreYierXnN3DcO1s7mQCrC/lIcp
UchUpcvTgFwk5V754sSygCyxp9ekUE4pkDqlBQOeyNMpjse3mwNPM6QzjX24wjilswWJJrZJuOed
L1eNxZah/W31Yppv9ZBDQhk98GZzhCWriH7b1IC0DH6osgjPoFfFu5SKYq8dNlOhV6XKr76NQOYj
PlWAJgPjF8yE9Bzuu/7WLf+qhCirU+gir9oLQtI9lF7naUud67G0Rt2+tfAkCxbhNSEAfATyCM44
U6E9j91CCeQ+fLXe07i2JrYESXHWccKbds80kod7tDKaAjpT4trThWzuuOQApAYxIZ3zx0GGINP/
WpiPkflwWaH9oM08aaFst61xP82v4xeVh01ZEho1kZmrehsgbgQARCddpdbpu9LlC8SPY0mKG7Gs
WM7TBCVo/nhQB2mBEIqJiAMsXsCR0QVDZycD4if1nZ7UAxgdvxlUd0VuuiudxC2Oy0bi3kka5bws
pvBHRMYqXO8fhib/8khyZL4ztkwUoXBEVevOqN8FlBG4OQ5FitRxd4TF/6TGnP4n2pN24V9Pbmi8
C7g93B30El4B3/z3ZKoKsZhYeTooUyQoeFVhcj+E7muTaUSw8WtnYQk8RU0y1uGBK3RO2SeYYAsN
K2j2gwPftOFieU8G6wdbBXe4/sDnmeO5i4+3cLm7+TcfVNaZFNHUvWueX33Klk9ecZk2h4uaiA4T
AqW/rkTV18JZpOMfy7ddqY0i+AQwGnAIh99vIiCXtIfxX61DQoIDh9BQ1D3nLB2qBKiuxpo6TSdR
ta6yUdip/Za0JYbfb4iEqNeBN3ONQeRMQAfT9UbZLwWkXfFh1M4vS4DtqgPd5aQ9llXCLXegnl/n
GW/C7DSwl84u+CbpWN6eJOBdpEASZtUsMT8OpZVpzRqjFrT0RmfaEfGnBN95WwWeKwfYdzp9DOnG
0twfoDUuecREnCpr27fg2m7zM7WOQybpL9Cvis5yLCXbzHDZLRnqjWkp8d+f7OEueQUijvavCWwg
FQHhyqKs7h2qiKByTVy+BP4h+4i3+GUde6nSMkS4HDrSVir7vv89TMMZ7qswsJLXn6Gl87zl+yJ0
bOPMrIqxiS5pIi5hqv1pi2BCxT8vzMLXvshfLcXk5VDLpyFh99XBF01iSvizZSA+G7fZC+DzAq5J
5L2X7Nl8sNBL6Oo777JaAHMObViZkrzSMP2HgNhb/q6c56BZ+2dnG84SJvEHBh1zZq7zWKRnc0fX
dpbMFF8uFBAxWEvW46jqus3wdkjVi2r/V5p7PEMWijpr27kYtj9JfjHTp5YW1iV6Y2J49x96j9ww
tSKzGE1q0ZIlWpt7AivYR+LGHagF2/WbKvDvx/fxXeVBrM5a53T5h+U2nxg9s4z+uGJ2t1uh+fmG
T6BcuCl48jmwwxa1JEI7S861Ve+2x+VNqon0R4i7E9wLCOEcYg022RLIIM9Td/xsBOrj30G5LreJ
fyWbexBmL4b0m3cWaaSHI3LH0A1duIhS76noMwrTFmqL/ogHXMLH/ZR1k8BVg3AFGLkBoNxNjg6a
0JZLKaSRkyE/dKRYoqZM5ZC1YUoBrTx5nyThccJIp9K4jTqSQVUmTLXb9K8jDquXRTJ495Ft/PYP
OT0erbnE0MTPvGGqRqAQqaH7i3/YCU24eJybwYDXvz4F9TihyfHi1tXZcZD3Bs2uEzIxm6sDxs82
TV/tFPoqXIkuCoh0/ExSgKKSIwl0YMsr3Z0AnNvxlixo8+x4k+MarTmtTBN5uHkvarYKT0xEip64
CKY6eRAKp3viarC7Tk32J4QEIz0b7aDfnscCHt7xUMB6Pxdtyx+J8cehgSonAEUUc0XEBPUk6lWQ
yc4bpl90a1nBtjgZpMSOjbfUOXGYC9uDsVZkqAJe78EKanFccUPQtRxw8IsORqQLLElEVarQERg9
BPvkZLp3fWoiL2l98JrJOl/EhPz9cjP3Y75ePfzJUr7tQTARDKs/ZWBKDLPC66UlsCvmHJSGw3Ms
TtOzSlxeHLAXlRKgeX06wvC9FD0LRZy0klBbF/94kDgc136UfOhq++yzTKNfLjuzxLqv6p0fZgqz
W/rag9BHNWQmwPcYVpPRALkrLG4V32azGMGKstB8mSeqOT+zgDmGbwkdWTd+B96PNKu5K2LLw7R2
60AXBzEc245rNpovXM4aQTBd69S7meI6TMAUJ3HJcuGHEYkBg655JXktJJR9TdyXEvFXE7pINdYK
u+j4eMdwoFHa5+ziSCDrf4hUxGi+L3s9OpTG1+Gc2Wnk+oC9wLEO+1ZEhVdH8BOxHsi55jVh14Al
2xjcS3lq3OuOtvEx1CDlosSzGw2xxCZKvaieIWPZnV2V9bU0JKNzLR1DxV9xyyMBRZ0J4oiGzP3g
TX+Z/UAzXJMqSo4EgZO8FnyoGB/ZYWx+672wC/cSNt/m11GiK5ACPrqAtQW/ovcWoiFqD8FIRCBo
L7IR7Z7FhEy9nR4SSfe6TyUAyuP+jtbdx4VijzVYHza5GSgEZWl2aFZGMX1hXubZNxR5i+AOYZxm
wwGPKRXZUp3E+oyb8Iz1YKwYvL4vZVVO0pvtYScoggYlcjEdt+jMVK6S7rqNhIevo1RQtSoINsQs
ugNm9wPkaU8wIuGZ8vJMhJ/lGidOL6xp9elkz3qmWJ5UGuA8yIU64FF0YRhVmUrxsDBnTaCmvmqm
QdAVkk8Og1ofv2ywB2MVQkBceYuUEYjWntIvIkeYfOrJKfZduIsbAbYKVbG0cfY2fM5d+qPVLaCL
n7gPpKDvvJRy73pL6xmFGpHbb3KHTqkQ5hY0sE1GzNXUqlqa0BesVC04S/ejGpWXXZFPur50HIPI
MCRlYzaeFoFqyU4+gd0IbRy5DeBSPed65pPMsJ75QZFSg+pbFbsuSPlk96XlCsE1Lh83V2XNR0RF
Prtm2YZUYBMnPpbEALEjb8f3Ol96T2AhU4LcYRtM37Y1Xuk8pbzHch+qKUtMD8amo5nYjJCw4Ltw
abMcDJ9pHK+1SiM/iI3kgzHfQ30Pxue1sL5VbR0hGmn4NvXVrgeOYYmrzHlwDFSOSj/ZDrdHiuOP
/kX5gNIRrYY9FY+lZTESC+XkkUdZDkaKLHArK4owfDT6GPlGUkTQMLNKgkOOeco5mBaFL5RkU3LI
FnXszmUfhECSQyFzxeSzQl5+Xod0LyANR5/huDP2i4iJBAUcVsjipSMDscjlgf9yW/EpEVB79rvX
5T45PMdO/0NIswQ6Om/L/AClfNZ8tBkmRry1g6HEL1UgZxoGYajqbcZvxGS89EXGO/LVZ6VNjYHQ
B8yNVCser+NNOABc74H27TjfxgnYuDeJN/uc8Lhqq5sD6W+1eYAb9leFT2+LrfXU/8bIb59c1epa
gv/g4W7GmnacSCeodebl6E9NvNXoL7MnUg0vdx8jSEMYTxGGalrmHuCjuoSWmBrH2myTXJJslWdu
OrjGi7d1f98WOw5BEB45rhFEj9Xq+dhwA0Uif2mEd+RD/hdxyXMXewtzSIrd3YQKjl+/zjZ7I3mG
DHGgsgAKM7jvivZm8Ma8d+7EzMLHYoS4tjXTL+AQzMH9uGU+GJVuUkPysVfP7wdHSsBZrEYkKcG8
Iibw0Jy2CWp05SpMx4DyGgFoDF7ZhSN7VI/Sabasc4vcM5itHcKoTijDtU82ePT7O/6Hg5b3vWtR
/8cHrCnqLYCY3gk7dwwg9dlf4SNuv+AMPu5Rv5vgOoa09a/cFAVQlf1QasOmcFdgeAnzm9gRq2E4
6Y+mlGW/GD851beXDDWwivIpgYZgeFVuPJ6hFOvoxXH7I1iL5q8PBvy9d1MkLNaXai03b0iWZYUJ
7HqnfMgUuvm4kLwL82ulTWdBfN6dbX/GpTiSgRYDgv9AyR4CsRs7EY1CX8fDRL28jWRD8A49pN2+
sfzLpb1awqw7EBUAR6Q92hj/Smr2bX2eIwXechroXCIyL5ZkfWGTqI2fkXU7pOec8qRRY3Bn2rPl
PVx3ZztZa3XOsAdu77GWzD/4DPtfIEg/3molzPLFe6jkQ2Ek1JwrUjU1msr9MWv9shsn+3Ui59rp
tckLQAnbJEpXHAs+94xnNsDJpT6jJiLpimnmwMJfTp5A2/3amSYqgexId2cD7DwjpKI16brJr7TE
TeGaQW7Ch/KG7tNfQE35r+pQ3hJVfcLDBHiBtlo8vO0IWHgdaMj6PMsREzH9PE/VPzu/xF5HbaiF
hp86AX5H8HXlS1O3dRnR0o8/Zbcmxk3ixu4ECnnMJn6BcjsoRQFC6UijtP+91b1s0GcHwaCdjHqf
TRSh1xpMWNL6TcX4zyJSYt2wOc2VLqJ93nNPZkGTHj3aW80KcikmocX8b2i54CwkcWLbJwaBC7p3
Q5c6tQTtfFgnTXjG3P4h20t+w09oU7NHQuNf0KWdpCTgNAudt0ZwtRoHwTzNE+KA5smQhMPJGDTU
88a6HN4UB40VBzxRwoJbRigjXEv2G8rJjF16b/fxXcy8wwlqtApksho4UOQwmplVFyF49CeSF92b
hZeprLRJRCqsGOBY8iJxW9TLpzOrWMNLJZsvzJIDwfHBEVOyzhawK6PAgehioEBSdlECVFQ8wz3V
VRQe5eQkVXV0SUnftS+ryfTUYGxbcd0/xE56tzr5eQdJJR5I2JKhTHwQ0s60XgjX36IhOODPrJOU
5nYfR98kex+yefhqzLbp+/TJvT1Ju9q+qx/uejQxmJ2p/hpXpmQBpHEchAexGo/gs14inR+Sk+P/
ijHwkldbBKE7BaHZHnfzb1Qyrp6Ex/5pafUCAh/675+agM9H713Uv2DzBUJtljnp8V+4IQ70QQfT
pfNFRoFQDmgxtoo5Tb579HRfiITAgMsNmfVF+u446mSBMBB7bOLABiPE0bfv1C4xozTi/M6GcPZC
rks1Uw0RL/f9VEOwy+KVt3ST3CcBKIgYwU4zK0GUVA90EtaaS+q0JjVGBR5FriQAYS00CBxj6pxR
im9Qhs4LRmKEHBT1gqH59Jd9r8ydi4i1qa7NQP0BWnjkMorjbHVDDoUHVpA05tGrn8r39oieRM7h
7ztfBsa4dnSFifSrXOrg2BaytYhkPJN9pNDbVPEDRttefpkys7lRLEu2Tow+BjbQcdRJbjTL1H+j
UctK34+6gCiMQNjg/xmS7nh7DFqN4APChSZbImEvyPlwEb/K27JbvoUyoWb/fYYBepfG3f9Elc/K
HmYwXkBansLynha1XOy5pqRM9CTAjRAna1OKgrOquj7CxHWVmUlCHWc6X6lCnhYdn8dMUhRrGWsC
ycrWsjVacLuThrf4vZR2ebYSNTKQnlqq5mn74E8rJUXIBjN9v27fNti+8TrT/EOfRqymxa+RLQ3Y
Ew9twtk7LGhxHwmGF/4PN+s8Pq0POhuFAp1+jzuvoBgvJBGU9XDDUJVQgeYaGeKyr+qblV3km6Vm
s/WeQfB6y9sgfhi2fTHi6lZyM4by269+VGxRdkaetC/bwWgYS7RNLqkz0W+eUU3dHw/T+JtB04pp
7bhIxF5ksVNFE3P1SZ0GdULlNV/7NSpfnpvF3MsiC7lI7E2CAlixnHu8UwcqS/sqALpennmWFEl/
xjRWMv+03lug87w7xsrAtM3A7XN+YoZHjKfUkv6A10gfhnI3b16qK0WGtj8vYPIOueoVJdM3UBHD
zqQfuD5HKAAzA3uSCl+g/I1DLw8Y5oDTU2MNV9TJ32GB6Em2KXpKwGgwoEbgG9cUP6eUIK+EFZL/
OAw2FeQneZ7jwKbim6iqkjRo/8BfvQnsw61MgFTTwJvYHTIC1UM4ntLqXeUW4tg++sQWB8ty/VGC
ynW0jlfs93+tW7mBUUqLPxSLXtR0epIAvExTQqxvyNMcwq7QGIJRuhjKgBDjnmJFZh4NRRmgnUxf
Bqx0CdxqdHgMBWkfBv7KZ7eaSd395sZCt1vXhBGko3RtZtD8O+gqyIseobpS5gaPZdpAgYSQqVlv
4m8ibrg9aBU9KD8pc4grgttWhFVIoE26A0hnlrZRBUz0QveljmbGwwyvRnlBrGcui5iGFd3c0npH
rLCezuX397ZwXnlfofSvBPGpE4Z+fjxAo/ObwpBYk30tc+7X0asdGTnZ4P6E7sEWCKScRO2ujmqM
T1HmU+/1tuPwACQOzGPsRL1l8t4dx3r1IMmVRkXmU5uzGxz119zJTmpKaeIr14ErIyp/YSKadCGD
hMVT98YoISQCtLS2h2+L3EyjZ94QzBPWzNvUeYPinJhbSjSDrXbDXKpo+ekWvCNDyn2IhcBL08jq
wjWb7Un1dqXZ/7wyCuPaMSpeG/2ZUruTd2LZPdmygjH6t1HtBRn2ZxWwkb9/tHLjE8HZAYqb0W1C
6KkM8C7FFP1nvQbkNGRXd8UEKj+PXea8uJKNh4CDizPb7vyOEM2NOF1b0e2pkoJRY8Le+ChUjyQl
B9PMDlwt7epkXgYuK0dG9cHoqHXw92oy2R7sW5qotwL+rEmPOuQQPRo7VCLsDYPFeBgbQRCEell+
rrO2CTNDUf7gGB1zNaKLeGu43gPwqhrtiaUce8OZePgHLeiY70oNKenXkLh+OFWoNQlkPQ1RT2UP
pIjm/cwO52SuxzaoQgTGwUCxwOkmI5Gp5DqR2OxRKN+UeRWokzDe5ICoEuzfUNRhcwYeKdaD1Giw
MF2QfpPcoczATqyHjC3g/CXDiHpzfP341s8v3zCCV0Vz0S1h6Woygg9g8UjmbP7t00IKFy6XY1zv
X6KeBt3hvowkURZRFgB3qLSTF4YJ96XSC3M+OGpnkhYRAzHgWujwl5FKaq0x9Tk8CcVy0p4fTF5/
BSWZk4RZMuINygi2G5+sMSTraqSZfAu4gOXo59Y8Tm8GIm34RaQ9MJLp8KvEuoxbFgINTio+dpFr
fQkJHmTIGV4v60t0LUfUS1O8FRoBDXx2LYvvW46mYykAYvOhvxu6bwJyzYhNKDsCWaWhw/KcgbEh
8ikJSRnI5ld1J/Wen40GUCRrgFgfKlU9V69hUMHF3XFB8Smngv8d0/Q61msR3s6NT9S1iU51MPLH
pMBQ6xCkfkXAAdEpxE0TrU/5q/CPT0rz2Q2f5vlUuSJWMVxOf7iV1PXmx7NyKY3jMs2/M2pH/6kJ
WZdY1ONXPTBYkg/sZnwIRxNuhEQ4ct4iU1PgSUkB+FVkzxL/IaPfaauSxAmTsSXUW5u3ZsyF0Ahw
L26CnS/q5T8aJJQ3YGy0xvFIv8dG/3hp+ZOlxKNyVwnUEH4mLo95GubR5UVk7xFebTSYuAfRbCMg
rRwM5GH+HSFRKWXcWLDGX11ucL72F2iETpG+ERxOGSGTTjL7VXRmGVWCYqRHy6aOSGI83DXYtRfk
i1kEo91jbLD7atkqaWlPusslVWzc4aNdUBdI4fDNvvzbexQaiu1Uqmo1lqwlv/azwI06ZU514I8a
k3mFZy2LKpX4qdSlKKf6l2S3t0gS/8X0rUj1MreAQPECnMwcyAd/4cgtJ6GSiVIFP0A8i8vcKBhL
R/w11f/nHIAmS2bk3hn4YaCjjZuybirgAAm31f994Sdr9AKNx9SoLrfMUT1z5OXrHk0f0ubb2DIy
RPxM/el8PPnawqLmu2uoNzJYSelaCCqRaHHxqpHRRGMKx4mMVLcPVjP6L96qq4D3CGNeH8onsdNp
5knRlEHuyaiotJ33p+xukJTyfCtfS5wJ8j/YvT7SF5r2HAiNOoGBEeGBK0D+LB+O4CRwr7EyXy8Q
IfgXDpj1WhQqjcYkl5zT66ocjR+WVzVHnkJWccm5mIl1aFlKdqnd4YULbQb+DH1Ap2CLJXRROFRd
DFwmHFnpLWUQD9foLg9iSXyQj/HESEkkINIz/ptsmWGTQNtcoN8y962Fohd3vngSw3c1+DIvm953
vcOG4vOdG1/TeC662HQjsmPqb0zfL0eqRTXb9n14xgXgGvIT9mnZEaHqjQGAvOoQcTsCwBe51uOM
lfDDwLZLsgc09Xk2eb6ZHYxiYgzBm6y+fNugKlFdl5wg9ODA2+WpXJ2pj5jh5kEW5DAteF1kddsZ
W1IDydkq5/YZJ9zGu/rQJe6cTbYhJFH/Eg84tQRA/J+z2Q1UQWsS3UN5SeDjE1qqnq3ncJtVEJKV
kbnelz48Y2BFSIX+L2JnAl/yjBPyCOHzHbRcZ44BToWaMEftaB1rBwzc8VDoGRUIhpN2aQdyXHXe
xo1O69hEIiiP3AQ9bcXaJlsop5LLEWVy56WrH7usPFHDVFViUE9MzfYDoMnTxqbw3yPpgw/6hfZv
R5hnkJxtyGdaCGpJezfGgkkmgdaUfwmr/E7PaxwC9oq87C56nSZY8NY2341IZC0n5HrZ2DIG0XN1
tlAQPrFPoFbArcOG4u+Mp4kwrfc8kzwJZwIHbXxT+/cx+153VAdqE5F0fHHjXebxRsfJl4LYBHnl
3+s+3dug5xF0GwYwpMBiu7hf6/QGAQcWTAn9BjrpAybkWWCvR6jLFmjq+sk/Vz8ymsA0bZA2Yp9n
8+fMtTFLlcSsdF5V75QfjiFhm+tKaeXaBL7Xnz4Ri6QRDT1gdK3iySZsE7lS/00kgqMgbPw11rl1
6EO2Ffrp56h/F8RNgSYO3/2YDMRMuidoC9LqGCYb9y1spMWA/mmKRfwR4UNSG/Y6BwVMsv8K0JoW
oM+TGHLeRZtm7R/YaJSsWs8LWuwE1S9LcYzGsLsH2z6Oj8ocqUDkJotGnI2DE+oU3128VlxvcQbJ
UTNNx3ATyT+VW5iCeBn6VfA0QfgkOhQjSIZulRKAP6N+1zsB84TscWGtYHY2Vx9OK8MDfrlWa7nZ
jQ+rAFRuWUOCJURd3UqPTeHKnCQ0mC+OKGQ5bUvtFjqNBQPHKGbE6GujLfFptp8lA+OK+KbY0yAy
NZmET1O51chZ39MZz4LomdjBiISM0cjSl5zQLjE9QQuwCTr5HYpGnpTLiQyy8AHUMUZtLDLenMkK
vWSJtaR5sPPLZVrbD/JKCJy/T6MpfeP//jX+pkDoofF4hIm2cOLvs+MEg8C9mKGbJTQD/dIs3J/q
E4HLBzLR5FCLW7sVnhfQSeOOJ2cildG8vwuna9rX4+3aTXcobQmnYzz/w4WjqD2S2cmskTff9QOY
ZpSC8OMmRfqnFcoZfRtKZjeQE4/ECeyGQmvvjqIr1v2p0CAvCYPKkUtwqymKlJ0krgFf2VaSf5sN
sDi2b80e+uzo9Cr+50YWZ1UbFg1IfkOzwGq0sMaley3wiQipfZSFHH+IFzD2VbVm0KejM629qP10
/liwAAKjYR1kGNIF5sWOlSETn5GmRJTvo6NbVt1o/M0/FSgeuFSPy+nTlApLzSdwr8A/aeUzgB+s
ypssqpqIBynln+N83jwkiVmHnQ2jl5D7CGKpxlu2mXLaJHSUjtMMKw5sF6LYuMWPoRYDrRy5R3ak
vp+wa06ngVEZKvf6qpTz64l5L5JZ6FVxpSXTqpyDbCtGMXr8qU/e6GAa1GEPX/pZx256Wtbrs0Wo
ep8hp2P4hY+2eiyhqOjNEA56JQ17rYp2IbaoTbCbNbCfgL/ScTTMHg/4SnYjwQrmBFeveS+dUv/n
EZkWeAzzX4Qhbez0bw+mWiJhP+yXiKHYwfgoNrJ28SNRhz6c2yVnkK6KCPmf5dxzSuxHuKXuoS0L
LhKLPnvltpiye0IG1yV/LQ9rratKwUHCwIIu0Jqbw95FJH16LHO/0wCMIY8woSCi7dRZ/DuonWw8
QJz6JzhMRe/KBR6IM/rVrx++nSmQ9GvoC73JYIq2l1E06kI6E0+E5ySEmTmuKjzWkFNns/FV24o7
rJrGjmYX3WSuc41jAzzzndr4r/IZgCaFuDN6PXLchnZ+Zt0cWpD8Olgi9HVH96QSI1UKrn9YwydJ
NzrQsgQviOZsjP1CQfYmoYTYqqtYll+XR3/k0Tezketna8+3JUfWGSCMoOIL+AHvnRDI7VT5xS2p
MZ2P25vLQKbjxxjiihJaNqVZr9TdiTwExM6O4y3rj3ywMLwpWHBtc31r13oqCRgoTmFWMRdo7ajj
ys1ILvSxUh2ITa/f2jVbXcuqgKtViXNCnNBNrglphFQc7rvAtWWSSfScQ08Ona30QADA68KXZ80W
Yn08H4Do7ujElIB1YaDMO0QaaChCP85IVh4O10AQUL0vdg8iS9FWZOHLPe7gXeuMvebO6b06/uR4
nIuaA9nZNIh+AU4xlsyevxSfe5WzHtW7PWhoVw8dBrjp4rt/Kc0hvn0hkW0fBnQkMg0+E+qolkx9
uepfF/B32aZY2rF1GuAFo74diri5Kpiwg2eul/Yu79hr2KXb4hVAzp4JKkhiyuLBhDBdDs9OmB19
CzrvVuUeOShRu8JrvYp31VOyVeJ1zNSHbWtgsvhfnX++rN92pMAnByXc+0TPKJJ/5qFtD9RwAQO7
zWb/ZjIPlkFjO+n3OP7W1x2aOc5ODYz4141MHPHm+WCulRNVze5TdAqSRSnny12CkqQTdAHWiCs/
2mnVhog+8vaQDxTvGM6r77XkLXwBa3fy67A+p1Ngquf4djvhlgr+NtSaAjq6fGjCg+6BuNBIkJ9M
TBWyM4Rv69XvyEjgK9jmuHgSoI/Kn/uO2b05YRayfGr2W6ckZ4m7WyXkdFrsgHIrVKuQJWQ2Aj9L
WV557HQnI4GF9my16SWTVojjb63tlrc66LbvZLF8ImpU0jZzAFjSsVL9nMVgClU76v+FlAujw5fi
MY0jLAlUfkh9hF+XjfiGbz3ylPJzPIwcrH0OQ62gqW377FkYuUbU+2+HVAd2uzEYNvk48PtOm2v3
jyhEl99leqUt0q1F5ZkFGXzzwlJnQl3r9VOONKRpl2Cbe7hLIyqdW7WwBvTQW3P44+RduvW0HjkI
1VVyiQZ1HzFUDOQfR7fkPF7wSRcjLmCRaEugpqU9y6fl5LZvmQCCGtfCgGurNTqdN+E5tvE2LKiw
LMxc20z+NDp/NAMBc/Ti3AuRAiWcW8Yd+I9Ff4wRmQ+S+xWrVT1HQKOkpEjhCluK1XbPf8/VGgLN
lcijEkupscj1JhZr8eVbeeiuJrhdkSRKuZvnyqxwLEpVZYm+zMcMY8oUsvgw8jV5oaBrRhjYwas9
zHqecu2ZKsIjii/TvUusorHumgT/4uVni+uC1u/swfkYNXeH5u7Ix2YDZOlMBjkoP3S39tzBv2BH
M91xbMP51InfrMrcihKsldMFv/55+M0lHQRBpGRMhKZJypvozprYXS4PBPU7CpJ2D7FpWFBAqYLB
5tWXQVc0Rj7jJnzBjJ+tN2wGP6TokOi6oaklXnEVtifKjzKhZ2asN3chPbe/0K+jV1nj3RXNJiPH
m+AcQ3IsjKVAsmqoA60Mqu5oGGCWkDT7Mjrdwh7RzFOObytent39HZjchVglsQiMLjEwEqBFSzdi
aO4pFdHAVwfoeoAsKUAT2E7/BO2zHN8m5FU1X6cZX10SdKmPHbSNQ7FClTxOuZebU6Fr05Eozo8C
LLKbahd7E86vqY1INSGW4S2RJGPR9016FXLY8+BpPIFPJ/X0KZopJQM2GGXf3dI4o666vPv1dMKQ
OSy2MfiUCHpypXo4AAm1BJmzH8AazifyQVSAPRE3SkHD/rOQSMmvYXf/R3erMSViLCJ++ohkKk4D
XeCN6L7UvAG2ahUxNe28NYIa/QhfMuu67QM7wPqiNCbketTqH16RjgyeIVJja+bk7uOn37pxAobW
ZN0jQ742RhWJ1Cw1ps2OLBWculoQ13p2F45ttpWFTk1Mx9e7rPRUF2nr/bLv4H+W6XMkiw69m4MN
yBXQvi0lshvVtKpqh77qJ3Ncr6kNBcvPua9KgVcvreUaBru7DOwPnuWpujxhg/WPVqBtVbGgrIFW
cG89hF2mupe+imDwGMawczE5APBd3I8nGOeB/IAWpnxF9m3N5Frj+FLZQTcv/Kbmj6w7Iqg/INqi
zZAKvPZ9hczWvNofTIWttCG5pzIzQmWUC1Q46ofL4+4MwGmmuSUqXPkGe4YK+KYzvXwPRBBoG81K
oCr0H87qqBun1E417eHIRqh7pW0wYJElVRuwr4HD87uC04Qpispco7LP1tIOGwCV7SaCcEPde7tW
/fxfuKJsizCjFaCmXV3d30JxrsaQKD0t+f+hN19yaq2nhyOCLcEg8IC4KT/lwqx4uKTEeic8DseM
vdGPWsI8GXZhEVy6Fg81SYT42/aacwOEFq3EZE5ol9fjBciUHP6EwxjLuP/qSnm6/r4z9yp3KDrC
ipR3Rj56rOr3RX+etOv+/XGjGTO4ZWwPkPVq8ok2O56oNevZGHVrGjR92WvolZ/XpbfGJJgNHF0+
6n3jZzIMOhJR7A2wxYx/2YP6EVyks27rdUz9oNrMURLDjdH2knHsb4mi+bSemXDaIEuTS4zwcZBA
qJZPPJ5dOAQShhN+mc9Q7HUoMKZIVBGp93wzw8vBbHjwGOm0o4Jf6WJ0CAg3yS9DUcLktMdCDtme
9+9TcnnxJjfO8bYZnbCN/ml2EbjNZBhKMlWQ7MX1j5jHzPyzab80SKEwS64Xuy9VGGiWh8zoEgrw
OecSSQdbTgDp824FFojAJwRWY57PweQTL3ds0nRNze8Yy5/xcnXSTbPH6Zqj+XTm26qipfRGjd3y
vd1tlGZGeJvmJerKDmRZ6DSvY5BaH+MJmb9D9LzQ/E7/KnsyzW7hR+H5Vdn//Z4fwJh7EEEQVMl3
q+YnIQuQWdCW3jd1NQ/v38UzoxziPdySQIGP9rMgX8xhlBQ7RbvR6aB6XyHYnBgVNDLEryPSYlJd
PcEGBxNHQA3GzQoBD4sFlZPcgpNPIsjNY5IqmsYw46KPjrb4dYJeIG6q8dmPCORqoFZ3Ly6yBQyx
EeFQb0QNK23+0BxV5Vgr5ZYYCRQSzfx7xjx3IiTQDhQDwZxxtW1pAc3H6M8MHc5bJIBdfvy2LmGj
Z7p6lNPcTt69ru5f2pIETYCCfK0P50byMpLgxZ6eSto4zr3N2GKca8bp7qS9OSuwVSk4TaUep83X
7JhPQwueexNskDHeSnN5+gRYOAMOOHHHEWenuBB9jdtRy6KoMgU2vCOFfpm4p3ewo0skM7Y7PI7u
slWvZQXwUOt2TZhkqNjPwhWn/k6kO/68UsB2Vikiw3WRyd4H3ldX01GAwhuGAnr1GthJeXLLKxpd
RkMQPYKce9Gf/7Rak7tknsDYRnvvsy5D8o4UV4DNFP4YB6JcwtMFEtNGqj6Ytn3rtx8KsTZ8gA73
XKsYG+mG+dHNCCcmuA1c1HJcAzv5BMawI1dSfg6uJOfJm5mSlSyNqPWghtXn8t8ioBoSiHJxerRD
IQUuxgTK/BO9XU4MQKRXIqzXY0aP9fPcGy2G2p0Bermk/x5CqshoDzuaHWMWDGJj/YnAMaKkNd7s
rLDwUIF1a4ZiajZBCyouOZBYCE5cdgRoRjM6MmT/+DdYLsyILLVLDmIU/oU68qWavM8OoAKCy9JI
YR0/LtdW6yZlZ8gkM9WZJ7zQ0niqtjHo+ghvlXimAknKC8NFn4f6Zu9I4fjJoH800n8TDxKiR0Dt
MF+ZdlmDkSgId3HR7aarZnTDzh5uvi1KGSDL7Tf3DRlXToZIWj5gmOjjE+OxnmbOr5Sd8zyX+2PB
ql8I+BeuvRDTtWhIKt+N83PJPmPXGS9h8Rh5HqRiJVDSe9GpAu3BuWUzSy8vZV1MyeqqhTklLzMo
6p4mPyDQ/Jk2JHLrKRuOq943Qclg7eFnrHxtUVMM3K0O/DEgnUz5nNNPnVN3wU4/SFJJfrKco+IC
jHp/oowuCUcb1KlMHRu9x5R9OGjXUmKI6JcwFI6kwWpKIIj2MxQ67M4iiWI2NstZCvwjp3fDVF/G
b5QqwKjk1dbVkIawxT3WPkj7bsOWSgGAd2AQWUdbOvur5bwRFxVUuAUUIfvonM22zheTFe4T6sY4
CdSTka8J0uajja0oL+PUZ+4zSBU5dg/woq8fZQaC7W6dp7pKVt/fv4j75Cp1U0tsloDV1EyxnI7v
ye1AdOoyaPXEz5/f/wWzSCyETsJ9X9bMBXgbxCa3RjipDD/mYeNmyvDy8nh192463SqdaxqtZVEk
6lxy8Grteac0x+R1LGSmGKpqtHsYoYR+bscyVYGruJXdEUY3XDftFZMoMWuz/7ye0xP5BmZlZCnV
6QbMe4OFALbE6aEtBwyv/OG7c5/X51AVz3HJOvYfO7gsdNQdM6nh8joqJblqe+hXexEFS6T66ePx
Hh7cS65QcFObN3xbXnz7rd4QVlmlsW1DsK/Vi56aNbpcw8GnA+f41EG3VdjISRA0bm2OJxF8xGLS
Z7HD2DiocXPgZhKcT8QhqUoaScT9S6blnGms27VozmrE5Zlo9oWx6rPQRM4QHrraW6g9O79X0KvG
4AlmXdzBrTbPyUWmJzCrsbFhqIMtOb5fQ2XsBv2aZXUJfC1u03j615oijOtPIuiPAEX1+UBxlsou
N0EST4SyAU1/hNFbf15Wz9Isty9s6UgpD3TE3yHfxn/p4hDe+NVpJjFJj2vgRiyk6YCcDbrzA8TM
H3xSywmX+qH2rCMqVAoS2a2w43ndgBry9k/u5W+35eMu8idRlg2keiDkGLr/wNInKVOR+Djszvd9
8+VIe/oAx887itG4CiFoe+U+r/MW50vASGFzQ0C53KdjeWcQZPn4tnDtZ91fAPaDak+RB1QJumxk
Ri8KTz1Nj5OhEwtPh/OOkH+PWAQLBXIuY6bf9juQ8Xgt9LQZRQTqHNo1Tkzu8YnJNp7MGLy3zSom
PMpHJXnkDZ6IOy7BgWO4q53jIoJSfbUzd/Xi9jEj2v5bgKUgOKofU14pxcdusbHBf8nToomhE3+A
E/hrEMc5lA/5TRnMr66mNxDN3u2p+DLNHfFuZXsgFd3MSXPFkInf/An9n1YdyFPblr03cBNsU7n1
bOcaUf5xaqczGKrx3QampszwzjMhZiig+iGpUw/7Nc8LH+oZOr3NRxTzEo3vPXz0XWu6IpjqA4cs
2bGlv3DhqclzB4PDGN1+vFJWimeQ/1PiGeNgPmhX6t9MfULWdI9SZozzaqgVzKJU+y0b572OZSgI
cpMxjlbKYxZXYz/3AgME1Vjs2zV1Bbz4+z6NwQ9BrzjthGchyMN9IBIkTnatjX/PKT4zIaE1qecO
u108u5KffW7/9qkK9e+aJ1vQ/xiblfk3TZXX40luX7O9p9m/n82Q9sWjvgcTYd4DMlJGrAP/Yru+
y+sGiehpvjj8O+QXaXfALUt49OwA/ZXj864gqEWOP9g+H8plnIkz0o31iQ9jlQQC+RNrvRmZPAcD
iC/9I/jkcL4DZIxjI+voGHw6AHHNm4gb/P9+boS0iNX06m5h/JuqLZJHe5vHOclcDUxqpaJiqZmc
HM3YoDmoiR4+6w8ywqPTzuPFAMS9buOrWNaK6vHK62ClV6YiH4XZC2lARR98U9zoOQytAhTg2V/w
UR1leFBw6Uaf9zNpo5L7Klajtl7GLxaRf3RaA8nBAmFp7jVNXxve1gQ/s+lWQqPGNLKtGhxsUk68
1LJeqdAeZD3nJJ18DgX9AN7lBGCuJr9OdrY+teNxsqWrZ9MspKeoJG/ZebSVAAKHOas8PTUSAT0S
rcg4bY1x3dE1O+H/A7N65qf4Zpck4zSJnVSDxVYfQ0VgBE/FunaNGLDLt7R3lUw3Is7wx4zhbFe0
tM/hmOdiIlEfeV4/nepk3RzMmWzy1aPIZET8hkAE4ygeCpV8jrNr7UXqRs56f0L+Xoo6+OmqWShk
EhNof0Btw/AEMbTcjCJesg3mZIPvAoXryWNbvuASOi1wsuwSkH1bP8aVYpfM+fmtYzNjZnWhAT/x
cL2pUEgDd1wL2cgf0tE25WqZuaO4bnEf1sKIkxXFDgLRLH/+rK3IAMqK2JImkb5z+9phyxcTZ5jm
5Sg0WoTfYBSD7OumVtmxiS9xWJASlYLP0jRCjw9sHGWPgUjDQhUSy2NuKZmuMplNnWFfamE3qVPc
vwtQh/m/0O2jLWkq1vldG2PtkiZAPmPL9qNvetcAQXnHltiy92z6nkd2BVl8M8B7k921VGs+mf/i
2G9tVMLBa/5kagZIVf6CNSmP8niwlmOzhON4GV6vNEzOPb9bnTY0XPJrC3TgAxh/Wjo823LgQvAy
hKqWSk6y6pRtlnGlETHT65Ns5eJUTdEdhTnD4W+HyQNmyxSQnvKZb9Z0sPpG5/pBzbM+dxQ8eJt5
RZS1BWwfN8F43HpLu5Z/l6IgGK9wLfBB8ptx0WgMLNvKtLZfIJQH44cXfTyvRoapsEcVApDv1z4y
36WQ6Y1Kf/cCmH9ia71UbDuK3RDXpNXcRFWOb+dGPW6PRN1h3ulIDm/YwB9JCPMFk3IRzVeYLWGt
DbH7rCPYeeQZ8uMUflklaZ1yQ5ZA5nF5g/PwcL1w0mSKRUq3/m1IrOTBm3iGhxK4JHbtsr0SgNlx
va1uMONjK6wRFpGkpZQcR+veSWzPoNWqkf/JDmcVd8eoFPOKx8mlWscuVOlo1E8p/okKWLpvQomY
kZRtr5qxAsSeYlTmT6gBRjf83CxShw8iAc82U7qO7kYf1WEtQKdz5nzn70iU5iIa1EMtH9CuzTRl
V9jKM10za9pbWj73ePr4An52Ufhz7LOpYjEHjosx4mreXRnv0UJiS41YKxaWP/aB3BOe7fGiHm/W
OsfjsL15EcZ7XroM+wJVKTZcOPyX3CcwjU0311Jbsxgb2nFyr9N7iY74EFgm3X38rPGo+Ui6DCo2
m5pelWDeU1oj/c/cuSDHgZgEmQY30OFQt2OmYFBbAIpSwXccl4u6Sj/mR/w5r1FfPsr0CkoRFTQ4
YHkmz1xi9SVMEQIPrllxBV1eWR6iEFlLNLy2in6dd09FfH94D/brf3zDlOckhO0aOYte/74K1vMO
opnfpr64T49+7aPRInrKE12HWAvvI7UtkEI6RyPe+qzZGfQ8kUOeT9D/PlLfunnkuhH3F3m0S7er
NwW3nk0OSAZIBue2cmM1Em2O9pkMarPEOqoj7X3LBJ2EDkI5fBkbwvW70ss9/luRMqniDgqSfUI4
hdrO849JbvMRl8pXl3NifNG9MzrwZWCVrgLWHHBDGjSJ2KlK/j0yQvWkKmNkKoNc4sLvD6VYfZrH
g+sYFfuxRC0wbwvZa+QhBIaZkKIg6nhg1mVGclJt6naktQDMecXepg6qdY2trArCXVXqng4uNnY0
+rOl8ZYQ/DtbdISJog+d8TKMqb3kHzQahvu5NjPfsQLQELOeuBDm6Cvnjz6V6P1HYWT8KpxhFeQm
/zPpSSddHi3pRmoBhkx3PzTBcoyyOywO2omeQN5UQ4SzusvRwAfRLH48Fmy1XwsUEA0Y3Ozz3X4S
iYogvGzOy2T3ilzb1eg26/Jtmz7cploDaKndiFIMrazNmHffQTf3gYfXsTrdyP5afz4rarG0IMMn
jwBclyC1kZ11sJm5H3wdwcwd6KASwmsVxM5UwHziA9l+lP29iw4qUlCcmeDfI3wk6xlDCbP/0y/i
BQ21q8YjTqZywtlL16iZ0Rfrh77wozwCPk/3evhJga9LXGu+qIVtKSqOzTs2pd+BiSXeEAIbQ51u
JFx5YgHjIs+RsUi1XVqmPl+va45gyhNobNLy6ex1h13jucuIsRMjk4TB8/JZra+IGcmpQ06QdbTc
/0X59IvWzk6IGX/XcAi2VnRoyxQ3sftdVnct3kf2sz6pqZoCK2UtmLLGU6AzSdQXj7bWcT+Q6Wp7
bN8Csj4z/DhDuCaFJ0r+g6LYiQ2DXf4zeitUStkV2I0fQzj5adqqJKMNc8VGVC9jHpB0TYYJ4zqf
qSuy+yZSMY0dDlRPy+uryKvx93DMXOfvfFHh7LSjKO/skLIFMJWFQK/xSF5KRBG7ZRAxGjRcHn3K
orvitdyY0HdrgNTTnwrbarr021/F8ZkFSfUGZ1UA3/+hYE+1hqmtTE2FR0OCjN7UI74kTH+juu6o
drkOjCoVimxxYdyiTJd4jN+tjiuSUZ3Vhp+y5S39yujFW9CgbLDicqHUrSrTtqtMuC0VQP6nrV8B
ie6oLh7QCQ8TtBndg9UKfHWvtHQFZfnS8qIKGZEcXCXwXiraef1VAE4F6Ehm+Qd7ffeovDi/6XJO
beIeR6IrN/Q45zp44WaK9hQsiGphU9SrDsveB+A7FYQbMor4qIBN+01TcFKrT3Ab9zZzs3u8Gpq4
gSsAeit6/zAKtkendlq0kpF6kIqIUhEL9jTCWyi0myTPDKtnrRKghnVpFgTK69UhXHI+cu+HQqG2
qnsf4xnDb69idoMHsaf3vIs265JOI87e6awp4VgCNqHWV67/b2Gpzz6L4sTc3uvGvMPOcZtp/DaJ
PDeC6l9ynF/+tLxgCFd4wc29/+YPPpA106DU21Ci7mZVLn6tMU9u3OaHdS5Ugo66HRT9isH/STha
h9FsSVPumpkNGWS77j5yzzZkHTV2EWgdJqh/yIhaxEwoVydrdsX72Klq9ARxB2FtakxogTJgD/qz
ZjDc/wc+oEvzRkGnlEDRxVL8JLjqXMPC57cfdBZ9yTMvZ7EL/KM3sDuYsuV9C/im9j1zQLOK1rsY
SBwurg69m+HBsu5kgGRiTPtG20S2CZTpdyzoXn591HSlTTlZLLpNe/+ODJ/bDisR564nkbMbiTHv
cKx0AQ1lRbs8R7MsnQCFsy8IEEFoiuA3xk5uGVm+x58NB4gvrcUWGcFrQBHzvgR4GlNd1JyIYUkL
IqgrGaFCJ73DWl81nIkJpj6Cw/L6B3oTWHa0MyTgFcB1VhQuMXZnAMvDJJgawqp/KFDHUGbTxwIH
mwzUImITr5Mity2wMfzu4cnkoZLX1jSHeDjpUorUd9ebKig0DIYEj5wUixFYt4kxpYOpqZIS6pT6
LSULCjBp4K195NVWtzBomAQObuMhsWU+yA+JF2SYP8NMzzCurPCB2wFb/cixhf/swMIGS+Mg4uTC
uaLDwTV9zrpQlZoh8a3zToT1lAR213L1VJ0+4X1Tw7ZsYbJ9ShCeiwuwtI1YWawSKnG7rCLazySE
vzYPNta6LYR9/R13xpre0jep6f9sYp6B4RQG0IrlAmCnTmUMu9NmzdefI69EbPFKhAGrd6oaHZfb
jAir8RbuVxw/7zmoDPCAXmkNZK/EidgoALF/hmf2+pJ2TzoLJJ0f0CeEA8/GWObkSmtQpkVBFegq
GNzOpdBp2Pg/kkjSF3wQVL62yHJPVHzQPIxFDT8PBlPddUX2z/zQd5E1iS6f21LRZsO4F2CPRjm8
HSbJPO9oLBTuGIVPvYXMUwlKHT526EHfKJzQB4gILsxjAOczpk42X+nguB/NlNDMjTAUtld7Kp57
5YV6v/LoHiUcd8jATGHl56mhOlI42Ks6dWVtkFHzp/5S8Js3MNsibHzTbf3YUpCg4wHMnuH1B1uK
hOmGOkSQlTS3aeTTrxbnwua0HMU5JuJ/QOQfJfZCGf88bfY411EfOMaq/eVZDoi+yQTZDMI10ZHp
vUz3ehHCDVoJ69WcP7EwdKiU17d08MKAVF9pchRjEG3ZuOOnZTMzCtDCdO1jogOt7Qu5ZxTcXnQi
dYfwVgqK5kKDRWqhEtlyssYenAWYYv+aCtjUyTLgL9EsfV+qRaFPZ2uEWWmeaYiVeOclo14ippgY
80xljnwcDj4s/58ogW54G12hyM+SmwjSMp7c/31/uk4hfbObLnNZYfYtdw089zlvjL3hwzq/yysT
kMCxVT2ZP0PqyDnIOHih+BEIY2fwdMY92BbFni2hqnyUxuEx7tNUSaiE1WqciA+fJAJkwCQ8StZW
CUj0yVuNZdCOKtkHp3tORuoI6Chs9cIVCLsenfec5ykK07pfO9yK/YusdhWsIZ6ePt6B1z3DyQxX
eZNv2+1MOA3/IWtzWJyr80kVnidb5t2LgUItAW22uunlThpXneQVb456mvxzNLAvBG817r6NCnng
gbcJh0jm8cOksE83DfcbbyT7/X8vWtfS/thmBqjfgmtLKpQ9WmffJuROuQKRrSJsx4+YfY8cyD6I
4Ca+FZABqIC2XDEtiTKJgtAVFx4nfkYsUv00avFUYnz7FjvuEnZD5exp3nAEZulU1XCkSMt+QW7Z
7nLUReEtbG8kwAYoXDn6FDClbvZe+yLDpCESkTx67Ss3/AyhoUwEeZqXJ0ptC8+ZimUV5kxB2NNR
Q+RRnCpTHAaka48TPQhd5y1LfxyS9pFlu8wfCEx2TuapvVPf+3DiV4yFRpy8wx2DskR7GQGQ7/ya
kRH+KU5YsEJQpAUebh09IBOxGlv8ZIlC1t4dlvUi+9YsG2l2uB/i0Net6vIWG3tmEcx3x0OImjhV
dGNmrufa01S1+gpXJkRzWVvKeZ9S7j8H2/DVIkGEWo/6VYxAmQWNRN+U+ZztSrixag1FZxjFAZJj
AgzI/wjGBbiUM5pp88px3AEuS9IoPEK32KL4KiP9Gq6uuNQP13rNY/e8lDbca2a17CGmzaqHKrCy
moYNNpvcrQEmvy70pxvf18pEa+ARPzdxCIIclxOAO1b2DhBiFvAbIsM1zdnDjy3DfI7L4dz+X/0Q
sqiHHRx1Im7IIBx5cHC9KSS0tir6kKwa5lzhqJIYq50sJez/5l2kdd987czrzrhqv+sGe5xPZgzy
35CzySmKR3CzkYQdMGcXYhp8P6890rCwAhtLCuRemFK8hwYYrexwBiOdfgDvf/pwrFJ5o8lj8cQ1
h6t7b143VT8ExpeQ+DBeT4Ju48GG3NK0AZY/hYYQR0fN72aExZbhxe9ZlGyT5p9SxqiNVJfd6weE
qdvsBev+Nzpvz1AR2z6gTPBuac0KtdxI7Tqk/bY0aERzb3L1fGT5Y7Z9Y9Lq8K8W/1b8Z1FPmc3R
1n3blNat+M/McAlbbVqYy2PtIFbkmfHyBHVbMIK16+/gan77QgDfvjksFO/Ffk1paQNy3M1V2zBH
Z1oCf/RD9h8kMZiZ2uLm33tgwZTc6b3mY5FliFdU9cmLUxqppvsqhe61uMOGIcuszevU2sPipbGD
0qWOeaGD+1EAjNhK2FjJzNm4ccGCx2T5yW5KWqvac+mXGaW1n8vT5d18/wl+DPpxsQljKo0rwCnx
GPlLJVojyenQ5VEAvk3CCiAbw/+1aZZ04ZIgD45nACFMAl5geTT4SLkHKgJ4uZX9MYIFhFgjvQs7
urg4H+eRdKlkT4SPle5SPxIx51wF6N0r7LQ/1viUnHPhFSAe4Ocm8skvgFH+R2jl8HTugMb4MAP8
DAZ/DuRCfm7lMdn4O/4ZFETpT5GllHZ1THXDfQ+GNRZyHZB/raYJhxvUWqo4/oHddvdvFAWNIYeQ
VbEaRdBIsKN05SwyRQ5BIWZXnwZtTAsY6AHUgWYPU18QOCzO8bUdLfU9LOYYpwJw9hxwauc0tdXJ
gXhUBsYuTmOY94QbtPMCyGtkPXOGpetn9SyGdPcLpXcdLEcY/SsMYlyMCOwcNtP/L3XKYsaI53c1
+10l7/Pjpn9lRhaT9UDZw4XbPbry0X2PYV8VgiOUIzpD6/Qszh+UclDjpuf8fVq3QVYuhXcYy4KM
ks8IuXj6gB0hBvneyERBljQBgXowfT1A6lZxPggpJJbH9aw6isvkFrftYnWFG7GkDX5HVO1z4zcZ
ImA9uDv+cbpth6WPyHSRrpdi7LbL58ppSt30EOePobc0QMU3Xu2VSFeAVtFbvudAxmQ1hifsJ+d3
Pc4PHET9eTMMrHyg43kuwN2hkCJeVRMOhIp9f1uO0Lc1/2kp+RIijY1sVFXlFNFVbrc2tXUg4oiJ
ohrfKt8QoxshMZfo4C40vCnbstpFhRoZK6JBc6sFbaZsl/0i4RHEnzHcShGlfj7QiLsXGitnwdyI
diYOXx8IrXUbjjzDp/lgDuOI5tcYrLvyVCBx6nlXkjTZCRSrLvuhXcsVlUlqjSFIbI3/o/4oVUNO
C9Hft+vc5bDsvUHj0gN0sikCihNzHhwejCYbnImb/+Pfq0ZVLKXmjpPDbloSna5gJ8N9HoyYtsBN
xpZu5gxCYLKNyTDxcaV20EbQ5hhwSsZxZhUCT8BBq5n6+PhVGPpCgNJXdHrdwr6aQoFecTbG3AN7
dqKud+j+gMbx6oQlCLowh9/bub3pKGQj3B9CTzP43iIGHlJAw/Jh2SGHbMFdQBdNRtUKhOOO2vin
Au9cnrAMx+vaDTryt65gZUqVwicNJcwXRMXECzGXV4QLxTI6sS/3GJaMWdYJG0FjHAEaEzz/qBty
5QPgJA9vziq0QN8hBirKF5WDTWq3X/KAfDVFXFCyPm6odiL2Dk4ntO4UQOQJR0gI+6mZaJJJ8wMV
4T2yfrDKqNoMc/kBpgEJPFhX3cCzDgTX83K0joER7m7wztt9ykyaI6vLneR2zX+wmH2ygE0Bk575
0KebcI1M3xE0NOHG6kp1Yi9wpvcBTBDjSgLUQYlZPYjmyhRYtYfAshSfomCjbqMIbsba8sXHmLqX
50AK//VtM7jlPtRu7QYsW/qLHQkrEHsuJrtZQh8vfJ6QEfpTZ7M03RDIyysY+7Mk1ntUjHY7ErhJ
T5MNIWQUr7sxdhWoMu+8roGicDBmvsFbwDi1285UKlD4kgLtdi9mxbrQVvvTqgOjh1DULTh3T6cz
d18r4OnYiAW7Pr6tutr1+jgUuA02iFPqDgpdQgoruKIlDzj9swXAHXoebJ63rJqvkO+D/iSz2LuQ
n+etIwOWgDAbN/d+EG8JGWQhSk56LNHKqF8L/ULNXJPmV5mw/lpAVr9B8PzlKgUw5b//HlMGKajn
aArYU9vhxk7Vj5COJ3uUUeBDq5s9M14KM8pvIQtWJZAlfk9ONqAKB5uXokyKwAIKWRGKYzq+YF9G
RBGPZ8zLEImd0SRqUnrm2ugk7NEYI39xvCzr/xIaSJVf1zT5iC86L0Sq9U4xCrgeiLbH4hqXRDj4
GwptW17N62nH1apNUtxczByhB7evheGxGO5DnijGYlMH6xprd7TbfySFd/f/eHhppYc2tu61nW5f
VKfsOvS75cujPjkuD0hq/HjvGW3D2dEU7z3ChsNsSsdmh6xp7Um8hSzC3ormRpf5ht98ftWxDuBD
jYATagjeOB8GharNv5cC7SH+tykruTVCO8ANgCdr5cN151kC/PRaANSXfme2bU91HirxzP4rF8vW
+axg0t91gozbofC87Q01B/miIYOMtkJS+Iqzi9HLRJ0jE2L1Vjgr/6HvkMTkDfiKfW0Duumkx2qn
EDIpYtyShePKneBDtIeVKvm4VIXmGYXOXdI8twFEzokmE8kzMqrEPcbdmJCft56lGbTVNo30QS20
X0e413boPKPcgTLCCSA9YnhPpfHe+Uv9Tu5nnFZE8q5jpak08JJJblLb3qxYhLlAQ93QXcm7dtIC
v63E8DE1qIEClyrkJd9IJai0B2581WsMTGt8Hc7qv1s3eWYM0urinhvMWUx+drBkk6v7Wg3QjuHG
jJ203N4hHTxM88YMbMXoDJhs8O8kIhxoOkqbyLEsV59j2KS2gO8HojSWYfEpUy3ZBXoB7PkBEwiG
ZFGYbi61YDXrOXmnJiCtSptCEkIkdFolXTMeUi1ZdDKn69xWXdSwg5Acn3l+ntgoxGsEIVY0J/cT
mwbLdlsiFZ0TvLRwtmADprVPLFHWPjiHHsE0R7ORAkRzX6k+2yXrqPwlSG7AIGnxBtj56mLYUeDW
YDGYE2y79jpnlGi3EkNXcqe+FVS1fc7J6mrpeYBQKonZtWr6djIM5xQof7GSF4+XXKjRcVoN6R+u
Z4Oe9tRc46gIVBnnWVruBuRcnl0oMAywSaV4g6i2TsLMLsTZTXMxVWq9nrxsuusZE1Qu0Ho06w94
ZKJ6ya4wT+m+8D5B9bLKxqn2hmhVLl8/pn+pxXHHhBykZuB6whOlrP2yne/Rp4WRPzMhePq2pOl8
wfwPdjQL9skOOFiurNZLP8M4CXDJPb5L4K6V+SISyz5ZlzqjHp1y5GQwXQCd1X/Rp/J20xEg/I6s
4mi16BtuUCE74YcpaAA+j9mOvyLMbeAdv+UPYOyX//oKHU9cxwp7De7ltEHEO8xY8MUPmo0EgFN5
DmRyfkYKlt6W76+eYjF5p/HEqLlm0GIt+JPSOAKuV3MJ2yf+epx16eWZUjGNLNdO2tCTo2PvQM6x
UxQ9iK8dnoAVWOhTLNat36cATpcneTpx0TedsfeNLamRWFcM+Tt4UQT8s8uNitgSzUemc58kMjle
XsZWwpelC3T2eNEwhuun3QY8Lg1BsiEzEDcl5bJbQaHmh3SZG3bwKE4u86vfN7Snh++JarplEf+t
szwk6pKomPG0ScKGZgcSkkpfHBAYcEgf1g3XEU8uutWdEL8cuegqrCLh/5W1bseJL7cURET8T685
CYc5CocNKSthGlrZqvRWICgJJx6gxdOZw+AZ4Pn4LNbOw/VCsJsGy7od28Hsn9kTv6ZdRpubn+oj
ioLE5buco0F6TkOPYXsTQBgdRpDiToy5QVY9n2lovgVK/e1AyGQHrnsoG29I6UVMuHyWp5gTO9+L
Eah2BmG3Yutzz/sKRIr/lWcXnHpzHziZCtMBDahWCOwRiu+ZzAeX7DXV6ZiBFMZjsqszh8vwIJSZ
bwI9C0DaxSPqG5G8k7OgVL9FBLyDSSWLOiYSReusgUfneoJyqBpK3ineVL71LfqzpxQdvLRfHOe0
xXK69JQNjtp5RGqOFlWaV5vFsZzb1eGEp3WKENtkr7CNc7VKf9MYv0SoCVjNFliQqjHCRF54iCH1
NNLj9vMU3hkUD6qAVZFtQgc5tHflhMLDrfqPEijP+HvoLcOFRqdGGUR3DMdu+gPZjBmjoVZ47OZp
DPUw2a0UGNP1nSSbz+/G86S6cCULIMTOacV56udfGV3NpfBQg7JeXS0p/N9J2wybXl+P1t+GyKTx
x8dP+aJhfsOQ9YA4OhnadhQPsU99JHLa6JL7oLphgJCCat9jg77c6SlFngID4pctoU+4lp7pb7Jb
9XIl7NyZ2PtWZLX05K2/Yldg2jEGOT0eyoQwpv/XnkQZxFuC4Y8bc9bM+42ydlgW2L8QoP1Yh9EW
Z6R2/M5scfG0UoNOUe+FGI3/Um87rPc0n0EwKzEpQSgj+2KWVMYY/05xoY+IxZpXzSkd5ypGM5Kr
ibLM+D30gJozez/0U9Mx6amfWPyJK/OKfX87J3aadQVQdqxd0W6yHKYbV4Ad8LRdHIgK5aOcg5/Z
ue2TbCZpALNaUvPiNmhZQud5z0GV8DZ9KMMdtLJ52ZMV7axtbSxzuFk86kImT0U6OyhMl5qycbL3
Q+0MzWGbZIpSoTzzXnN51yBUUQNPMYFjhDj2v2S56uwZQL76kta0cdV58c/hHUSUlWr0SMiukrDL
CwSn03qNf5f4d97YjPu9VXxHFzr34sA41z7YgoU4W+9thYUc3skkwVzdgyU8eCOnmWP3YsO41YDY
bJG+vNuqKNLxM2vxkUV9CTFwH+pnE5xAFAEfcNmnvwDp6iHr1+dvCIsmTSoIp/DAQfR4Znz3sga7
xBapmO22ZoNmeUm3tUsZfcJU8pjff0/Ka7b0mzW99kDQJCuvJg4d56u7wjdkWfIrlKXt8GbsRQgk
wFpj88cCoufzPaB2iZnw71X2QcxXyDLSFKkM6iBDxAcGVmB2c2SP6upMNqX5EysafZbMfVEDMO3w
3O8Bw44kQTAE3aztpn4aBRtmUWj0l3QuECvt5hgl3A1HBY7GldMRxJceTOrYtxxGWthHaBBRAxgq
zxrtITdxAlYep+V144OWIDomK9WaehshiTLTRfeP/c0NyJfHJeA7Ss96Jtpl0Q+d30ez6uwtuahM
+JK22ebszbougkY/KtA+bSsOI7I+YwG27HDtNlyTTmOPn4uvWpuB0iH964RN6yv0i1Rm769h/eLX
jmUnBVgz+WDtloA1+ICy4ogG8DYQxg79g9SllbL4942llmIsHmdFtLq4LKPVXAUpQCUKhr3KbJge
Uy6xnsOwldZ6+Eu6dDUSitGXm7rPrf3GTR5XwSetq+CdZXAP3SBZuK62S3/8zc8wUg+1IkXac6HK
0V3jR2w0kZ3YxcrqcBHCxgD7qtC+tEsslevs6+2tfgMX5jUHeF5OCv4UYadeZM3YiGZ4k8xuI8P3
30PUVEkdYYTbFFrP0VlurrRl9JI8wMs+yt3iTl+EZousbDBFeOD7AGl9jARffgjNl1oqoKChPNgq
bRIjRrofbbwkvy8VtY5uUi+YsHCPiRqRfWv7wt+KHN81Phyqdit02va+TceASRy0aq0kpCwp+BaR
mXDdg0JV0YZ05IVKyA9R5I7NqrupLv3NtraKuxlq5eeYaDFiCiTQti8xMyssYfNINVugKeD+9+H2
NLynQ6PfPHF7Ib1lj/lCsGIu2xZJgt6tq68FxECwrFhBm6BYbUL85eS3JdvuZpBVqeDkfpQBS+Eo
mdn3+XFYvLTBzW5UAPbtSKRd2UFm6vqblK03f8v3OiU2DPfD4xxzm4poNVj/X1YGLCdKbu20/0Vq
nMbl8ZhardqGN/aaXScLkkAOHiDtOJ5ovAZSh2xPXFfOOWYrNOq+QHjuZ21nBc5iFcMK6ePAou4c
yBZuEBDMS1WJlujxDGgJPGHynSWkNEs/wLsEoUo+8V6MEDNWhSmW8puPBPH4fosoyqhcFCohY+rb
1t3XJevwww7EyhXN3Ilav/rMKJlnZpqWB82XBwnnxeNR82QkZLXvaXQp37R2kk36yq0JPZhE05i8
9yrjHhWM6506mcLNXrNwR/n8QysGxSmWZBCtij7yxrS4cIRChOu0cp4I+g+ArlXXZrkiReWZ4KGv
R0jIjavbVokN2riOXFkXsazmZIfUBZ1NSQBgZY38JSa+GeWxOZMxCRsUC3ABVtFHuJx4P7QjoKw/
oQYka8N15fFrhagnpmXMioIXFnsDYdVfHhIXs7HTZYZ3hTT7b53BVYkG+qy3KO0oI7Jp8DBSsWgX
52IuBnyydxTbF3mXaM5hj+xhRFlryOEUxD/ITdj9+uuZFf4q6FMB34a7FcL3x55MUOijFPI46e4R
q7TLK+StAfXAoS1Q0AzBi+ybAHWylozEa67PHwEF9NFpmNXpnz2bY7nnC2KEg0MDUuy0Zbwera6F
sc9x4kw0KzJzFUfpzFMOmqWpLBoKuYVdIO3XU1RAxH6yG5/HlLoWFf9AnwFuMyKrEheFKlfax4cC
RzpFgQZr+MBJMQgiLhr1pIzAENJawhUVRKIUhnIDRVRxkcUcVC2Rhm+GhnZMcAb/cAzNlWccmlg5
mEIlklWJ2uFITGw6RP+V/aPmXProbJ5d83GoSnJfbfvt8675BN/gYWgQjlTuMB9wqCtEReAT4+Yb
WtIEfv0FMBLSWlGkndhwLvJASJ4wdjZ5Ax7vvk0Arb1uHc15vk8xssrKpsp2gw5mil38yuij9F57
Z9+HFV6iJp62f4NLfR7UpvPJiTAJamqrbm6kh091tdY2lm9qI+Q3T7XcPMTMwn7/Xh9jvSVkuUyl
SyL3o8VnYKM0+pm+pBpQhYAz748QAcN9wHjUeE7dt9nhMqC77ouB1Zxr0rTXPOukTb5I0SkLicPJ
nSQbLtgeIPCGhJDzyGXT+45y7lEvtuA/VTzT2IGUtdOoP8hbmLmt2ApDYi7W2vpb2wPctXp/tKwF
X5Dg4q4Nc9Xqs61iPdHOHllouHKiNVfEM2gThtZLf/zrTX5q+uChDTeqhpw/Wy6SO9Eg+nKCTkX6
2UJYYJ8lBiIp6idp8gFuNxJPx7eFY7Osjm7zSkQivNBfzufYwWcxOp+nJU1aGrQrMgYE1heNwhLN
UnnJRqe0fP/iNqjZJjG4BLyacTZQqvTowVrRGdwB/isxvR9xfjpmEz19pp32uy6gRyuZTOmUwoJt
kmm04zz2UU24NwBnyWucOMwzTspoS4HVswbfxa2T8KcRjTbZf6IdLlCNhAEFsfOkfDK5W7HclWtb
JsLtsT/d0BxmV60BCkzKIVwRxN5H+HhIKxDopfb5NK03PivtgrMYDoZBHBR7udAt7UQVsvhXGneh
aEyxLq9De1f4PlzcTFNHDJAgPe/QCmhzutkrL6qCedz4EeOWun991LiGbkWTFJc4kMY7dMYGM2yf
UxOzxLWy5nKg30kEMryg5x32QajJlh842Z+Wk6CUc80SyFKLdI0Qxc6pX9VQr4oQQIHfOYLRB/gp
FToHZLHALFQKJeJAdgqaPUQo4ucMX9yfhuE1z/wDaPZBaTfXywGiUyLatmdOunT4mnp7KAHalgKN
w3ITYXEvwPspbvI0+CFeM4xh0jrfvYi/zGc7Fq9EtEOXc0sWqSDs7cdXxkXyJdafwZA+6G1u9gm2
UE3e/P5URQNXYf6NIUASx0fcC2ouDTWc2TbgZC3O02kjPc4A4sdi4zmS8dKUdi+yfEuzsX8icstW
j9dK4kmArzDbxA8opr+MjV4VNyQ5U6mC5QBAUj3JEH/HJEmO2udFTpFKao3gMCnfhvrgnB/5spJM
bRKCM5b0q4eGbW1Mom0iok241NwmCqfoqahUzAaCnz+1BXtBCYf64lF037nLRRW8bFjh+aY0G2xY
OdLP9Ckoh6sRawQGjHV3BX594taEmjTUjkNIpf4aqoTiQWYKuBcJTC7scyjk8eoVJsm9Ut+KnxLy
s2on4YL6C4EwpGZ5iVoet/L4v+TPHPnuh0f5LXXv5ShHZUJ4axkUWE8JVvAtt6FyqI0ce68ikN2I
26wb8FJ/1xCEb8d0iuu1O8TYhE5c/OtNPqftJmaRJ6vrfGj+5RBqNTAz6SBYCRFXkxT3vrloi4Zi
kmNgHnp4BXhyE5e3JtKhs8r0ksm6+78Z1RXc9uibALt1isK0GdlUUnWJs/gazRvlYS42HinYqfjQ
imAV0FIErWTCoWVYzFGtohYB5QNO0tY40xmxaL3aT62NQPW/qd5m/+L/9d5i4D49s4yinyvvhmDu
4oJCopUysRiuZj55SW8tDdTqNg6d7ru6YPvmgGfyK9YyX8rxhBYc795w5n8SzGKRr/q2lC7LU9eX
eiP3lNy8u8bxCDMQxoirLMmONCnL40MpSvKqqUncirkVdJcgi6De7w2h3TawoZhVJOLV3JDszEm5
WwrYsNuBo2P9MZ65IKwRULr0OgIy4trtllIt5+3wvKtR37FDUTJoh2WpHngxcZjl6us/N/Pntvtx
dOfCwkIourlqvW5sTqJ1DnOf2Uep5o6qtU7bpTKkUQpv22s7f9Y0aZZpSn0p5b8hxc2ntA1MIo2+
FepALuzCVC7mB6iuC3WHaMVKXJ8Npt8uyEaomGDRvfEqilDawSXqICMzmY2OdKAZWqwKpQEEO7Oo
4heCpMO7HdebtSBxAubWMLhxZC/oxE90gSBENJRi71yIZj14M5f3GW54yQzuUAmcdE5cJQUg6h/W
bb83WDl7t6RL2Gjl6ZXpTc/STtdGBOnf6vSFddgQmttpUJAxrYGaxnGVp+OCR0SCkT1KKpsV6IKK
HfTds8Mp348AFmBadF4zSZjKwIa00JtReWqJ9ZFZR5uzvWeR7OGDWL2iXko6ngSFrO5kuWb8r8AM
8Ac9ktirCyt+kXvj7YU0xOkm8WK2MMLh8Arfr+7rH5bxxHkyE14DnIlD6jSZa3qttQdT9dRCVBMi
FrebOhqDgW9WUJJ8ulsI3Tf616CaobPQ4KN6pbmXArmV3+7FK5QqiMm83GBrB/Eijo5Nxcn2vinc
koe3Aa8tDApSO6iV4470dvcst1nwl2sdbLRn3c3riQSeXn0h1ZkJsxvBX68SMR0unCz3gZgy9z95
46PqZxfCguLFkUgXleaa36v9Z9ji836y2kUzFAKQ2xKKbpchoaqrBEdUXQtMtMvfNRp84gDDBCHg
I9kzQNpKHQBV0noVGj3KfXKlWgN0LY4P4c6yM6MMrDYPbVf9QWUtFW9bJaLITnkHJWFKjWdiooNW
8cM+Go63UvGnOcOEeyW/fSwPMYvgDyoP5sXwUSFpKqOuzUoeOlwAa8NzNPlySKGq4zyu2EZLP9QZ
NaIIqY/t6EBu8BmbvxGhhLIGfXsuDeadBuP14hR8MLUJzt9TCNkg1MaODSxU3tI2XSUJXbjMURzO
IJJVxG29f9eOxAWV1IqaXQl2qssihkNUnDkeaumbW0Ozd2OvKcQHPnYdpxh/6C3cJHRrjpkkpefr
VbLNfwZQiETsruzowZpWMhgWD0PH6IsOWFynrh8BQssnxClPD4kr2RaEPjdHJMIWu0o5z4QOO+w1
an0ZN6dnCeAXFo+BZ3f6vbvDtvLeXRdnFLPwTFzHOv+lXupLE1q6U2yC5t7HYv0yChQQFGLBqFee
lrTJzyfid62FpNIJDs+Vsh3Nii6DyxAcSY3GroNJdrQKhK8hwlB4UCHzLd3AAR/oT6GNSnxF7Nvx
ekIMvZ1q+hXZM4DeLdRttrtBYCfDnNMriQ03JfGZ5+sHbOf0+eZcqAaguVhnOH+AHtBe90sMfJQN
WEkNYt+H36tfwBMrRDWoT61KVfVylJVMUFg4k5Kp39T7HoEjx04nltBp/dI8fzgNX5wEm3njeeKf
jAbXoashhzCI7L/q8XQceIBGphOxnJCntWBbggm6jhNsgb+Iv9AYdF/nfBeoEzZtP6c+hKpjf+d3
nEzRBDL/q0264NHyZ3SJZtfTL0WI5CX8yPoyTXlMGLeTdsfIiPzxAZsThSacZdAk14zfah//jk4N
irNgnhGFi9dC0fZtOgVeGx4UuPtv2qVHg1gcE2QEGGPJDFTbiaTWxQ8e3MfqbmnzB5ku2BlCXgVT
ghPUO2ETWbb2prhOj3QJk9s+njX9hVkrW9nM3N5fMMz5v7qDPbzZczyqq4FNBmNysrMUFHEzvQbf
PD2mTi3OxchOhetMdeigE0FrZgQvGUOB70XirWykefSPvXHBjQ3WC2aMduIavVsWXSfS+V1O2zgQ
NIOnplUtBO09sot5meUHdTNc7vX1AkCyYOtn/fSM8Xamz5EO7D6b8EKV/9FQFO7mBUAauB26Mfay
+8Y0fab0BOw/Od7GlljKCoXQn8kLWQhR1oA8UqrqRUHc0a0fWjJCSiHtgCUIIymaoLnwN6I/16np
hWAoenC5Pqh/rvh27WRI7gxWZPUZVwL4LlLYfh/L5KNgZWip18ieA2BuHBl9NtwxVT9Vz80drDeT
ZC7qEUq/Vs4LUHjCvibE9uperC6h1y9vCIvvKAMAukpbd4RAy4vDQd8utNT1h4L+zLdAL/Nre+fG
/69+2pt/STYeoF3Fh/Ht2g2L77akl/a7JaK0TEbAJSogbuPSLeTSWyXMuRKTi5py8W0QkB0HsfdU
mfHeVLRCbO9kdS1qjlgjj0sZmjCc2H/3JSsfsIHIMVQcKif1USAvWaVoORxvDm/9xbME/FcwmMny
qfKrft6YUQOPYJUGV7Jx64aaam06WxHfIhLaGR9DV4iyE98FvdEldgSEqVs1cfGlRDml7p7jd+JZ
T3479AQ1/01AFdZV0UWpsclAlRM8Z+V2w+YJzyl1U2sJyTxfc9hq34bCY1ohQ/naA9e0zgqYaxsE
useN56jzd5PEJpS0zGU0fuV2KfN5Mhi2Y17pc5oeesGc3prjvEJmeV7Tl0pw0Vx7kqoqWDj1M28l
oM4azL3NoMuZgoEnG701spEGSrwhLJh4phOFZ3yv+IiRTC/3Si7RxMTsJBsPHkAGmMENc8+R593H
cIKuHeR6UNe/sPA8AZPVduoffSB0kmfnaaAHJZsW3o0EJqEkBhDVPDa840aH/vVCOgKi5HgVGJbN
tvGbgu4N1Ly6vomQ91O12Qb41sxjaEo+AoOEvFQT73H0Be++rKxAaagtpU4D3wzUvmLrF0hugviP
ESc9nmrAJdMYBXEIozQ8oukyUeXXF6QBqJYomGU4fbs5Jqvfef2zl7uQYyv2vcIhq0DAzv1vbY+d
wCbmUrY3Xf9/UQNGwjmv157sOJJ1AX+JYoow3oFNuUhgvOR5cD9mL3xKKZ7OwaWYdT1RIAdsqPDr
NlReyztR2EXIPWNIOtLBqe6uBF5P8bgfr+aGQdg8SKdvR4u3mkWx4o6giM/5WTn8yW2vVfUCcS9D
OVjXRIG0GbETYEsQVOOflIyshjlDVzdOgn9EWMupu8NV+UxzlLDK8TSDNk2SknzbXpQQpI3DKRB4
S3J+m5wvIrTpopggxH+5gYdVECWlIESuvaFFXYlDOkbjkUloIOippL8UZVveqMcWgh40PuVhZiPF
nRaIU7L0xvB662wlcYEatNt+S+pJhQGU1ziUAPRhceg4POj60ISwubE6yiWTsneAfWSeTiX7o1cT
UbQVwRtB3ZUUTzH4/Tgs2PItHqBsRVd5mqV1EYvDMsWnKq6fy7Rpt8ofoA7mtjCCXXFnl08NdaWK
vEV/q/wGfSFdLl7dfLpJ4VZ6xCrK4FTn8gSs5g1z7jR6Ge3emqn8ipEA+xaS0e3aCAJWBS1hXd/q
ZOb5p2wShVtCXps74BxZNkbi2zXBIRqna5JIobR6C9+MYa3jp3JQeHcCv3ojRd7YTcjouubRvmcd
6UJVL0cOyu/lw2oU/rbl1uQnLJSmaJvo+k1wvsOmt1eaZMHjXUfU0nqfAj971Ynb5M+uTldUHGZL
Mzph5btOft3J/RdWYRc3GZSPzEoTU0HrZLlg30iAV95ZMk+XkQmbXv0OISr23BCgXNU0tOa8Ws22
0nSWUVsVOauKGNka+pKxrotvIp22kBk/fhDJnFb/eNwlwCqtcxkk6wSgXzZIGWG5uD+z0g1GsVDF
P01jQHDIEtmX0JWuuRHkF5CAiEXMa5XE8xeBdt+CVpnBhptNKCeD8FtTbzb1SF5rSFPPgHIBQo1K
ayhFNzrWcPb4vJccQgDEJBMVe7cIzz/St4KWTUN77nkxvHini0x0aHZzs1ydXDnZRz9Ts/ZtH9h8
uXLms4DNm7fdDqB1eYPI53ZmMX/yKjy4/Ieacy1wi+aEJmulp+mHjSQUqNEWbIqorJZe3+2KXJlw
yNNKK++66Vj6bIzFrj7RCCPpmaBRXg18hYaCbxhNgfHPTEbImqotxSI2LtRro4u42qklZpL7ZsJ8
8vAOqhRYHcBfMmkL7As5qVbRnkDYO43H6pR0Yt7Mg6Rj4EHyJC3ilKLdYkJnfjKSbREsLMPGlJzL
Pq8CBvLeihKo4DrLnxvgqdkdpFjjYAAcrPc63E/cAcBdTRJyeyUY0zUDaEtdr303M/b+GbBA/Guh
Dvkoq/VaLyah5/TA7bO8qWO2/dJ8m2mBCuJlPURkiExuRPTSTNqbUKMJ4dHRZcDp0hxbnYEvVjR3
Dk3wrpcIqThCQwl5wNSJ4tNOYh1zDt0WOCUKO1ddnfdVQ8aO1jXBKS69BukYTVO7Oo2ASUOmEpBp
dOyYmF6Ruw3MLRBuwh3KKw+0mkBjPxw/vAVwPWHn3xY14k7IKU5IdJzBnPgJ+skW6u4GSXNCBv1p
/nowC0C3Trc8qng91eU7DcjStSnKV5wG+Oop3qg7m1dNgiztcDb71AGn0DhzRRWDmo3TNB2+RqH1
RgsAPNS5jnboD6utb56WCamxEhRH9sNFpnlXJtlGCi/jL03L87Fk1piwcTb7hWRIgvyQxyxQN9fU
Vd7ZznnTFH5k9wyl2eWgttsPXVqJaLcvEL4fExamjMoFLmglt6u6ZlGmEJDzrYBplY6HKi6IfmIL
1ufSO/hb0QMi15hNqzJzt2m4kLWbxVOcr1vdZfA/+2AN1ByX/XU4yqBiRxHK4PaOLVGtH1YcKE2j
cswwraDWntzODACDsAFL4yyBByXqEx8+ekUiVSPk5/NIONKIDGTDFV7Cq3y4Wh4mIXbBk3Rci1ps
KRzjqRzo840pSouKU7pNU8+Cv5dZfyiZE8aETZsv7oH5b7AJkls4j/WKtNeM7K7dq4ipnHBEOTzB
YlpJ/2CPKFgUd+wyiw7yCUBNxuGJnQT9IhNAwIbih5N4/vptf31VlxjeNgVvrsIYHg+rHqkLl8QY
4nD++0d7P+PCNGYbFYdWl9IAmB1rXuzYoSLYok2hpEyp9KWrKDHM8WZR1PIKIcqKGCN4ZN8CB6Gl
WJz+YIrBcBJ4GMVPIoDGBXOCPQAo5xmrGvQ962+JlnHtED0qa3PjQI9NdEEMc3muuDy+Q1UFa/Jq
0K9KPmErhTY/9ljm3QzJLEYjtlPAvVPjk8grxDerZP01rr+W7v6qCz+iNpvNBRcTMYOW/Gf+CYVK
K4anVqTqDmbJOFA2qEpUroBFsmw0z7i0tW6IQi4wwQMRb586AbJKo3JMBaLPZV402fDwmahbpikl
G2dEXcm9OU5962RKatjgdhrLrRqieA4Sq367j68tQhR/h1cKqeDhj5AAk9hJMQVoBbMDkJfHo9aF
bjJNZ+sNlwtxKDXPD6qVhKxFYfpQPV2jeenhx0TX11qIgW7F1QlUpooXHklnZ9OfqrlnFbF/ksFX
lD6YXyFTsoDursh+NEsbOb6E0fWkwYu2cd6FrvL33pFDGaqo2hacNgs3HA8cH42+lSX2zLOIxCVA
77KnZ9eLTq8ZqHGGkP9+qk4v1vZDiJT4imJxGXNVHWPdRNPCAYmTQ36b/SSvDwkYzArS7ucnTfEp
1iMe6CyJo0S5y45T16e17YyXx+rRqaaO9Ery/EnhmO2+fE3gNpYfc1yucGX3wqHwCOpgdRroOY1P
CKe6BIi0n3Ndo5CQiSDHuOh+D3u0xAd8Vk9mCWtwxthBnzczsC6epGEkB+/9y9nsLdEOnOH7eO0Q
Rn7TFkhn3kaWl9Pzfjmg/JFG2l5+5AE0EuRlkzzgTrEZzPPK0SPP5CWpUnaQEQ0zyo54zfTOpDWY
VZa1iHL7i+aZlqHBw9d1P1qSrjv6Zjjn6T5CZyt3U+qSu8zxB0Loj+L9Sl07MgC0xUHaBzuAXrjw
Mi7/nH0v+DngIto8JXl9W/HG29yuZW5c468ORvcL54u+Aj9on3Y7EA1ZuEUytAlFktvh9r7gDU6K
futgCUC2Llqo5TvJ/eZRIxS+yjZ3+af2Um0vE0kSJu7gEneU+Q+aT/MYfvFD+71lxyPm1YWknO3a
ni/SajnjTF+UcGtTP2CZ68nNMytr5UTr74lLfByogG2kA1Dnp4bE2P07AChiaxxx7O9toLn/HrH/
P22eVNtJjqOgR/3MwO07U/qR+e96armk/EKdC9v72+hlrJtl3FZwE8zTA1gQBfcoe8KuOzZJXGr5
12qgRjR/CliUWAxhaxIVKsPf6ABSfwv2iMRM9WH/5I9QGa4fwDDPzRMwgx9IaXbINBherj4Scej+
O6YWCUZlTCuXT+A8W4w4ssmczTvsuQNXCnk/k5kuGT07e2ZqD+OCC3pmXl9DBhNbgv2OcsvQc3mM
sXG10QwJ2HV6XPF45+JCr6zfUN1R5vIeVzO8z+/Cz7U3kRs0pQxzx7BM7ro/G6gL3uG8CGINTzuV
pwMEXUHHcgAuHAkmzLUY0VxCDLx0TX7f77wLiI20LsGgHDBsEFdOowCHfa9hM+/pmRfb5u72jWO9
vKCZ7nrDN9OFTXmYVBaILpCU/s5bRLfxjGxjoqsceT7wHmQvV9oPqBr1Rd/GBDaSKadLfC4H5DE7
k2MxqtBZe1JvAQXAqh+jiG8EoYumVCSTNbi3YXWlyCMlZohn42+pM7VY5po/+wQiOKTswmuISvV7
jkEdvCY2sW/5NGMrNLZbiuZR05S9oKfCNomxoD/9A+LUZ5dgqEXEaIT9vNT9CTQZj5V6Lx8LzjK1
Jnss887rcY2/Baq7d8PV3gMVXVLyYiUuJahC4kn7mj2uKZAYVnyoCytmMVrDpkaiHtM8l/vwJqup
4dHPQFHm7NhV6aJoo0epEfoIhLKVEh6N/B6xTl4sehTfn8r1SO1u9vLAuSSigbCr019Vw9O5/raZ
P/Qmoux76wLonE+jWuJ2OVS+2G98A4xC1y5G9IMDFYb7fGDa9mw9olmm9/JXJhcM855JnSf8xYsP
GZGFBLeqaX090Dn4P+ZUy9RXCbnpxSXtbBGj15tSDnmx2LsbGuLUxA1ORD3a53/I5RMqOR/+KyJ/
s2+xx6pmpeQDPzTcwclG6vtOozdbK/VeSUxKrXL8tZYXyTIiYtDidb1sAGgjXUhhZIafcFT///ZT
SCsJ6S5c/IXYyp8hkj7f+IgcjaHdGvoP+KVo8RPnkKtuMMtvIeJWeKgU5g45Jlrjx5lQ0WOwr1dI
Lgln2PhZ6Kq9aGAqrsiaKfDjaQpGwBLTCRhb5Q2o/NWCCj9nMz1cbYx7nOUElTlMipca17r+fLTP
wBTi0YbLnEB0w6iF9EFVwJJyPv8hVd/b6AvG3Xbl9AWspr8smX55bHlvt0sR52nxcPveUOwtWKRi
w1tm7TRq8gZdIxr8F5haUSrfRXWRxEtGLLzSbMSgGdLbafmvw2bgY/D7G1M6YqzAso1idjhBQxet
fwwxC8TgAbaAcBRYzg83dSX5N5eAYgAvofDkYcZ9vt1vpqKT8FF5JOfmV2uF+H6Iw+FvINhxgW/M
0CLRJdin/nw9nO0ZUVIZ15xW/lSSjpBZILMzS4SvQP9yswsaHhfdwJz5uWJJ9jk47uqRUSUOiDoc
amoIK5jt6Bh+P3gS7XJDQLKWwEeOCDMciStIgzTdeNM0f+evTa6aW9U/sdSZ8Cm5YqMTJsNK+6ip
t2rmvUS09IptpaJVubhrZzGM6kO0+QJAyZnJMdZvs4rp0SlJjaz2raKp7rKenwVTey3MyTn0NFM+
1XrTNeX/TLxVN5Nm3iBnZ5TYlFPKdNin/fdjzhYUAqAzpApyWzYhGwHzPtoQpP1CKaIdu45J9m39
26/E+YUv/bncM1ZahBPTW923TgPSw/EuPksWbvnD1jQTRj/cLaPwLact9fu00VRwaI+Ff6nV2YzL
HrbTQXu04XhDQIIv+6yycn1xsmMlnb5CtjCBKrB4+yXyIbAwm0WEjbIPzaa8nzoR99GyTxxIvW2r
j5XKeAugZKz/0zmh1d+opNYiTjE2gGse4UMZhnxjgzpyIZFQ+Uuh1zccW1rTQVRBUGdf5FrDRi0C
4NeQ8cdxCmsDbAXJ1+FKaRTC4t83HjEbDM8RkXXiWXqHGhC6HAcjR81RR7j0SnrhJRiIkutHAeB6
stgvsqWo54vMCUqcVlNUPI72sVJ7kU1hAi8rQArF0DrpKshyrc3ufuu02pQkz5gCCoxJ05g9UM3y
VSqWofvznZl0bfccYboaxCIOcDD2TFpSA22g3N+PXid2GkrDJMJi4QnqhDRcZc4e0gOfEJvYIxgD
Fl6INKZGAssTN8eGJphQwcivvt2akwEK6c7iz3l6xIxH5DwYX+exOl93yM8UvQ67WarWfV4GM1Ks
0o5+EbOu/Gih/ZqSqwQJNFNOQrUo6fBlGTKOVy5q/GNKePUDzQjWZj1e2I30OO4QsNcHwR6OBZw7
8KY+TssLu+UFcoFNTYt0D8+YE2whJ81N5nFV+3pS/BCxmqGH8gY0RdxZEb+4aPFZukmjdayhhVFg
xxfjOSecQDeNonTHlNYmQUL8kCUIMsOx55pQGsVv87I2Rg0z3/h15STiOcTbTw6I/Q3/QzuCwuGs
IaJJ1nWQ+E9ZroizUyAataV+Q+0xiU9TvHj6nzCAzNzIlYbI3EG6lhCeZmU7M0zAe0Xfnkya8NJX
JTNnrOhlTHUgROigsChFesEOx6VsQaZOXSueSl6Feh3piEsDlt0ga781daPR2FT+TD9t5x6h1t5b
Whjc8rz9APqp+Qnwacw1/5CctD0JNMoAAx0pPOjrMGvjJro7NlxoB4pXbW6mjr+71DsXknhvfCHr
RRUf6M2zfc27J0G38/tNGvHMMLX36dI1pfEb0hUvQeQEeh0Gvv6Rq4WTWk5qNjz/T/pyXBUZBvym
qpmvjK25mEkzfMGOCcKs8Fiw7gZ0FutB4aLmf+NTcHTZ4HOTYaGKk3gSBabH1f6ulVt1rNbfeaLZ
sNWINFk/xstYbsZmjezGK2U2d3ImjfiOzXM6BaQCU+1R/coXS3Q7KyoK5I6l9p5RJ0F2MKBLv4+I
AEMcsA4HfV9CY1ooDCQADlhjOL6syiNG/rR1DWpsyZnyJj9lND46lnRGOo9A21XcKj5jNI2M+fpX
7+XRhOdAzh5yPlI0h9TsrJ5xQ9LwQuhewm/xg2rr4SJwWSuTWyma0B2I084avtcWTba6+IXAEFjD
1/wj0tWW/ZN3uMGJXFDy1ZqkbNU3cfsLjA17dugF+Zs6xYo6vSPXBKIO5ZW5XLMsDIiFb1gA4DUD
Gbuj4c8fdyZ7LWvTGqizV6lmwRlAgQ3MoKUg2BGjfXDHvWqsY/7YaW27QE/f02ai0rTRbp+KlEA5
Bp2P0gNG4qanEikxkyX2ogJV1fnwlObaBfy8hTpg8I96d0a8QquiTH91+bGDxB+W4iXav4ZtHc5w
laSe1l9NpccwQqiD8cO+k2kThUAdkxyeexuZ8mdXYKwCNMqGQbBTaKk3uAYxAz9yrj/k/fdBdXB9
Hb9ctpPrMoWMkCyA6gcOnkOKYBXZ/uieySaHJf2RQ+T+xgf2UCFGV1iMK1lNKfWNrD6flIUeOjrL
zV59mRICxkPfPinX3ruqag2TKc4B2FlzBc0RPZpsTZTBXjSNihCm3+aDL1gfD+iFkyvNeCfu5ueH
/EkxuGv4s+crLJMePcqhUYYZUx+nhcxfNAaPKiho2nTGq9jV5aZ/nfJNJ7wBTYjUJbNGeS2yETuU
w2OJXotw+KLMg9ZEwm6jFVhsMOrmqlq8x6oEhFd+BN2v3ybkx7U/d2L0vJnF0m631uEnGgSgBvub
L5+cn2jIncOx4lvH5WlQYjUf1dCP9IV066XOa4xPlIng0WQ5Ei10SmTKiaPG9vT3fm0jFiIh6LXw
ZtJwrIE8tEk9FQLzI8p4ZTUHLUDtjYFlT8oPPa0+QTvnBfI0ZkCT4WxwWpubPCAVAhAqHu/UKiUL
41N8bVUh+TUxNeTk5Nw3R7XEdcL+P2jaJUwrPnY46zeNMweTUmar5/DHYn1Psa/VedCNjpNFtVZg
xN/kvTx5QOh2IrPyqIjRPqQVRcOMnBxdQncwH7STIyLsFBbs9+Wt2VVbzRqRH9AO2VSpil2nQmVf
eoOZ8bYAG+o4xytKM7Ck+QRULh2lDfoBCGsqhe9GpxJPTyX5/HkcxG7ORkzn79eTuBE0Wzs7w4Je
pzm39J2nK3fpxkge988/3Ce03bQbBbG6BSMJT5l8F6keWSMD5lSZqN+ik1QO6pBBsEEXxOawtq1X
tGudbV6qjqyJRMi/wbYw9QmGUsb84u0sFdh4vvDPKA5jYPBQmQKav5uPUXd2A38ort61M0UAm+CT
tI1Za7V0+TQ4aC0Kf1fxWJrTVVG5unIOcXY1rzSL6biG+xyPc5Pkg57qP6SH/6JuNY5Pt9bOzD7+
wDDc6Krc4uC7FXvgwNzCK3eGhOTmGPfoY8ewp7rmwZOU4Cb3BkCJGbihahHQy9vzJdrUK1TYZgnz
hJl9af5YkOzhViO5Q8nikYkSWZdB8Fl9KpyiyfIHPys9zVQ0wRU/OIhtLib2ygCC0Kit9Um97iGH
MgyxE1SED/DXGIMipcZ559j18YaNX62xNuKFM2Z9Dteq/LfxXArv3gJzv7tLLsNqBZ401d4Ld/dp
zq6GVqu6ubpTXIw4/yXU1TpXbf6QOeWDFKR2HRYHUQiV4uOvhVLzNUayJl4A2E/88yhd2W2Dhm24
b9y5MbkWTWnUE3ob50SP7YuNmPYIn96yYXk1tyLrIMq+Oj9XFTyHR2SI4s9EfDrnGRi1jc8QUC8x
oybAWpT4Kv4j0TcSqInNes0Oib+7ZcUU+NwVvsHEn0wMilO7PT/HXN2mT+QYaCLzH1X/rhratcI/
Iz3XzlndseNKOq3+VwvUNziOZgU8kbuy39pkrMifDKimlTda12BAgL8Ew+zT0ut8j6gcG1U1U+7m
yBrmyFWJgRkl5Scte3pr3YA9dlJ0rL3LIqpKp3VL/8AZU1HGTNg/V+JG8piDHa8++2Mr72gQg53g
FYqX1zba5LMeQ5L6XGCOaY2QtflcTraUgmEL6/O6ZtAem2K2cYxTZeSLJsq61OjjwCuGjYImAaUL
0CFg8Ik5qbi9rF5u6K6Fn+D8hk0VWHAABNiwYsjQ0E88hzQ3KkncNOfyQsM8vegn2ZTpQuXyBCoi
dUKBG0IsTXMRgNMNBvdHjpcMcLlOlVHff92YcleUYupuQhNtHvGqrRQc6Oc5AQp/EzgAyn6GpkYF
pBX62dONwnDLYA/cC36dERYbK8q0kxU7AUvljWA65zhBPni6LiHvJA8Q7jRru2qXwbS4/EvggpJt
wyTRP4gtlwT/U68BJ1CQvjzZFQAIOAUMdSYf1u5u5GBelYEsVDgzMNLbEr6UQCF2XGrKRcOt/rTS
8ToS0JY+exWXca0WUilp5xhOymnocZFr6wc31JKMM9R69+kIqBgZi3FSLq2/LXaQ4kq27XObOnm3
vfx4B674jQjzmps/quZb7h7qfhqCoXeqrO9NHX7lfK4GZJ75XTgEyPceBD4SNEtjL9DflnrS+SjT
NdaqJr62+e8NbET8wRmDXJB5iIXPBp/M082bVH2i19zCaUeAxhB/8V8XvE8ugboJyEPglX6pzM5A
lJDn5I5sVJZd5ffauHcVVO6tOgMhZE84xE+Q49MVlinBFGV1GVJ0Ht/dmed1TMwKHaQznFrl5Ntr
F7wwvPiUqtMKA5CY9Gr02gHZ505acJclQQIvAHyrFhpOA9t4+r57WwN8fWukvdZLYYtMgoyuZAmG
njTctPGJ5B3jd76JtBg7N2B3PtP7AwMp9VelSy5Nhs22LQH66E5eT32dNJA3WWKMrgx0HyGWgPM3
UmSbeICDWN716K9BOAAP5xeJ7hzTpZ2ZpbIyGtH1sb/agG/cDtqXM2Y/8zk1PYWRsGOib8kKF+WH
65NK2uVBMeG8fJNG8eDbmeBofTZxdz5fixig1saeE61JOCquiTUs9hO+717hq3Qi96wMlRn5Wfn9
nlXDirSUWmKaZaaCYFSit7p/6xrGUZTQbQ02ULi4DKu7b6e1XpL8h2FF8rQ5aYfqrpZSZQGFMLfm
T62cResq2sdOJzF+zkvfq8axxRJY/nBehxcXhGZ+NEH3QDQ7EEsCP4df2La/9WuHRbcBLdU/ClYY
ePRiBuI7sdYnkgnUZ7yLYfmLCXB5oL9UX1QgSljlprFAT1/ooAOKI0VdH7yvtJcEkuQIleaq9Twf
P+3vAc9msDqeBKoE/+BQAaSOXoaAU3zNEMonnxvxH8wXmmdmomK712xdjbuATebAI2nU5GpXU27v
hB6llf8DPv/UCIz3OMBXDrLQ07ZR2x6l1bNZ26BT29wM25mI3hzeUFmiZpaDChv/rUfGw1ZbpO3p
TwGN/hzlzrD1YBZEgm9FPOC5FG/o6bKP6JpzGcxwKOXFj1vMSeCxbkmZRFyJoghB9kCFuzWajNuE
E5/pMBSqJ4ekOR0KRRoEHs6aM26XU+83d77sCmtSCS9upandNNWOQGUTP1Acu9JE8ASrfjZztf5s
K/XtT4dw5AuIPCvBMhbcYDRjMK/COR9ySm8CMEzhwgPjWOLO0B6byCNLzVEpGr41oG3Y08LwpSSg
9pyHV6MI0X09Sue4fRKlRrV+C8mJ+DAdlDrPpL2PpcUrPSqNeU9Ucx/QLBKKuF0XclanE1op0pc8
Lv6PMtV/GL2Si+HgxgkOWiy5aCcpdlyKriUzEiALsepwi/PVwrKULmuZXHGPmR+pnitfuJtJyY2H
Fz7evUgTaZcDYFMXvLpt2eHI6Y+lKGyOGpwQe3dYlihQCUC5yl6lKP+wawBZ0C+0n7f9MhW9JN8s
hR2s/BXdA0ZQ8Wz1w2wUb18OXRGoa+oNou0Bd9Azd2DL1UzM2IyyNBGQsZqeVWOmT2D3ilgL9Bql
phiF/zIEMT7Jx+gl6BbkIW4At1pWoaV5wUpNGpwGeSQ6tL/7WrXPnEabd238LTGr6ecosEAGq164
SBTKOKGUbZrVSYBwI/9BJebUaGcs0mL0Z4ayFyG/CimizvmRdbmeEBdWztBxOa3mPZeMr6NYOdwB
pLIsWCH9VczQATiVBMg7zNBISr12G6AaxueIAP+KLIWOghR/kyLyaY9tJgGCyy96zxJgQ2Ve/5M+
d3Dyjri9Ftg2wxblymEEcX+Pi6+i2RCjC3Mq2yv7rgBm6aIC7wRXTl/MWtpcrHoodxG7H5bF7Ilj
alpkF/DNRdvwiQH1OVw16DWg89QnQbCN02CUmozONHzrGjXH1EkSnCTQX+CR7PZFwUMRGVagFAZL
HA0ChpJ4NcAeVEcQcPn/Kk9lg4p23bOuIXNFZ7BUlIiKLNARHeOaGUyVD2BX83SzywTkxRXxgTit
NTORGlTTiwdquKdCy3AWtOY1Evf1g8vpZiV7OrZcRIN2irok15UJkZ8qQggOzFGp0GlUp7f7mmlQ
3ny7VDk+k0eelaGkmkRFYFFNpPL0ihDQSatQNIVOnxCl/Ui4u3jZscAyEd05prXpR3px8aQwNEY7
NvOQonOEiMu0792ieSQlfrEcP/fT8RLqVKZuZc9eUQgnos/76RgM/PwODU0WpugflSzPGF5c3SRF
NzZu2jXqDb2oKb8N7vxc2674sxIbZ9luZ54FQwZFQ/zrIN560SeujctM53GiZ6e2FHJI3NEJWXTM
gIXpJ08ypOYX1q1hW5AnNJDbCGQd4SRmRQNF0p+Voa5QP9a/2zggL7VTcXPEF2p6FiHwYPXKOHZG
75DG35m1kE4UcRSgvLHMIKRvVQ3LHiBg6MMCrLOeN4LMK/SrkYksUlXKxCSsRo/wPWCyYWGJXo04
uqEzwhx2QnwoXxtLugV5s1KKFIxEmUmwCY1jtEB8tYx8bYPaTlek02v4vxnZGkrci7geCPeNXzPc
vL3WSiXkt2GqBeYzBCAqVAw1Qjr/zFWAWkY5kI1KGbog1/FnKHKxXfWHnC61x2zU9SOKWWvyrk8n
w2sCWhugiUb7/tr1S58wPpF9tU2oS7qktBxUT16U+izmNLLf1zQ1GocC3HgYLoYV22MeYs/ILWKA
7pYnQnG9ywBXBREi8oAWhP2cm2HraajhyomSZX3ikbtHnOiv1sSFnMn10cNcZ2AnjLnwX/T4cV3i
53MUgPJY2TnTZM8uNALBV/6BCLmAXDgUFd48jYeWdlXDODuhjp+Z1f++WwY/ZBcWvjcOHUuWCrW+
q/pvJwKitCbthkI8YQ1U4hDet9Vcm4VRqoF+RdFhbkbLxwqv8hlBbkE4Ov0SJizaIgMfydZo0MCf
zkhYIaQQYksjYN64oCtgqLeW59DUJKPWttg/VlJ++zxaJk6nvBecWqk9UtZtoUi09zOLZAjaO5kF
EYTTl43/fej8wpQ6QkNw5kGEHPtrVWF6JpulkNlUjCk73vvtijgdt8dVBKCYwn9gqfMwo9ypHicP
MpqsdX+04hFhuEkvPR/SfLaWMTiRHgvGawrdtp1sb0fuV5beDJvEjEuKc9jfRzKZqDGXje/fl+KL
bF79g1JIMsYb16lh55PwneE69ekM932nRjLiBthlj7fycs0X/AabEPvouDvWM6UTlPa6dyKubyoo
+QfGBXqonOGjcz0zoPSarr/EOf5D06p1AlmIajjVbkbMKsoFbukqnDpXGO8kItZkRyWxWiNtr0ax
/sf2gART2Zt5NsBQEhcM8y/6lX/b3Gfx4nSg5Jby30vMPqh/ryf0PKazwJJrbair2U3E/iImBVmq
7QcLY+uRDYratYCUP7P7Lh5JohgX0qi22zBT7EaL1gf+HJQ5QxgBqjtuyLzFw3psNAbJcy48Kn1D
FEqLBl/r5h+ysEINnh++T3qtGb2AjXuVmwmtyAllDdnmp0yq1znf2znFabw1oh6mzG9p9CmY+vYF
jrtS1ctP1owypbNVAcNJoMxBIXWzBJpWEOBtt+Y0pfe0AcjW+FySZNCU+g36sI9XAsSOi6WwtFAx
HY3Nx3OobXD0BgpupGxNo8h0VwgN6J6W+MwntU4HQog1BGoXMXzv4sYRhdevB7DpXUKSW5OzIzJ2
tDPmbJ8Q/CDEE4BYpA3IJyFN+gze8yV0Gzxe94FeuhEObNzGTm4h7CUkfOoEeEB1xXoBaZpOJ/D4
y31rrOlSwxQMVvG8XHoV4CPHh856IXfqVuU0JwgJvVKONgyuWU8skCX/XB2ZO3kKqdBSBlxqliRn
04jtLRw0WxxqnFeF3AfcqQHjlvuDccflgxFdCUGb3/C1zvlQcdsPts0SUA/wlfqjJ2+lcJw4cywg
NluTJj/JPeaa/XRdmqD18g+E4qN4n2Q0UD31Ke1sXnb6sE7Ajunp9UOlcrOYx8v6HaQ/ou9fgh09
jS1CUjwpEWRhIIkkZor5KuMYpvHvq7mFwsndxvELv4rvE5uFnSZoXHXOJUEP2eZbvqvyhrUjGN/q
LltZjTURsUKEi3mDMYmLU+vsLfhO+HvsOxKkl3YAHVPAywc/jwKSv+4ggyPsmBUQ6sEF4ITNSowA
0QETLTzKc9UwHEYJy+il+7toUDXYWjk3JSqaYiJ0dEQNq0rayOBe8gUCLDtm4puD1Oh96XLSDk+I
K3P/g/y7uQYxIk6ifd0AlKqc7iQLm6DuyP95QIFsREtAbiFMO6LM06FWqTHZJOo5ZVThTmeAIqG/
r1UPPW6D6cED/qAVXnknBDZfg5/eTvKMeJ/6PidKvJH1g5DQkh81oiI+fZ50hQeaiLH+fTqzG44T
v0nqmNBxZmIEDctnsUgHVYP/RZuFeSkeW0NLHIv/oMfESmjiUWUZPRBPBPQeHzwNifmoSX/1GVV8
2+0DZGv1aGcg9oP+XPVymoWzlP6Er3IG3r89OxkG1jCUC5/+9kVCIPb+/+QIRv2168YBmMk5iukH
99VtNSGzT6XzgY6KPvAWbWE/tn8M8elM1IaOEoDXfQ9pWx0Ushlrc/Aew0ONGCDVLpp/oYknh4YF
RCxpvsECwifgwRNW/vg44RiyghV730F1oqn+nhAxW1IBPW1I29pAc2ctbZzEdtgkkig/I+w+m0lr
S0D8DBkz4z3nzHECHbaFIT4DIJWLy57ufGqTCY/8FJQE/b6RRBogfTMMB4S6BedgftcNENVDgoHW
n8LHy15kJcNFx4gDQbuCQd5vvOoiDr6Tq5/Jo4J7rhIwloTr/f21p3tOFftWcPbB79qDdiX2E7sl
G+t/GrqHOLzt6L4jay7Gvtqm3u9t4XYzcy329sAP1gGRLtytuIJvCNxje4ysaHmZ6E1M7o/vQaMR
Mp+TaaBN5X/HXuC2nThlLJQOQqj/j1CXXthBM3hEgVankOttXa6CyR6vE9i2JWBTMecFEdwB1sYX
dtNCc7RXSdBOwaQ/hqKmAwEjUuYxGjXnXGULAF/egoTEFaz9z5N1escKQMbwqGM9WuFZZcVuf7OB
rADzaCQeh+t+7gT/Ul7oHc6l5c+seG9EqTmyC8wvaDmcCPaxzO8W4bhna8SYMpnz8+4j8Zo6Zfy0
NYWqBQt0TEX5DcRgeDSeu0MprkQ0ijIx6VD9rfSY0gfZykck9aFzbr/4RMolXspWqJjWOjbomjLm
Yzow/O9PClWtsziRDc9P35b11bc4hneYEx0zdAmC1H57tz1GebtH236L5Nk+yjPCd+P3PdCEern3
0oCUof6Rgp6LkXjuP3towvtYzkuUHtIjlm9pmQ6R24EM5NEfL29lJrGidcE4oMSjXp+6jBJQnbqE
FHJz6yfDl/kZg3cNDq9MxktY4LmuiuOozKv46H2UJZeRYbQH0sfxL92wFG+AiHvpLo8ZEUPPj8GR
6FMnAnxIT6CvVXZr0okXWYwP6CfZqqhLS3lKIDOLwY7OUXG84i2+h9JSbsFgzIjGgGhzX6Neaa35
T23Iae1x6gTkUOpAyvSectwjT6HHg3Va6/wuaAjS3TJVCUUkY84FP9UxDXwEfISwfTLNnQ6k3AtW
ZTa1hbTkZkqRTqXTrJbHIYu3Wjix2KlwqubgD8X+UHGQ0qMhS7L2qeYj8fvkwLTbfWkjoWBPyUkg
Z0eGj5WndK8m6mG+pCXoC7STzsWRoCZb38ufKdTt4tHY/dbjRtSWfrPCzWN8drBROvQ2zSJI6h2N
ANBZxVWYyNf1BB6pgaFIhLRXoScHaOB09x0Z71W93IYIYumWomSqPpvo3hFPegvBEXV2Xs048E0O
5/TlnUn+tYiClHs59rNaMvUQ754zMxcruEm2vOzaWTGWf3zx+ayNwvnLQXBT2OKS1jzGJGK4Z92M
NlJBOl0rwYVxZScYUmG13itOiVyjRLZAlNJi2sgbBt98yPd6EIhNhEjR3sNApkykZKHMlWVs0iJW
s7BMlXf18n7Zogj5qP5TRvYVik6qnnKFygXQLmN38HKpVmsE1L3jV3Qku1vgfQii/Lbc5LpCNplb
UrNiKqTUmmsU7pfudJjYajoG0YWU3vfPoYUvPnzPVO7++sIUZLBeHxyiUnTlFTjZNl1Q9EU3bvV7
YwWLeFCjXc+m615+GRcLvQmYDw3NK986z+tn4AxuuIbxDCZOZFz8C7aMlbOsv7NZz18NYLqQQMV3
YuKem09uQS0sF4+2V0QkLUeD6aAzT5UYejG9pQpGbaxUdYz//WeDBLHp/8xb73Yfx7T82dKKhN0x
OfeIaUbi2RjWch0K27jXgXeH3gwgJF+th3ABtIZXuoKRhAHwFwhLMIcQ/VNjOQmeagkVZmQM/kaZ
IwurKzZIDHtX90ZES0U3PqS8lkGiDiPf3esGJP/BFySeCeXUV0STQX/yx36Xo2LGmuSiiYg35kOh
glBRyeshQJwqHK5jsq+zn9l0wRiUbeA2Twgwdk3LeE7oEIoCnw5B7c6LRf13qgj5sEnXNhjD+RXj
Epn+ndGBQwDw3rsl75ZsenmcEBkrziafuP+ok2qQ0S+9fJSThFsrJAaPpZfwl3Usb0OrsWdJfAxs
YMWHzxH8ly4pEOvgcy237CQACFcr4KOLImUt2u7+UzNbxzRp89D3Zc+p3pfvbh59IcWWtVUu3hip
y+KqPO9c1N7yHxprnr1F7jK0AlZpR8na2ooVa1WPx22jQuq+GweJDzl6AtMFoJqNMyezntERnRS/
dvLKxlrQzYiLJcxoFLo+1JiDeX0oSqyjLwHi73tm8ay1qbvuZADcxRViBzYyfwkkitWZdLERBfVg
lT/1yzUmYYEH/bH8b47RAeJqrOy8B1y04uwttwQLrx9ocjN3QQunTaVAQfbu4N+QVAGn79Zi1IRe
Q+vvgfZxtjNTZZQVpxuFfNom0LG8oS7ePjy0d9Y3Mz0TDWW9Gc3cvhMzWDxQ92krS6HEPXwmEavM
d5LDcYXrRjo950Vjirl0f68TCAZSAWMgMYdNLqfieOgItJwKscbiLmD89fwynbno8dE+wB2CGqnY
HIWJFXemwCM32p4zr+a93zv8fnFc7LT+6dIKl4dkq1XLgkzsvGlLFetTNvqenx+5nwEeq0cdK3He
MLIyd4tTOmzdBBjh0EVTP5/X9gZQq2OZwGbTx+JCIesVUahFhuhQ7/m3dbzwwroQE1KaV+pf/qpQ
EaBXPBzeqc/qCsZWs/RizUvl/unqn0EHjmPGSsWP6JMsjw6I5U5oQI7ZS3BDXlmHFOKrXHF4co/p
fDGPcL5mFh+04Ft6hkujOxzncHRF5yh7+yVfcK3r1QXGdsI3TvAAPAKprHmM6zpldEX09x6xjcw1
UEV9XGd1cqLeGuBuz3DbiYb72xLpex36XqQa6qfbqqTyOg0KBCrkCK2WgJGqrr8/wc+CSrx1J9PU
dtYe2R1mm6hZuGztjhfxQcbq2M5UF3l8lOVrRZQy9Q9nMEk9FD1Om2OCWP8Ajvqt328SAP2JTvWg
3KeIijilHTsz+B8a8WQoq3fs1fT7zgAqlz0Y49AUbHauuRZQEJLF/N3eLJN2SGqTnUun+IXfJRkY
rdENHNTkBwC71zRd6VY2RPx58OBAW0NQMqJ2pUexq8DobG0RS5mhz0ssWwkkAPHozl2ZIhSdPhr8
LoZTfPgnpUIJc1XQG3psv6yk7Ir0ljRJQXJ3Fn/piIwWtKzCbdMbsht/8TRPjV9EYtkK7n3w2VQf
nK1ZHcBmvKzvdxmyduoP2HmDMfXAoxDh+b+BIOQZsppasBtFJQe8nrV6HdzjVc90of24sEVrBowh
TaN7ru9rl3YJyR+Yj3wQIEJhfMU6Sfdm2Dgu4jFumZYdnvRvhqEukyzj9AyjWdus96gKmOHWFJLn
RhDph15WQFavApDyD06UcUP/qfZDTEviJyLxcSAbS38uwUuK0AQ4BcnQ0Vju7lbiGwv7ruQILEyo
Nrs1S4cOmpy9GJS3PYH39ednH+FmLaEPI3emxFacWDwNM01AoRpWJgZj1p36zCcEf7QEdvP6xi0u
AagAGu/DVoCL82lF0JnzeHMEwhI8jIjN78Ov+j2FhvVOGy5Bc6hVYSXqxEEHkIhLVhCN6f2k2KjI
j/QdR5EjYzg4GckaOkkgO376C3G/iuw2pguuIZJbuk0maJj4V9nVqrA6W1feaNAvfFx7gQz8k+mj
2cqVoyXmvPwm+Z1XMLu0OHCh/S3eynn6uZ3Fk1EdvcHNwLrn+CAEEYo1RswAHi0InPHOx8aqtdl7
rQ/2Mj92MJ1xMa8GRXf1pzhAKTs+wKbVaA3JnR6P+5zFRknscEmKgnP+Q9c1H07XZbD6oDmn3eoZ
qTOxzJjbvoiiPDEQU51v4kg5CE7ymFM8uJp4g4iOTPZkUwLtvSh0kK+pNi6vsvtrS5krCn/nW3rC
sSMxXpA1/3A6kPBlAdwDIxAIZ80i37RMMN4JMLWTcgg/lLRtq/kFoTDcxG/5S7tfbY3Y5OjMHbQX
IHmjVjiwbL4CR73sgWmkU8IaYBJAc9B/WtZ5CgM/7wcAYHG/gRovAUI3ikclGgl/4K8qFKpBa4Fp
0q6TgFNnKCkIcTCwjcFcTLYuFs3gE/APogKefnRS95B/Hdi9Q3zuQMcaOlX4vt6Xio3qTkG/Y10I
BDmofLk+wq6xXQ/2VqyG7r1yPUoG7ucEdHkUIXZDy9eeZKpRwHssQxV0yEe1cjjO78YCElhtCmAl
w754xOdbcJqSiuG8hxBgBs5Uke75j42Hu5n4nKNTnQy1MrLYAGXLQk1Bbvf04eCdt0SPM0s6r+1e
uCeEAiwPH6zgB/PzJwH12pLKNhbW3F1caHdxhQHnN9yZhWP2DoMwPpxoCE90tkHXFgR1mhPLJvH4
5SH+d0hXEmC2VFCiCPmhk36ITUPhYiTCAizl1z+R3/SwWFZ7p8ZbTSGP6CSZh8YC8C9kJ9n+taf9
P6YNhYhiUbDrsQKnO3gmymwUBLjn1UZrEtUeHD9N73RMZYMJ+xuleY0kAnu+2cg6J+I9aSwuzQqh
B/h+tb7RSivTGvjGarXwEcYEAxm/Gr/cvS300AV7Zypm0eD1pxhknDGtf2VVM3h3lPullpWlWN6u
Jh88cdsEFpI20WXk1vB+xDurEvzGQ8NuM7PGCZDC8zuOex4Z+2dCvplI7Yb6o5m1D91c7uNJzr/7
xxO65MTIs42z1Q3X8X5CQlW6qNU7yoFStfuh06ZpPiLxw/kR7mnW1Tz+9Gkw9ShvWyEhUKRt0pKK
sXJV+VZxdXE7hI4FJW+/138A47onJa5aWKdwHxlLKapga6f9oWaGdpZAIQdr18IQIKp5+RZK2+cH
iIF+FXsTggXikTS+zTP6V2B5kpG0yoEM5d8mMEMGKSfWKAXP0BBoTbYADYsUU7ZgBvY5EtoFaKzQ
G5ws80ou5e2qkFtwDeX+gaDQ2m6OnLrI8vRi850Yzk8gTePfb3zIhrE61XAfPXfymu2i1olyZ9oL
wv9KYYUqlzxJnvXRrQqiyh+9p7V3m8RIDOkMBhYETZjZ1AYAIgRwLFyROGqQGjCpiHfkUbs0WPhG
oO8PArrrTi3UGbMzcOmekgMmREl6j6qd6vXCnxNq+Oc20+PUrxeOcsmqbrT99uJYTF6YFVUjOdsZ
JfOmLPgW/nfMDr9XlBjNqwNR/On5+SlmMzcLYjLa+LTm92RhZTAVARSqbxrHNUm569btdSF8E7+F
a3qhmXjTQyOwoasb8hxU+QbUfIK1NAUHIKWsnaH0cCqV68WKg/iZci/2hTkY1faQgJ0f2Oiy/x38
wsl9JXO5F6bh3D66719HJY8SfNJhLBlyuIErxTaV6hjEPG1yWANCpYX6TCgw/6pUUeoQl075Jp8v
Pipg1UB9/5qhJJlhmynFMtGVPnlR1UaTRP3PWAPRaheLV5fmtnPBCvBA2BJYs6S7Q7OrtfM1JLKm
YpPD1coKAGuat8Of2p0p1Eq4PiL2VKypF1d9qFMD4Bc0FgBtBTAqgDFJqydu0tSABiE4DhDlMSnO
4NSvV6+qoFQRwjEfJkUKp0KqWKd6OVAuNBLnoh0DlVNMJ/fPDoMNbAnZVCEY7ejfW+euJWCpFWwJ
BMdC7IekBpiysB5EmK10JQRLSBTW+QyQwS+9K59cYd+avtIHbTqGhBaFgFwQy41ZRH7wNGApLEDA
BljeY4/6Secnc/gd2L2PIgBcPep+M+rMTCK3hK+Njxn4ZGNotnSmh/7/hWTn0e5cebWYSj4XAAXL
u6kcoHpneDgjsRNetAEwvnAGFawZLbm61id7QJ1/vv9b3nyJgs3GYBZh/XI4slCz5j1f++m/HiCZ
eAx4gpdYAZIo3Lyt03ZcIAXalpfMlPhcKuGFasF2SPlD0a6+nbRApdbL5zF01ZepkTl7aF9DWZ7P
849/wYBw5gs0pVxbjIvKUQJ5lWDrltMP5ipXmKHpovIDO9xZiqFtEuQ34MKAvYvNVBiSpAtiluZI
FBuBuWE3Bs5YSwu8GBUfMLCGcx+LOfRlFmLYNflGGiktOYU7FsChEX0svYhRsnc08kD2jwNsnFnb
Kz2E2hGcVVZllFHXQzjLsconsQEtfMm6eALLr+jXFoXY2VzfyPYMnzQaVMnIZBfc0LVCpYP6cZ3o
ugFPRYVmgxj3rha2cMl1RGNG6XjydKsJlgX1QLX44ripQxtk/QSgLJ8ZzCuBa72WwEh9xCwfoqVS
ZKejVf3LUFq6+paWByG0CPh6vc0ZX6QGvmAcuyn/UOcW1eDYyEAKUgx1Gs7wljGiDRfO3IYHN6tw
UmQ68ockl/a8wBv9st35rfupi/focI3nZDZzI0JRwHEJbgemSpRYWv7CX3WFIsmo1TthgemkmINn
0tAYsfk4xwXkU8kNvKSzftipussuKLkRU8fEcGP5cEXASjXPQNlX1w1zgjoupDwpxkQTOgL66G2r
7LA4TXgZINbe7lSdUMmt4lEvPIV27qAgUnsKurGwS1EM4GE3hfvx30p1/VXIPI8FCEbWCfbXv+kI
6Ah1cypjKMWsS57AXr8FE7DjjxCVuDAHuSKGf3wTnla7bStx4Zrt9j1AjiZ+cTeHUdN+Li2ZXv27
f410wYVMdMmCK7fUxZHgInbaKKH0ssdpMHXVqXN2GUS1cYYob0mPqhAs1PF1wIY+7IYWdt9FREVw
rpl2AqBOJiJya+wy6YmPC6/FF+/N1LeLQNWUbMThnqnX+KvQBzDgLpuMpzKmMjg70yu26mIj0/ts
UQWgg0mz0DAuPDMZvtyCQCiFFrD5iHvLzqKU0Sfew7OGL8TJaXaMqbaBQ/Tq3ovEWoOTDyV76KeM
7dkYe20cG76KWRBhSPnXDCMsUTPitarZW7jPfDP0LrMjUMgb3sk89d6eZCRPoIiop70v0GbsMCnS
SAqMthEOpaLe/wRPxpqiJEm/YZeLRHUbP/4i32b/H1TT9+FPycJeyK24h0OvyJQv7ARUSzNIhG+M
m3IRd8kYl/jxs2LrQhZMzO+e9JFNDQL00XUws0sgcxtRYLMQSgWU0lTvqHcU7q+Lr/P0d7IfnSpo
es6hhDg8Wr80ukvhwhk/A7XFvgdIOjyXaPTWHJVOItG3CxdrctEcsHY/HdUVvcSFSk18DGzjShFz
BO+l9JTOVVPhYsDGfIHMckjmxuCYkfL7p1b9cChUW4FQM4Bpe/muhyrqiQSElD5TYHTB7PdVUJ/o
CTGEEFQltFYQSA/ynj3AUAB99KGfDm+nn4HOYaczbmqJLrUsAupNcmAQtgM+Rt/ZsZCJiTMG2Gf0
1uinhfIzrYHQOjyVgccupDEuN7CXkNY6M9O4nKH+keZs4a1B4JyM9UFTcz2pSjsba9yPUSsDndoD
lH1/Tsz1kgoaXzrwXupYIvsZR98oX47rFLs/lqEsDYuZmxcF+e/YOuz9aSzTPXRghs0SQZFp9WGm
bsZ6xAacRTsa6YwVE4RgIxHn8fC+bZBKqz+rns5si6TnwoczmUDUmqYdmncWCsfWcrb6744FDNqO
QZb3flvizFm7saM5GYyDoOy7putvf2YJH1unB7A0l7DK9oZ+gRA8JMaR5iSFxWIFtOn5611Vn9uf
cqDO1gYqhy0MBoKjAxyMhMnWyOwumLD06ejY/d5R2xFHTM1BSKXRXCvSmkZW7qoE/6IL+PmzLC9W
Rp1AVTltqjdHA1fk+GD2vV0XLeQVD6M27acIdoPFo4zyOUCMQkUfGr5+NRINqOxMdrKZhKJrRIdT
ErHHsrpsne5Q1Ct7vYUHk8Be2p3khHWU2hMN/DjjKFR1/p6al7PYB3FytS7n2HEywyqCOFjnD2kn
AGXk9aa2N/Wujhiv2pF1mliPYCJDBsto6R2Dz8OsUF3i4TILl1vKnfC6/i/WD0wVvdh24zjPSntC
Ey5ulAdHHbqqeY/oxB24j8jWlpwH3o0NUmrByZ2kmdYKe0ZBEIankRNKBmKGudqEiUq3YaomSyfP
M2rGP+ax7+3gPEWZIZZWo2Dx6+DCJ5hNud2qImymOiEcHFO82wOjVkhM75a4+drQCKfPqWr5uUN4
//BGCd96Eb6ASG8d6AYlkMZS7x/FoNgy1aM0Zp+hPWCybnTDxfUYHDnjbTLC0fJApe+2QK8FyMnx
miC6r9aLz48WcxHpnVFLwIkHyO27biLjSvL0eL+QmWSmcpijWTY3YJLcHnM2jVQLZm6OeRdPdIUF
TfGz4otkesn4NDKQwx2coLWBkS74uLLPv9pb1bIiSVP4P7UBuHVQFElIqIO9hpn+3BZzCbzbhVpa
vtlroFZbdVN8YNbVdpmS3s7RbbtkAl54BiT+MGJCYSfte9lcBx1tr/GljMmqGLizjdzpyt37LvP1
6FjXsAAZlTLbxwl5VRTKbhCjScDV4Q9G0XtK6S/VgBhqciqAPUVssVumRyT7tNI+9+1c3dtm8Yng
bL8fCvkl+dCIBzaxLeJ9NVtqg1BIikct7pXykqa5lHxKLx7df/aKVbMGz5OIHZialuwndAhx6lCt
M3veclvp1GibLNdXOJrvMbDt0IvrXlgGf/ies6FUGogDad8Y4KBmAqMV4OtIDaNEXWYKYp4ilJCn
I6muysS3jWrFqmr9o86z9hsR4FiSG2BWL7LhDs+a0Mvy2o58b98SaT0QQ6qiGhDlhbssBFZ6eHTC
YPs3eYGqzzz1DtzvM00xbVda51qSB7ip9jxdRhFGeMwWuL4lg7dOq9YeonsAlgBwnXlpbzoq6RXO
yXCb9zVwesTGwKOut3JAfHQcrZq7+xvnR3aT9VyIF2KlEo69p/0TZhQgMyfro938vYOCJRt4S9i9
eVppmEmM+moK5g0+KhU1iYrmCM0lEuGZTnkUb5CFMjobOxoNLAsHxdyYrmSxj0wr3bJBBRUrUMXP
OBUOC5UvXWb61RWaaLdAQSJId8MvcahtjJfFTeCdWanalwM9X4kTifFeZlJT+CCp74pc/t1h06NU
ZHf8k91KXOxMGkcmFzzbuFskaMStRHx7AZqC5kAEQfzRVbaTUKk7SloLSdnDgNLTQ1dn1V7doT8Y
ubaJiGnwZYbGKtU+xfi0s/tIYPZRqvyizjFmix2LzgjKB0nYpG/bT+mCGSa4YaZ++eOkueksvNBQ
4satnN959r60JHJFBxUHLSycOqtjHqO6K7vIIR6O0l0kFF1wd7I9izs2m30PwKhBSVlwt/V+os5H
cemgr9t7rq7xr7qRCKOaFGSw1YlIC72NZMr1sQGOYxIlvyvJMERdKunzIhg/GYB/JO0ie+gqIIKB
IOgQlP4PdUZTgUymG/3CewucWTsFdz3pOrY52WZGF0XjtWlyoOZ8Oye6f9pz5TXnykVyEk+llPHq
/t0lb33Ih66kIVZaQbk4Bs41K+afUokb7umVRRJzQfaT0etCaFbrRVce5A+nFp9Nt2uL2NDDg+TT
RQS26o70o9FTsqgWzUUfqeaWgHHpTFKFKxL8EQsXFa1iRE0xF6MkH2kFctz3KK+EhYQS60HSgcxG
KQuRzJGL98XmEHmlbu06a46NNF1e/RIrUsHdlw6XFUt/ZpDw9q0we2ePjMKdHkd8hiJZzOaqHQZb
xAFeFEmMrbazadcYJeWWbco+ISzDLPFDiQBb6oG2v5EiNlCn6qJPVtgPSlvDiXYslpIY8Mrw8j1R
3+ZBAoPJYhAjXPcpCK/TzKF/3+sjOlJjIpakie36mtoRY03G1wFhO+Q7EWAR4TIuqAB8wKW6GCJ1
WhKrSL8ls8Kspduzs8Li37Z3h6xHaRR7iPPzAIVQnVlJk6nfxKM4lA0J+9C+KwwtyKyES4x8P4Gp
gi4mfWqmHK6WFGpEBgtPZTWrKrssX+7nIlWc0mO+PSEGnPBnoft6n4J+vB/2tZAGypIv6W9K2JlN
7bxzWDKnAc/bvUYBIUr3YXmqKgQll5+biWyAN+IUPkYIDbmkg1MJNNGOESzqjLiEV7zaQMx8cf1l
ZaJs2Q30SLBJJkEBPnW3zqf2hvK5QbbOUbm7+vCFYFeZhutsNR4PYRz2XjJn3cHQCjxrTVZI/PE6
1e06nAlT099A50s35kTlzssBrCE7GJBNc2Fccf74Myc7oxUOZeqP48U6kR6WUur+VyAYUWaS6Ocm
fQ1KRxwqr2nOGzGk6bJF1dEP4nIUMt4k4v8BT1PWHiQSHS/eiYKo07DTith/nbAC2eVAzuMGkoin
92VNN6DNqjSeoCIE8HcwgVlDWWnjptHyX+PxWSIyfk+x8jnqCFgy0TObl3m9bE9QCa6Zn1jwsWhu
EEoKm90JNst5IZFqvlGDytJVCwxukyeCTcCRRk9ipAZAj0LfggWzJXZh3uXgPVvQ2OagNeC+e6SK
lu/C9vOUUfBBwWZFZhzol5IbvKYFhi9uQrzsiPqdFy2lhCrgLsTVMUiUzxB2MrRILBbgTKma4PEK
UqXv7Vw0ZQC79QgA4V0Ds+1bsKSMUUUnU9JcJA0SH9Fsk0eACs25/uGYDuJQTQwhBL6gWVdzCWxz
BofMSZJLpxY4XMVs2e7u+eRDcmZbYLcAHziT/+GFecsa15guZf45CR2KoRE3JqPS7m5B42jjpjmS
F0tOyI9Q6bsvEH83vyO/fX74YH3uDHgyhIv3brLOX0mUNLGZoeyG8hY/s/zZY3b/d1TRHhOsxly7
SkVJeD+Mf4DBmowhCWOy8e24K4HX1++6le+o7zBFZ7Oa4FwlbYPJ/p5O5ONMnez5qyqJGkdaJKpj
7GN5PGdLYkywURJTrq+9JQqD5Y8ZVPGf+Nk1KQ69im9ZT/BiviAu1JdRmHoGUfzXfaAdzamo2qHu
yGzi0b3TuL+UaKefB2HVrL8nI2zi6nFXOJE7a1MeQLDwm7snBYhziS6jxskBKjCy+nGrzOvLrNsS
RcSQn6YV+vZ09Tdx2A5Zood1uYO/c01W33+OjGWviGGF58b3+btwp+JA7wwOoSngzDy7YMn9kvN6
ncCPGgqEs7O6CzE3fluXomylAI4cCmW6bN2XlhuxPOtfPYTW3LqnNJMyfiJJ0Y1ltTA8++CZi1KN
jr/PgPzUFCh8diP8yX3vHyki7vK5bwPZn0zgLqfy4iqV1jrVughguQw7a8OidX/yfoloX5bKtG/U
XdI3UfytU5U8Vhe4QfISPpYM14uG/3FN681lubI/qYmXc48yoyg3ZcVoELwUwzrPIouuj9p6yUU6
Ox1ltERDuMz1nBEMO/nydk/03mdHebxgT8x1FsVYZdDr8IKQSUkPGqx5qOHf/Lg6ST/uL+7EfmJs
AChMkrw0fOlcBNxBnD3nS/8HW2meglQam7I9CI7TDReep7qLPWQq+HGsrh61Nrju7d6CZtajjyfE
nyib+5BMCZXEZgm0QrHhNbf5RHrv532ODvRuYgR+KiML3IpSqrCKvl2TyAzkWb8cOciVmkKOyjms
cNZlbI2rwfZio4zatEjIWKlFVx1BIC5UD2PJ+EuO8rkiOu/NJtjSDoPDmsGfXR8Wkft8pucqiFfE
0mkV3xk/qxrBAFsiVlki2Mt/WGznYqicEO4Pjaj76oTbsL0um4CbZwt7QkBqEJYR0O5IYouzi2fI
4HjwGRzQTTTwyIg3XcaD6MGQugkahB/uKMMGIix3WKIisVQPk8HBQFXCLEw+MffTBgINGvUk82MR
hEPLRuvNAt3T3Xs6a3wD28rbEETn+0KYT+di+2JVPtGMvCk2kezDRoKSRXoH6GWzk5Y/R5I8Oev5
hBup3loDYBe5S5UJullL3KabVQddcp83HTzbMcU8mI80dRoajzWcZczfShZgBOX1TPnuk1yNlg7I
qIYhJfaC2xP1Xrp4V7Awu2XguzAxl4R2qzfJ7+9mcof4W/uddMTwAXNt5oBvcyC23B5c4ioRd979
j5WYMVB7xu9p6pbry9YkumPtxzkh4xm0kPgqL8BrHWgE+dWIjRkvN6q7cVlGMvTUu0x5nPj1P7hj
26BRkl+2ssvfqPNhevEpJO405rIfYjjzAqIDWFYgUUlC9BCJ8jWHdPHdsXPNFemMM93wp67mPOqn
vCzzsJ77Ywhm/lP1zkqKveAyO2Ki4j3WkCuWonpeSVQU4KjnyukGYcC7rOWsuPnaXRd+c+cKEU5+
aIWIjfWhuNgRYVJL66Bba55emtVvaFY3O51retO9aiyHSTO1exIGAqyIKJQhYjfAMzx2EIe7+BEV
muLCHVrtwTpCx52yYDHmz26eiXOs2v4tpLKAfBfnAIHmg/kLEVL+S5XQ98dEpOQIKEip3OGTgczJ
kZYFDQ5saZj3qM5m0w15Gg5mDP3xnm7Wd8+q5HdnZGQryJgI6iBpoXvX3I9oStLwLu1jLjJvTlk/
rKtnxJbM8prfcWHPxtHtt9qxxzVXBp9u1a8l8vw/2C0LqmeI0bVZwbRMepxOdmaUWgjvQzwqNgH3
zjMAVII7cNu9wM0zrz+zsim2LYwmUzrm+nq06PGWF4weVowKp/+oKoxA40RqzwKBhhiJVTYvP7oC
x2NdMcX0djw5QsHXKZh8TFBdMZzg1rShzOP7kEgic6PRwNFcrwP08Jgf+LcgWlcXTEP6eXayYmEy
UM06AtyG04tIUK21wpJkhbRsWyEanVbpj8gZxpfQRETyRAmSf3GHq8pAZdWiN27qob2hV/78Bfo8
CogXDalxpShDouULQbf94pLutdi2/h4fvtHM3zqhLVOa4N7HWPp78pz1xIe9L/uT70iBiAFI+XJV
uUFqx7AohR+6MS9KnhHIM6FkISY+Ew97g/2dyGFgNE8ooWbvGhGvqFjvho5IVn7Tv7Y2L8TKxZ6a
xIumBv2ekbMDFzLLci6Qxf9R+l5acRkJBUod2eZ6foQsgovgqyaGcLxLUSUOPYOksOheUBJPyBEb
RKIXVUsJLAhJ4ObISCXH3N0J47aclxVROX+aTCvLXI1bSzu4b4sDNUulFoucFI0IcWq2rMaxDbzo
BlAkXL+rFUsjHvV1cs8JcNHXFRAcdchy9jr8LXQgyv/lUiOE7P1ia8uz6mTBgGBH6yyduUzfOlE7
hb5QUIIS5aOl+E0LsN+GpEJRPmxqgpnpNRPj9+y2v+PhH1M0VfxICuBM+vczE5wzlryPyN0vlaUm
ZD7wa8mxzmqbaYRoe4Gh2mc7eymLVwX7zOMbyn8A3bmOVTrMTUeyJUotJcKA7wNHs63n5jNMD9lt
6Hgm7+VA8HaeCLw1SO8m0dUG/LInQ68NGKS9+PesmBqz+Vq8gD0h9toyVV9inVaaNhNWyLB/UxLd
jnjwnzxvXf3ZGgNS189ErlkBe+U/KB0l9+BsQZiZx8ydeXJ45eu7cBd5jcn/C6AV2LvFOK+zNoY9
4Gl2pNxpGIJtqSLslNYMYoSxDSX9ZHqgSO9YFtuQ82z1vM2F2LuEZbrPuLzi4vh3u5c+ubJ/6yf5
LIZ6QhzAcI+8kSKVLMfvTG2RPcT/Uin+yBsBlHighYe7D0z1qsIrBnFdDXaSw5p6ZCcAqkquJob0
GbfECLcn5NqSqTbLOhJsAHxCvi3AhO2jjEMM9FddbU+XF17/4iAwB89LRv9pO7p2E8rJJlaAPT1R
JJb1pwYiVVAcpOIZbY5k8jusPOKUL6/L6UZSxRo4CXIjhluBOBaHfdxtuEmm0ExzlpNe69viqTHK
map7zOp7Rv/Vdfv3Cdu3b2NmfZuu7nniCttJlqoargqvx+42oYLZlMv0aQCuyDChvVlprqXvhIyi
CUG7oxmV+Fkpk3s9IaKJpA7+BatGkgT9iYUnhJI4J5XZi0h/fRrwx6VJOYyXIK7nD//vlSAMChD6
LIMY6kVEjA6dmScR7XHeBbPDqiTirfN7ez8qAwSuGn/uZly/fiDPmjP9gHh/e7y4Ay71+XmYDhO9
kUopUuQeQ34cVfdCl4mrNyM9nFwAJwyFAF+c4vzNKGjw5tsBlGawR7GJ/6ES8Z2rrRD2nf04v2Mu
RIbtZGFPavhlVE3JWuNeiglcrOvAIC0HAUulDJleLwauybMdLCBR69hywa1oIR4P9spWEZR2o7QU
ZPfY2Cg6Cjp5VtZhDIDx6BbFwKDFt8ECqIJLMoCR/pIpcdPs5kAMSa24IfsDZARIjouZr7gf/L8/
1A1Y9tgYvpgrqu/YqN3jVyskiSdCha5bJoXVlIeTMxqxxMgxruD/gnVziUEtkOZdHA4COVE1k4/t
fiC8l8CkHbCBZTneesw0/h9wyn1prCw62qDdLDcVbNw9VZxqXrE2UcQJdyqp2jkcTbxlCxq5P6K6
c6jWUw+PtKGuWSq8j7nByZ54qVP/WXC3jLlD1w11IPICBa4kqHmypzbucjTFsnBnJ/Ildy9hJXiW
X9K+lIscn0mYB0PdUdcwOmOPB9LbpNbbRZ5CN2+g+IxVHEwiQK6rnNu4Z9keBGYDls4JLt1ZW3u3
gfeX9p0Ru7mhtBY3wpn5s0AoD9TMiLRDzhq5GDvoQ/z5/ayo/WMTu2w/QA2+GhRTkBPpCdC8bP7j
tvCzbBUYkufferZzHm3ugge3QTH7MDWcOf/Ax0PZXHMaiQ2ina4F/KEvR/scviNGt0CqIARE/3zg
giQw+Xlbpx7/HfbfEC3khItR77Vpg3Tjm8vsRN5k4La2Nak8UzB640VJbKPhawOOUI3ze+DL4et8
DnTaUe4AXu5EEZN53bfnA9feviJW2oYzW0vdecvS8WaaNvrRMs0//OSB8ZBwicQrYVzLdkHgWGop
nzKgzA6LvgInBtkEvTY2XtwKhEsjToYpOijeZHjcvZWDgSmyRNbPf1tBOMd6h/ha5uixsfIrnu0m
eJZpr9inn12AR4zNqga6W2sNCTL7Uaqq1PJKrHdWZAujlclH2nlSwN1yWvbAlFECSBLXaK/enjVn
hWNBKNPMaD2XQ0iuMeTgk1cKiTd2+MOwvcKlhK7POrQXeeeMKfJ14ob4ZbYnUdQh7TXcvxirTfCE
aPCj0zYpNMTw9dXp+IQ/M/l8ZhdUVu2mkkY2lCF+6ak5jkvVIQ7SUz3MDOd/Bb79EJPymC3yzLo5
Y5V93d3rzP/7gS8QyTJoKetUXBW5jgLM/YoUCdYvUo17yCdcb8hKKaDVI/ujtQtDpoVEM0SEyddd
eJvBc4H/xSgw8aoia3zT4bzOvvZrqYuMF9flSweq4u/ct3ONLN9bHX5X9PzwsddtCwH4O+GrfAP/
HB6YeigyFjvtqIpYA2U9v2H1MTIP/x7Y39hNPtuEVoywKY2VJ6s5etfuaL7gwcoGMZa823YrPV11
ZfN/7lZSxGY6xQ5+u+xuFPxo8JAYAgEUhtq6OIG9FTZgKi8sw0SrIxDFYHqBqnZX2HRxLm3GdmLE
p+drXcC/b8HKfD2+Ww0a9bqOSEZrn/NiVKfzbWDI/ZHKOl3Xwjb1XL3gmK39u862lA+Ah8gdJf5L
8LK4Mh0KJNQCP1VAg9b3qqbYx7VG21WGJFYv+V6nnQa5ah5zohbB8O2dDq0muccJegqMbKZ4lVtB
3P1SYRspkBYtXgfKA0+9fckWOdZl4gmJu7zf8iH6i4m8bp+j1FapXxC6SpQIQ63bDHuCuz2vdQgT
+sjobZ89dCKZEg0RR1G85tmmh738lzGc2qykzPQI0/oP8PMX4pj9qZq69vLJE0gMCmbEP5dcB4/4
/RtOYhGlBGFI/9/KQB7Zn912dSW+AepsOmW+wg1RVq+juobgBrOuesoniNDw6yVHfXiKIxSVMctg
GEL4AkrnK9jm0JMsCLr0mcSAKixI5XgoS7hgnzwvEsdKEEIbV0ZG60JO1+wB+9IcVtwSxqYT2iVM
4NJGvwuRFw7ELhliRwyXZ7mwM5RpfrHF4nSeKvMlvWG+XvgFR83fj6OrwCWL0eZ5krOMumTFnlZw
paBxcsMQKuNTFyFHLuTkAYXRgZWZqrdBki02QNwHYGXWyoJN7ChAPuAyWCQePKDby1b4pjrelitQ
2dFw3vy/TwkVo4nd9oDhCiW7q6RCP7geoJos0IdfZ9SK1noyAfyQQ5tI5ul3xRjL5WajJbmCoEuc
wValTqRANiPyxwUTYrE23DEtCzPRB0/EbCXXN7/0YTkC4Cc14tXHi6I56ocHkVgr5yqRqkGeb96H
gCVVmDj1560BugYnm7ZP73x9Hjlg+s0HZ6/biHn99j/je8qG2UKyh/FulNB2/KI1Fiwwe/Z4whyq
KkqyURxlr08TvbexQu0SSjo3MCne9+y7Mq4852w6ztw3c9qUgOToOH2uUNUrragvh2SWs77MgYKi
rQZeHCkVOkfu5twHRV3keV7ASvjebcjHG/Wstj4SM+CYuFlZR36sIAY4+RfLy+JuLh3NaUtWZrH0
sIt2jdODAYWcIec2Ukkh7bYsOQsQ+j2eCUa/o4VREno5A0hmsFnguMYCKSFFXIkjqNR3yneBQvlH
lySP0OrHIUTYWcD5WrQMaXOEjhe8vSuw8xybWydG5PjcHJUFK6NcXZ8vPnkwHTsKyu8NDnrf8FAi
9iRN5hgmRtpOuF2b5IZuythXbKvPFlh4nbfA2rXEe8foZzfl5zwiwyvrR+87IJ0wvPD/KMmjDY94
txNFG+MBWdd45qWyJh1DoUoJJ5Ovnheb6xlwYa2rudjULreygUtWaaifwKex4UPEVfAMJt9XuEUh
G0dbGiusTCmGiQUj/xeEjCr1CcSLz7Ex5NYJm5a4rWKi3UUBycxN551fPmHsGSc56MlRIZPblMvE
goYMqAo4Tbzm2YgK1yX8aRDpYgNy5cm+cWcX0SmcbxKwxG/COF50fpYUaN2Fx6/i0JjPFNsoldOb
UJwR/16Kc5v4tuR5PugOJKFPannKRqchGn63QlQhJM+YNaRhR+k8hh6pOq9XR3cqRknUXUhOvDD6
vTLUelaUKX6j4SOm6rqOJ1d94Bf6XsEBW6UFKwMULLhYCzbSXH9els7LATpQDA5F9vUeBSj6TQkC
gQTgTMDFsba5URuhZpSMek62/n7yBfX/s+CRbLJFXCYj8T4kMhI+KMmYwQcI6tSIOiz/1O652uci
GVMWETb2MJ8CDnoN0oe6nhp+SsQNQKBG5kXX54AmCtNJOdux7T4NvlDd6of3dxde/DTQkmynpY7/
D0TYVnNkrKIY1vk+ok8D60r7lRf4nla1iSjKXjuoTEMIMoMqpj8MGrJk8gYXe/XZnaiwyK0HEVLP
l46CAhTm23Us9KVyQHXzNXzv+Zn8i68b2BxjTYmBY0J4sThcVLCzoPgT4zJVLopbUj0sVDmt1XHb
ywT5UW6WLpFwVsIZjLeAHKQEWH9E8pWOEK7ha/Qd/zvRtYssmelWakbfLyPWZjHM6lNukdMfS2PN
8PmxlDlYUfakEqogc1xsNKs6BLnoTWmEvt0gzK3QgSc0Tld7VIdpbOBdA6SDB1GB92bRB6l6iDAb
qOFOa2nUemNMtDRJ8HthqAo8KNKeHMGmySg11Y80W30sT4iPNswDcr93s0Le7sxRT843cM1YjAF0
BppV4/t1MCJXCi7X+CAydCeD+o2R5LkRt0XXoCiUsx1nt+ujaH2TkH4XGREBujO9btEP4lldT/bL
0y+p/lI2+KlBFo0UQnQpc0knBb6XZnh5PrAMW2cgPb+FCqKE46QdWopN6MFHGY6NkdLThchSW/Td
vuqwaU9N3RW14eTgxz8H5Lzz+YwdVm1ZWprzhdgO8IbR4CPV3qn1yGpc4cxjCoboXRZ2wHMSeeLd
n073e4dBdOVNQ/4p9jaesQtKPOYa5yq/H7Zv73Q76qoQwrwwQ1/qfcnKKG7NdJ4L+ErwHpWabuam
skZ4FQjD24z6PsebLZzONSSfgzkrdVjWz3G0nsLX/XvR6HrTq6B85rAB2Gnm7yQe8Ena/EkYg5uF
Aca4AWlQ81PQ+sJb7jiasnXGeysP2o7Sbt68ygarnRhzps6qOFQou38RZwJa/tzJHizYGZWvQf/H
1X9MxqQ7H0+zVp8lPWlSCywgt+JjZsZYhAFIACIhBsuJlylUPojWiVulNsJTSPVJWO+OOdBoN3AN
dV31IWtkFR4ktvYPRtSzjQQQaXb4p/OOy+nU6UIqT/EuN6NdeQaJC/sXFMQESZCiMSdUesbtxFmX
KqjgJUdY9bG2HBYvHNx3TW3nCaJVx+lfuhM0aYw9deTOUjmOW1pBHjfu0MNWerGC4j3HR99D34gO
dcqHlbR/JudiNZD+OkGxSrFzehzBrHrkRTCG/8HxfClvVUDStAdoew0YD2lrG9E/GDnSjznXfwPz
nfaheXWKCtvaMhysh9XXcP/10+/lcJH0efDbYv192WURBT0hymd6aT2jQeOHM3rU8wwffGhv3uV2
m1b/6I0Acqml2sjk7DDLrEtvxMk9niyoQizUpfIMhUGESvNsTcl4xk/um/TVagttnDh9s3Buz71w
aGo3Q/ZWL/cw4ymKRhD51OacXhx0VEHeODVu1HS7hHMPBZPn92x+VJLpXid+kCN/g6rUKJGYD8N5
itljbZzLTjc2mzpX5vDfDk70XDKfWRtIs+XGUutT+EQYksVR5tG5Gb+y1c1A/Ct1+NFzMoKxs990
MKVoCstUeumS9eiZAuvnXLLrZG+eZB94C9nEn5K9Ou5atCDpm0ohE+bv8oZPMDBr8dyvmLSxI5oO
8OiTQTUQfAijZ4mNhU3clE0Fhi0kvESDzM45jSxLqhfvPzOWuaHwHbixPOUFXAVYdbChxDMRxTc0
BArqSM1Y1OuyVDOWJVC7F6b04YsFSOmqc8rQsD/dvVh/RxIfbzTaxXEYq6TP8KFEXZxo8LsHIJcA
CMhuqjW6lLwjGGhMvM+4mZ2x+RxwdogugOWuKSjPdCaZUDxcKtdtlrT/+K0p2mGntCtW1UITemmz
CKxTfB0b1pLABv9DGq7StMQe3JELLIt/GIrj+nNPs2PUxEMQQW7Ae8KiqMPNlGz5/EeUFhHR7hQM
xaLbymUSejo5Cqng38NSzf66+m/wM6KqQZKuI+crj+7ScRzyoR5z3+ydqV2zrLqNyAqIdP4ZmUHF
lZwIOe9i5ujgQ9+ENJz+yOyOtacnvuE9ZPyv3lcRN6pI/RTvcVcR6gTPoeQwMEUytL+Fm3sb1sz+
2upmG3KDKc/Ko/Bl+TPr4XPuF17ouVsuRXr2/VJMGqlMSJDZeYB6d9WIuUWyqiIlyd1EmZ+/zMdd
YIu8EAc9UtdbGzedJf6Eh2Lh6ulD9QvUlzMXs801Y6aXzUexl3YbxQOm/TyOtsucyxaXphI9yofs
LEkStFUu8vSjf7WakvANXjRcqcf4ZM3gTMIAoCVVW+0AP6d/0O8JMMdUQsLsNAsw6alAHyIoHRoq
xUfxGTb2yLlZ8dOaEJ1ZrR+SmWRODHxDDjjbIBbSx67Lja9+WC2V2LxGJEV9hx4sLx/TgD3Xg3EO
fKC/yL+vayuT5g8FBjkcq7GTuiiJDTcXDcM2JFgzq9MpKjeucKl75Oz8HCmApzfgR5NvUzoX8vJ+
dqUK0jfH1qdUgTe5bvVaAIZD0EnKn6u1zUgmVuRKj8yfmhDCfLQUnRgS/tp6ZPbgu3kqBwq3P+CY
hP5/l8/KiZ7wRp7gfKZCJAMlwCsOeIRcUpP27lDA3ZLLlGOHaHGJwMBfZb8uCKEvmP//l6O3au9V
Hj8etzuygvOyj5tUVKZaYWywpn4eYjNVul8G5fh4O3KO+zv3pqrFwvilXXLvxb4zpVIsAuf2L1/y
kMy4z7frxfHdqKhy4gWF/3ODHGAjA/Q6nT+Y+hMNiw+NkJiRydU3zRTEFjvXfaezWw23XUHQgjs5
32uezsLTLvslcDXQ6/bC++/9W4iG6rnKbQQlaUA4gMP76EPZT3sgARWTw/5EBDFnKXowbMhMwmgX
m/i/e9bAMoAa0C3Cr1rNrD9F3TgZJwM1nC681UNhkArgkJb2nTK6MCbM6K4ZQm4x91snthwUq3LI
wm/2gKYIytfPP4r+B81nIBzIJrZInHYSYDbaocMHBI2842eK+FnjKTdjdWJYtMS0t9Wq6rPgUKtO
z2ltdGiRcaN0WoUwe+6nlqg82518lKx7kpfENhUqmH/nkZPAd/folhyAHXEPPPGsTHDQUPBxV0gc
gbSw02wMo6RIe3Nk1/sezoiuWS1zU3zzBQlcJ/6917X05T5Q0m2t8NRdvXf2VmOExC33K0PZ3mwK
O0BAs7NzD9DJe4mVrCo76v7/oYEUV87p5GmfHSJ/3j+0U4XQoZkgPd6ERGaF4LVvdAua8dF4FCpm
vR0J6ncivN2WcIjeksRvIFFdOQjMBlSCYAUPYRxZbO0K6ywk9/V77Fi2doFWGCRDYTSyD4tudZBe
FKw7b0h8lrEC6yb9InSJCg4Ra+gGhmcQcyk+ZxNPwSMXSf/R/29WRPjBmVUTQpajHeYRS1ypeKxZ
EXeS4XE2ZUetd9tyJoNurmD0F41Cx9WWD6W/szKm20Gb0/kCxZ//CiVHJ8tf8+vqHCkfBYpcYRX6
SJGc3TXnV5z+3poTXsmegEEGhyDi1fBS6IiE8QbexCQ8NWqG+BUd5jgb9nSISZXEJyA05bpoYrFD
DhoBZAMa780nRN8OJnf0CQhwfnLARCd2Dir4KqkAPKEEVqDikKwJhc0z2SUoVpW+Mp6fWqZUaSfz
/DiTg1ltqbvhlwyZrAwJ5nEYirWkkBWhjR/5MkEWOG/y3P8kIQDjstsaixP3SKtzneCtUc+c5yXB
qc3k7ma8KXvsnpz2Kaedv8sTXz0Vxx0FDp0Rw+RtcOIsOMzA8SdePcuNYTTdHScJmbDZmAfJ5l81
WfHqajFDNa8bGOO44pzQYLozu9QWxPOrcv1Qa5oKRTXHtuM4+aRoZihpieXRuM5R0HeelDstQ7U4
wbToHqdqcUCRi3O67SbT4T+eTeE3Ws7fuQ2KymBywtZOe8UGuEtbBYHJldhjww8VJeIcliEHHc0j
hNwssyt9pahBAGfsUviPKUW3ZUuiKoMbXIA3ctOPfwtz1XZ05eeOWcr1pcEpRT+XwdjRTNj/LDAM
lPuIVlZ0IgSYSc1B1OFEyqPpv105qEHIQHWxa4nqi/HlAx7b1CQy43uKoOItuCxticD5WlHGkF6z
P/w8OxvUtjWxbW64RmLo8U26v7Xtip0BE6Ea5pIaV0MWriAq6t/4VfruVY6YdUZgbqvPymtggT26
HYohTLd3OtsnnRO+xyw3AYtmTGIbKCL57kkxV2xCLaJnR9jaJYHmO5YICCr3W1Xmaku1SJU2edj0
Z1PdiY5lnRfIPA8w5CMLcqjx+TAEwg5riJNgAqa75/D9yIMUePh7Ra49haXhb5u1b60VFLesB+pK
eUPr0v6HEqpOi8n1Jh1sw8nXWGe29oSXZG9y9ktFAs0Jwj8cPchxHlR3mu3oa1CkBeAMUiPWl6E5
iBrufaEbQxcoHbJZxvqG4mmFB7a4jLBlJJ2Vg4qrYNWWgHCUpkuvolO8o4XueeG3+neQ0wngC75+
aE8FpAp4Gs22nIR3oxSuzKJf1U2gSR2nhkM+TrOgnAy/wX/7dKLg0diFyaSvPQxRNm8ykpKCE3/B
/g5/L7/W46orbRYrpYJEyBsPw9Fl6S0OzZdWCdpA++RL0p43ej3fKXNvPuYZ+Gn14wdehP1FHADE
wACCvoUh+aN4CnQhFPgAeYGHHAw4JJSP1HM+gZ7r7FTG9ZpMcfd7DjGINwy1anoLvxkR0DRiE3wO
z4F7Yr1ihWJrLRZsngMdNxmltQZYFCD+1zfblySzKrlp8V3XRm6Aum8CY8TR3ygdHzfasJJEB6Er
q2vnSZSL13LycT+qr9ijLRle1vcEMV9FWVSF2uSOHPJSzKHfD5tWkhYTrGF3hBeVMjNydS0N+MGw
1z5977E6EWfXazhxkzrru3S9KQc06W0GTHQcmIbUBCLrjaJD1GYZqSHH4ON/xvA2gJ2Kag3mZxVO
bKI90cMohzwPL3Qvc++/PpvfJg1HNEsLNrUQLSRjmlrTo+geqvdNaGF3WN8jUjdVyddyeFTzYxLR
mHjmwMTKHhynbZ6L9/TTytkgRfACQ3/XNlxRUWBJ/oQRChlzXTLAjO9+72Up3T7WOw7/cDCksTO/
z5YJYiWKgUecNH+ZpVOjyzhYz+/+g5iTgAVKH1/T/dIp/cXTdAcFq1pLx9zJxA/Em+U+Luqj/ou9
bVu4VNQQ2KXYKrn31sar+JZq/JRSfWAQ2qL/QbkMCSd8RS953mijpN1+74apMKW1u2wiIXBDTL0I
0NFM9J/lnV5CXTFJZmXqgDHaGCUARsxE9j3ZjWqF3KohQJJdBfeBI2lMcR4ZxPKLDg3NgPoHECMw
SxBrBUA3ZXXN3/izKGpPuY6E0hUiDmsaDhkyU3ozZPPLGk+qftC781lEHutyl0BJWZ+bRFnNn3Mn
q+UDc1Tfid4YtYbbJc4KpNzdBM/btttPo0ICsk3yU4OzOESnZRz1ZbBIdM6FGjgKr8oMI3OrNiuS
mdOyG6Fh2GbhQ4rpUjR6pRKfgTG79NfNabITSrIrj/QbrXyTl/EYxcwi+xYFvhB2EKUaRBDO9tHt
rJCDOcfirJLcB4TQb6vH9OQ/O+Au5WvWpxyoIQeemtLIdJ815sHuSslh0Pvs6cgFACSWyEPZAU82
RpU7jWh3Y1OePE7IpbNjnTF+gviaDdFsDRGrlkUlLEunOCnBqMLJYvTmaxnBBZSs+7/ZP2wsLB++
kEjaOSbBkOXP7pvM4ndjx+tF0ms44/psP1/mjDeu/o1/H8cOoO7bwiyc4aEOnA0hx/15ijglvO1d
rqqWeTwx/POGw/fIMGvswbLm0GA6k8BpKZupjm0HzqqeBX8GDzgrY3Iu975bnI/0llMRbVA3AagE
YYKWdvrFeevXkzJ3ldoYcZl+/uIthZYFBByVxRR8l3orHifspyYvvFH7+97sXA/If4lawR2gGWPX
eAkoTSbFhncXrylKrvHp4HJhCYFB5h/ny4cR9cfEFFAmTFyWEkEJyRYAXXizQSjBGCziTGZEc06x
zKHYa6jDJ4Nmpr9FNgUAtsf6o0i1TnNgTXORE89cShceZcRT2E+E12RbyhkUTHN9lQYbNnd6JhwE
ucLldskpYGM/rx6+Ow5hLD4W2VSPh+5Nx96BF1R7M32QzsmZd6jlaiZ83WE6pVIyqzmxDxPuM2C7
9NTwpiGnRgAKvWCE5x9jSVUs4fQoxSIzdrE44mBxvzkkI+RdqAxHpHGAsqCB5AZ0facml7ZukjZj
xF6dEingtxCWjBjsI/6+79VEetlFoOrhhbitZfWGPVD8T+Dwn7C8oh+UYlDItnvZlxyY6deyk4ei
wO4JfdSTTtTUvXJXev0lCfyzRETPhKnP9rwpK90oUn/ObIdirXvQSQQ+cNNeaziRjQlNXNeJUwMx
0gStcpxZdxx1A9N9+p2Wvka2qPS/b7lVtM7BiF87/6I+Id1XNCmrHANcywsW08a/S1nI/q9RJq5R
T/FMHVIdl+kg/fAEmW6reyJrMYsANReuIgsXpiu4qhKvIwZq1xT0L6egp6K4d6QWS9vbi3jTwyev
Fd4cDNr5JQTqsQ4GYSHGa0YItvE1CM94gtN2Wyv+OHmA7GpT4YwfdQVG1TZ5sMOAoWjs5qJHgIoE
QwFNHhRfKxL0dWZ9vXO5vXml/c4hRZC3Xj5yUg37C+BpdwAVT0YG9oLuyg6y+4UMicYNZeu4u4Z4
Lc7G4Z3aLFlgbZD+c4vRNpbQGSk83fRdfjCQ64zAzE95cTAzSx90rLv914/C8UNVMfJq9gyXRtGX
PkWEIJKPYEp6XRXGc0fbx+ppHfesVx3bCYRy/yOTmevAHgGNQn4qUJwo7mlTXP6NqpQvLFGpqZOK
JAEc7AV3W7MSkhj1OVrCToEmEsvHbkvEZmL7Ktk2v70PSw/NnldO22Ei0BSJj3ZiH9E2IWfoFoUf
YvCmdONZs4ly4QJWErMh6xEQ9i/xHxfRAohZHwm/TUF8viyemh2S6TxSeMs8nuNvau6WwGclhCjd
5D8JLIThhaRdSiw5JaRK77uK6JMS+b1XrvnuLjQCYCMWj6sf5s6w+69MdPkOeom+pRxNVcIxtHU5
c/S/tMeM2u9nAZUMsYzLDdl5PU0JO6UgjLkFQC8S3ggluNe7bYgmZtulONZK7TkyI7umdeXFdH3J
VrevOLvGDZYPXLiAhN75wDOv8e+k9EfTXwEWO4aoKyS3MaiN/Nj4f3weK8Q6ZbfyNEocIiKPdLLc
3QM9wiOyJBQhg9LcWOo4EnKApfqOZ3lRGUqZsQPtuEbn2JqBNbRa1RpeQqNTPv71hrHS0FL6Rg87
M4httgXGBtxDqW8Gb3FMUsdqk3FOHQEgONb8cRwG412t48+RTMLvzd20qANuJ3zwwsEsPDV7Wy1d
Nqdh+9g5iu3FxPNWta8GCvjmepGfXg7VyIrkgsR5KmnhyDHR1vZqUud9rRRkLGJrszcOtYHGXGC2
1lEloqAAdCmBblBzrnEtGPXNSpPqNxVrXci73t1x5hcC+9QqObAG2bbB7U2UkAGSZfkchLm37+KS
0pKnsyVceXjD3V0jZm5QYz08Oudsbtz5KTHjcD5KGfnUZJiRpJMOojugcnfZ6/+1JIjyFSOcjPNV
xcnOo9Mvh35QT5Fm1z+TRGLm45FQM8foNpw0BAlSYYWIdtP/3ZEpOpWl0Bln/gX56+oIqiGeKKY4
Pn/Ldtyb9Rp9DHjVNvB/wIjJJM3kXNTKGueatdUHMEwyGcowOJQ9qnuYQRB5XEmrNFZc8AOSJZ84
FUIOaHKHyemJnkauZBP1v4VKKCAZmmvpwzInbXuvoBuCik8v8h9r24Syt2U08gj57nu63i/KJ0qw
zqNjs13q9SRkBvlKXoxK7/Qb/o+Hq3PIXpIGY2TqtfPvitz6J+d8/nLxW0V4eYY6S7bk5EqBRwZD
D/DE0dxlQCpMFA8fuRqeOjOudMTM8+/EyLH1qKaExabGeSgJr1ds52GhoKXATbDb46PlgyHhx23t
zLQhXd6dxfPPPjJKAWjLo6Rzvf8eF9X9wY6cfzdjMwjIX8KLuDLK4c+dICDYmBKrBT4uwIJdK0HJ
GklRXjlLXJxZMxEMocDEKqa7R+80W0bUIW9R4LdkoU+kCYNJpqWRL0B6mQpygiJGgmpFEreBQ6Rd
C0n4wFh26GjUehMopra8iFkOZPo0cOEi2iHejYGELEel72vBZYrk5yIy2CJE/FXw/3UeiGD8e8Sr
jZ1AyUN328rcIdIJ5VRQJ2CALTciEmwqUDEWvYxsyOu0BEad3xTF4OaWJHXnfp1jt7u9Oe+Eq37g
BGPIJZWwG26VcFkE073++Zn9Vz3WFyck596Gvt8safi0Xp4N7JGBUC7dm8jrrFIr3p8IlhRVc6ek
HnLV8Cr7VKo8wQoFRj2/RX0qHqZ3LBzyQk0OCawhDqvYYFRQN3kKHMmBgPXTCBp+cxx2GIYEA0vs
/7ipq5SCRryMVJ69rahRexyDJYXBvCQXwCOgi83t+8RkSzC74OfoDIW4ED4RLfuv4m7jBKa+I53k
ZIYmeLn91rNwHpmpUimmRLAXq1bDhuGDEu6/JEeb05NX393o0mQwBNq88paj7MB01bd8BQmTes5f
NEJYAEx9iMazl6DGyUTTBHDqwWQUzsw7mrU6Fux9e0HNEi+Mgn8KiPqlqtRCrJWZRDvVMhA8N7sA
/PFlbQ64YgIUuKR0Zt1OfOyZtZiPLV4NGDfpnKrACH3Va8F0j8+a93Ne4R2JMUNVyzxOrktHxSpM
JKv4nX10vpymRHDXA3PbYt4JPgykHXDjI2qXZt5uoFd6eNQ1rqESAoRLHbkzAAVyaujXJjhrQ9xb
pb+er1c2pgcbFzUpszZb7dRYtkbXlSxjU+ubTHtEExmefhYm3NPii0q1yDckc0KBVkZuWak6vQ1X
GGu8cacOiiwJRJIy7FLUb3zHyxcmXqjE+rymXmwCYF3txmsrO8JqQENhNvG1JInoVX2d5/zeSxc3
YupaA1Ptl5KXSWSIhotOXnu4mQ/EAwlcSsUr6Dt5eb28pHh2IiERpsHJy1jAhtPaL+6DeN1NJS9H
mausyKyPgYrcTCHpYuXEl/GohVVqoiIyMaU5zjj3lWlLFM0O9420yoVedtFi3OlT1IF+dRo1GE/a
QEGAyXweiPnEyZ9azZBr1yWM6NmWnPdTLH0QdQTmufrAFV2yHK31k+jL/Ss9kXkJ1k5rSew4+NiL
E2y4pe+eyVLbmEcqipZg7FXWCsb6zJb3Yu1qagl/7pkwGcGZZKQMMqtEX36sHJJuwo9MS0/yQrTk
G2QkYgfjWAaOq8P4AzTkL/Lyw8ME8qXPhTMnIejHiM3Yydah+HoKIoo5WHbdLHSKvtc3nQraKwr3
ORaDesa7iixPr7viVJL518vSifWuDDR6aq3mvjP8Xml7P/OieNKWByyhQfcyYLs30smB8fnlsLtu
hYBW6CI2aH/R81igMGGO6pTImYkqJAvvEQx4nl4P81DnATCW3RKf9HxAN2sJM6N3BdPz6ZWTe1ID
y307G3vn77J8cYAiI2B3A8A+N20vkDwAf0avrRLCS1OlTF7CIhe5GoCorBR/l6KAf49guVTT639n
pcR5GVTUMoiM+dhyO9bQkt3YmsAguBAerHAd+HdeXMqR5Xb6WNLKULAR5bHahnqlQIhWfl6zAzYl
F+nwPlrJ6JD3RgUfKjJCfc7CRiSpkqFWXR1aHgBT+HimBXmIbs+T4gsMvl5MX6875yV6aWWHIyyJ
PHd7tPg0fPgcP3Z0+CYZ7Oeo9C2jRV5zm8Olkx7rcpGIec5s/nRu8nnJui4g3nFAy2jwJfGZf7gX
35vg7xDV2tOUxZGtlQWBFnG4PZpCEoU8Id15xz4sW7rk0EmM+SJ/TXnYyDBQ0yaUXs+Lj5+7XTtF
b/c8QIfwtEFe/kuTUD5KhFbdoV3Jy+bY+xT7E4fqPwMcm/tm2Sqed9bLtPcnp4vOFh9c25lXAjyI
DGuZwGj3wwOP8U+SkNVkT0+ayi/THB5gNtNx2kuNFlM97eDSj0sBw9398n0MEI28pe6/n+bGRozI
cPX9hguKhm9G9GcxXmhxK0NHMqGGs9bubQqwOLgzohwwiHNxg8ov1qvBjMl+Yqf3bozETu7GvmqF
eBqkoqm0Cv8cHd8H5/PXHO/NsWv77hi7cC6t+upDSvYXpYN2UzEwthkqCppZdLq6sMvp0UAYcjsL
/s4NsFkCek45KToYIpwf00tXe3jfNI4gQgg/YXAUoYdAWxseL16RnJF3b467WPU2PNtZ/jiTCHH+
ROu6SNKV+g+mCEHAQqlTSFlxfJihSrh9D/UUaGDdQObbJ9PDMSJ3iYntfymbANNGGaINaunrLdxA
dj15FZ5nemMOcFmJxR9VbTpm3B9GUDmyVPwT4uqKgtYA/85JeljMVOhtWJb6f01bD+GsTo6+CNSF
9n2VDpL36FDlT05Qt+UiebewG98eyGE//6m6UqOLTq3pMmLfOzKTa365b7xvkqGiHvSaYfGocu27
DB0GZiqEDtNSykIffAUWPLrpY4HYXiNML3Bc29qxFKOE8dbP0ncup9zuAs5JTDteyUVxRnP6K6dd
z9JnfI6uQjnIeSkRGCg6hASaFuux2JQCPpW1DLPLYEcc8c9cAwsCyoiEd9hwxMWfuZw0QTJoQMTs
MWe0VznYjgu+brZGKoCcCTqdNy5SCiFgQjtpP3mvjGrvDwoXRtPFUdDGfzU07SiENs9lSNiclY0i
HJf/J11yZ65A70wgUzHxNqHdAdkGPOPc4BUbD5P/R8eaVnJssscG1KiUJQI8nEB1psdf+ijn7V4C
epaKnhVfqkK9typ9SpT4Nkqhdr82PTJILDiFa+mHdnx8CCvxQAIx1/34Jqczheb7DNECpzZlFeXC
oRBSflK7Lpab5zcWErphQ72uY7uKG99u4LR6Ri5/SC61Rani2E54Xe8h0ZsYWRpscodDUpRf7Sld
ArgJp9fRqHhb8GkVHrrQzSepRprpHb/ShmhNANuk3dG3tEsn+t2jSPsXbBTjLlWKQgBChFUaJPky
ev2QJuI3TjxnQTX32NzdJs+aEepLoWK6pf5otsC7jM+uDqHlUwG/Re/kese8ZgNZ1MgStk/89+Tx
R7hmmYlaNCvsxMNFZX6bEBbxHX39LJM05nQt0JDifuWYNC+K3jAwbjv5ZU+GEKbolGwnvidNCLJd
MotytRvCCOHXH0PV3XvHMVCPdvVCJ6zcXSdTlmuBeD87eegSs3wNTgZAyiCscsuK+fbiyDK+eqRQ
bf2mO583F3+1fNoA6KzxpWmoLHTVX4BHTb+bOA0EPmaMsXwhKC0/ticR7KdX0tcv5L7C5Jcm75qi
cnlmLbf6LEj1JAv5oWhenyMicn4VtKiCXnyhro81TBkmiRJdyFBKMnTvHoa+XnRuiTsfcWX3nqeI
OgFiL4yAEdyraiavV64MrDQ0Ce7nvU1EUAArORJQlRoff77uV9LJUzF8rz/FnSwKKWnLyE14rehT
KlW5nxs1q5Ja7g/0yOMAu1B+LMafIsB9+vT7DdWX1sYDlpt/WRDEN3PYBnGZpfZLBzo+G4GLoAF9
YvbWWqsTBsdRg1FpWfltaaeqEv+jQ6Jlacx4eh5qLIpU/6Bmr0xJRUw/7jwZSgzPJzTlntn/QKCR
NL0uNubT8e3BI3JZiyM5APe+7TRysWofS+mvMMyJTp2rugvJ5nED9Tg+Aw431OJL1B3K1tXYX6HH
aqShLdru/gxupDsoeI4o1p4tshGzHBGJ7IOvUuKkFir8sV2kHIUkoj8IvuOddJy5rKbVI2fDxkxG
eQ6K8kh3RcguyOQ7wCCIcKzHASVf/lY22RwHwlZYpmJ0/Jwq1UinfIKNcjWg8Xk9RPM1ene3pr3W
5jxNnhUP19qF2gSBPg0VwFHeHFORe5IkTUAoxxzX+xqIDxm8oOuqjpSyLZU6ve76j6+7YHx5+sLd
42M93suaISZ5rvKrIoFZSonQJV8QUzUbv1Zpyx+UN6PLSWGFEQOA+JqVjJSIdkYK+ZDmUFicD7q6
U3rS3gCsFjzrbL/WICghdh7VhXee/f2xsMylkXTH1txYqgpKxXeYmwu0MuPQEOzjG6ogRbACaC28
2aztIVM9tNGNBePLwr57ccvPMXeQa/cznGHrR+lv6i748ERcj2D4v5R7OOHndtGEkPbox/nxqQEx
ZIqWGZDXE5F8SJ78ffw/aqDJmwDB88WtYpekBofAPjaiN0YKJYZkvY7Qh4LuEcWA/XNnkx7YoucE
enbQzuWn3PZ/vLYvtq/4lifpvUeaMGbf59h+B/LUHgdB6ZL7RTQ+P3zU7ln8OfdZfvLiVNIgMyBZ
MS7yre5+pK3CuEcQlxfqEkLTurF/HNn2UvS1P61wWYAnDd6OMu3Me2VLjrSk7haI+18d2KxsLFDK
fyHyNExWovt18IVdgey7QDaHc9OLL1DK1jTWzYzK1dE99eMpE2+KdOcUMMWO6c9Zh0QPcOZxXK3c
l2hMcE2xrCSNgGVO7lpSaeu0UmAJTdrWaTP0b3jiHml7/UBWM0zP3EtECV3d/+3K2LE7hhBPPsK+
fa/Kldm9+b0LU3sFo42rT3n9Iq4LOure3lnvV2eXPV617IzrcrOwIcJ37HRAfvjAUwKjUy+gapL2
eH5J+/D3Tzthn3PZ+BTYFhOKtjiHDm4XlQc6eZ7rqTgWEHCHskGkNFJLO2rJ00CH2uDyu0Zl8gR8
quLMnk4dp/5+6u0fKzWygwFjNCxkyCqlXz92lxDzFRYDYfpM03n5RUBrBC3XIhIKXVGzb9AuciwV
u+tA2i4imlolaA/qZmqkA26yhepwclxCxwIaViJa3HZ1utJl34YAum9Rip4kEM7V58H1x+JJttAS
1tCXwfOfSUJfpOzzTlA7V5XV96IuK0O/fOLBZ0BUPd5gbJNSgRU5uDULjgcmfXtNXNKgKBZSfBQP
zWVuTqFaH81xZ9Ha0hmnKmVki3eRGW/gkklG5CqNWIAyu809Qb/9UgBBPZcFdf7KNOGJCMEtPIlX
HxGzW5/Vba6ohZ8sBgPb6rhQMBYr6O6Q5Ud9j2F1xzHyH6vhiHp13Ys3IS445/NV+9usqLIvIQKH
XeSfMFkSx9Jx/yRx/djFbJeZ+/1S0eBoOUWszef1q5J7+hWGio1t1WPC7OLetIwq4Juk4ONnh2rL
YMkQswARmJ8bs4l7oV3hSWiMP51P0CBV8dQh7MAtFTuDuVUEjVeK2oT/C4NYv+NHPoIHX1jrGEDH
V2zH8QIJbR3QUM7CmINcdpmeYvayorruALFVuQ9TGe6wqub03PA5wq6D42wNsnDpS0c469wDLpIE
lubDc4DoOSw994c0OnuFYJ2HqV05Hz1XtIhLI7q5lenNrAUzLxKG+EZiLzR6q8MUwVo7THI1f7JN
umhOxf0yPxhuJL3Yijqlvn4spV1OaT07a/h5s9UPyS14dMlrkG8ISzJFyC3yEIjURUILQgDqChN5
jn9rvB+ek1BCdnDQ4kXlGtwSvmqLSscFZWT+eAwwiMr+BcOAXsQa19w5rgBICQFF3wiFhRpUpAko
HByxfREQGqavHHOtWNZB+pKBPd5IHKv7XGge0nxXXJ4THlANKSbajrMumFtWQ/CFBrtZpfAkZQdK
lUVAXWZiJnXFkM16g2fu6BA6hjIXCncIAkNKbyEB23b2+lbFwvFpNLu4j71LXlSaEHtsU6MHbtNf
BLACEAfEn3ZTBc8XVcoy9/UywZbcCDxvmTAA0+V9U1T7b1VP3ZEMavERU7CpOmJDg4id2J8WS+0S
OhZ/W1i/XvPK33D6305++vSYeNaJJ68dGwiKiXXon8MXQgLiNurCpcnHxpm4a+V60gAL1zgz6g6E
gWO3992HRkvA6vpN3VP68/5Bx9goXqeUCKFdlmw1UMGZ58GhmtGsc8vz/L5B93HgUaK815bxIo20
Yk/Gr0tNC4InYq7q72qa8haNBxrtAb724UOFmi8Y4fvWhuQ1w1UVBPMMd51DdFxbeKJI8xq4cKk+
DE7gHlZnrPBE58kEhKDN0loee6BBlp69s1vmQwbh6uWJY2nF7kjcA1gGATST4aFnE0L2FIQVSmHi
KyM1mGioIsljTATLZb6FEe3lYN3Uadd/MfQm+/nfWmWdnLtHDs8OHeGH0V5RvAzdQxnl4TmcBSff
aQ0gwdyttxvQ9cXZqpnWH79tRYZa1YczzZrCWqHkpnuYEG1817TI3TW7tGqoE+b9PQKOYM/TCOcg
RTF2BX6yfKjaXrBcuZf/7ix/RqIKh4d7+Z7+fxqAZLJK91dGx92b1k+oxC+T1p5yDy9YSIsL77or
U/qkbgT5g9bUjdMnzPsS8zjBwVLVbddCmugjvLRn1EdztE9Pp+6wcdbYwiW30w/59+HTqyuYHl2p
eQ1vMnIJKQKAmCb50VBvVfsvgiPJBo9s/ukVOmei2VRZq1Dope5sT/es6XZhrJH0qe71M9QnN7bF
zkC7Ajw5Bn0px9gNptm03NMIQl3kA1jGKIFELHKldD/z80JI0HveoUyjsbBdKhsrIhpIcV1c/WfT
qcMXkXd57Q7AuI/XpvZSW4kv3PARsBSIJwYd+V/bKFI2DICQFZhoEA9byAPWLE20TpcJx0XAK1LM
nKinbaFea+kCr7zzvH2zv40G5JXWt6hzRaNX++achaFi81rP+EbfOep3hQWobNAnBuBMd5o+4FOv
fLM6KOF746ymTlsDflKLcAhS0KFi5lUehOKkYusshjioWmK48O3BGC9adRbB8tHTrlZGLIsKimqI
SW3Xo6sMbCkFb6uwHfyVT96aRf/n48Je7TR5Bt6X8m7pGnx3ukDVF78CoX9fz/M6+uGJPoHVlVua
CkW5TwasMOc7Gtgr7FHwAYe8txiq4DYibhr6HvdewBJlC6OgjIy0VdqaSMpTqVAzgo0YSkwkjgFA
+JIwtB46rbyCvUEiINNOi46hsz6iUP2NemRoN3pK2y+l+OXCfQQ3QTx6hxOqL7Ixid58ZBnvjxlR
oSfPPpvJTp2roohUBgoYAq9JcTUIs4CfFyoA8Kjfo3gJn83QUokNhFgX12Rtcpm7yJ+gYIe2I8g7
9TACG8V8dOwHrG5p1HZGISG3m4nedWJIYYMd0G3IGK+1XeNW84NlXK36aUejhlp2v8S5Kb6v1D9q
oCXmRMra70PwcmXyBlWINNFvCtMv7+lslp2nh0nRTwfOpYq/zD5nKJHmW+QuMRk+8lFoMGxczlzy
3VVd6OXbSHZUeNIsDxF9UU4uw9CmSxUolsWRE534m2QhnmY3T1+0eUdzr0rpXnbTWuJg9nldXECQ
VWQKnEPyUZbsK4vKkmPbUYQfLt1PCl1DXtITOPC0RldT86fY+3CyiZ4KUXqenxBa9MCOP6dTi4yQ
macfA+jhLVwr7gX0XP5qpReSTe4UF4WrUGpcolzV4aFrMD7QJlja2CMVThts4JwIxe+4aSAmuvpd
GYmM7TOTR8rsdebJnhNgdONT45LttGnHAhVY0+rBVYuDd/18ArL3DL3zy348w8sxAm96kyNoSHMG
d/plbhakUxHwM6Ma/cqO2JrgqjSbpwBoULnShkgEFPEXkFrBRg6m3EGyumWVNUJLmY0as/PhyK6q
F+M0nZbE2Kvn1/Xdr8Rb/hZLX03L5P6z7zgkUqDe19beRLVECyksvoNlex/50vU0sGlxi41V4wOG
H2Up3W4FWP5+BGH7r+kgArOP88e6xrCozbqOfSL8OE1om07nqat1d8mm5AVQj2D7nIGjrujxMaIS
pYRfaDGACE9sjjus2KkCKh50tqmN+8i0petgX+1+hCuvtMxGFy/p6ZR2PAVTVAiLjkD0pAkzEbyt
52j5ckL0Zc8SKBSk/wXOJljlCpVW+u7iM1tpfbyxLNLWFq8aUhLJMl+yygAVuhaGq/foL/GHhvep
ap2MRKoAGTPBdA6NazqTcWQI3Syd90wgwRegF1c01I5SFWbbO3U0I7Iaf13ZFpd+IbfjXKIVhH8W
Xbi389JGwLznWjrwFPNe9gUkc54kSTd/CANxOvHKm8+8VKHpPm8eit4QvS+A9aIGSYAFmV9akNws
0qe9+e4Mym3i3dM8w5A/8S9iy6aVzqy9p7LdLSwwb7ICN8+icjoMrXFl5BUgQqEdA2pR4tIslOR9
1KzzgPYnzZOBmeBBBFKLQZSIF8TWEVARVy4tmt4dRJQSms80rA6P9Kf7mU8Z4M1MHbrN2AcUE1HR
h8+magv5iuEQbEMvCRx5pn95CETEZHGjIlKbqkYcDFPLnfoVc8AZnrM/RXKpzjDSmuL4hsEOdRO/
ri7fJr15SY/fcf4Jwf1V/w1Vwly0/7rGiGG5qugYiJQ6p0aDOhNCcGAUyURypkoXa4kWwumsbVj0
4qF1FW52Wn1q60nLNl8ShV+xQprWjsBaAVmJl3oJbf/tPGnjYijcCYItNW6c6Oxlp9XlzrpA3tw3
L6M7SlY0Ywqp2U6ZnFs1jpZBTIweVER1AWEVjq/4AxrS+ORebewYN0+3EWqns236zlWYvFg/x+BR
RKntQwOr9iL0jy8QQfiySYAT0tTdWN23mIR2HAHhf7NOqM693fPSipU23U6EmiZRAT2saW45NWq4
yrAbMo5yzVjpKt9/Zo0qajkTSo7w9IjW3APITJDnj4m+xW0p6f0bnX4cwG0MyQ/etBOr/OnTJclD
tqXMyMcFJey8v7NvrYztGWK/L7f94zT8GatieemKVTXVhR7OlYhYfDVPF2VwADtHp9shgt20i7Xs
ZozXmy6RQb9EA6USmcD1j/AQFJzTrEIOMTBNUShwaKwJkjBLFQpthCxOQDwvcwkXsDjBEa/OtmrY
S7SpR7bnoRrBwsR4fVdfDaO69iqrikoxDAUVHm6+5zeVK95J/q7ckK74BGlKXB5KEP/JN3fUWslS
iObhnLpfFjlRDyNbvKXf9NXiVJNlWW1lox98koT8yk6444S36adJqGjdz80rRbwWqwcLn6bwKGDc
6NJl4NYBDQbSfTEa9iWnlcXRuKk4uEKOqRaAv4Ini7SED4krfg0448RgsGiHOUrrnK4T6zW9jjTk
tMwo4LuFZwqrgfMRUyUFZoecUllRB0CEm9VOJ3maFN0aJUun77uiDZ+et+k19smXu/mxjOmRoLkq
Xa/z7ofY5tbXhGBRVNv0xDjGRg3e64UWsD1JUsVK09vJg6tUfZgSaV90Vdqh/+dHOlont080mAjb
WhUuLu6ofw/D3O8sIDeVwickOvaoT+dXcl75OMWJgkNoAYgfWaDgJMQvD/KAPru7Duy+s6db+xnF
BP9Nl46fCEAB6rqbcXbAj1V8WCaHKCYfABgXgq5GJh5pzh2iYlCR3k9st46PZ87iYqvAORp5iJEn
+WpsBeL8yl9tFo09lOBQWH+rWZj8yGpuvXsnrZQLnPSbl94bXTv4VAROgnZ3HEvLQyafnCaJKidt
JvidF0mANCShSjPrhwZS+wnJ3cK69ClvGuV6VzvAY7SWYRNnrKY6FlslWw4OsTOHScuq0q1wa0LJ
aqP95+MuQLyS3e5eTJLVIXxrjVRTaBJOMDc6NlJZ4j7Nlocy2mTxIPKg47V8bSiPZfZZSG7nw5WT
fksIraMSuEQOyQT5NkxkonKtcVulox/oxbIP8GyZZxPPxX93Q9Bf74e12FShzqhCw1RA6X164WGs
OIFbrvqT8drHj13Yr4+oYMYr08ke7A9rSaMp3ME/hb2kPwX+EoyJ0S6qF2yhUOQNl1js4CCRnNbL
i8kfO+aXs7YWIyDoQVTMTjVSA/zdfVvvF36gji6w6Rnx0nB/FNR8C7da7Y4JiWYJa+anSmtfi84B
DmZzbfUKRhNq5snVhlyHQvrCmHA8aXdyLzkDIrcaM3BvbKZLKR/AMQwp0/mBFWEdgQBHdDG0jSNA
n0/gQZCkUUxLIIKnceiLrdRMDXqvZgOPVv/fAKrMB6ckh7utDnKWDBl88pD3ajo82q4GawO+IzjE
9bTZuR8dvdovv5QcAzCy716vj5Wjga96W7ww7D8i9kNQQsN2QKhyMr1Z3U/Z3wpFpkay6+aYLZf1
4dTvwhyaaeMjojIQm4gjQ0T6oLV3U+hdTosRt64boUlNZyk3c7Cz+rnvUS0dOlNC07WruDcqkiSs
b88acrdoWV6wHCEi2DM+UJSbTukQXTvI///WZU8T+qxD8XwYCUZFfaI0NZFmJb59rfxdm7i5E+aS
tC9IgwYun8E6sx1Q8DwY8PP1RcdKowyPx2GgH/0YfKjS9MQxgzLK9NFYPElkx+N8ubDV6aupO+AO
apUYqIg3qn63lZ1LRth3fvR3QoLTmuitkLUMV+qMOaYtdyRj1Idn3QuNYsiS9InxN5UgBbN7R3MQ
WuAlugws8qMipYUy58O0SgZS/fStch0Ci243I6RywaMGJpog/K5jqfEtuNGK1Vok62kkJhaLTZsM
G8TXTevCEneTAzTDPf+VnsQCjmFjPHh8RE0yEZbffEoj39tK3fet3Kh7YPuTaif8gwzCwnaO4CD6
NgAIhRfoEedxuwaVuPgbLpKa5fgfSjWPqFDI9NhD/l5xnQcKIB/Rr5OrbXBfllRge9tj5QFfvhYN
+LPs4zDtH8GwJ1wB9IchRMP6kLZ71uyYMq+jXeAi0UNj392+Yh9gGfrieJJu8pvUDl6o7LlIzcuo
da8uP/lz2Kjr4AkD6eR+l48HIZd2PvGxfc/+ADuGmvfHDi/YIBiMG+wjK65KDoglQ15ffXnyBF1J
nI1htIWWpwy6uUT2wy9/XNt+Bx83AxagNO8HzyoQQmqoJTM1OpuDsqFGTnLskC4yoIm+z35nJJQU
fC3uOuLmC09+6NyDCTxpeJ08/72Lcc8hpEAjAvgwRHEdknRU7YpIWm9wpRRUPHUyM6ojLzny2BcX
UU/l8jqFOfoetJmrMeIkllg59IQIysTjyogQHCe7+ZqxdSEWPFl3AhpjCWfKbG19+mN9viBpqf9j
abw9dTb45tQZaM2mf2VV3+EhfbYMTLDiTQC86/zIyZ4jX0kSfu/EOsh8Avx/uOn55KaslzNGwc5F
VSwhBkWE+qaRdp50Aq+lCHEPx9APfkHk5DIHkvdVMSFl5tu39lVv0LDHgTwPwraMW4I0Vb0eoxZn
2k3GeRnGlHdkdWPuMuE0T//Dq2BYnVEly5oPTDcrzAQFGUvlWS2VzkfssDvWBLRZ4cSuXFaDsU2u
PTyQJ6ghZcPqH/CWV/2n8gRD/6NlAJwH5Fla77hIVmdBYpWpojZmY9Si5TaOIgbY8rqnh9UIv+cm
nUIqMaIRT/6+9YMExDG5P7LvrwFVe+UScSLHMtxSuMJHhwif3NSfFdYBueC/60BfxvcHZrndNouZ
aqYPES81E/5FKeCFB/Wooutq8q+EnAg1zHKVChSte3bhFgUecmR2+M7amDBWODzN97oBCkTFCySs
Ld1ud2v31E0Xg2wW8LoH49rsg2kalPNlbcKzp7kaw2xHia9NOKPqrGA9Um3oMh7Fo9y9e7t+QUBh
5qZLWaMaCdrGmSfdJ45cfujzpvUcoDFp1mOcXuXISElIe1So7si6Y7OIjZx4D+aemqNR70x7Bwwp
dhn0CprezQEu9bIsRWn8/3yT8/KL1ldrpx5ks5nHfwPOVnmpKBc5HPuYssvzBYYZjSE3asuoa5nA
CQLTyNFy1zuGBkY7fS0D7W4FxEiPjk1BD1ccosq0dPk55Ex4E5J/PSdv/pmBvBGZ3xdb5EWhFcvl
SiTvIXokFx5BqvxzMrnFs0w7m0PW564wSoFAdb4UyT/WvsFmNMo76LM0Sn22XABU7yfEa6lWv1Z4
NZ4rZ5AuRVCqUzEWv07uUeTkl5o6RfRIUprU8LznuNAWCpffBAfzywv7NiIyhpsndT+jMoNSgvxZ
idCsBEe8mJ12kHGBIhmAc8fiuWmBxRfjVH8x8aXz3ri3Mp88eP/onKMEjH4ldIUAHrwjVlwGUT+G
XpBUPxj0x83d4CW2j0jzlkHnDiE3KbP+isywN1ioa7WlD6nqlakcBLuC8VFPFmIaYMmshvidhEOs
vDXS5AOn85LNbM6/V1CG3qQtahBh4RqfUI5t2Fm7JUfC+A14wYaxhk9fgyQ3dyib+RoD5c5/tAT8
nW1zftWlOxM++7GVAL8jY+ailxw3IUc10qJHCBco/M5A03ExSa3rPItN5nfWLHNF3iKSWE7kwGsF
fl2wDIuBiuvz/p7WkH4U99ZZSR/saR3wxZRpGF3N38Yrgzj4xnnVbLRKTIj1sSJHCxPozuyVHRvo
LOqOAlG83oAWJ8Iw7scYqkHuTq1nqoZaMXbmMlrV3AIgykECS4eXbHwRaTOOc3X/t81x1jy5ozm/
8yxMhfZLVss4jMJaWJIrqvI05ZMhonMHqCMIKpPDQEs3d5eSzDN+Ulu6hftZE9fXEDwfPkdxZB+3
KNbrhJIEKVggJqCaT0/ROcPexLzEg/MJhE2uSf7G+e2BEp6VJZgN4mW3bK6nFOJLhdIa+81GEdvR
+AfnfIJfZa60r3fY/JnNgfRQBAr3cCDVa95lHRaQ1jCBmJ45gr+qPYYbD0AZpLeIiXtNdbT6u4x3
T5OlNQ1flIvS2EyGwR36LM2tJMMaR/p+6jPEurbjo0OKivDu7WzO/+Vq9SNKrDbgG/tJGL9wxz/E
kq9+GRkKXuejremUedtmriV9eEIVjXXpQBznDQ9XEQp0Gk2NJotHkz7qkhPIUAIwS8jjq0OyC3aY
Dk2VVqhZ8ThQDLrqZSXBh7h2z1HwFwioP78ETLwQPluS0C2LwxZYI+fEKm0CpsGeQC8eKkqLiXC1
z311Ahgk92CZlBOCCCoVGGiC+IGC39S1JPI76J/kWOE/fP6ZOqp5lrLngCmvWqnYlHi3bGJo4WAt
V7tezhNCdNPNIASg1EydgcixNf3z7x9gi/3sFvLXKdnyPxDidcS0dbCs5v1eFdHkd4bOPO3myr3h
15cn+44rmieW3sNH5Ri1V6xfwjyjvkIhUZQJX5t25+mg/l2deLwy6oi5drU8Sf5RQmynRaGaSM62
ejPBxPSiV/bkNmRkhkMHe0G5uSMpJXVqeB8/oLlMp10tvnPdtj9mPxKjX4EB+ePfFGABSCIpnLHQ
/ZtAS3VIUR45HPjM/GGy41YfNmpEnMmxwPfslVZ4G3a3ymZhdw71y1Dxif5rQvYA8ToieyTDoZK9
Pl+XTi50HjlNtI04TXtKHIaD0GXz8yuTNgVXxi0J/2lsstK3dIFBLu4QDmsNjuVRsXfJ4zc3D2Ov
nZM8OCcdGN4sYf3qvcEkr7CcopSEw3GAxocJ3rawXB1cG7s3tTvt3t/ojL5Bx0gACaDog6O38v8Q
OxqYo4dyHs+iYLLUXvIH1nHHOEISq/s9G4q5eG2vr9ZT9gGcEWIAO005jpuau5EQogFYotldA8LS
oWh6FEyFK/ICB1zmHkki6W6JG1LIi+/7TDHlTz1tpg8rmCT0NmazbmRGqwkYhKjpPlT9GBbybSp8
xInTBGdTs7m2mKOmsEf9RCC3TOYWE5oOChVexV04+u/gCDCSWnkx20OVMJvoxaCZLGgMKL1w/k0k
I89jcl/FCst/+8W0E+2yKL75dZCwOxihILN4D281wd35Ow8B4vf4hovLh8Mvn5n+A6w55o3emykw
lfAPjy3Q1vG1bvQ5FF4IvSuud7TotjVE51sHCRLZdOsqEAd1h904CqljxW7fnGxCftzHciFwJ/rA
QbuuXdRkv9WzJ1J+navK2qPRZiSMqbFhyP0gMpnzlWap6yybljYHuT/eMbj7kUOI9ylDKhbyh2AE
uCYVvTEteDcjDU48P2XoTb7hvKjUgu5zi8a/eCmaAomFHvJn+ZZiJPcNrd73FjWJe4dFy3ZTm+4j
tahBUUbTCV3+3XOuiWVNw7hG32/sBdJhotLRIL7fHmSGxuj1pTrzlmvgDDHow9W0kXtRX8bbPZZ1
uVSCaAEsGFBpjlNAVEjZa/oTRlt5pZ+vCmLGbEhvhHS3SzC+edyJmH+P2iyWYKhrvmAnk85cpOBq
nrxtKOP1DTgpDEzd5MXCF6juj1j1tyORV06hZC+h2fDgy129ocQdR45hYxFHhrUNbA34b4SE5XlZ
Z1EX1NPmn26jX8DRkbatS4H3J44VkrfONPPuhqFYvF0askoxkkDyYWXLM7UMNyZErMqN/jT1BAGX
MT588Wx2ZbkA6MJf9dZ1J8E1Tuo3yDQwZajIrLQO0PY8JZuzrPYd0B31VinnptCFfIrvi0fbXarQ
/z6Ha3+4fi119W5XijpnXubztAoZdbmignhcFGejXQqm+i19QFOIoOIbuns7kfN8KcT0iyji6Xe/
q3kEgbnJ9c9kvAlukSWLbS3RuWzr8F3h6/EJZ+xRwqqxWgbv0m10qUDMNBV+3YaM7ySRB9qtmA8J
hrXiQ5oYhdEj3U00Tj6k3YwfBwbnD5xlHFAlUnu1K9m0I3Z8vJW3k3MgotRpC9EpBnJjskoBlva0
cHgoxehRSKkCPkqeHCwPU9l3XjLmkdYrtWeTN7/cAZlVIv4M1TMSM6UK+g+JSM2lhB8H6GbdS6qL
nJS2LH5WmrmBsIocI0A6mTbZS/dzDMXYQ0LihVJge5vOTT+WNlzZ1jR7ijmCjPeCvsQfYvGQQbOq
4OAOso2fbSf9IAFhqLYH9qeR/R/ikHdJ0pOeIvMhaajIEFBbjdQOVTHSBg+7ju8WX90w8cps7p3o
eZd06vzA5BCPSRAaLUYOwBdmFm5750YqHfIOxkZPmuikoby53Uz64QSzblRAdx/tT23z7pTk3xc2
n0djC17IXlb2A8D7OaguklTu9eyU8Uf7ddg2vJIvAZPGp3CljvELywbsG6ICQnJzvtV+B0eFl9Sh
Fmkod3Kzsmbk/Q3hg0hDKsk9jctNvGwPmEjwkKtHX4nwDuIx4iRGzi3MkdrIiqle1UMPb9XvJgyr
1neSdqnmeHkE9bK0UIRoIaCRxApj8yHQN3n2Z1D8XPB9NnDuIFFqEQb5qSJ2nsJXt5ei8hHWeJXN
kjPFAjMpoTuLciLNbmAggKWBMbLfm+p3JCc3njstFN9UJiF/pgK3NWSaYbf+NUUySxURlt62eEnO
cC1uLYMWWRngrDD4ogFnCbmNAT5u3EsnbZ2PQPoCTPLHL3rY0Dp+4EryqxkpA9sPW/Pf9EbkwRQQ
xBJPlso5mLmqKFyJtBe3Fv08+XRYD12LW4VjnXQv8VPWw4sUiLKCOokE9xQRfIBJmpl7exTiYYUa
9qQJcpW3xBBADdfu0OCGuZVxogOSjyVWG1470nvohYz/aaJP7vGHvilsn5t/gZ4b4b45b0pQ/vNL
gUnb+F0gPqWXOt5r2RshmHie/BB8h0B97CiB4q8GH9+mybsyx1MqwPRMMN6brCNuYb+IUgDjVSbs
G9cIfAMfQi0uWOHS7sEw4evnahuNK+raUIZE5Qv+pfiUaUS2ZgDNph9NcQDu7s+RqGKsXqptNr7d
l7bOM0WDj7apjdDU+y4Q/EsygUTzU28zwkT8M0Tfnj6G0cSr/cFoncO419dZwpI0JGhwGyY9Ps64
KAWIVw/aZLdTJd8UOBuAjwDPmYQrtTjAaVSUJZLU9QddXdZT+2v83RyIr/iVD1GOV5jDo/es8IJC
eVVlzZgQQJIsuJVdt1QPSWK6PlVoUQloRfyQiATgoxk+J52kfXYZQKehAcJGJlOpu3uCflgtYp6a
12SEUewNpoalL2kuUCzOzp7cMyrejm4bWV145zW8L1+Z7BGiEZ5ackVxs9ssNciPl4+CLQiwv318
uEFzNYI0ww34V9qx0qE8frSEzw0DQHzKzW4bNqFlsl1QTZo4I7TSvz2bbiToSX3+DS6dPPEmkSm/
VhAfxuRrxJnXAmhS2hV/a+99/0Wo1Orn5hjfLw86sJfgOYulbyNJwpxOEcK6cu0ofaAN0ob1xoqf
4uCUVN65s9gJE+HAwQ1QXUcP6jDDBGFY7k2DjupfLhNaKg0ceObHUClVutAplLIkC7b02GOXHFHh
F61HJpHLw4l3tZT3Y9BCtFBtPhTL5DxFiwweWLTfOEp6d+y5Bs1Qn/yw3lR/b4XINqGrjsi52d/b
lktDpQAuoX29GWLv0warAZx22mTmnFHWeo6gaO0R+uVJ3XVfHX4eWpRCKxkp4r8sUz+LyvIooE+L
RJWYntPP1iFSKgFDcQ6uUoe5T3ca22MVWy4daNP6JDE4szSyR9Ne6H79YkZkARR8P/esHubQgaA7
cD9PjSw2xWmswgEgLXsz7R6zo+ar3aZG8EgEnvM76uM0AnIDZD4bykEVf69W9C8KiHW8a8RsNrgu
haBLQKk7Bp1HOLaWmZ+LIRPmRGqOPfocCjszHYBJQsb/FlfsK7tYubDYJAqcOZXnuOb2VoJfhrad
ZuvfDrURAwcwhiVzy3f7IEu2/ACjuW7nVYgOReyxMjUi4T/m71gG3sw2jP/cWE/o6JfhVYtQNroE
S6z3jrm1+4Ci39pF30fJf1Q/+a8R6RsMSo9X2ujnuDfSd+X8t8hHze1x9Yfy21jg5XykqDWiVSNF
Y1rhHN+meyXGfCIf6zXp5QaZap217hToNgGaTRYUl1K5eoR7AitXTJTABbJTQ6LVlv29oEdqZauy
deoz3bi2OxcP0MSggUPNJS/qAnQNBiFFZ4AaQYvzAQhtFWLBR//HmGDhxMwH2xGPoFwRCeqBMHnF
oibzQFu8jTrANnRM4jQxOuecca734/vkhyzlcqaP+wAAzan5HOV3dsS1xXS20fPMJFkN/W4hYd6S
fMsg6r7QwgwJpOCGHeDrDT+eZKyA2GgdKVALzC1acJkD0jlnEARP6hupjb8du5h6OWkYDplr7w8r
B+tFpd4YUF9Ueh5xS9hscXvZrV/XJ4TsI+WoZTRlRQqSkxmFwQaOjvK7WqWirniEenyb+LZIv+Wv
9Jt5fuALBKlLgGG/GGH6TypKkZ5x5Oz3J9PRkj0PT7WCvnYUqSFBngT+7DE03avehplNug1+GzwM
ILJsX7FIRjfoKq8Ca+m6NjSV/o1XMqXR6KEpsyKU9xjqu8GiOZ2gVwnAhoEQ6orlGdgFQ73BLPgT
eNmymJh9NkyTp9c+7P83knCcEc5cN+48G7tExtxYjq6NTlgwZUg83gX8EonL+3HyJDH8KVQaAXGv
V35sInWDQGACjGHrGWnrjy+rV5vzPaLgecDAka1Umo0pUAv8PxfRhWEJE/3xV75/dm+BEr//EF7y
cC9hEB8h4bDxaWU2T+ZFBkX9UiwXSZgN1igOXOwfQOQpEW8KZv+5oLg5P8BXG4fT7LkA9lQlacqA
ptP6mYpStZuieCAuvaBoa5sCReVzj44Jiqcqj5lb9IiY7hgxmPIFtKuKt6autZetIacH4vLCW+Gf
HLgfhp3DvB2yJUjiLbab1gE5fL8L0tRMMkGCVxdLxaWx+mrz7nJ0cUVEqPdTdjPPcxTN8AOVOMz1
U5FZxm/M7AyrQ3J1G7xdnLyA+FIvw81JZ7Ei6KYky7RROPILnsNfaE5UV1Cu1BZAXbfJHE1PoXc2
zD8qHvBYYqUMDiB2Hd3wLWfw8Z9EbtgqpO/ApnxgC5fPaLBFANtrBbx4cRJ64zfOAbhz+KLQ0JLe
hvMWDt9mqRgxaECqU2BFCpW4h6aBsLr9/+uoq8NNTXMb1C8Pix/2wleYsUt5jdTfAQfZKfm6EVc0
JZkk9GHcUDVgPn0umYD5Mr4HEDC4hPl+S24uH2Upq3RyTQyCF+1vqVDhDMCavsFU9gGTCloF2PAT
u66zS1SNHbw5Cc4cYKGCwa3xdt13O8Et2SuHG54x1TJ/SbfMmKTq9rNScpDBwXOhmifMWO95Iyjw
i9WJxeDlLBzcr2kCUI6Tnm66rCMxxpqmAcqetnObZORE4gYiTa0YpAdGRIWG0Y27Qg0M5BtIAU3t
VLYJSkxGGjqunc4MGB5qOPZnH5keGxsYckRA9s+laOujyBXWq1nEyTqAjygmnCJDv0cF1T3n63lF
RZpXGNKmKJWktz/PBCf9wu/mUaOnOC69IyTPc5tWHU5nyfD++mIAYpOxEYsx0WQQxFLa82CqZZrD
eXGojpbQXAeU2q2nLUHcccZ61FcjNsG/N+CwEBUFxaTOLn+onhbNXDhBPapsGE5JHtR436oqM7IQ
r5vpR0IUWqqBFp0P99oEG3sIn+NtIkiBxwICYJ1+1HWAqi5NuN//fi0riTUL/+Kr4tf2hXh4AWcf
K78+OvrdZIZy1VArJHfrGwrgIwI2cI6z662kui8hfnUyzzqdE3OC9ifAHVYbKABaE0QS4OEqkDZc
sseydrtX3a/VlVfNhH5gmagmixahLlBeWrIUy76CleUIS+jrV7sKHUzCI1Rgix9HFBFnCRxu4nkB
OkDmAsX+e/MPC44SEJEFIyQpVkvQwl0YyuFKmbQi5Q9W4RaHur5/n0ulw3wymTCQAjzb1ZFVLdE8
DmazLu/LDZDDnhRyOmyikQa0YjpbMm1To9eER71h8gRo1UZz0WTc/dxskYru1ilRVi//bbo8th4f
IP5akHA54ZJ8HgMA779VBZJvE8/QI73V5p8ZXoFHqjpsx3Q1lyWB6OGT7IfzpbQAe7lKFDord7PT
MkUqH71ptSY8yvzN72ZnutzJO+Ahgkmp5ksOD8BdsdY36toYNDm1anBpA1Rtfb5bCEjuFK0CzJCq
m9iTVAzC6yvpVpLzqS6pok/pHEbVjccYIWJ8Dit+8lWcx9CGmzJk3U08bW9ynTWRpqZK4B98YNwY
6Qetyehk9/DYmUvSLZhtlEkIkrRNZRuJLiwUIPHEPeyLhgFGpkLHSFUW++ZIJuGDSy5VUOZXANqo
iXfORTr2ts2cW1rODk2RBFcFNrEftWATS0qQV81GQfXqazsBbPcPW66B5lnFo7qeHWTLW/NCNjnE
Cvs5NwzVpZlQdM3UMvOU0pYoITSEkAl2kUg8DobHRbvXY8mWSb+FEnorCWzpvuZfSK8dV+lB67XA
V5a0Gn1mBhh94ao807YrfZZLR8TLFVy1ZLsR3YkUbYX93N0GZUlN4XEPFPOldQEwFwVk2I/KJriV
mnz754uyz/m2Io2t4Hu3rba4jKwFws454Zbn8TXHVonZfi3Vwzs2AQ6EpBauj5OBsyXGpXf8L7GT
Tna3of4j77COSWYXfYARAAn/gmxqnAxM9lNDAsns31DZCWVpOPeLgMGRXFkh+b3bgN79tXHMDgIM
0QfLG+lMfT+JUYbpsQkPgOrZ2OdQvLAY9ktYwT3U0IoF+gBumL0WuSP6+/wylSxCqUG9+rFaNI5j
83VNZuvvB51hYlaHH1a6aDyfqRBt3IKxcAKlaln2EzZXbksTs4EDw9cVhT8LxU4z54+bqHOH9bAq
CzTSb//GfQhTmDeE6zBiqS7KqlohO3ua4iKBL1Icli74vP9F4DxDQS/EPZFL72qdekHZGLdi8NRQ
Ih3jwRPegMxILBrFSnjfqMlJiqeS7RVyu0OyN89qK5bZ+VyZsGfP7hnXgqpwgKu0J0NSvhWHQwel
HY0diAQehj7v5RVdkZU37qlxMXS8NZhDwm5sDZR4deRZOANMfK5/Vs+oIti3SpLyyLNLXIiY22Sb
LGyn2i9AX3tjPbpb+oTm04l1zoLeuy/8pS6en44kFZiBKo8/5JbCIzijt9Uohq3spCkUVjugps8h
4PKGPYwxrp/ZeExTcCKEchQpLjsrF14dQfTlwRl7CZm6T36NyBvxqRzsU4c2i64A8fKVO+BlFM3W
2T8h78ThMnjzP0xgy/OsZg1xZk0wFgtooRdfRAFyNcADWcYxywUiBW+IioCXsl1xlvuP2VDnw8U+
ZjJsJUAT/Mt3QfkFim8GYnVZnADRDT2vYpuaV5p5CINPdAEl+HhwHLUKFAiGZizXMQDDvUv2rqQZ
5ujCjUvhb3PsDw1yJThejnqFxBiCeFhdxC5qapklS58Qv5kPmqNZxB8zyCaocuYxSHljXD7g6GIA
fM1vb3uMaQewQgLU7RdzHTHlhNRA/wbYXdhdvI1LDJxRNI4buYbjczyur5tFQVFJ+25z38qwEOOx
30SSnHzRjp7nVChovaJB3fXL8IpSoI4C3+j7wiGYf57/AMN5kPxPArkvAaltBcdLxR1bl/ZWj/lZ
La9KLajVrJPQF+IgmNknECdXnc+tZ1/y3s+GU+RXloaOd9EExGRSBGialvlSl5l0BoTUNUnM41/y
Ce1BMjj1dPD4XKuH/WIfh5nrWDWQZ5Z8fOE7PKcWyaaXsV4+yNltWrfYxrC0knx0vqwlh6Xuheo6
u1I/lV1U/eglikfT8o2xSdMBeC97/DBs/EV8n8CPkMPS4Z/HfnxcQz5CMW09jJbBVV3xlV10saCg
IHn0tC6AcEPGzZpnUYEaQB3hdaagz4LM7VH4t/xfdQMaGia9eV0C+QH3H4uFkNKj4H8DB56rOo/N
mKFefWB3TDEyS0FD1eUbGyAXiqUthoy2m+OYEZHKlxlqOEW6JBNYAl7P/dutnwDggZHQFQjzUF2s
oalDFkuiHP4QQUdT0F4Q3k/rduKdCVWUO04jPu8mNVbjPpJnUn0Lgis8zhTr7jmVApjpjvxq14Hg
MchDvXmeevEcX7ERTdhSW+vn2iqStCojqIKS0MEnRUik047DnSSC5Lu0FsDdDk+IrJt6nggCJx1/
kIjlr7NWoZUBTGQIBQM+/xBVXC1GMgALzIyC7+qMvD6U8RndjOjZI1G22XWrXpjFkRAQJfXXKyhB
3qQUMtlTU7+llhPVau8eY3FY1wI93GMDOozt7d4LuRntAXMAh2/VY1Y+0KB5hARCiCx5PCPSz/qN
oLdCLz+ukw2KJRRyrsD5pZdOGg1mrxRu+Q8puYYn62AZTDvxe/9QNHWTeCsHcxaO6105/p+/7xpr
ybmYInWsfaBzK/i0p1AK977XIJLDA2SR68y1G7iLVdka7Am8wTpaFAvId1HROu/Y325hYKOYDy6R
64uTvNfEa9SVK85oytOrJzUN4iDsfudBJcv6bbg92rOCvosRNK1UX58gylRlXfWmNsb4bhunGVA5
6XtzUGnt+xQQxwT+OlekGAbJ/QYB0u63h8+cjoZxCu8bk1k8LlXSe0qU+rguXNR6Xz9pL/8QqvKJ
ko4Os8ySmvaq6kgw/GRqSGCWav35Gd/Yydai0bA7e6qOrgcjwEYUcYZYwd7a3A5fADRSXRAYacbl
odrLSHfjV462f7stNsU21//EiB/z8bT5rBIJ+1EBZJ3BaT3MhiUCCFJLwav2J1WFX17PMkqrsfjS
AxRwpdBtv0ziLpPOa7qNI9BL2SCwqcTGVI+1lRpuDsKcKRGyTvzBwXabDDEe88UKIPCUerv0ylEd
1W/6q/snGQNo7eSUB7OJ+XTluzYghPtMW4+ALO86l50LjccjlcHyaqXL8iiId6tFmbJwsO6Sbemd
AN+fnoU7afhlZJJuJdTgtpu4CMMdmeu5sVwEjxmch+nkxWdJnD3GGQV+akGi6+Jb6XG6grZRUrrQ
ZTwsI1sWRmbkQickgIBcBaHDSwMDOi0/FkM8oni56zvPnxWLD1xpTztzn0HZ9lLjbp+AEEGkAKaV
8fdZHhk6gIryOjNfMsMqvBZfGqXjAZbIN1IA8XbKCBZ9XvcOQwk98QKrslEw/3HvxdSTfykINwiu
POffbi7cLRv+M8p1tYVzrMXAyaTyGKgrMEnEENRmkXy3ostvZfupPKWwC3I1T884d4Ws8v3KGRMb
5oFk4klcdM77vwVuDvmumSEFMjnAYNo1MPJ6eftkFRnqoeJkNM9cJyqmAUoTCpMxN+Hq8NB9NkIk
Qx5y5GLnZT+Q2HrXHaSoG2ja2yK2XoWmJG0WpygUwClGpMhuELA2ZY2vAJVq/0XnukdbBDKFnKvA
YgV5Glt0i0vE+8DJ3u/iAXX1XYyiB6ghIgvNskSZAbHQbuTGyMgNhSNOjejWVVP/4Wj6UkIb52yX
h/w4R8AUmzfbgehb6VEfU4uaceW2QFbF/rynT91CyYupVVuznd13gMUgB5MJKAv2uhEGSRN+e96D
aodyAhPpVquTPVr7ErV/6yKZcfdvuvCyWX0ay4cnDj9YMIP50vjemD7EAKI6gvf0uZeEgQVSHd4F
AORERD/XIuce/LVbcIMdwDJy7sek0JAeDjurcgPQb7K0+eXeHJBuO7BJ9ygG9MVK9VH6kTBUUQLd
9b0zOx9Ow4in75FzKU38q3NneIF89QDmggNwXYyTAg7Fk9WcIe95r8kuX5LUIwA77oFOGSWbQhNJ
GEan269yUdrICAwvygWy67rISEN/e0Ry84C1lFfU3n43cv0VqHET81tKSxSD8W2uQq1BfGu1wPin
hltYdAO0G1GYSTtFIzLW9pqcj/q3ExKajAzZas2PsqZRGUURqkGGgUxt/l+sLSTOPeIBGPhEicoS
HjcGGOU8KRHbCbVoOnusobEZQPLt6EXMnBbZlFe6fHd+HkKmxSgegOl6WiYjjIaNzeOJs+Gt1MYz
fCYw6a2doHLbdxm07tJU9kouG0RBrw80CMDM0imTtQgdAWq1qxPDlil2b2xTuJUtkdDxh5SmnwaJ
EyG36JMVCfWpa6k1zO4oferh21hGLgVfGtQsi4+nwFUEd5kzuyISZbx0T0flh1tR+CKfcPkgcYfP
pSBnrAmKM3UV8VZPl6D3BE5oVI1rMK3IYurcS4LShugkPi8EOSI5Yk2JTH9N6VQpTVR39w3ntVzw
d5WmZ7jaz8ep/nNc2/Uetx1WfOeGeIDidVfTCM/HDwK2ygW8gvtczmSpehdFEbTSzfBonABntKDo
ZJmxlDliY1bn37gshvk6CxJ6ARcpZlnRr4dnNPVvqo3dtalI/hPykbfih3vHfmlQBp7kLTDrEp/2
4UH8Ef8FRAi/3LLdQPjoO5qfSDotKjvvcA2E6X9l4zIRhnjV5qvsTl6tQab/xCem/S5qyrBcBCVi
GLOIoeviXzuQ4+6/oaV0pH9gr97DUWF5h34diM/HF3j00Xlp4L+6ukNqm5/Xx6LvSjKU3tu7q81H
WmDAXBoRqkDAERVO3Rqoc6IVn1eoGYJVVDH2zK3AC1kvyFKi0wnY1kVmGS4vtkjCzGyThf6rTt9z
GaY90Kp3caUcPri+ZsAr1JUPdnw0nxWpICku82UtlLzOuthAuBgBLgmRGPDKqAcr6edkEseKXWKf
Fqz4Iqlvob9iNW04rlqHLx4eF0h+c6BlBqasH9F54diLxVSTtuEWOugQC74ChnYN2PzDgyZviPFx
K35J8TiJoUa0F1OTeQpo9Im7AM3JF/1Tk7xZPHl3a0gq+sBPrPynVyCngIHU4jrwJtt3OOBP54VV
WnkphDGK1KUacB/uhmSQQNNQ8puCR2gNJbe1TH9aXnKmn1eEv48gZk+EhSixkDkDfCQPXC7LNrn1
2AQ3l0b2o6PXBWSiGP2ibFnJ54LVDqc1efw6PH7Q/jyg0zEuuQ0TI49S+Wg1f9ZiNF60yMfkLxPP
VjbAB/rsY24NwOE7LgSY9mK86rX5i/Vg0M6vahm0tcS86adDD7ovtVqNIGU4kFHrzvVG4Fhu5FfF
v9zvhSah97sDPCzNgquy6SlpthXp8iMcnLjacBz6tZ/XjOWcuBT8Mf9mxjQJiAXirpy0wl/u15Ng
qQyuFb+Dm/BeNfXmhK4hAVDqyNg66j1Rd+plu5hvNJOQDf8QxpNO7n0dpC6jsbHXwVHYXgCwHYjt
sKwVhhTPKXSs7gfjeeGmfds8uBCKcjsf2o57g9proWCn3gXgrKXBXiei4WKOF9omDeWMolHTll5s
BEiwm/S0SfWv4z2T+Xp+l+RjBBCq8CrJNoMxvB+4m3etaieZAilPk9ogl/PooFtS444nzkOa6D9F
v1FRLWKg1jbmDyV2ATPOaoxH6u0wJmmU3zP6JJBoDojRtkqalAsiBhePmrdr3ACbQSHNryEfaVt4
OI7cIT1mvVJzxfkuxloNXfzdY5IgLiCaC/5XauWz85s0G6rHRTGUGWYQ6m/AERJIvpNoVHk50r8v
aFEMCPtP5IJljahQ7DkFik3Sybb446Fk4vnDpyQ1PUaw854FkaKdVenU9uIRp61EF7PEcyxdWZn8
foUL2XaXDmCr5tUAE492SILkRbDqM0z21bmNl2X/cy403FkfwzBH5yvVPXVcu7Fki5un9p5Pjg80
cYtIBEqBgk9hFBSyDr4KVc1tCuQgLjrdEPEzkhhI7lirXeGDDKKy28tw2zX1u/CVtZnCEeEBE7pz
hCCUUKigjGbytpaA/mTJqCVEOp8J9OVie9TDZky4aUtNHSj4Jjcst77GJunRKYTBMp9sHadzhte3
Kz35Ftw3MFhdUuTzKHXxaG8gF0cmn2lbXmLnRvA75J/MpYdsGczqXW9U4XeeG0wQuRep+78RZy1K
5cjd5x3Bv9TjkhL2JPIJtJUJ/pIav7acWRqS95kGECvOAhLrGMJ8WwtyufMOhZlLsNww6ltw4tlG
DyXEdgH7AbqRw+mf2YaylbMh38B3iBZzPCQXw04oFCg7S4CZ0Q4ne6QZ549VKBdSPwQ8erg52cDj
vzHhroWITaut8AdkYSZC41YoPuJoC6bshUX87sgNSPZBlpbwUn+/Cv3HSfELZSbpUZcOkIS7/nTG
JN8IiZP/awkU3++qf9TAGWz9ljYrzuooAvH3dQYsPtr+viHjnRdmM4Nhy3jHGmuDX9kUg6Ax5kgX
PPjelN08+OvvydTiQQJsN+e8FD5Cs4yetnHLzOrrBSpPtLg9/30hHkgUMWMnF/kU+6VAr+N3IuBJ
qzTngJ49MzuiW+bADZxqpUcr9qioTIThOP3TQzae/qh+LPq1BRSe6I0YqTJcuc5wSXjvWJn/zZ72
gxvUJORov+q8IMGbogTWUszVb7c7AuuA/UwQNTXRScLHIf7VpaFkJG2u8TDqwp717OjtB9KDBgUb
Q9RPvrfcX7r9xg3u10zhpafz0cecJVj5WehnsbqSZ+Ax/mPrUatwHlLREd86/L5we5CPrg2Ej9UY
JtJQyck/0ib6ISEjDrsUxtbcYknVgzAtZT8fdcg9pe/THcJsgwhSyp+fLjdZOUurzwss2nDnXQuB
mB1PKHSRk50q2i27Gu8oaI0Z3f6wMP4ryVK3IuikPcZDzXJaBewF5xc/qEhlSGzHKZlTS+2S0rHr
UrqoC4fslzwnomKYT43LUPUMF4Khmt7AJkndrs0S4snoih6co9s6HVFOmtwK6y+vJmROyv5JUusJ
5+IuL2s2W7U7/LvRyeV8QH/lfWxlCscaH56aKa/ob5PloBFPzllqpxMf3KhYcrJSnOPYpVg0dieb
KA1lL301JXPSGpeJXHbJtl3QSoefkJWsqH4Hau6m6GUp2RI/vjIUSrj/mwdUe/fKeSjHMbMtReqv
0t9vVFVw5XcQWTCCarLeviFEWZ0MDWmdodjRbTC9MqLWvTgVjdouRg+xpzsDzMZ41ZYn2KmOSN2r
LLgK8w/91+V5kmPY9H9jR7bE+M0ZFTPqesqhya28oxVy/XmeVn8nCs4eu6ziE7lq8iNpoHnACjxu
7Icu+GpjuzXnOwLnKOGjV/+LC/Sf8QOcC8gOyMv/R3obQ/9S8Pw0DDUU8/Dedl0b34RW0m8/hkmD
qfsieaFLCejOXqgOrEcb3RrJPtfGy0FncGHNVqsxQ0AS46hO7D5QIlhh+4Iha4rSVh815Z/4mbMu
mPp3l4WEH9T3U9+LlyoXW5zIAfJIb8uXg/MebUaC9OxBEOh69vMlYGsUIavypz3pSK3xYdPSs1v5
aSxUkutqmfm+ULLcJrgNjM8nBMjXnNexLDXwqgRMJvQMrRut3+LlXV/CmpYCL6yjvsZ+MLAhbBW/
zCmYoDfOxR8pPuWaMcKbDpCV+QTysFISyVKmaMUqfl66Q+dvnzTJ1nQ1lcARD8zi+s9dcy2Qb5RF
IfSn8+vrdvZ2MRJPcIwqikv5Cy1KbxQcMB6XcJu4HSaoC23P5J1tBFQecPmnXWoukp1JWONTLnEz
p61Z3P0XwxrgZ4CmH/RUkTfhyvz+F+/qPpKgfOyzoRXHvripifA5yyOX/DjagarVz/Mka/lDi2cy
XbfApzwen26BEHGuWnOSgQN1akX/UaVSKuZLyYtmCr7taICWAmHD1a3wmtU357Og5NH/1hTJvfIJ
Pa7tF3bmke4Lr4TzmA8MwPPJMSzaD9FuuXSEdKtuOwErKpObggK/jMCE2YT3U6HVIUXOfd+ar6YB
tMjJim4Q/4dKaWNLACAceJ767larD6wBFISaHIZ3D5Tk6ZUOZJTK+a9DYkQsr6tdeF5BNM+NUXLF
L6LJuy4iUJxRMRRNFW96t8tM5esSa7403nKgY4KddE2hVo05R5SJOf+G21NmyY1p/HppDoh084CH
yjNmg94KOTEB2XsgyE5TZ8QwOw6kkho1wh4GF2pWCnuJxV0SKOcWGotTlICgJ86BT7RcC1reRYSg
be23tzNbTjb0FyvSx2ygC5CxMXCxp4gTaNDaTekP3QKnbpm4uHWhaOgnqoO4G5uZa34V2kXAoRg9
yWcfKk+Rypiv0/Nq/p1C1yn2kyJtfguFMOj5uTTY63tv2kq3bnajPGmPbUmYDOxgC6jaShCQ/ROJ
460bq5DJ/ENhvaXZfNc4sI44Vqkw1vKOhX21FGq7XVEv/uaGGD33rIQCsNYBrig4s7Qh2yfAvirI
gYSirCPTM0w7ke5Bj82A3hOpv+ly3vQlz8bV5zUZXEyNYdPipPaEG4itfu5lERVP5J5Ffw5HvulU
nsvrd9om4T4Z9Y+mLAerimp3PtuPE/C1+3cXbRzhbpiS6bPoFdxTvlbUyAMpEmZhwRlSqZcuCtAX
DH4FA2r5DwFMsqiPF+q8iJmrcoPb7iTnhvt3sD3YV7UDl/orhG5NfiPoyB3wPSme3zSLYvwbZ8FN
66NmA4QHUEV3+YOFV/lIU81eMe1OhSpMDoAwvkItQimbG5zoVmrP+bM28YclL9t08Q3bB1k+WkBL
iROGGpcfcKg+VWEcfzqqimDHST8Zv9SvMPhASUl+QfHkrNVDtwfW0X5GHUXPIu7fjZXtrHFET3PS
kOdnK7jrm8+XqQU/mFx/3XDVElMyfqn3ADhnjC8QoX8KY6BMM7hIciHoGfwM5DXMh+0SI8OOxiDT
c0xZOor3GxTN+cdrjlXIcRTy6QLXjgkApnce7mNr06DiCUw/oKO/GL+3CGlYgzfzdQivP+APtVyY
+4KqtyCjooSZsODZCNhDLMo7lcLqmdm0nhzjy8ZSQ2WdEN3b0x1j2me7U+t5cm0nwavsl1Vy86y4
3dB0kfjno/FjQ3HghgWsEnPdXSTAgikg8NOfbArzhyh77OjeOvRCgcwFRgfRc6+XRwsNIpZjnZ2a
CfpSnMj+EHGJT16xj4rK2zElvWWEiu6L5jqyN49YeYvtfVgJzA9KZyXrLRZlW9tCgbdtIKhvVAOZ
c1NsdCXzhLaWCmjTSJtytx+wd1wC9MB5zeiWUmRfseGuQErj5Ar12PUutr0xSuta9vTJLFBHi+tU
AfoLVM0UsSQCoEW+uxVdqNsLwFmiCQshTUGChYlHPOZoOfH8pbkSav1B4rp2o4ZtG3vBRt5MWFyW
IsyfV6C/yxX+Dl2IRf+Deuclmm2T2GmXyYaVwqphbihKuEBbJrITFwHgf7MKSxh5RygnObIC87N7
SbbQFtNDZzpRB+gpcQRIiWLvqmlzg0XzTiS3gDgku9sNx5Di0nfWtdFATt2WfomFIr6fv95MYVl5
zy2QzzwQi7/N1qYZTQ2a6LZ6SeeytQnIg+fOo201iXJNdmuWO0CyjVhyHOBHRYvA0Kexhpg0fzNO
f1ApN76MUsFGYjW3i8K1jnAZibcGwqufmhsWFYlAMM8sbkGSKfjVx3khPMy/+QPCPPi6hJuiHHht
D0vXvH2bVCKWfizMgsaKL5RDZv/BlBUXdzMZbf7rBtj6E+H0URLLmp9QrbNZSSkRK/R1uoYNcSU7
J+TKClH81DGy3y5GjJaEYly/N6bWBLm9asIloIvCyJCXDvl61eshoJbsnJNbP4hJpMFh3K3g542U
jVXiMVxSkiUXxH8CKpu22f4aGypOUSJGh7sJVPBwDSyT4Waf0CwH08yRQ7YtkwpaeHxeXu6fJzZR
BsuoIJ+OXskKXp+jMrWen5z/YBJ3u6itpP5aFqE7m6726kpJzr+hWfdTTKbCG8Ri8SY83wTrmaa+
ufpIdREHLjKF5ZTMdiCN7hgOboWeSM6RJbUGTPe7F5S4fFBsFVh6ERUBVPCqJJQ6esBZz+bJ3E2d
QK1hV7QlAT0VgwSEYQ6vDsUKlnfCrs4TY7l4G5KLJ2i3I9hwuJO871KzRC/mlbzV/sDs5jmAR7kU
8/9QpRg/ZkTCWd6cKQHhqLy1EmLT14pMdD/GMfRKO/uTI98RKXvvijOvyoYrsmYSQJgv6nsZnPwr
0L54e1Rr/Qr688M3PHo6RbtdYdl2LgshuqNJVTgFACz24yYjEf8xyD8cUCOnemYYpT/yyICo2Eno
DHz2ixWfNh9nx1hy+01FrN9eudqe9CNBjTg5qagFxTvfhfLHbw1QgWK/JF1Pt2k9t7qCpJzCYcCE
a/kN5dkGaePo7uIXqBP/F3OS2cB9nZQ53dL6pFKlvGr4oWBOtAfJ0j7TL+QMO2icrIItwmvfr9ke
viBAtLU3gsjYwEWfCaLMBHyZtKu6rEEP/JRezIlhPE4kkjCSh8hGn1HKeuU+/9k1A7GvUApp2OJp
k6u+MmEeegmXFY1x3IS69PqzLjgi61yi4lwwersEdUmi0Jr+O1JZi1QJb3M/XaGUjUI+URsehJbm
lLKiczb34Ll9SBWMAsS7zC9oCX6lTEOD3wDhod/r5X+nAw9Dx7ogPyJIzQgVebVfNkQl9VAe9SQO
r2mKkxrTZyCCdkOSn/KO4CcFJ11HB3xsreWUUorMEUzu2SlvJAncnVyYDYH1oVEA3uel02dkk115
ma2456OAB8w9aRlWQe8zvmd697tRafTJFuaFD7V9FFBftYHCYZYqSl+qdcXuMKjDQ+V9c2t91CUA
Sd/plIcf6qazqFnXC2UYKUvZ5YNnZs2Gt9Uw10gyE+s6mpSWvLDRPmZXYLO4ewVfEYF96OhTkf2R
qSkfrBh6HKOmQzK4mmUsiY3QP9zKRbnSOYQHh8jnG0YAoyk4Al3k2rfKIVUhWjP/zwadtIkqnFYY
yike1krU6Jg7idI1s2IjEFyFkb3i5szBplvaxsGUwroJ0gCheYJ9q0XBmx6tznOcG+vjxSUbdne5
BrUweUdqPDbex+/6l418/GxOVSHJkKoDrqsz9p3lIr02aqGVR7pa9wvVLCpfjbssRk85Ek3hoZfj
aU0LunGfbpbCHXkAHFWG0I523/9CaLHMuyARr03svAJ0yGgsG9hK8RfOWGQ5Fox/BGXtb+CUwn/e
Z1qcoyPPOL5Pt22q3Wz4n/nlB5CNtK8jFyf0zNPO/LVQtM9sJNOmKfvxXkuwtvRQ231fppoMojva
Q3P6/wu47iacgR5MWHzyL6HrAGlygdpf6SUOMYWskh1hZafNcKDXO0OZKyFU4+EyY3t5HMzkmOpm
bKdS5TUklfiH3XazANhf0joGK/fcVqRPbhrk5R5zpSZIGIQjxI3fg7TVHvLqcph+1AuQtZIPBVI/
IT9vmPJ6+s5giQoVFt6I1X+pndymRoAUqIFodmyb8V727ziQnbTZ7x6f2KcMFuLp6s1ppaXLGXDo
zAXajDt4Gno4NaIffYDjlKhyBFu/fikiRk+dGZEc26e1GeXvGMfYIEEF25NqOiej4yIbe2kFKMH+
tkWqeeIOb6J1VvI5tbfIl2O4HnTthWrlDkd1s8B1Xt21p6D+TvbdSeRLWM7gfBY5jQVJQcMPwdGI
I1vGNpRUYPKjjKKBDl2WXLVJ31kCc6aLGxfCzuOR8lVfMbsytaikRfxLjBBOSuEjFoNJFEAs12EN
eaaGXvjZvhmlNkKnyt1NeAghfArAUoAS3+0bJ/DqDaswttuwy89ruqOCbFXpbw08aaX9wgSuN2Sh
DkRu6BzAuGX1PHJYaiGHz5bYQpEOUaTRZtUuF+FKK7mjXv12UHbO1+lg2a9s/PZzgw5z2rsynBqx
aVwwSOTqJn1WDw00FuO/46oJqXnF85f0iMAdJYhM1TQNx8PnJ/diZxyRIJIQuKSuWe/AJ8lwcNk6
qEBaMmtEI6NGFCAAwmJhQanC0MDJqUoudERgVZajIYy69eFhfxnU58QA6yOegpsN7AZTzCKPxZGc
x68BIZAZuzpyjrQneLobrnP/OSNTLAUF2NmcUvrS4hNQTQvby7iagyHbb3/QeTTu7ZU8sgL7zlhk
JoDIIcwiArd7X2/Nxga+zqYY8vvMZXGEPwqV8RvSgJYx+IE1wkzL9yAEue1M7J5LbXZXdnePHr3I
/qF7aSZXVuuW6EghD+L21gL0rqcNRXLOLs9Vc+MKw0FwpHQa9/w786OUicjIH8a+MGrFz6gDhUXx
HxkcbQhkbCm5KuW6/0SEtfCys3oLbwLgJhtR+TrvIySxXyalf0LsU8rGp46U7AkzVEd0jd+W6eq3
kq4tulfvjzeglBqNHNn8lhGsTMtYLquygnAedSxm8IXkh5JTeCE7hRHh7ruTvq7Q6ynsalHgCpkL
qPa5qa5r+YaC6TUvJqLwROI8EEcuEpiJ3d+Z1NG49Ug44dS5AH0u9H0CgbHhPIoL4sVir0/g2PqJ
KMYV2Q4HExhPs8OhjFNjNcUPZbXg2mRNohSctXVumdcKFUgVODKJU3/PcXXoZWZbG8Ht3MUZ2y0R
MHi/nBF9WNymXwhF2RNhgk/ldUCtfS+ZPeVYa0ftYRItCyNHWfcCr3PRx3BcIxBhPQtgFPwBWnyv
QqoYmptuTNlfqTZ5uabmwS8hksxyndPiR1eBWXkUo5a3iIQPyxvr9C4o7zwmPZ9KnmFlfoyI//4U
8cV0kQFrahdhenu+mYBQZujsFChIk2emEGd0RX3lPgueqQfLhN+Z4tkU0Uzcs0X9lxgzft+DrRvQ
JRAIBjfn3WmRXv2Fsqn/G0mAZ/ATxtn0T1fy/Kbp114jK8jFg6DfafiNWwBjW1w4Jid1+aXhFeF0
+wrqBkYZIAD9KjZqljS2Pz4I2XtwJ2bwzjbvTtY9DyYCK52gEXSWaetm146ER5mWOHRx/DELNZE5
er5sfb/h/0Uz99DdLAr8acxJs9Q3XIAGpmRibubqutFiiHUpUtcv1ekXDdx/5RPzbFHG1sjA6vSi
1tWhQXI2f1jaKFIGaXNZ2u5xPHirCQQ8U+zmmC9zzGypPzk8oAf+Xh/kZqcOGFoDHkO5Uq+I4x/W
efn0LiQnl/cWuSD1LfcNJ6RpEx5UKvb8isM76LB5i7Ulp/g/VxcGGG21ykUrJ2+cltKmM/ufueK7
sTF6Gkuerof4Ysmw0QVtv8fngj1vMme2SRWO54iPsq4wgFNXzGv40RE2ZtcKfvglx81QHdythrJR
hxJd87aqldjhOeuLvb4ZNetqK8DeHgKKUF5oafDHeSWKyvJloi1KWLBFMT7NW1ZwAM7RuF9RK7oR
RDIV1D5pX96dU2IiEhmVoSaPFC5XbsnkhkPRg5J2zErFYEHw0ioP939si+v1EewRIcpSg02WuGK1
kTQuVdv5yEO9Moy00odJ0TlMO+AGvVBR4Jy0extDtdPJ7zEm4WqttxBzcUfwkajmnHSJubtPb5Di
a+grVHfyM5K4zTutQFq8H+4TMmKVeNXhTmmPjZ3haSwb9nl2tlsoxC9ONp0ERYngvQs+0q1/c73l
WgfDi1RG3v5WDBGayy32AShBZh6B6/GVGkSH5opxXbH0P+1g8DkDFzYaoNVYHBTP0iiBYxIjjELj
3B2n+TZB3H8AftiYCfsn5NTDRxa80lrJ3dGPIBLGykhlXV1ufIFdlY2rshG/Npc35cLZZNR+JJs7
nIFVasHu4DasXIWi7UqnCqci+NlRPu5iZn9egRzp5M07KM2fdWQk3OQNWhvIbtSTO9kpw9C4SF0g
BRvlpCpfBvL+ynGJruD0T7lJsF3p7sylj4XBA6med/CZE1mhhsLEDUXrJLrTplVkDpjib1paQUcV
sp80tCBdW9yog4grjUBAHCtyjbJQBWYqzug+woLf21GPNV//71TBH9pXIJzjhsBX8q1gh9BqzutS
cC3NVGY7YUvR6P/T8FLsdoj3rynJfDth07/l00iV1Q6xjnHXy+1/WA0izyabjxWvcmTWA3GMZQ0s
slsizcBL3+lex2o9raEHZCLm+yWR0uNaKq5e6C1XGQBwGKbeArPxxXNRqIHQK+d6QHn0QA5QIX7D
JlcowyckGNu64q5LPDlHiFPAtZNMKCEqxnXF4QxEWM6rXkS7KCWR5XWba5lYB0hhJZeD64XmALmL
CjGj5DI4SyHBxiY8LpW2+6Q0INi3mJ38vPJ6USBK6mrGfuBdvwwoKTMmC1uwmpkSXwYyeBFATfu4
pdQrOFk1+Jd8LqT1nNsCwP1sOQztCHvwW/B9vpYT9wnHlnTbUsnqoW5UVtk2miDCJON3QsiVyJmz
0/Xj2SMfdFEy8eHtWJuxss51NsrQ8DV8wxee3IWNcq3kcE8HTFQTYKYYncyqdvCe8FA8TjqhvaoM
8v5bGxb1+hqdIldeCNbnCf81AFOTMXU8kHdPSPGSlZbSEs7ynYaVbN66e0tfKu6P889e0ZjOZcp7
o1Q8k74+W1JHa0rhr8rWX23wSFQXj5pafn3/TGtDFcf3ylOxdHB+jHsIp4k1IHTxX4TGu9u+sCiN
L28HkN+h4QH+/woPlGCTNSMe8PHQazFJlLu2FNyYSmCrsJ+ilgsABxsL8WHKUlk7nJ6+e73PfKRQ
FfLOUImZ6RtkAbFhSmJsLZyuru9GFCt3iXao2vu6uSWJgqP26Itpu32xuJMF+AtG/+iEsBCk1wRD
0twpOGmUywnUOukhLYVY92+ADjTdi3dZ7kJOO3sbuSzKqYtCJFIjeoqKbZM4P8EMJRho0eewhoea
TPCkHEJh/s5zeDU5naIxNOCTVA+6mbAut7p1rIb/grsfmnmfIDwGvSF5elduf70pl8ptXRTTUK0+
k1sqoYMO5jKL0Py9Onfll/LwIQBDCdy1ulfx80v5chHJjZZnu/dC19khmJbz8Cl9mtkFBAsiq92g
5fA7xm75N7YBE6iRP39XBL3uc3H8LbbfHFZ9UVZAbFexF36y8jI3Sl3BoH4Sfl+eYP8ZZkUVAENu
dVubDCJgHN0m/md37cC1lU0p5lCGc5oFOcvxU/5dqOKYXBNpSE5Zw7vxN3m5sTYqaVVMMrHyUL7z
UvzQvF4AKglHDfl0dUv5Xuc8tXp3lqsGeHO63xvi9WXq2AyzcNes6wBJYKL1yn+YAT3z4xL+WB9l
vGEbjxAMnDqpqk5ouspGnE6u0WOjhD5rsARleHNA0ZHMezqpFV+4UDUos5SKT9CAlGj6QyDBe0dx
Nx3KRdK1myhVVHVXTy28B6+Dggv73qlVf0NUlDsvKk7PLb89Sesf895Ja/anGSyIej0R3x93w1cM
Z4uiUNsZxjvJfVm0NXJusOtDAOTV7D3OJBguopNb2ByuB3WYtXqqCfelWMFvWEPFurPv3pYYMLAj
Sq3WpDqOReQQpJc/GFZpnWufFucmDm8ZN3fb8k43d6ImlywnFF1YLZdVLe3Fm3NOh4wz0kGQMDYV
bl0S/opCNJTZ8fbhfzTYECCufxqhRzrhCXbUr2UVg/FzXt3WsZycsOkxlaUCor7oXGgjkiZo/kvY
z5OWxTvSR4VCMDfRkqhyfU8uRB9gIQP/N/gZC2rf05rRsxD+sPWOF1h+7Mm4Fy5cvOOT24d3GNAR
zihYItdlyDDjea9KCpI8Styv9fD0oNp0P4OhpvBVpJENaxv0gvkHU3RbRkdku6R7jvZEwIP34Il3
j2cj3OMlXbA7vcyKl+04vFUYkhESnQWEgSJ3z+4PGhYFugbAeXcN7qDYAkjigxyMoztvplkL+18Q
FlKzZ41C2wFcPpfBsqeRT/YyYfAba2Bsup79D2DcRZQ3C3VXd3uOI/Y+Bu9gN4hVyU3epTfR7onW
gq5uy64M9mD6+690iqUxjY3D/Du5mzXxJFqW475c9PB9EyDdvaUqOqIKDrkCM/Hh1hQVx1S8XNvR
ybqRUsmS9yQ7q6uLiDaBJbqqr6cJdrewnWbdW76tN/RluZDCc/yn5Im+DT7pLlkag0EFgPFI+FAT
/vpotDUbEmYkD1Pu5xuXScMVl/39r8hWjEU8gpDu0DMjnSGIOQgaZALzhpqbrFqppCGq8v5D3Wh6
vzaU6afzU+Qpb1EiQI78cNaKMkytd1hbP872yNf7WCi4SQGrRoXsW+2blVdrXnBn1LTjwTqAYdcC
wBHOHTL4wtL1sjPdNXwMWra3ZquviClovDGX3bPwgVsRgejhF/fHHtSeXpkYfKh5RuNM4oT5PlWc
kFYMD8vxUzLbqVCwq/Qch+8q4jEU8JMF9HEdA0DxehQeO+QmSTlQ7jd0+GxKAMF7A7LAfycmVzjY
TLC/+OCzm8XWfNI2RKuAOoSKrE+nuhjTzSxjSgwLYHvxbagvXlWUMwhlAZaKSoR9X5fyFKlS/KAB
Lz887caHcxsKzQkEtlE4KlLFpjN+bjfDXJyqf8MloHs0CSePayC9u6VvSl+HXCWZ+xAR44cWUhkk
bT8+S/53AN4fK5M39xSyWgGAIoigy6hlPM6frirqgA2+1g/a0IEdUMQ6VdOyT8l8OguxwxQ7vDgI
GANZJlz0m1xMUXefF4JwZY9Z1ahK7enGdCFswjik45Nf3W2fzX+WdZJjiWrGDupBOoOv5fN4/Ukt
oevBiel5VfGO5UyMqI+4erVvErdJpkChC/dOr+j5HGIiH4+a0sc1uth6dxVEHAyhHqiLfkAgHl7N
T2Mv9tVN9+uByYKOsD/Rb/hktZ67nU9QxZfJJIOirBxDIpIh4HIJ0T+RQM3WSCK/wDs/W/WwHrzC
2bcRytlpMg7/+YucOxpSRD8vQVreddComMzsHuC8di1rL7KaB1JMNYh4BKURM9iDllKSF1/6N68a
eBhWDo02LUgdueLdqR3acu95SRiad+wK2C7TOTargIHinx4+VKTMhOhxDWUjioGnf4TfYIYzgUT6
OVqWWzbarFj+zQlxep40UI54jf31oSXqakxVynLETDF2XED/3djAAcLjnvE1lyiGbrRtHEPNRgSR
DZlz0bysUMmroO8RqUCa0RJABwrGVeKnveOhPqmWlFWtBEqWgXeTVdA7JjQlQZfUjAwXDLnxVZsO
XMvb5WjX9aApvC7GlzpksqUmjG8zqEC6TFucW5aIQUucfJ5zZb1pbC6FXSPStT5sjU1iul2dRx1d
ibte6hGpUT2KRxTfM1DBgUflzht7WfBOfb6JdficYEtbRvGygZjiPp8Y8NAyhr7gJHUMjCXzWehD
Xp/Vm6kKDInOhImwxBPQNV9NMGA9KUALUYL9Kjd+21jPtKfvS5bhz0ZDmeoYavoNi8E5PcH626UW
hykPKV26VDX1YfwyM/rivuY+IamKJfZvpfvc4RYIZ5XYTU4HVoXiJn+gzNhQbi/3+Zuj41Hr0hAf
Vl3TJNbNkpfmBHRqV0lr2cL7T3yH279+Bf3AJrCMkZmiXAYhHzqUVOLlSTbD0nRq4Btxehz0eMPz
pdx37dK0Qoxk6lc+OQXEUWxB4ek4spwJg4bTpFUf/FVjabYb9HPxyKyVLn6LUru8baoIgL5g9x5e
DXaS6+K8SPE+mNRotxNzF8NBLMgLUY8nn/KaWKCfHG4tfhKQkODQO0G2mAiUSvtlueyrjFdJXnEi
AtAPI/KOIhoM3ZtB6xhMlBTEGh8NCnYzos16EdsTsNONT8QYRxNo7OO5GFNDaJYgQzQKXdBke5wz
/Lgx5kVRhlLZo1BMNLEa/AS/AONQyRFFxnoDfQm8/gifCKTSCjgtwXN9cp4zLTIOjPFq5zxFQu5r
a08NLlhVpJXtKXXlI1JEMSIpFaFl5N/kt8x/Hl33vuRnIM9we/iSnIfNUUgFho/XDiccHQv2cKNl
c9C/RPwq+gOfNEwOD+rHGVy4V/lMY3AhNROARRwTUOFFRT8GY6qjScoaUq8hPRZc1CZYTATfIue6
okSFHjvVOad0Yjl+MhZH2IEliCmsHCABhewndnJG7W7JhWi3yckBrc1tGrZZS9h0CJmgAGnOYCWW
JbumUe4aF9ywjUcMvs2b4x0bvJjIUo8F/1qBJmHgkfisTnEM0SScuVVgihnzUvJnUhJRxfLl4lUJ
NmrfFcbhgJbB0SgkJz0MFImiWpW/7bPMXacqMr1qO559KSznPu3Yqc5kChZO29jaLH7DLNpnv6CP
KiGwIPvSWoqmNLQ0PHZGw2cZDbrbGlYrDc8MlM5Kfo0ofAzoLTczuN27ZMu3AZDI+27DuVOMKqDs
yRoBeN6zu1zsSmnUBbtHSRaxXtJvG1iOUW/13nFZ7A/XamuPFm/aWeEYdAemOgaAUKZuM13EVWng
/2p4Rr0MCfkLkgwLd1gXVDwjY0gfbT1BTqgEnZ+QnxWRog0YzyQ4q0+zS/PQZCyB7uUeyIVjnSz2
sYj1ZusL6NcYZ+yKZ8/JQuLMMy6RPlhsKpJ0mxXxnvHuMHk4nctVygHm4ooFcMxJSJ+iQgSYcuwG
bORdnZjkVYnu+TKYEWUUozxM7t+mllzMTcYv59qf7+dNSWsdsekZYFQtHb7oFktNIE8rGX3NGxtd
ndZ957MGE2ni/3oj46f1JA1lDxixWFPhCE4rjvqxHtkOff/mwrRoR0Rl8YG9G/mjVPow+I5+gebq
aJVLw7x7IXdRgrPZ1t0y9hQjYvGlfLp8rWg06PVuuHaAboznwFWJjEX+mSwbGioCHnQuKfDqahxX
7bKMiL3mJf083I/sSIViCjr3HoJiGpPqPW7GTb4sJJ4woiPWFME1Q00Vx5jVGbbmozuYwGNVUJQB
xDo+RpiCT9OBh03f8NTKHjgjeWxJUw8qR+mZaTyRUOF/SZadVirtSyGGvc8V0brMlq861042RsFM
8WzjELra6u6foXGQIJeorUrPGu9kbQ9piq2dp5cy6gODRoefmhLBl4I9UdUmpqN1jGXl48q7scgd
UtjtB+YZZmpiYeqCDIMBAN6eHPsMayv621pnMufg2wlHAQfztLKuj0ELtGbcii3NW8Omj9Z6uezG
A5pyNrVXhPT25pMujPjlQaYSSjvGzjugDlf0SaoOm/6trph/soK8ePCu2oSp1IpsDEXUooIasYo0
IoRtZvelKAET5ty5BtS5JRnPQG17aAX99e+Ep1C/R+nxtnqsAm/CgkAjsRdU4IYqKnm15fR5cqry
3+kmv7wYZs4bswDeqH9G40NuTVikmnN71lJNuSsCsMHsLtS2UiiU7jOXlkEWg8clATQA5qekMDzO
roOAVFt57MeLP6b6HoNmc3yfB+x266SKsdB/SXeKNU8spqxydh2PWe5hovYZOgJwC7SdgFRIOhmN
Oq3Is0rvKbPCDDQIrx43FwA5F9p77lceLNBqlDHdxJwM4a95We5TRNAnxjQ+/ISSvAEFKTKQNv94
lSIgorSbisE85Od3vO82plS8rOf9H1AhTfy2YXcY9wRLQqKV1usiXnPfDWXtOHqlTGK1wlekTPna
E2D+VGwKDToj5BnoDsCw3qrmJeMUiEfaofl00UkDz3v4+mh1bdEwfxTWXaIdy9ef64P0Cm8XfHMp
qjpWMe1RC4EVjtQZLyRXjkg+/khFHInVJvR2SbgcgLdLtTny0c/0jISSCIFrpKslLcVR0Vh/nyMh
qW5uYUFuLq6avit/I6+yYlAsAIMBGzK2BsTMLSHRayQ7QzXgCMAO0aWGIuPINE7JkMa0a9oDL/3V
KixQoafE9Upz2VoB54Tk02VfzvMOr6UkTHay98Qc5t+sH7nqtuCMD9pAE1uK4Wapwojp0c4H/5ny
7e+fsrEdrLg+QcHZv0OubvX1rR1F97Ws9ZOvCWr0YGHuLLc0g8PQivMpOmSlA+N6NrfBANPTjiA5
qDJ50TFFut9pIU1ifbI/MKrhXY6JVO+IzPrVxbHSkBEXNgqA31AmnJlW4uT2J5ZnDRkldzn2LYbC
RgE1Ifi090d2ROpcwOm8loNi+cdrR0Pm9pYIhQ1Mb9zgNR6Hi/sacQj1cMptQhfzIbHUhprZkXrU
T31glYf4ybuDzxVR0JQ/Hx3xnqOVEsvb2HfQXiMhvLR3Y3XpIeYFCr+jHD2/iveq4aWtsIFRqSG1
t7P6oSQ8pqh0z8I75UszDZjtXDfXQ2Ix6d5if7N33a1Zp8NwfVN7nWC1Ct+GQ0nnnQ7PcssQR2ry
+nW3iqQlvGIVh7XX80u3N//Rjwqrw3HKaAqps1LvXyAeGaa1hcphP/nchoojxY+ba6GhhhIYLy0e
eJtBsrOnRziypcZ9sfBd9FDJEwhOAfXQMr2g4h6OfC4iUb5kp1D74GM0OPUt5878Vi8jBOIIr/Tm
joEMrI3LtrZqVmZB74/HoZ9yZg5AsztLmpsd/AIb6u5cMyW1ClSf2qO9BxFzCtoMagkkONH4tBkb
wTwkJM02s/4Chdpk9x1CrRiea7GE2+DpZkQ179j1aKGgs9YvsU96a9sXdnf/fOy1g9qhGBbWWP23
E7u+Hl0h1t15CBTtilXMtMlduraVl2Ad3rqepQazxupgd6qzBQvlMxctcPB7CgtBwuuGb4JkBQap
uaqFxdmES3maCAQ0mRSPrvNbHCWgryCPsE0i2txmcGS/VimlRktvdgIYuOYACP0QtuhdVDotrPo3
9d7RHexVA/kSMQIZpimXW922FoGwZlBuekIBAI/La4Jia1Rn5g7L6r+sySvQjCUG/Yzteuufpzl3
0WxYMz6qI76oI/QXsreWlpomfEGzaqpIYWVkEWrz9cQ0wvt5GqOfUcdUlIaqCBaYr/MiGdH6daFo
fpRHM6DL8ah4zPuaRY6xGHx0mDzqonCpKASopbg3+pWYLD1jY6Jr9wCTF9wuQFNO9DrceZg/h8h5
5cYqqnE5wwhmP5yDCh9wQ5X3CqmCsXtM01XhUFjnEF587+V3BIvnXnxOB6mwX7P2/yHJ7g2jJwsn
c9MrVJxKNJhiL4IM6CHCphre5bx1exHZIHZFHV6zzfAk0Wqi+HmprY13zWosDgJMLar6ZJD+HCTB
Yv1+kWwY6cR89Z1fOqE0+VLa/j/qwCiHykEl6m9iWgImlHcGTKZGP4e2FwL9jZ7i7FosM9cWbwQ2
o5MmHyBM4BT2cUW0lugObGjAcjDWh9AZza870FqpspKTNqnMnOzrJHIIO1FSUF4yypg4XPa9PzVa
tM1nT2DhwSAs4uTYzb3j9b1oDba/jLYaP5j5c0B6XtxwYIiDuANzC/p93+1hmUzAPYh2LrfFS+je
rGBp0w32Fm1BZXP+I172+trH7pW39e5krD/mJeY22Lx07un6BiCSzMYSQSKWO9vu8hc/SePqJecj
CR/2CgS1SjtHoUv1PC6s9IOUPkCA40x1AzX+JG7Wubs8ebO1r8GRzkY76DG60QhhmBTjBownpTZj
rpOE6EmD08NgjrfwNRDnmRf9aGOjAMT+ANa9sU7A8kLLITA4/jzxpCjjs+EvVhOfvmJhXOgw78M+
C6+mXTXwOqF4QSyu2IxRxUsLAlrlPBoAfDD6y5M1NAhqMLL3KqFJV8lWWSuKASXEJKIRaVtVCVER
mY9bUYPk64kEecJmE7Dv3NIPc5XWXpyQ9lXmDdUaUn26pV8Bz1JpfV0ocyIfKNgrwrdbmRgbDvjQ
pSMg3M3E1e3tpMlQpfUlzCNUiaX2o+pxQSKJabBbRI0zpWWogMxc1sIYVxjXTP8adrHrVCrIlQXl
WUH+D45Ftz+9W96WaDMJjpGGfidbAnnPks4hix0Vmnonb4O9F546Oy9ItPNz1a7YWmr3dGbW7SzM
DfoDwsDRMnVmFs6w6v+xIf6YxWBR7Y1bsN4Vt7KXIGmyt0Kjl+LQRGcC3rCTSuFUfLEBik+4jd+2
MfHgcMANTXVIwE0n1nHEy+lNqXK13t70ozwhgxysInSDKLqPc7ZNoTG0u3WPXEPbtQRvreq6uLio
GPnuJrWUbEeubS/Qz9t1SsF++Pz8VmNnuBu3UuaJWr/Hfi1d0UUVW/xzaeqU23p3ivoHdpO1LgZ5
ear5t9FVU4JJYqe2AonNrpzg5Sdsv4lMfclF7JNZDY+oVskt8RusYEFVgQUOVk2RGhwXqdewSkCf
YLuzgSUGDD07saML6BVMpFm5/SoTdqWc+aJqLqLsRhMKq/kSTXBrdHwDfo0U0JQ+Thd/mVjBi5cy
a6i0SeUcBgO3ghv6napZ219rejw3jAeEfYiTg+9FtOZWzppaoIoalyuNtGVNfI3gpiUL+v3tmzZT
ggLZtN8CGBLlanYnOmDbro3PraDEaPrQtwJcMquGuBlndj0YgVhclGAdmEPHucdHy+xuUyIFejE0
VHtpFiRS9tN2/fYL2MYhqPi1WVEixxOzwjsMcxKBQ80WJxrh6Dyfd12y7LLZDq7f8holsVx6xntG
MXRAe+uHaFdnPZPB/6R7Ij9rYbYCuarATk9w9hF40eTTjbLSe3hjl+NdBBhwwdKfW5AgaYJO0Rtw
kCcNs9GDVJxrRBLMj4tpBPoruT+MlrYXLdOUvl7MjdxHApyIiayGDGVGdYl4IQEi5lulzAB4OcBw
A5F29SqCGP7RI2LZeobQwwZOjeLRe1otTw8vq/sGbQcA2SMTmBDDNPgSURCwsbiduyQcDyNV9vC3
rWrQO5bolbHkdhknS9/rhNjGMrRmS2U0tzYI4M7Tuw0pF1iqK/AcqiRX4ai6iGBEDnOelYab/SgX
nPqgmE69xwFrQaXK+pJkAJdLX8Vx969OM4T+zVAjygPY0xSZT4PsaLs97oyq6qEZkkDeyKti0Xql
glIvnLZi14gSwtGN2KqQlyZasfmdcetQAu9lZ7X5RTMy3ax++Eqd4XcTiMuVe/ae8FSzM5BHkthv
gnr6ks/pwhoxacEOTjGnlf8mv7SXptz8gOHTXZ4CTS0t/mafTTcDfKbeuLIxFKO1wtj8Ir7zzNm9
c+tL5mDd+CQ3dQWX+3iShZoaWM9rt8miX9nKD5zj/ycgyeRsSPJnodhHt4aaebTfiD0h9VdP+aq0
oBqHAc/c2rgg6yHI7xyMj4rxKpEHlO53hBIucefzZ/gdxSQ077M9UzDhansnNUuCjZmMD8isTlzm
iArOQ5y/d7KMxvxhKwKeXIr95AtW0K6oYYVrAJzLIT415mdCME++JO/IGX4bk2HmqiOo+O83SXWm
ey2z4r11eKL5U6RcCZDwQhbn+Q/uzRJKJaSMn9l9ju7D/WA3x9Lgxxu0SMGkHYfp+K1os6Z+jIVT
DEhgJNebFLjoSVYDxGAt0vAFNH1nu9Q3j4SgHeoGVYdGQ9+zX3urtXWhLer6tV5T+MM3pgWjpH2n
zwrNYa6KMUeEWWq9JfRQP9uW9cghozE5K6TQW7lWxWDyAr6WkJpa61U3jy3ri9ZF0LNqHX1PNYVX
mZmTaALqnYjAkEgSxS7B6q6/ygGzdqESEmcMktSSHcLqlfKR2lgwG22cmKsdjwfEJWYDypMQIGA0
lwlParjAHXjo/w255ZKyjLzPWr06+Z252NpP7P+qUHYsZsmJYSWORz2bQA9w3fEp0DzE6nGJr59+
bnZfYQA/Y+xxUGbFCjWpt/0A5JlP/e7yBsT96izJw19lRTl78F8Lrgu7YZSY0b0rH3IIekMi+bGi
mvtQNEVWpYVp20OwMy/JB/UAtRuS5cO3c+560QuMzBdukejCslp28nBtnzBwoMLu8IpVdfBSuHrs
wHnupYBuVCYw+drjNFdr+s9QSh86Lq7qpJWV57hBzxSAXhK7JC6XaITmLf3GTr4aywDiHRPzUBn0
d1mHT0QZXJdh+Rnj9VvRI4CCQFFf3OsqMXATptPQPsIU50i0kNtzfv642GjNHnhJ5sjP34A2vviV
UlSABstltrcQLdM7iRI5CdFrdRLevqMAulQXLrGhZ1mE4QPjT2guJSibPmuX1cE/Gb65MLDXXHQC
HEqI4t2Ikwh9mTMycfehJhwYP/YCaOWkxSRIMqBB4gUEn5HBiso9To+7mBE3yDfj49xs9KxdtdZy
KScfFNNPDbEwD7tvnUA/IWRimGC/iYheB5L8SfVqMFWg2E+AmzhyMbG6D07m6ABv94lDDE51BV2W
yJQbrkW8M6pvXd80hYpWqDUuEEagW/ODt9iqjC6xWg92GHrlZqOBQ/G4cOHAf2SZ1rQjEBAPOaNG
jLpEtjZsQNPS9pCK9qSKQfi5ckVOMUrESpEf0sfFTNNH+bZB2DwPyLAdDhQKnxipthpypQJFR1km
8VHeJOOZQOF5u028X6FMlbf95w3S/BU/q9e1b2Papa/nOOfMB69utCgSlhhLGmsTtp7WmfvcY9ih
hLOm3qwYVSFrNga4Gv/Rckdq44tdSzQBQEHerkSH3oVgpsnBs8nPt7Oi6RnlzRzN6KlUGaeUqoEJ
Z4ZAtuHJH0gFYbOpPINq4fl1zwmSTLmo45IcMRLlsNpnRikOn1hrxHOPvkXYHVN6Qh39fmcepJ4B
40g2gzVG+7Ioxi/jYCpXphIYdk3MY8QnyXhmq3rQ5S2oAqS6fFa0IEr3uVHqBqa66vk8g2n+O2+u
JOfbdPF3n8gMF1ZGMaV9ucHgm5j+Y+s2QiQmJxOzIh1d3PxRyRH9DoBj0zgL9PDfYbvnckCKETzc
EB9eEr86NulUcXajfJJXARINLR0kwVKpTJql2FBpavZdMX7qKoieZ1+Dz0s7yigDY8ciHt8G2MVD
WPoZd9TX+dMVb9YnfKQ6EEO6DNkB8HZJS1x5Xgr4MH0oehCJD5+bDNk8Ez4N3WiSlxaO+bk6+UrO
Dw77E6tIuaPfiWIbmb0TiUlHLD4J7gzpKhiDOszerayDJssj2v07fW/tgyqM7OzbcpV9KUWVQMPc
MVeAnZo5d7P8IbH6tI8YX72LeHK4tqLVZj1CrqtGwlRcn5oWps72AuOrdQDM1jAm24pjS8lq2gvg
1jRGMj6sqk51Qh81y1z5xAlgAtDzsYRD9oRttWjbwGtE3MU0fN+BszI3EG+isXq2VqTaYpUG27ja
6oRn5YMRG1KmH4utMZrHFzp6jie1UBgx7asz+Z6CHcL+yFpXVYbbbWuBgJkijLW31n49xNLXNErz
IQmvVGZU5HrP1Ev7eqONQyU5wk+IYZf//mUlEOVRXlmIXA1wE9JDohHe5QRgr9TJURu79CU7Sv3I
XpKAg5jYxq03qaLMBKTIkFEd+DEh7EbB6zoH9EGlG1QKhfkCa+XnUwakDbXJFic52A6Afb2UMVqI
NW+AUxyDASltXk7Dlt0uBGLnkOOtYpiQTSSJUJ+L/yO7bKVXE79JsOq9dRU5cUFTmCyXC0aJFwLM
/wpS2oesXPkcMTPCuiK/iBLXt46DM8tBWqzoMw/vv/iurBe1+sT+mCUKsqhEUNIv0xQ9zbcFOjv7
5I1NFobnRgw5iCp9DmkpZ2ztFahyLUn59dLyPqx+wbsu+2NFbOBI+pfWjnyGz6b6K+5TsEwoWEKw
FqHcu0z0BtsAwhOK0aSO4t5cs/0wPzqMrbb59fgdrobEqGI9/R0+CckEi1e2Fjv2JNG9igBpkXdu
gsLUuD+OVR4V24204KHfuVf1QNaOu3CJ2tnOG/EmFxpGSB3UAkjTMpi8jvRAq4vt1Y8IYQvHhqXK
+b4QuE+XUC5e+bwUtLXQFaC4yh7fpT1WxntTmRdsdnkJPSh8ghgoRJMyHpSh+UBBn+yoX702lmlW
i2VHJDXn40dOR23+jABBTWb1P/bX0TekW/La2bUGRRyiV+Jn3ZyJ+mjeF+PLrkKxzGyhx1Qz/P7k
GixjzeX47OeMASuyprsL7fXCxzOay7ZzR74eJFaHCepwxtfai5tq4D/FGXfbeiFUNrwVLEZoZ5l3
msJ5MqO8CiOkBs2peCG9gdLjR6+gGzu7ePSIpcFS0hFVp5MSrZR+FKN3x76p+8JBw8tVJ+YcIjiZ
T6JJJkuyl4OWaNDGRdhqjIIYO3oQlWlBWbpWtexr/pOVjoXECJJ9y6dntAxFSyRMlDG2ZRy7Dmlp
HkmwxiL+/812rj3xfl1MF2d3T5dOUtinwrzxm8qd64+9KwY/NvXBrsDN5uo6P7+PMOAm3W9fZ/SY
mnOnnYSKbzjJle5NubbCRFIVsH1HpRjhsrT1nSJAWQVIcMG0lr5Xs0UBmoZ+/x2rSMCFsWRf/tLS
WehlgqqBtYu/enQyTDqBd1amWrWE9Y+5Xvz0r+TrCvhRbBZFNtB/YoOKlOJHh2J2ZyVaYTXuKQJq
EhnhP4+9TOuY07p9Ixn1J1n0K5qfeSy8IN8ecXJZ7KdVTYq/ObgZOrU2VXqkR0ZR2HS88l2/g5ZS
w1JMVzEoyu2oyJK12z+26n/MEA5tm7zTzFX++wtTbkWmv5WJRWQE73wklpM94Tf7/saAX6UN481G
EicJl1Kw44jInOk+/wWGYr2/yeil8EzznR9ezfw0ISdmF/F3JR4N8CU1gLH9h49NrxsoM+s8Hn5d
c6VfPIc62lj6Znr+dZetaQcvGke8u6U+l1ADPxKz5Xdfg7m3ICnzCnvNnhh+xcYKEbNcP6vMdnZw
leKMCMdjhEUvv+XLEMe4vQrXOeB+2jqLB258231xZLxVGL4OtD1APGkKGgxZzRhJK08SITkTf1Oa
HqK1UczV7tAq0xf1hVJj0SSrtfwJMcNxMzq+Vn/hLLI5VPISiQ20TgWfmmQIV12f4pLb54c6OjxV
YnRlSbQA8F0fhgcLsFsYOxJ9jSlLtayLSYXzgKd06p+xcOO8AoMDIEtEy7Fo8kX5ZmJOZi1lAvn7
9tF8QpNSKlWwctXCD2sHPt7diaTevrdx4yt4wVX9kRL6Hu4Q5kLnH0RMUCXFQM9pxdboRVWFyM28
8sX5PqmB5GVWbw5amBuUgD763ggw7FAb3zLMefbnyLZafSRFpymXosFdhLsh5OSEo/7SJ2PF7Q3a
ge7N78JajYsmFu8zzbs6tPrS+jLTRaxFnJ4r/6sSMHvWIIAPjP/X/SIzgfniv98W6FK9rQSoR+wG
7P1J8l+nDjcq/6JFKndLZfRQXCcaSzJ+UyWRbmcOudLIddzkeUBcjmRgRvMLpgXKqnOz5PdvKmYx
Bb033Vx5ieX9YAwU4LeGJBRLIKX4faTkyp8kPBXkZistz+ifBht6wUsJg1X6buyncXmabB96lx2C
XrMCSqRqVLYDXzKP0h3jwXJZqy2P7DAvchxmzS4Irqs0QJq8M8qVbn/SxmiykkF5G1z11bj/njmR
2subyVm2K5PYZ3OSYvvWzhlV0RwVARnbpoWAMDGmk4r0y20NOiDgGgjFZn0kjMNeUwAShMN/UCMz
AldEl7Hk91Z8RcSWnXj5Y8YWBVNAH0h5dEkWF9WIyc/eInYeOJQls54YDNID/webVwndipgP6lHo
tZ8n3bI5gFNtnp7wucmsLbS4Xata5thOxsS9IJORBdKTD0h3FKopoEPcNMizBkmOMiHOD25fNz6M
pjLuNn+7IHMUv35aqVFv54Ty8UYhZ8ItSlOqdHcM7HFAZXZIM/gDrdQ5Lm0l5nVyYgsqL/qe1PtA
hPhJAvrgeBpVV4AU3KIcg/tvqkglpUR5tDbj8Yk8vYswNKcciiYvgonwx6Nb5YBjaH0breyjsoiQ
CqSfvHUj34mtz7XKbpxnwqkMT1pobcboDYogktRmBi0T833QiTzBs913WriVVd4+Mk4CQt8v5Zad
gbrolcYQguruqnK+27sCSyqbIQ4HzmwVygWsNv088wk+ocZxBynPGcfotx7+B3glUdHVtCgzFz1k
c9L5U3BwzQmVSMYTRYSlAwIIGjrYiCeAU1x0+JVz5GqJp93XlfS3BPqGenJ1RfHuGXQm9RKJjAGB
y7eViNkDaf9WILY/7kbfqO2ws2LMQDrx6vEe9H18/PQwjM8/hVzHs+mJYbgJbTSrgR5lwX1BqMCA
qMnc9N06O58ohf1qrFZs4lpyZtejFdH62IVPcJm9gclKncEpuA7sE/g8J+nHiJhBOMPn16WEL46u
oi7qPKcswAX1pyrm2pa1vWAAPfnopXPrj8zRw81uhawIgx+iKoiE5zi7wX1lKEAfH4xP6dB7PWFC
jnlkWFmKk+ie8wkX3AwW6GqPGGTREyS6rGEz6JhVIzJcLKOJ4+buGRWn1Qg14zfMmS/Qc3lbcCEu
QHADIJ7p0qFIZE7g1A/IW3zsIpvpNPKeiVcCjvHmyvf9ovKcvSiKJQHGSmmV2L1Fn1TwAj9kfscO
zdxb+IAhJ1s9MCTuzH6qdfCohz3Eyqx2vHdSIuP+Qj36hbsMCGGBb6dv5oWc69PXb5dfOcOWvkCp
r70yh272BFhXff6a8h809b8U+T6b2r9F0r8yq0kCPfwdcRyJtuBxK7ooDMnpufUNbihzI8MrRydT
1Bu8xhU4q/L/BDG5b++c465MGQTBqPIDTdRjB9ax1SsuRFRvEZWTlGLfekqrRPKtGY69TzuiV2nO
DQmOG6hWzsLWZ/qwkPAHoTLZ2xN682PvrLKYVgpZ72qNnl882MENdMNa1d2FSiQ7oedvSTaaeiIA
elRNnXa06OTzc9g3LAgzTSeSaOTTow2QADyMSwf279p3Bx2jTBH54+JnanWTjVutXKRGAd3Nq0C3
U5Wx4mywNybSLuf2xCABKGp2TnagnWhIC+zm9dg+vx95jYs7lVZ71yD5wfaw6kRSuylYxu4mTzOV
mE9WGOiiccLfjlTI66yx0WqlMIAtzOweITixACW/eUGRO3P5xEI5hP7CNvDy622mtYKtD/Kgs5lD
LSXDoU7MlaxSgdzlG+m6nHxDEom5XbvgUmeEmwjd5MGNJKStIWS/saHpVXz36IgQ7mNuHcHY+sUo
0QujtQEbbPE3knJkGxhME431KA9oWXt9llrnQjxljHLkrQMBtdUMhczlvwK0/mFmccEQ40wiHO4b
sdfW+W+ruV8lSnTT6C907btsmsYVi1xWGUHmNavv0AqxfWhYEF4qdHXrvWkd2NUgsgx2lygd09ID
rKfBASVITXdnvlXMqy3zyvrK/q2p+UTxgQe0ipCbANP6YRGrjDtZaZGmwUR6GjnD8o0YXWXMbeKM
w1dy65vEkWCiP+k8koF4N8iRhXsbnnX+1mN40HKMA874Gn0+MkFFgeHit8IneCwvlSVE5FsPfkLG
ne3rHYpFZ9WusSlAEoqCelZ1eUyd9Tu1CuPHZ0fRK8aRdip9/n6W4ZnJDgtXapPhM4Z9Q+vptGA7
vF4vwGRARxSMcX9xmVDOOb6roM+whmHRShTtY5A715ndrOGMzhh5FMIN6eBL0UOC7vgaYceY2ovu
E7lo4u/1aqNO3FPoMLqfjS1KiasW/bGFCGPWfGaf+GOSqodye2UA9gNrOQPmubZaziYtrnMVrUF9
7G5+Bqr6l7p7E8+0KHt5K3HSjJ4Jn+r5nnqiR7S9r44SkMOvZ+lLgrex37KfslCEo3qTaOIFGb7f
BNbquc4hJdXzzC7JX3BRdTl706jnTYbG1YFYnKd2+wEzq9DWHAFc5A7eGkvF/A5utE4QvGknT05Q
Cb1wwXuzS8WVQPR5vN2U3RwToIRsAR4PDi9RLQpnyxd3yPlWY6TVojqw36OFrwLGE/C7Y3DsDdNo
r58yshCO6R/2f3RfWhJoy2SzUZ2pGmQeMcwAgv8rKNk8vX44/Kuo/A3CWqnaTUrnGiZoB3o28FZo
eVh7+p/xd3yZ3ouU/l+gl1nBK9BR7Rw0MuLxEK+WJ1Nunj/PQjxFvli4Q3jW3SaQnjHZks5ARvuY
UE3jiWLw4zQwV98abjmLF1q4ETiE3oJaIeAF+RGGHKATWe22dhT3f9AGbQb0l23y03+1rZ5dstzY
mXXj/17DE6cg+3+M686hP1Uh3Ebj5uzssWvEaAxE2M0islxhzSY9r8k4onUVYPuCIFrqtTIjlKJf
jrd3Dlv+716KN9FYP6Nj4scPuvPdWFy5NLbibrHfrv39k1UUBX7uHT0TYQQkgGQsUqsZ7KWCIZQj
nVAtPK2GNANTtFT/wjfnSIezx/ffs15Dd5S5sgY8QrpTIAsNfjcg1JN4iBhaScKf+4MLx2QT/zp3
ybxF1o5Z8ch01dv0tgpJGD8rHZbfgtbyVFLwBUy7IlrKgYCsqLu+oPU7tcxId7cJNhrqzMwZ0Rpu
MRFapokR+iRqxj12NKveQwZCC5pXlQejVD5jP9fUEKEwSl/5daD9d/zW5yB4n0OvQNM9OEZF67os
G02DHG3Y+D1MIXGMYUa54HHGr0WgXCnBLzdpVm8gsTE99SE2lYhgE7J9IebAizEuer+mCMqZxL3k
xX9Axb/fS+myOicTJdYJxik3MSyYuQu4PGFLkzW4lfcuBeCS/Y+jLkPih/cEjjdV5Jv66YvhOLKq
2O0TUa/8eBZHwtCp5whUdjCSIAbBfoWzPjc/RkzCKW6unPQg14sjwhiPQYPngtSyPqF1dP8t/33Z
GQnGBKGsW8ft1zu6WQYe4ueDzEo04dP4juv9WGw2MIO8WhxtKA9r6R4YkwQBSQxpu/BX/1mGymfi
iaXL/7RT7WlUlmKEvU9qJPC9ImS+H/7+RRavAlkJyQLD1S3GV45wa1s4u0KTZlU20PgM1b6LVp8q
iTO2cU1/7d1E+jFe198gIlW6Nvyz4x0zatx14xrIPO3nZFXwTzyItM5gPZnKBPaqIW0Koj1CSHVK
rnqc5zXww97BbhGm1w1v1gwBQRMenJmfiC7++jBsMtsU0rnuAnEiNCVWiWV+aKQQojyjDB4UDdQI
Is8UEFbDxm4SzMuoOp4FK1Cpffv7wrs1wMcjIKv635tFUbY2/OB8IhgEzfn9HrQm4XtrpCJrMYU6
nkfHc1atdeldLeVrR/zdX7B3+jcnA9geSdKqphOKvIW2oOSYJ34zq3GvrvHos6lsPUPaWLTviKmh
WtRKImetyXCg5dbXRGuAFNqsZKbR2s92U+FGJYwu5fX8sCwKWIf3FoC9iAxspwgavo6TAaSOyIYo
Wb4ANn4oa1Hvoj55sPgF8T0SD8x35+XmtmxVmB4+fdFa9IKxdV1ZFEJIzRROuNIm2HnTG57oy+p/
RyEISFuMc85gLGP3Ysw4hNsu0QCVKwdMEtjAbN/Li8Pyi/B7rgP2P3QX50xYQfY+SPEKTrbC+wJj
N5CCwXsyxW18ifwiIRkYChs24jfnDTYxgeg/whKR8QR1JLgmE3/A7W8Qn+XMGBvlmkl4zPitBQu+
VhvBwxPvRzvFTSgcAwDbIynq5i6oMRXA6sNJh6ZmVhnLDQcVG69E+uPxbM5VcX0P5sSNTssU2fAb
6OYdZR8dLJFXxPiVJKsBrMCGo4F612IzyVvJCMwWqKBKJgAusD4kmYnJuatqBbjmlHInm8P12DGU
rT7sr8WbOXtAbyO/TTTYjDVy9LF5ltBpLPnqPnGhmvBDqEu50P+yzYHvEkRzno9PzETnAyVn/cPp
qiucr7sbGZgDsxsbFn+mDi8QK9PbKBeriVtMDFk0omePnKeee/z2fcwcB2SOoOAQUzaI0PXGwM9I
PI7aXEDXe3WwL7F7hrb3aoqrgxoMJ0pI5IzqH/hjpRJscP3l2//phJ5T5ti3CR6IR3yCADA14pJD
lBivACBkUXir0Fsi0JbA/zfUgK52DFBhA0ExFdaPirPPwDJrpq4ZeeoVe7W3gp8od/VL/PgIQ1xZ
+hFlnej1x5Br4hiNRx0Ltl2Wk0Hep7/2eRZ5y2T7qZYFfnx1M8mzpbkPjp5W4/tp/jmpJDN3s33L
6fwQVafCDg478lIwUrU9g9SmZW4NqWSXvYZpiPIW3FjrmkQR6e5CKU/a8IXDant2nZ7mjoYW84Dk
bfP20O93l/uJbcrD/Vcw6z5sHn1GtYGG0CXBIXYn93qwHlhXOVcmYAUsuMPs4+LjQSJBWBJgbLMm
FZmDMOryaJcISmSukJn0FyNAKM1rGy3IwKPmlPVoJaGUnJtUutg1PxoiILtyH/HicP/5Ybj/eqKV
HzwqIb+bwY0hSEsq/C0OH67/fB+Fgv/xGwOmo5l/zKo4Z54Bq7EfEy1HCDcHhfEO6Fs2YRnjABHH
ibU8kI9/tJYSe/TGNx8trtXov8+r+W3NuBIYsvyEz9ms20p7AbyaDISd1EAIKi8RYk4K3aNhnFa3
d+zKLHhkQKHb3teOz+IvdrPokgJ/jprgNPwI0Cqi8UIM8jj4uuY5VXInSuYYpu9RLbVfxHq8009Z
hen7bOLETLGKQPqYP3chxvXc16XP9Uy5SymFlJI3xzXo88QXYUQyv3ODHLk2GvT/kmEhcZ7a8L7J
/lHXjXyS2Bt8vIJMLdQsXGKK1+tclUwshoRm+QNmhVtIref8YrJUU50cJA1h/5bM06mEa1/gwalM
g9vh7NsZyw0h94HApExvLhGUcIbC3oLRI5ktJ+ph/Uhkv0YE6t+ASBfLfbr7rcz0BIh9EwertlzK
YgkN8u2EOqwH9fsAtfJaHWOijs0sod3DiBDepgdDVoasrYwpFQV7XqthbT3Yb314m3BMn9pusclw
g7UiJDzNGfrDryCmeLG327lIosPTDzGp8j+SuJW2BtBykYhszqgNySi74XYnd4lb9B7eCZuTDMdH
E/gcJRzY7OuCqI1YHWWufXYdeK3EQXmun9hsMAbmaIHQT8KI0tgA0RaaLLxO03jRRuMLB82Pf082
kVekNzIZZmPPyLKK2j2+WKy7jrPQaSszY02sSzL7c+RzGnMm4UX0sC12ukJlVVBW2HO7y32M9YfC
fBRWPWFrtbEYCKYDk6vzvS066jc0O2iT1neCpdfu2Fut6eAHUa7ntfyTmFCyJx5r10TyfGrGe50Y
0p2BHjyufAGmNKRXpOtOWOASnxVWySYJ0RRgxwX7q663knez1tMg1m+2B5xebn2s0NXg+c0JDt9I
Bi6e0AkGO0VEtqG4Ur+mRZ6FzH3wiwBj8plCBJPxRwrnOl4AE5Un128OJ+xs2ADaBcdyK6Z/E0ox
Acui+eVhZAxExTn2Ku9Gpfw4+GUEt3mXhVQpgdGsOWtaTlbzhsbyhO7GDKH7AFpVgF5+cvFmXDeU
09imNtpHGu9yUwYPd82d1qO8EZOYSMoMQJ7H0xpfNvq/odcwRUvBpRpGNJkaQHOQ+MumrG5nbFZx
pYU5S7WAVce5h8kbCgbdk/beeIBKeMwP4Iw5EYwIcesylFnkgH1pmW00KQbjrZuJ9kSq2yCL1hMC
TQql1yab0uVfO2b0ArS86OcXmWwOoGNX6BtpD//y2RIMz13KM9wiXJyndd8vzShe+S0Lp/wG6B7Y
0ncFFJAJaO2o0C0AV4yFhf6+3Wd2igvchtd/OMy6YVwLG3Ht4BaCSZwxAcohrDn9mPmwMXO4Cusu
ASI/A87qrbko/R8tXoOvviklb57N1kJLUC2zQvDGBCZ++kWrwdp8PY8ZKutyyQ6rfAsKwiG0VM04
sEkY8aPsUEsIrL2Tngh0nj7jlZI7zJGg101/u9zH+SQBTJLT3AZPDhS/zR1xN2l3vTkosIn6Ic/w
pZut16KUde1lnxVXEm+7jwGEMZIMDkY0Y7pE/TRvpSMmc0P4CBxSDbz0A8Qm4IddhaZREghpRy5j
OkGuck66WshMoAaFMmA6hf060tMhVA3DFH/OAeqg2WzXTt0/BZcnAveA5vvWDZVLjVIC297RR1KE
08g/hPIxzXc9r/u9N5QFRt6Q6PkEgJ4ws6x5fgRK7jaXvWEovb7xKxR7zBg94NbC/d1aKWCbRywY
HKTVRQ+YHnvoMjwXWfYLtgxF4nrzEvy2t4CYGaTXakbRJyNSZjTi8St8d/jrvJgrIxUGUf1FJs7x
q3hczKVsMiSdy0flpfSX/8qvqVORqA+u+xDZ6/JOcPZOsLhcN6eTxKvROXMSvCtGgJaxEh0a5lgE
uAA5foidzWaqnDWf8gk5802TzdvTG1uOK1JO5iH6w2tpbi9ceNt1yCAtMTN5FbRxpxE+3wYr/Gs+
03EFXtNMqNzsOpw+twEiN/Z4NgEIDP1zpwO6XXeGchSZo4Fvnx1D1aaeAkvPSvZm0QxwWBH0KJaX
S+BKn0Nn9hgPqHf5hYGuH1J3PPX84CxtEEZvhR7wm/R9dzBCs0QNMxfrYNYpeV2ZagLFowuNQ70w
QG7cs0VeD7XhX3C6BscS+ndS/HpngbRKC2d0izG1iQveP+3MtJpRNvcOVo/WSIwMKfjimA+7Ca9X
SRLwF0H2wKr3BMcNPzMv9ec9g70q+eZJa9aXTLwJFMz/ryve0op7Az/FoXI+QGb3s2p5MR9/TYRX
qyyuOxGoAuuKxWYYTLJNEXKo0jc8oPBr78KGStziK7Yh6g980dUgjIb1vxDfQM84lUX41XhQngua
HKG2gZeWuytKO/K+xVKKyv5fC3U276vLs29W4QWPYxV8IXzS0gvTEkwz6L7DvIcKSg+FkuI7ul9y
Cn/8qRR1X9YU21fUKSBAkzcyxc0mFq+O7kebJWuif5RxXJgX7sbXwAExgv+QhK398/jGoPos9ZVp
7sjiCLkOwQQVX9QZcLx+DZZTuv6gK+f4bio7zC0p8/tSqK3rBrhrOB1Q9dMyExMMQxOHCoP+GxmA
V7s1y4fiI7IPE5c8IKfT5Z/LjqzcLvhwrUzqB/sS95gkAU7gjygXq89GORiFBVOqFgY6gd2HuZUb
/TaQOgfk04X2Op8kKY3ffZiXeZTHiYF+WU+mmNgFoGtC13MEKp3uuJ9hhto1AappY5/mw+ATNUvI
uyIXIaPX3VB1BZthM/BQw50+KINMhnjFzkLtRFol7g16OdxvOlrZTQGa7XNQbWmnJ6CSJ56t+wir
SYoa3wx3Jfw9U3kMwkgcuL5Oq9h0xq7IryQgTcga/o3W1/4Lxr6gFuaLAiWiGQEQpRTkmrRbM22K
+FXGz6+Q1/i4YGxW6PV7mRWmGkU4m7JRMXBO75/Oe2mYImPm4TSo+lxHIHfhqI8OVU1Gt20EPlIH
6Yn+hiy8jgZxeqAZcONbgqaQ3Fi0luem3b16ZEO5LJA+mVeacm4UEtJSObZhfhalMpkvC186Z7u2
9895MI2Sg7dbUvEV115WKP0nMw9SF7sWIDVZX6J+M77Uy5pn/HKUc3LhLBa7ibykLbUpfBILrXzF
Ag92EzSd2r9UkCcQBRhiZa8ow1SzOfEpn6MQ51eVh/A58RJDCI3WU0amoChx4/9GtAXOC9VkbiCV
2Ufh+jdbkNbBxmAMJN2MUQvs7D9EFiYK2U3INTSsAF7IR7siyYCC3WY3hozQCLPS1NMfVW2RAHM+
/H7Oim/WsLKf1mFY/8VDJP2aGegAUQimXZjKOxdGXcIMnXMnwch8+stYW+JA7l31PDcW/XaNE6Zk
Oynj5zLM3tr2wCp73zFj02thS6wFDR609xuu6R2qQHt8/pYnPd8Vv0eKAe/mPWSXy44T5KwkngZY
1VV/aowcxSuhWwzVb2OWURwpgsLk3uRs793bHAgLOA+udj8jTmfOFCvmlstl9MZTWKwpafPfC2oL
llUvBAdvdjGou2PxfF6hA1p6BSq1sp7hVZ0sWdNCUKV+Hzgtqmrm01rb0TkI7ZKrdd7llzAYxxGM
2GZRxAQIIeANJ7xi7B8diCD+3kueCLlWLe7Py6zy/xUvDj7HNA5g/toAI7efnqcHF+ZOhLdfL//S
/SIDK7/MyiQXU+dLJwykSQhqQcj9b6FpvdMQqE6NJ4xegOEtIX0SkCmTjzxOW6A6mZfsGC+avBpe
ah4NhGH+IFYEnqohdufYbZpMOUJtMrhy4q3N0mMWWRgNEkf2OwXucLBeCX3BloDfGtP3TlIYBMdc
EDdxxG+jE3OOS4tzsHxVxy3AAarFpdLYXklOzLtjsoDugB04nq8RpwlcdReCU/Fa8Um2abftFE5j
46s/4MjoWThC+J9vONfpwQNtAQ5BFmIHKg909BGGXrtmyJe1H+m3xiqirpYkE9onLqCZtn/3wr/d
w0O8ARG3ecmE3J2ulZzEv6rVnUVpxL6uy5u6mwHNA9koNA3wjKvWFRSFOQw/wg8ci93Y3siBuGTm
EdtO0pDFWl/QXPq0mjZ3ZhnIkytDgWyUMRd5rZZv3OuYmg68FskKf7xOatJfWi8KfI2AxOnjy6u6
+NJQFdKF/ORvv+GOKgs/TvbUAMqCL+ADshS/eNrkRBEamIEIBr2aSJKN5bmbtUIVPXb3j/IpGDPq
VfYHRgzP7Vhat850cPpEghx2hMjwUOtyqR/kJQUSTrXHBFnEkMHzKmbOhhkeKHhXmyTtYx9h51kr
eNf5SzolyzHkrjHN7FPaRskLckHTbp0yV0oWWBO+yCJhQOwmh03qTRVFkZzIYMgitFLJ6d/GVCrO
1PCOIWq6tjIkKB41Hlllgm2XJu9KAINMfXo7XDQm+9zWuOsXSH3sLdSsLKCul5JJ2xSgOKx5WkL9
ubl53ovgf22yBjGOVXxhRHvM8DTbYByCw5Mj/jPemiTErlN4jnqjktbQAxWUj+2HBh7vAroL0PsK
hSnbit5PwpeHQX4lNLuBus32XerEfXEc4bHX3vZIcz+VfvnSxNn5jfCT9dJI9EnCi2wuRk5fjW2H
sNplGvzBMk0oTc7ZFxabUE7RoBc0j/pZWHbBgMozpQ+oup5svBEBT37xNmBXuYyV0WpUQtrouJ6S
p7jYL3J26fpWflNeU2Qb8GKGXY6dkdwKhvATY7o1aBkgGk9v5ahSV0FYjbKXrqYzdsLqhoCptySZ
Ia0Y7k52g/PPvHlAiG4jeV02iSNkyhZB0U0oD1kb6DXjiu+oPeyWxdYTke2O7wJhq1hM4yPnq7+N
jgBcEQlISwsq12SvbubBnTGRAVLRCF60EBEh9Wscwpdffn+vsb4MqLkzGdEUkJxYCdmRGjZokORp
wLwHj9oiRYMbZPO12rSn6fSDEYQfK5qIbiwvUF4zmAng5YXiSUjaEfHNFBNHJPHR4XwW0O2XUCkl
gVunJNWIOOeMWODaZmDdcYDtRwzm8eoQkbg+zBJCGQwgvCvLlzEt3nt17/9YBklGGxRnYZtMHZI0
XS/JcwQLcK6QFT1+8oQ8hcKvSJvKXRTL+Zs1L5lSsNmVROW5e8jT94z3C0+Ed3WDJJFBqPkoapWs
L8l95Hi9R0A0z/7hR1MBcqTGhc7VWLyAvGx570CPAYbBBqMmwUrwxm2nhWJU7FPkxUfXdJ/wh1AM
oBNnrSuX16/h/t3bi2Vdt1+gGNRhQep6HSMjGem4iMFn5leGVRFFe88G2maWg88MUiwz7rElNOPK
Fx4/sHjtNxkpxRFUhPmMUlJ3FficQRWZA+09kmJORRKr0a5IruQbsNlD/0t+tKBvF7PkxDReq7/1
6xLNb3Y4CMU8wzR31wML3NB+t8pjV/kHEgePj4bZ168gCPnOdtfM2IuL+OtSlwvkrk/aUI69vbZa
gpIjtKcepllinusImzotTrcSGDBUcd3OLZ30xYFwztpSBzVBKAVvOIY4bqEy0FXvbTExMkQ1K6Er
0DH79VwVdjEpjEeTXlSbhtxPAknmRWdQHC9izUEmeDem+Y56BfTfBMxRi3lIL8oF1PY1qQLuYrPN
M1nS1X7sx0m+J6S2DfQ/gb/FR4mHtVLnGD5fyRqBsiw2egvpvr1yD4lO5IstEhsXUSr+PE9GL3lH
txIW+HtmeyPVjQKqaKtdfUXDIx3gauD6E1jC6FE72kSM9yIBH30rjBGwnQ6UNgiugCkP9cdmkTg6
EU0nijxwabmJRAdIOUj/cF9sSyrHLML3Kg8oR2cSBDeOlf74sGauRB6RHm89nHC6u5lhKzWhNCZ9
dXNcImB7JYo8OqswgzZMvsG1FFht5WKseRwyXasUQPUqQg7Y1tBht+yEPeyq4WSvAtzwRUC7Xmwi
Pm0ysiWi/cT3DjUvrhm58potcfR90t4NZfnyZAMIBN0vcqsoXPFNDYnXG+1Ep/OEEgxfHYNlrfoh
HUrSe52pcNGgKA3MN2zP2WKtZqsc6JcBOKvZdNcKUdV1WS+MBXflqTzav42Dwqup0LZQ8gjxsQ6p
JLJt2pSEeiFktBVsFg3AhEcLRsIHljfIPymIhrnmEgmwTjYGT5Nuro2JIf1baFrBAW3yJsRiLgTp
d7d6m4WA7TNS3MEZIiv5RqbA2SzJaOQ03Dm+sRkp0A1M86XT48/uCToML7VKlgDa1JPRLXc83a7O
ONv3EI/H+EcjApp7lf6Cjx6RPQI7lFYtY6hJH4wSGKGFe2MCDCLZDPkZVivl8uoCuUFvS4gttHjN
RbSE2hfNP/nFa6k1ApGDxQApVNvTZFx/iWsnXttG2O9akRsP0E85RECwOu9VnNH+tGGyHbpyYGXK
pgDne6KiEv783DzIqq0DqyqB8n8un5PYH8xoZpFvlkJZUvDCNDTkCPaXKheV9ikezg4JdXzs0655
kOzX49yCP0IgZh5mGO0ZvkJouR904qHy57lmCiwiUqQNmLeFZdfvVJltMw+clUR8z00aj+XZZSUk
DKzVrhFxcWNubO000r9TCg5qjSZk2iuZhizqvHImGdL4AJU4WthXrWMHvxGqldmLQzBpw5LVX/wt
020XE5RCn92pOwNTEedjZMdpdIqsCYf7W3dW0KDkod+y3a0e76LQpPwGJWnS1/bULxP0+JLFzWFm
lfzDHeeH11aisnfJtmQgXaBm9gyp4udnaCJvmqJyqTs1o5zu2dYDBqpZ1e0l3oWkOtXzrBpLEBUR
A7zZykyKWKlCxnJtxpU73HbAch9ANW3NtApXgI+h+haEDqgjbxruLJyizE487dR1E67bpk6zW3LS
kZu/3082bDmdMCI8Mi3rqM/QtxhA4EpJw4MI4z7bOvrH3GO5+Z/FjYJ9tt+vAlsBCvaiyaxtrILY
3awrd6RYhF71sHCD76tf90ucNfQX4U4nD5iFQKckprmYB6/eD54Y+ZQm3rApcG5hRgbsxwUG8LiM
+LyEdpfIHME7QaKaZq8AfuMKN3Zwfp7m4hRk81vaUJS62fdZXN5ExiIFXXmDwpbFvmdeT9nkwVXW
vcj+r04e3F1CaNCsSCGcrFoLXmt+x3SInK5dJNlsCi/JWplJExjKDcdIZb+2Hxw9SyZbplWoYwMJ
3WPQ/mS7hneN+aeB9Jwr+9mKhhjLGXIuRRoDg+fNHYnhH8Mv7PWNXTnLUP3ZOEfxzPmUUXNkD3Ij
BCvmRPO3m7OreLRIJOn7FGTcrR4S5mVf0YS9QQVAq+u7x2hUhd7byiYhZjjk28PZ4XXtobQgyqLr
srX2DAA0vC+8YwDG1kAN5SwlqQV/uXzJpbxRorA698ly0so7knQjOBiqeWmXl6W39dfwE/Rhgr0Z
w+Ra1kVv2nKx39w+9gNAK+LzKqme/XPN2RKGcGEBBUaF9juLM8G5eP52TPpQPzgSo7fBwwMi4lTG
UAikZNwF1dpitnjg41ONDwqdcfHFihbdcS4ss0J92wN4F+1l0Z3BsgAlWOmP9tCNrGd6sdJu18kR
0oj3YYU3Dpf3UrKPoGYB4f9nSd2/q1gDugwWRrA1o1yqkW7Z/M1cWZ08+EM3lPANe0yHrlPlTWXX
tmLZ2bVxyUUqYpiC2rP4BRHqXRVuMrrrDUO0ttXBkTNxObPA27eNyo9nm4wrSfgc5JkitlV59dvi
r4V6N+g+ywYTMBDSDJOmKdsd6a4jJQWWdUusdfpLVCNQvnXTvfZ0d70gZAgNtgpHHvtj65Aa+W8m
HwrtZTgzvPY+gKOzTX/8ikzQQ/LZIzCrkZZ8OlrXAgN7X9toiDY3al5N0RY8s6QUyvZ5TsdlPzUT
Pqr8BMOVe8QnQeiISupKi5dJAYv5WRtQlHiEXSkZ5XAB0nXvXxpOhlkx1MMA3i9quF8HEX2tULoH
dho4/8LNLLn3/XXdxEa2/UJsOrvm9AV/pB1qTplauVn23SNvTyn/8FyEEbNXRTj6tkKKA+Cdw8QT
lGb0lC/YzdTWJFfYPdborU/92JQk7PEuGnzFjK4Rmxr5VBSdahg5ZoN7B2rj6QbC3Ly9tbCyiG1W
DoYIx80qdz0Jhf+tFhpmpQZ98xQJsvYMEtmQ9bFW4++oux83MyLKEKWtPHgGSVKJd2uCPl51nBBY
HRXxuCTYZEWU+Rwe1I33AG2F4m7aEwHk1sl4poU9JH6Zi5jOUFj1f22OCPRCg79o6FDQf52hjk8Q
W22vcI008qSC47monECBRiHgUi4ia4BT+5YPAY8HwVpbNxxqtTLsu8H/e6HLOlEAyX9JLf0hdT0a
auoFtNmfC+FBoMI7qLaO+kjEtPKFf1ymG05JYx5Yo7i0qvm2EhRPQ6UbeRA3dVWzx0Bj91a0PUWW
+hjx5ZUbT14dxxCoGS0K15ScEeCzcxVHAb8D5kEw4k6S+hWaMJlt1mq3/4vMAfoOoT6eYbSHherx
/MRMbZfg9Ix7DeJ8lp1W3luXbSwQASX2CzESxjeQQFHuwgSENo3qn0Q7V1CHpyvN56uF6TtIPMJD
kV3Gx8Wr9WAcrz8eDrwFWeF3sn6FwEHZvcvKb1gFLhNVKEtCPMTklvUlxBoDqbRNLil6knhYJQ+a
t9b08aNqSl8MM621Fh0DV/TZ1Tl9dV3m+b+wSBZNKmlXpwWPBKMQ6TBJCKU1Ah1/CXpFLNyesA54
dNp7LrllCH0bfNBtSb1WxF1cMIkgr5com9hO5ZrSmNvFrYfL5BkuZGHeFz5+aahQ8Bfouv41IVRa
hpWdtwykPa3hDBWkHVLgKnXsaXa+aKVIYXS9N/dNcC3tuIfjOxEYWJpGih/9EUxS5+NkXXu9Bvv7
z8R3CAUPShw9THxb5xi4Fz+26aLqCV/EtofXNELsrBde0yPVCUVSuNoqrmGzZHngVe77OXOhKZJa
QTZpF7Ypg71ODz80/9dz901wJVRG889e5yvpRGl5IMTPYwxNM4/ldrOUaVRdN+PEAMIhcJ4a5TBI
ovCaytxUcKv9m8E534aBBcpMXbrIshPZsz0sKPcxdaLBBGKF+sZnaCMs4IUFIVm3U65vfXR+enz5
D6yB+Dc5fRowzhYY9AarVvG6khEBJm8x9flV97C2sQx6yesT8P+aWpg8a+v1HgB3a+O6AupH47+s
fsOpw4+lTlTNlVXi7/Ayur7L+ZJyiqKmMOsDUvLWSPDkgSg7GvOzkoyYTKFi8xg2SxLF1vtydA/e
8in1hxj7VNbQtG5TEq9ev3eqTZ/IEBez8KC2+DnQ00UWeZJKcFiGPUReH5/+Tmq4cQnaqgISHDXX
E5G5A1IGraqq3YPslCTMadAf/RuJVhVyrdZaBjvmTi5lf2Y3doRL+X7Ky5sP1DWwegelHQtxSLXC
oArM+WNvB1nxhzJ5IZQnTl7N03QwNhYRu3SL4zkeL4JYcefh3SY+VnhO0b6wyGKXuSL/W/RQG7nd
9O4XhtFZ9EpVTvJ0IpJB4Hl+AQaCkFXQygPTIBTBOdeky2ndeDk/1bXr9i1eLrfenQj307tTnTih
eW2AGJjJI+TYPt4hKy1P82C2BNAxMIPgpZir/QktWHikKjtC4GN0A5sFXnw3t4onhuLrjT0RKMIm
bFaoVsMzyEENpC9ELR+EVKHKju6rGBMSbhMVR1rAiMREX1uld/0idPpGmcWbiAHSl7m9WBstM1RM
fH8rK6zXgTWJJXPZrcqrI43dzhz2EQ5HatzhX3WUFoy+fGgf5cWnaOVA4h15b8fiAxBPTpL21xf3
UfERHquSY2bBaxoHPTpJxaxsaNGIWvx7AtJN7Z6MLytJ3iLK5ADQlRbTL9HrT/Cb47O2PhYmjdkD
Ss8NvGo7mu6p3B9J2n3yRgIUfrRRipOZfLnGa9IVjPnSi2L9/VprayKw+M2fXXnU/iS8VVMapBhJ
LJOk2agviXIrvG8Dx+xlw1h0sGySRRqOHtczDvHow3XztIHoSQFn9vijQpTMvI11FJWg9iMyd6AP
dnpzu/REgEecxCZieA/rlk4PQKp733iWaIGcL7JmWmA9Pq4GrrmvbaVDPFCrrrkIFInLjvNhNIsn
VIr+iTe5/YYZYxKdxtFoz4fz4bwD+xtKmGhEabScqIQcFU5W22QqLhJHpHWSwTdhEPiRVwLfvoYr
BGzK9CpjKy6gCKXNUvmeb1+CkbEHO2WhON51oOOsC3UCPwRQgppRvU0C1od4PTI4XY7c3cNNKxBR
vQ6GW7+iawdP25kTKMwfNB0dRca5c6TuTTn/1dFcS+ZEcnZ0lJk3jD6X33u4QQZTXzUdFZh9Bs36
vEAEMC7XsuQ+qJnaGfU0IhtY4WXHmQCzqdffdebzVyKwCOFSjTNqIpMglEaHxYZPie2c9yz14Ubq
1G2Ybx0gFOD2zKmHfCSZofNSFY4ZwpPb88syfwP5BZnpwTeo1aS2pYAMZyi3bUTnmFPKWOacEc9M
ljbbwz3oQgFv77rcEAwHqm1iWi1wtMFpvg1aCqyQeTlTjr2JU0+a6JOV3r7hz3iFMlCNOs6zVK22
dchDuvpP3tCkvbGjJEUGI4qArZ4L3L5oO+XBfjvpQI7/0+Y9LQU4UVWcz0g2L10kj/TaIx1k6dUM
T4hr6XLdIruTruUamIvW+nQikMQeD7uaKscZ5zhecR9ppdE3Vk4SU4pvs/9kovmpfhYL5eoxWbpA
RBgKF1jbmMWutnTHgY/uyn2pq4LzWVnwaRGUew0SGbICnJVMZp8lBLrORUvO8jl4A2UP+qU03S3y
Bv8AsexkjBSFs7wBTRwC+BHAh/jpG3T3xsS+8Gt4C6yrAizjAibE5NZWLBs+Zrrrr2OsLMeu3L5y
kf8tJ9Av1xexuEKc0nLpFR853awtv5OLNDRNUVDlARjxruoCpSY7Pp019g8JUciSInUx4yoHkt/1
ZJjlOr/cRhZ8t6EN8fvAh0BmgUktbaXb2St8Kit2/xYwYpJuXXPtkSntJYB/HttpZd+dh9Ncei+q
Txol7C7n0Fel8a4Bma6k4Yfh/BqZWmHPtnBNdgaMYSef/SV86MZuhjSFmvsu7Ur18gO4uAOyZZdr
UUf4tzPUYXP7ORUGQe2fXOaifaqHSiOm7zVMXMurYz3sHUOq39CeoZpVKaZkXZwNK6jfarIZ/FeF
ay78BjLbl+QWlbl/kkc1ZpRStcxa1QNoC46zOv5C2x6/2z2FRrg3uK+8oiHf8g/FaJ1/tCeLtlj/
EJJWSzp6oLPqVXFJFYBd8tdrkfpVL8+aKD2EmL/sjy8RlJVCRCgwbPCMqp2+IXBRe5uXASiXIJvd
smFucaECxLNzye+U0XvkGJyV/iEPdA+WVxW169oxucSJA2IeOwXo2gxonKSzjVYbrUSyCLC3wxa3
OeD3mEeq04hAsWmrlbYSUgJrlIFSwiuhY5FtJZoJKN5WqXHf7v50YviahpDefGYV90iUx9m4oqr+
RkYVZWxvnqzzrSlFePd56azPebYQzushI15+v37osAMDeivLe3xnvhUI14h4OhbvD/X/J+BJpv79
aJZ3zzjqeVY+gKpNHcvXz9Xd9kdAazmx9MaDpN6GRE9KN4alnUhyllYMpS0Anwd1LHHpaV8M7Kd0
absUIR4u2Lki5k/lK3FrHvl5LMSZdcp5hSB0wP+tRP+WDqx5i8IhIpjZtMH6ov8+Xez16UvGBEKi
4IwXzDhfjTimUjLQgKcltOuGGaa990tD9CpwFSe60q1XiPuYHOtmSNwPobuWOTOMzQn7v1cRmM4D
khSO5Iy3+ywXW6nKA62y21IDSMku57X+7YtIrOdSF6L8Avt18/HgXO5hzoHuEY8grSdGlB2khCxa
a00PeNjxF+EOFeU7uD53SyunhlkwUw9bYuwIEFVN29Z+Q3T9Nmtli8lqO2gYNKVs7rThL14AZxvi
7rCvPxca2Ec/kLTA/+8188QHFscaO9rUyv/KgVAOn5g4j1X8TTrHwDX58c/IwjI2afggXPNZd19+
glYk2OVahST/HYGyKSNrBLw8Yx6eyjBQTXcgqmhyjC8T0zW78s6fY0w944O+V8v4577u3xG6ahGZ
v1Nric61f1orpm/6PzBnFhCnbf9lomETK62FWgMOQzEoPsQWJUe3AU6NRsVUnOisZS47ej9NSoD8
c2D/12Dv+zA878oEGtzZEnX2lijjC+wrI1BltmotMN6dwE+sgSRnCXuowMOqz1E1YGkv6e6Y0BKC
13aLsA+4SYz7mhFIVEaX2pnRKQMdInBOnL7kTZxFo2VfNsOZ9InYWUbXZRx3/y7pqBYElUqfK48D
keRo5dzB30bUiSeP+Y984VVLpKoLeIc0N6MAS558LPSftGVd8SQFWKjXfNBvLkZgeh4LmdjOAQZW
RFokXMyH1X61rehK8y5ALYK8BBUNEe3WFEMVgrNqy6MD0cWXBsmYQQdhl6/DUH741nC7wO+yWgJO
Rbzi5zhYcQsP64XP1ubaebXf0PBroa8F87sFnC1IYLwql7hjjyxJXdejRu6/TrVbCiMhStz5btXI
JAFvIUCZBusY5nido47Yeh5V/7n+K0rl6yS9bEOeF6kmOpBTThxEOioX1I1iTb/Mxl+HXlc6RdA3
a47uUqxodelco1F0I5LBb28W4dWZvfWV0I2cyqJT8v5LKeyJlGM3l4a+nF9h09wPldFblKTlIBPp
7EEKCETaGTh5U//tFL10ryuw2bFIW0S/BRTsPJUarN+MezkePXi2S3MaSKYCiDZr1lSIuCYe7DvD
ZORc/BoEJCiuZzIgw0NGXEYVdYg9pQVoIECqz1SCAswufWZ7FgDbJiwCchTTtmHnTTGhrrTkLpzr
CCpmbR6RAwJx7NVuNs8xgy2zhU27C2LaCzwwJguPT8SnQJZK99njkbA7GPdZN5IRiv3wSbYixUJe
yup0lzcg3P2g3/y7u42EwTyKVNM2n7Y4EjqNNKyFBdFYCkW/FYuNXYsE/avGdMv6mxHDGfahKRXO
j6vobPzX1cp3L3UeHub5P3oUPkafiizpL3vHpE2o/FZeRskexNEL2iICzkRppEk5tEyni8VUUWDR
WaVSI6b7fjR2go1N86Bd6w8pZxwxpQ87g90g5QA2RUxrqrxws3WdMXkFhXjMAzMbLUlVHDSi1VUf
mpmtBWIulQlJcicRXHF4z2mECMDm7i6I9Hr8OwQFqCmvaBKWmeonPuIarRYxS0KIJXvkbvSQFERg
SRVOIzUBJ7rKUb5yweRRzbnr8puPBPO5/wmUPTqz7m4vuEYYmZ7BaDuiaxi0gV5bjasyOg7YPaGx
BSBmIwCqUNqW28pIQyVX9hCWGlWAu2qn7DnMgvm6a8MJyL+7L6Yph5QienfZDDe92AHyBgaZLTGP
AFPuKok+mHE6+9AMMz0W/MjDQX62hbxn+0A/r9RQehnaM+ZylCMLiYAbzoegbGPaUxz2gsmnQOiv
+oHSEJuX1ltZkvno5Do1rRJnoddWmnsGmG7nhznfzxz2bCHYjulx8RWTiy8tsJOiEVb5TlTzZkeC
uijtsHTBiOz6o/KTOdavme10vYx0toznTsbG17sVe8TiiFyTvZRSIbtApcAxjtCze2weWgtd//Rt
nUoqQ2TaAigzOrcrgz+2Gi5cpI3v4YGhJO2+WNL+ZDswL/zZqc92G9Tj6EEdSkO5J08z427Ryig2
DfbuIP29qZQZT7jW3p3+GEEOlTTaBXq8tIHKSeV9QixI36IsVrIMzLYYeGA0siLM/cXaM4WcJZqO
ZkbSF4/Kx/SXsfF9WzjW1EUPhMHtYiDtrhFCIS4QeFsKGB4hjVc0lJ4JUh6G0nAouj2MXpx7yUvj
6QYZnuqhfqEmKxF4iCF2Jcw1V+ge3xROggzdABOWX3Hqvvwr5EAgPdxLh3dglzyV9rZ2mv3RHkq2
HCiso8AYRFgkOns29DA13E8EIQA7McuwGFs7u1ogHUcIj4XaOOpUBSDz04OwRQ/NTquglV1FoTMr
g9GEfHOJEJJyOn1Y18bxmums20ja7BqGrUg2PDqrTc+X99m3BPhhvw0Gt1Syp8D7Xs2XDhQuMF5v
xOMTvA02gou9U2+3Stnhknp/P4xynOX1z57rWaXGfkLCrFeD/cR7EpuGiwEZ9OGoVzHDpkJ9Xn7y
MMRySp0BugAuCtnBa1p/juBzP8meyeV/S/mBV9nyRdzLQ9uRGQECQ089oKu4KEFxweNjTiWqf8o2
XLELJ3G7vPmTEYT7kqX7xSUPxG1TLYu/LFcvbIvHAbDdlK2Y834Iz/1EtqkJcghSCKwhSCwC2K/i
u1fHqENPs1bWklFOpqyXm8m+GNmqobn53Gi+XCAksWNSMqlHFp3aZQ8nb1DuTEvOwbfuTEPNdqrD
ARemCv3kA3DuUoCKNgbDsrxgi8QM3rpGyVX0Gyrpq6ZlgKaJf/Lfzo8V8wLKCPDO55IPu3hU/Waa
UYxPgpT009bE7mUP/utTQ8yqaR5sN2QoR9p/mkMp50pyw+QXH9htBhFRC7yWpy7GHcucN2AcQBRO
5R8B+cEf0WHwBU56SOeT4UTcZQA73YT4mORICN9c9xtXGHvGpYxTcElgF3y0BdAId3OJtEoaTZKp
OBba65hHd4DXKx6BtBHV03ssX9HBPedvxN78M/rvXogKP6+Ytokp8QCX/sNWdbotCaL48+MMF3nH
RsAoyH+jAYwZc3Z/I6OMcnFT1B9IcRZDLUHBgC8/J/8WF/9MKQCrc79/sHrpOzXL8Pj+gQCwRf9M
Y0SHfd3v7fgPmsKn6aQaiDaSq6yusUcpFA+1c+TfXr3ZAbO8M2v5FbMjd5q+7BcrKzOP5awbyIMV
JsE8YdkWIMR8e5kwat10oA0aD7toOc3BUPloj2fec9lb+EVEMDjnH/0nlVYsbvi07c5eor7SUPZE
yHerP3y6+gkhYIGVLRmZI424AReST2pWMmFMZmdqRMKT2AURT7hYq196jUiPfSAflY20mw6myZpn
ctw3nyo8nKpLLFjfJ8sGNrRDg1UmEkAb8OtfpDpaqeq4iO4WGteNzWkXCT1Mrf4BoKm5LXXtM/7f
N7wXLbfioLL3tjbMHus9IoXivxaBiVxv89qJ3p7G8+1TgqJBK4Kmysx3mNTFMhJJfTSNCoAP1gv6
dBgBtczv/73+5/WooauwFA1uptpAifLsbqdiBu/HmLgEkoUejNXQVLwpRA3j29tiQ6Q6lm/53hTV
h4wH6/+R3kifJ2JE+ERKED69E66S35Hr1Y72s1DxvmZB4wjs7YjP8P8XYsOjb5vH6jqtSnJYmzhz
IXd2gAhh+dB3DKdOKR6qR/jzKNYZocrw3TfpDF0/nKCY0nmEiiRJG+seYAywugrcocT3SISBbNy7
+qqybzHIncq04rjh6UTqHVlLb1JhXn5lGvwgtpMzAiHKVv3boIgDVMN3dOpJW8Br2weoM6D2VEPx
/BlXzGnAKsppbsiSJ1lP51kGoPsWs3yVb+SFmpCCTahI8ktXqLv6X5WlLcYrdKPuYXcHc1qBn7HZ
J9wM+SMPJxIvfcW2gtdoxJ/5Fbzz6DBQ0h0Q5kfBfgOEz/XjpKNJn5yKbcKWdFV6QZdqohqGBJm6
gUNPXKapHNrm+yoD2VTP0kU+9rypEmSFGs+Sv+YQLBVIjYTEQy1kJSM2aeO4UjO7NLoE7U32WlLu
dMjZjHTpWoHaMljX6QVQcUiFcinw4kiTPdpypewqowWz1Scvi2mjR6FZj04gdxyiZsI/KNBrFQVT
jYDFxb++mrDA4ZV5yH+A/Zukj1OCE4qH9hXcpghaqsthg30VF28WKt2Dg5I/XsZOp4E9bF2ETLQ5
wd6qxGy8ySL08faBmw21VFfuKW3om8cYF5fGjyMwTXL2Q/tMzykDSXZlOksyy76sLUoU0fySMmUf
pZb2krvLP4X04mqWemaoZ8wZhvgl3rFqvwiYCPb8i8BT4Uzd86rgKsNo1OMzn3N2c4C+SkLC0bkX
/XD7rBkbJBv8c3v46+sQY84P4wWzkyK2Skbn/yekhCkuq4U71dXNwetoJl2HY39mVnIIKoFeSEvz
PC5XhRJ5ot0+YEbJo9GU44pk7Wl0G7Vddj/FlQfsLNYz2AC1FY/xCZxVBP5CC9RGlLQCdj2Hd5PQ
XABV7vBHwrng/3udrvpjtZFWVHPl/bOv1I8FTh1IF/hABdoqE43Zq03K1QFXd2SAnYiIIbeor4X2
fU68LWIwexaVK/cgCokitbO7diEKnlJs1UZtM2BnfYJ9OwbFJY7ktGut/++m2AJXBrxH9jyTvAL5
/nPKmB4nRv1+PiOYKn0I+aiQjFuCcDw3qaKQB3/Rpq6PS8BjPrOcaTL5UdOQe7ZZHlwNWGeW9ylK
chnhdbhHZegv7MTSE/qyFKFy75dYHaDxjSgLm2FC6loVDXfJGYAX7PC65joBFFkvq9X3bOrA4mVm
hYvMjg5bAJHAATkMkV8/MGvgn3zDDGmNBb74WiH8ZoC+6pzo96bXrrMhfn2eNEF8ZAFYsu1wzz55
z21qgRTrjVCO4JVRnz27R4edlQxdclKvyFbqqrfjLPYZGjD9Okv35btpxY96KnqflAzHNCf2sVgF
OPoz4z6vwCMA2lhua47WX1ClNAOwOPvevLgAqbZrn9urRQy5z2uU7CMy/kMa6S2N57naMRpyZd08
LRq+suIJK8RNvlFoUFVcPe6UWJs+INNVZcW3oP+oJXjsJchhw0lLfrnmiTig1ldq4EkRdo7YmCGp
9UJU9t7JUxhjxjzSl/gAcGRk96yurgWUq2DdiWEonexBeTl6nSJ3UTcaSBfoecnpALFlJTamXrD3
yyK1cXHYw8ZqQ6Uf3J1kJFYn1542B/YCGYFJXLZM3KwrSCozbsn/uJL42GdHHeoPHN1yY/xYC+42
BNYH7kl542k0APSF2Cr74WHZuo/ACk1/NhhwI5jQhkCIUAF9s64IQbtWw5QN8okHoFvhQzh/NkC4
34oSZt9BONupypW+wf6b5LNQCYOYdhFxBfBuOeAoT/E59q8Ol66lMcxK1tiDfxqK5Nq8mkX20OXm
iF1yy0YfGBrCpfvu+l47RKu54Su3avVGdnVPkEljKhNUKmY+AJyi/rbYLx8+QUF6/wO+mnvQ7TOK
AeNiyKTKeyp9HfIjCKr7ysBbd0i7ZUrsq1Bx/9o42OV7hzxUap5EnSg5nX05F8Oq3ah4Pa3VwtIP
PoTOrHi8AsXI7xh9i2zoYHzfdYNO/7IrAxxmCJIo8lVPniJggv911vb3j1NkEg1F2ICE341gG/pa
9mQCTwRwLUmkb7yE/OpNJsQVwE1aGX5oXkq9c8OtvXE8P6OaK/n22w8+qq9ibZXqbGrSzirHzUo1
iBaTx6mEkemavws98FwxtxpTFfwl+1KtFyj+J0seU6lczMl1BLdkv9GXW1mLQALFKDRWtixNhCBu
oDQuXIQmtAViNC8LI/+3Akq8pKq1eS7neGTsXYSy4mGtnAaTF9BINnMcAMi12whNQauuy7cuQYB5
IuiA/hc1aJn12DRsksuKvzvTRpw6+ryJQPqEeGr98D2QF0z9uLR8I98I4P+YrpQy1nGgtUmJn99J
GRi2wW+BISmuJeOw7RIWtJoYjzMPn33CxAw7Zrg8TAHD325I/uF2rQgXSG9eqdBPEcQBkIqh7fcZ
ztuKVwPNrb0VH2nH58V7+eRyWLnQDsjo2GgmEOaeaYKCxt8G2atSVSeI8/RnWO7JSc/W7fvwfag7
76Iq0c+joBnoz7MaJGsuqNd41Lb1CuE1UOoJfSeBs5MrhhFn9H5Yaz5NSB+YPICoEG7QDUwh/T3z
3kkkZBgz3W5TuSIL/Xf09fMSk43X5iuxyQ9NNhpJy15Y4f7wcca8ptBZgeavq60KwAt+gj6XNctN
gcxDIWEtplwUhKmot1h0QJ1i3GEcTN2R7rMVq/u3gXiLY4QSSqJOqHoW0KT8qYNNzfXJONFWmq7w
8Qxx9okPsYMBVaMTMAG/64KqW2qEB6H6LYfVLYfDPULZpItzysbIeOihnpnNFJRqlJ7P7Z4aZ66B
RbVLfGZ6oYs8vtcvAbmdrepdrPeRE/qre2dM7eYKUcRN2Yduai7w+Eab6D55io0h9Wx0gdrYWgq7
kSs/6THb+3t8pdq/JXjlVzhB1GngG0A1VUTuQsprUTv2ChkjVAa41Mj6egt2h2h5A2cjV98mJQkO
1bzAiGAU/+bq2zEm9z5ahg6FLWS6P+JluiwFLKUszPDl+qh25s0NcHzkfh1X0lnU4cz73vUy8coV
zZIC5Flpig5luQukrevOJX8knQ8SsLfgBeyCrildnOXnA1PA1Yc2t9VEgKNsZcC3tZflW4y8CYAQ
zPjIrgt5zwDNQDP8ZtIHD8fklpDvjykman5UCRK2JXEU6wSLVKOnt/NTtoLwtc2red48s76bpXIM
0WuqQczLyMQHWB+ZdJdybzisy2FJ+jZOOn12VBvo+kuw1M1AAIHgwqq3h6ifj2n7SEoG1MsMl9V/
lZBWvp/v4SgnG27ND1CuvQWMumRRSt2HP//P7XUoocmk1VNtqUSZMFsxh6C1k90Ue5BykRfJfAqG
AhHK2Ixe3d2RD8vUJ36ihTtY9/vYwrr0C7eZLF3GlZY14x9a0nxEOmZ3RlpMvRisadKoUph8sENN
bCTdgh2jP9ZDmGpS47PXVagTWLlM7xRWHtpdXiGGGDqy2rxxHTm+imLpmVa1K3By5i0XK2Aglc/U
xHFuZTvGiGJ85jJ3EOmV65gkNNXSPyvI8sPuCtZCNX35JMTkAZ4DVWTnPuuiTHGB51oOemjxYVlq
Weo86owZwpGjdOE0S9vjIf74Co3Wi8su6ioqYB4RuHy5oNZZKs9m1jyckRBKNQAtKAdA9kWKpTnN
dtupWBelxvJ9wCfcUydf0j4vmjmMIrj0qlDNE0SFDWiDbDBbDMNBXFKKy0xfcIU8Vfntu2lcltwZ
nfVX9wsKDQKYuJEoazkY4t4uveVpp1KCGg+wUUQd7I8meVNcPNdVhh8yp8xso1+MBJ0BcRj19XwS
6cyjQl+nQy5kXQSt5X1zlIsPtHSqC750QCBUHGSnrPhPxgQB+TcajDXCoN28udZehYhryNgtFKGx
0hEmMNqlaVIO3E7Gsclt4aJy21bzIa2wfZy7el36/cCRBPiCEAnj1F3eorQ8ZPotoBfTLoPRT7Vj
Ty4OX2F+skikMkUsl+G8vpFOHVUOmuNVa18tNf+LGriKeZdVwhi/0qBphiU9Cw9Z33kTgw+L86Q+
LVK/llMboymxH3PARqR/oUtShNNvY9FtNtHinE/ZgAMd3b1rNsZ0XnI2ik9Q0EwGyn7uoGm3aQA/
enR23S4KnBg1VnPw6Jcd8Wgj9wtWfTYqh7H3PbdkLL3Bu0O/L4bG9pnQRvNzNckSQaR7jyt+YAWu
hiTvxN2nZapMfR82mp0TdqfaahH8xDnZvQD6WxBvmJYi79x2xGxTDlWtNxEwfDuW0YvwggtG9iAy
FKpjDlsl0uiMCEl8ObvPhKCH/fLERqJNHeeyj7nARx5Qv4ipG9MDaYfRd3Xd6CtaXw5QpUdAHs7e
L5Cii9Ztzc8Nsqdygdgm7iJr6r1QVVKUcAzE2Ud1eUCSmXhS7zf1G3zHceqXrJOYmfBZDwfCJ+Dp
NNOZ8qlvpLR3NauNMX8ffxIIrR3TQBubrEm79+O7THySNH8wL5X6IZshXDbFcJLS4m5fKjmFvblK
BubNyxGkBdTEoxkMQdl60pEj+Aoe6hlazviXrET3iqpVbxDQ96fj1/1wHmSscqZCzcNK2xts53MJ
NcqiAFFaPaeBWo+5J4+EGq37G1b0VH6YJEf4Evw/x029npx1l9AwNXFMfRvtizP+mjA8Gr3ZZrOg
FFIf1CbetF03YHoZqsUc4zC1QSiA27+79xE0fsBVUajaHyOx4fT0jMoaotfoCCSAkJgnTvnSIS6W
7wzmbexNmLcT0e2cdnMuFdBAivurQGImLU4Gut0BlSr+h+JzuI1jNYLSH9NHHmaBTPJ1Xg1lQVqQ
IXdo/5T4oZ6Mcb5P0Ro04fwm4jUVXv6P2YfXYy5cLfvdgooei7kJjMNstBT6pARG9ihhwbyqOkGA
3h0nVAM3YHjMftSE35kQiK0/IgMJ6oodZ1GsIvVpO5MaStea7mNB07Ibg1jWx+ivXHSTasHL7EDK
Dm6HzCv+sn1WDFzyvt8XFOTkLNNGvz5OhgMPEfQESG+BSh5QPE9XkguW+WLTQaxseC004Jk3NQQd
1Zjjhm60wX+DdUpGmMr0wGcW47a7c0BnI7PWKMwHRnt0VS/oPFfia1Aj+HmSV91W1AXPLsAXvgkJ
VU6zGldJQh4tX12k4bcagpdBk7LcRGda4O42Lff41YU0AeGeJHB1Q/te9ISRVJ/9siXWzoF4Wfl1
6kO5rMveNrAqUe1TK/GWF5KrvcOavaKOKSslvMiil+VLnG4OKEtSnNc+4nt9hQXgrxrx0sCjJJer
rG2uzRdTgHNqAOM7olZakyPto0Z1P04xn1Yl1b8tR33i7gJRKwd12/TSy8uBCBE3oqFrqrZNcINI
bLB5Nk6FcHrUmfL8ZwyYuviek1qq3ohd2/AlnmQ+8gPhFlzTWRsSxse1ZR5rQ8JmxEUD8z+DjWDD
oQdeuIKBzOJVLk7gNVmYhPQ8jQRaAYhokY3xdwzIxvF+E2I1QR7H0grbNg2N9UzzB3fGWqHsuFqB
00Dkm3kXW8gPt/ywNuUdzbvktQkNF5vTonqZFE9aiszBPYRpSdKNmbTQa2YxHcLpPN15yp2212MF
bwA8KKKRVzb4s4kXXzg7XZz1/6qOf+TCzBObSbEjIJJVQ5kPRLxik3QyjtXRmNwqJmIWZ7n/K4PM
ZVb6LHZkMeVzTkQhA6oTjxBd1zmBJQRrbHn/gRSPSFHlarnpflcWxqXFOhiGTGixQEmBCudgDHee
EuYjRV2cPfJ6wU1t9lEPU46bIBLmsQcjAzcPeSfiW1A5IEfvijVqwC7WpAYOQQ5oYab1EhRVENuL
bvHek6JJ40E11DbuasUWZ9UVs738UEvH9J7eTBTLLvErqq8wPhzY4zxoULaqzq8q+NOqA74kqdR9
9p6Afu7s81t5bbZKJ86+L+d9Aufl0uF0yRNrEnFg3wUYGcHae0pbaFgMj+RowB7RE0St0/V6k4TJ
5A2Dpl0D+XETgN+Qcg5dlkpkqsu38rLRQ6DoFh7lv4m2DA4HFs671BQnfPu2i38V7DHojrd/P8Q9
nuOXF5SI/khq1tui+r/Il2VE6R7PFkpZOPyHcrVRxUvmNtFpaJkFD6o9DbmyGGeDNq7AWTtzKOfi
AldbR8MD0iB6aNUANkvZY3wuP0S9bmUHZfwppbwlDbDmD2bZ9vhqrX/vIiLolkfUDgtsbzxVGPOU
tLVO5wULnYsIGXKg4EC+9/LYGA314Ihm3WNXPhZ6nBfJnOYrhamMRq1xqJ1jjzFs0XClE6qeKyjg
f5wquR7feOfvOEUZSeY7HIUzeeaULj6DxlZxLvgqfqnf+GPcxSApXIojGUATjbe17YSqoHehZgkN
PJ4DoWaZen+lnNGjzhXRvAaFG0WUEoEPsXmRwHOzlujdvgPhh2OiMAoMX1G9IUkcIPBn/BQ3Ur48
U2HxEWy254QwG78VR5szin5MjacRYloSf+8AIaAU/RzF3XCtiI2OxV4CxObpDAS+XTruaH9EzT5C
sucClLPshnEuh0J6qL6xfHFja5XXUhAjasc3SLvsUlCHkIykF3J/kFcvP6PK1RFxnQzvuUMXTQ6n
+XQJDnh4H/vOV2ffk37UHPjBlhM5Zho/9PzXuclwyT1+QTgmjHlcBdRw2ft4vT3BwOolJcauOCxL
xv0bUgAaXqsxT33DBKkS67iyNbiLJIxyAjIsZRv8VcHbSNHbpXBRsW1Y0gRXbOiUrnP95yesDNnP
4LTyuDzQRQRwemvTZxNCa+/pa6x0VBHIfJLkvVKzyQZarrtGybOxAb1wlzW7uxBOV5leg9EekiX/
NdHviiOLLSgAHXnbG2zGMFQI89fVedH+rrAB/xICOFnD2jlPv/uVXNNHFyJWz+E0eVss0l/xhrtC
cxXmESicDNzpxNxAsQyMBPFqkpGzEUviUKrKc8XWQHaSE45KzTtve2htnHD6/GPRW80X3Zd7kQvC
5HupZlDckojqEYSz0hwzXciUSgV+lipIlwefZt/UdX5UlajTEzz0HgTeT6SWhPsVG/5upKJ5JJ3F
aj68bfaLKmrJaKxKgO37Xc4fBlwiRJ39yZ+Tq7Pi3JvuT4ccowok6kXHVXSuq1qx/vxTcFurQ1+2
ian4Rm+PfLkQHwCgfrNFl+loGdBFfBBvMLQH6ZVuG83zk39pWfR1B6VE759RRIrnOj/vEvE6jGzP
JsumHVZJAAeahj8Wi4DWT1scpLqtjtzcOqF3xO265QxQdSckrFykxQ3mlbEoSYVoRID1VAFPoO88
HB2amSm3/NLcYxG0tgOAr16wSibMU7vM+sh2EwM3FEBZZ0ACJhTaQB9OHHzCoM+f22ZPFJEB/xHw
eDafwDrUK+IbKdy4r3RuTcDBP8WcA7a3A81gHlfPS0I0GZ+l7UbFoNHwldrs9HNcbOZhsp8Ekvgk
TIFRDRSh4wMry2i2OTssZUmRHcKLyRHkOn+aSBqT+EckJBCXiTsKiTATCkaBYW9x2EbHNHH+6TJJ
IljIkdzNNB+8plfDNNmupLsbzSPaLnYRsl+3z1PRDkCEWUWsMOx17yy9+NtZl4LY2mJQeOLHaP9o
IaAA+H8Z1wgkNbi+QVwz16FnDBmN+1F+SeJuIaT0uKnjfQEygnjCvA/GxklXTkGHxitsKfce6BKt
TAWMoTIGqL2Hk9VPD69cDKcLXG9qtzPjM184nIc/LxKeH5ddm9kKJ77NsIFcj0b33VvYKNBqCay8
Ny1UjLqCVSZBLjKmgzGfvnLJuHIZjgnYVXUR2tyL0LxXPcs7KySJz0iNgWm6Y4GKUMkSMUz/SSiy
ZQ+wf+KmKZbaqW9yY0yk/IbtbaJKQnBQy1Q8MuyQ/zB8eKzWDANcTHKHHjg1zIap3cSs6FvR33bF
N7pBjRbYP0if3XsiWzeihXubow5g+97r3EGnyKBJl7k6PBUCvmMLDacAsw+U42v7HBOgrJqbKOma
5rI9otfDw+gP+ve3Pwn/B7hVHrW8AWE6JEP0Ahh8ddePZNi1IZJPj4wF0oTUkLWGTXHsC3yLleuD
n/qQwwOMSyGREgVhg4dnxpn+e3Ea6B0GPcwhP7c1gckw9t/fh094gKCZnMd98MDVtmRjoso7yqBf
BsJUYKmz5JSHWzofoogwiwuIyUSWpqk+yPogPF/ADdmbfE1qiKZ7+lTdI3iEBTMf7zkUD6CBK9Sj
+Cpqc4iGRtXT0Xvi7nkggr1Ep0E4PxLd1jK47Bm/BV6ezNJ/hnJqrt9vedDNncscr2iyvSyTxGuj
nYv3HgO+s2/inUTu0mhFPaaWO6d6dn7qG59F0W8IGgB8pC299b5R1cIzZQlg4Eu0T6Xd6eUrZr1a
4BYtQPYMsBtP6SAoCh+92BtVhbCnuv2EiG/8IvNK3t89wPxhCecb8kpY5hFDuHpOFmBGWn8KeVcq
O/0p9p5zhN6IWVMq1X/W//FecnYRpPcCP4JY8GNfvvg59XdZI4PMTKb+2X/niggyvbV63Oh0FceB
JZCi6IAywqjHMjrLBCA5/kGXiUpEnybKEAXYXVnsAFXz1d059q4j78/KrtMz+rmyEwO5T8UmDiEc
sV5ZItLGFcriccQTEp+FzaB7hNKl8FXhCHdJTj/w7G2lF3YO/vutSU9FoW/ITt2SaXEL9mA4Xror
Gdz0BABH30QDcePhCnadr1YaipnYzhO6xXbFT7lut2qS20navZzGt2rB0IpLAijj/S8gmZZbU83u
pvrDPNFw4Lyvi4xHaBbqGRE5MHytOYJn/suYteRHFSfltKFMCWhfNi78O6/VHR/PlSt0o8GbnbFa
Nxu+2bR/rfLXmnqfRNhXaN2qk0Ri4RyJzP2F4x1T2Rmems8ScGjkaTIxLWUN7Uvs8jmoQ9tgMeIL
M+k29nH3aa4wUbH1qcvDc9jzzoK1/OGKuaRhEUn02PSKQb0mrh1IAyAvu07bLlE71/LJfEoxCl6X
dYkCHmhGwCY43lCeP/qrjH65WMLXOmNtR92DLjL3466SCUKFqw/4lpd95MXh24MqchB2oy58FJ9V
AnG2H19WFIoIP3y62IyA9FoWITvVAt/kAxAxhMl0oy38A6a0dHEQUApwtq5C8Q5nSTfHqPc+0dXl
/CNLkXTmCXHm6spXob+sn6luV6E2bVakPP8Dp026Q6HlGL5vPDq5Nwszr38sjGl2cHfxW3RclBjj
7UR01I5MOUW1a/Nmx4MSyAZai11L7jE8fobcXltz560bvpF2X1g9Y0TSWwEPqfTqXDHATpRRlnC/
bsrLq8enugX8avsOxSxuP/iCpUkciFJ5CFNUKohEVRa9ihuxE65TV4HGh2X/E9mzLVcA7YLGE52d
fk1tMmX/DN6CeTJDY8791b3nW2zhwzOfoMXo2ZukFt5vXkYgjVwuSGldmM6UwLxzD2k9PSlOPcoA
93Mlyimuod665zxGdbj/PBKxoP64YrG7xb6E0ueyPITMu8SB4nT1eNw/0K3VjGAvDdYoYaMl1bOx
mjWp6RUjloiZ0WbZ64Npqo/z7EFY+sS5/wo8LQuaQ3qmvzzUjsonxqxGOBVZySpZ7NGqHKpw6Lp3
l3yGlRdyAOhuWkkcHc04OaOpEEY+isR5BbFfFpThGc0NUasKA53kG/w/l53FpG+A2jj0LU3J0X8e
JH9y0Y4l8ohFpteqzy0h/l+7Edft5cP65CYe0vN77KRPSeS/GcjPPOgpPn3febIS+pUVsUITpFNe
ulGevo7eDYrgocYNLJtiwb2UwzgaIO3vlFpAumkTVf9c09ua7SfBvnsAVYV/tZ97MFgbDnOxwrdH
XdEUjnk3UIp6SjoqLlvwTfXKqR1YFTK9JRq3SEvH2wCvdnMscUO4GAWG4kLSeXRz7DON3DOuwfMh
Ysls+aMg1vE/O7sMaHkglaVldzKbLYEeQtnjO0HD3U1CP2LZUwVmx7SDo9cKHRKtBjV3hq2PAVpS
TJREhlE5WW9Z3hvas5QzElJc4TtqZDVIZIxsTWzVAtTees+hDX4f4jqA6VoBmKwVsRfxHpnkkoUn
iaUQBwf18eRFl2zVztdmXR5v5c5jL4XqDzzskfQG9uSYBlqE1yVYfDdpdOoqf+1ecXrtqOl+Ra1E
G64E3CDgIPTVqhGtT3Z3LwOvbj6AjVYIgLU+u8VXVG5hgq2187ITLi7SaXYCdjxFdGkoH79jub6V
wkyk4OcIsU1QBRm+WeERr/6DYUeSIZghJ0tHtaA+4BQd5AZwSG3mRsF45Z0uubm8xfZZK3nFh9In
oDKXNPFREJO9fmzLKYbUSGRw4vK15uKniFzgDcdVw0NN/D+bsoeLPLvDQJZzImUIbbs7YU6+kVPy
EfkWzyJmmOHgcL7bagwGptdup8SReBhqTPxjirs6YBfAl3K7jUil+hCzGZ8X7033YY+GKBq+eIMy
7fvKi0syFwh2mQzwkkOvBWdjtHut+harOXEYEItmMyRILTfye8LPK91Mnn42/plfSCSdrXqUa4Ky
g0BDbVrlV53Wu/QSbqyNIUgNIVraQdwpx1IxoBC3EB0K+t1LqDsbqSp5coXqXooS8b9lAxReEISn
czw/ZlvkkO4Z5zHdTPRQyOO77b/S4aGgiRVgLV3qjB8UoX94hSmg7RG/UP6KFAiQdBIp+DBlOYk9
GfSmcPpobv+P0oojQo8T2w0GbCSW/4DsA9WkgVb4L5EloI26fd5ePLTRz1K6tE/TUEre1ttwlZY9
vM0b38hnW7c4t2dIy58zwU6GmlrCAHRi3rO6+hrF+yTxEAEycxsokQ8K42KRbIxjxYomOFAJWIQj
KkxBjKDX+KXLFUqNKQ1L4dycZvizhs3uFKQW9NXApu2G6V5et3qNT2E7j1Pg0APjeWsPqi6YEty6
reQbvFILhGn0KTDtiEE8YJd0z6B3cmaQpR+amiuKYhz10depe2d6O5k4QyG5wSNa2stuzqW15nay
e2G/MLLhuurQG7EMvFGMv6o+9VspvINXB0J8Vp2GVMnH1ebSLsN9jwd8q6l/B/EcTTqjPbS8OD7T
G85wjzkM1IRAhivWslfqnD0ZwWN6XVvQ+3hfVzgk8khNWmSVzYv3m/oLMB5WTpq3Tsf7bOqU2oEq
PpoD/EgoPOY+VmI/x0cFHctDaUuTbJq/w5Ll1l6+FpzRn3WABaWbsnkkyKT7g0YLVfRP/X2UopyW
QGUAOwb08IztKdP/1SSR4SWB4E/giMiuButbaVaKVictaEjTge9Nts3oNcXJOb9uKK1yiIMXUrcR
MKlqx4SHaHMZW04c/38ZtkAHqMeKeabBxfyBwyUkPdYTPECIkb6KYu9vryk4gs//JfSU6D8N5HY4
AX5fJcHmXXIHYpm3oJ69ENYzzJBGMXzIrvUC925gCwiEM0mLELvZvwPTviMAt597tjtnG3ArKDwj
y9MDJ1HMQsE3RIN9d0jn2JDnI7SREjChPM4Dspday+68Gpndji6xpFXmquv1dxr8p5uPxYtbGXfR
15OaOAydpu/Rz5SAv6c+hFGE6B5ulPRXBQ1onIrOkGaMJk668+vWuO2xpAJwddTibUYSAIjAh5d4
3ekQNxrhdU3kQ1wnjPzv6jWv6in4MMIzAOsvxgwhkrJ17CpAsSFGBjco8uRIU0TnHEGY6ytzgeFr
eIvgR6BaJgRZjY+gkc74zPt+8BDZqpphn2WXxx2ZzZjFE84Q9Kn/IO3Xf4jXIJffUwcAF1ftsSlb
r5P/ifLqc7Lbn1pIDCJTo11J+mcOvuThicp841xFgDUCcCj8sg3Wj1WsWflApDc4EUvNIxkqgeJ7
AaPlY7B+EIcjIeJAY9dFFgzc0+ZkPQqXn9EcrgiXoWpUdNVMnj99lSRfY5xClQdL++rqn72oQkAp
Rzh9Bee3gQuRAyYOzY7T3J1Lg/P36a2OP0zS6z/265Vk9hzWSovv7Zx5BXEz7vJpwIl00QRpk5YP
Nsrtigbu/Njn9NPbkQVxF8dbbZGXFGej9heEKYtBXRhqlIdY1M9VZfSV+5EAcsYUd11IKYeECfQC
GA1uyQl2HVUPTtjph5oZriA5mop2sE3ng+auIgT22h62r6IpWgu79d6UIwGjADgbUwj9sZhtGWvu
LVthLNwN5eww/1VmiatpOCJfeh6oWvvnGoaVSrcXT8sSF7MNFruqKKwCAJBUd67bM5EzVzj/Drlq
17zdj/RXh5pIiHg4Mg0uG2elOOEJ3LmisY2oRi4sKUUqnOzMqfcSfsOXqxrwjmmm0izgPURsBxhB
gFAgcqT6XZqQduhlxbTd1wSHxmam8CA6ME87VehZ07rgBKLnPi6HhLbr/K86vcoU25oex5wTkLps
kkM1e4TTq8xGIew6CYLW3eQKmUequSnhUxQb0si+ugKy6K/vTYDo/SutUIoQPSB/iCA7IDYidmrN
ypWKCHyFywdoZQXBnSQUGrfWSvJgiymi7Oux496MafD3wkpgKMCLaIo7Td04a4q6OYqo0obhRWl3
RJRgHLW2EMibsrZD4IF6MeGB2AqooA0CEgOidbr1QDIxLHMI8WxzX8Y7oHn14QJUbCiBPuWNneOA
Looz8LWklQt1eHWN3ct9bd46Bz04YTjGNtOgED3DCXufITOJyUS4/VwdMC1CMdK5XLyr+NfT0q+Q
BXTRmnT4ctoZsJIkgfE1YG6fRDCHfSEAOF0rH31RZ3NFuMmF/ykgSyTdXln6qP2xVwdIzxQhUr/d
y6lGHnQTXJDTpSX8wdNE6QFo598ji37sNCmWXo+FfgmR17MsUevoCvsDRFNPsaDz6P3Kbq2j4+md
NOO2MC0q0YYPFkrL0ft7l35xy7+HGim1W5M4IgCBZEDIKrqmzUh+z6JeVighNU197kLKht/sKfac
HvhoD2tO2KpBhtmhn5poo1UIyT2kb3xlYtHHtItE5KhYV0yUEQIM2ILSV6h26phRHJ4KAQZ+Ng/1
CUZTmTs0BL4lvNJz0FYNCXoAAPdiOltDPo5Oojcd/tueJAWr/G/qlIGuIUphEC0zCWwfPJOK03ej
j0zknCrwCynOfsyO+DhvpzTSzDQZJP70Dq3t6cUFOdHbKs2oSP4KjbJcM5Wfok8lHx+9l7YcBu5I
Y/kqcfOHcs9YxyUfJgPrE0Mo5VziMC459j43BfeUJZO00wF+wL++gmJmiAkhodqjVrGcqrORhINZ
A3EfYHWNoWtp2ny/CWKCUoisli3ZDQbztvbz329QvUFFs6LDVdeGgUOyvnHpmAYss8GeIOwE/2+O
08MG6OIbl3DdxMwsB13GpiK/ubuNM2Fac7xLlNGD0A5aaINDHZ9kCSxbjg80mbxICURZDMvFhKwF
h6llThq40a2GOmtg2qKGsErv2xcaXDAdoMo8Jfalv+oZrrcMSZV+Y6bbo6mOS4HUOvawIK+foALO
ubxx/09t5F9+5Q45gl5kOURO7ChFi0cWl08DDxn1/kKOuRO0Ro3YA2wrxBy2UDS//2VROwnpTcQZ
uMOIKWNzejNXyUayn7yQ5IV6rFm99G3iKwRe6h8DMYdZtKh+JVT6Nm1pfHsHb2zHlnXIf07sIMGj
a8MGqWjJPHGEjnozChdsHbY1sa4ItmY8u4/1/jkz6ASBUaPYEopydZcIUt7q6GPMc5hoji4T4c6s
c71NeUnSALEOjZM2AhEs8hlWJeL5S87W3vM8NmnfaTvymaHtFTRJtF0JFR0suwV8bp4928dxWBZc
Zbutf9gaQv9wtTn1VeUEFgi4z8aoRRmtdG3jcRlQ4Oy/UuYnrGtFLxvUpf0V2HPEtggMXQXsOBNK
e3AGrmklA78CgkwcKAzkFUK0+NLtrOT3t2lpTxr85IdOTd9bZle0RlYlP3H6CrznFKqD3J35LP1V
zsDj8tJknqtqdy+kqzHoUdAldaHPxsbSCjBfbUUHwizTdaolGMfr+p+HCvAwt8ta7agD+kcCx56S
UfSMs11j7rnKlLKj0lFaSgnmXXqOvuZX28ocJOZLTwH7roJ9I/fQOrNhsWpi5zdh6OdkY3nqNz/m
HRV+myyRLWzjcZm96Dk2qqIu+qWJy0m6Tbz4Vbwlb/S8XdYIOIPKEaMtyJXwCEnvLuOdwmeebMEL
92eYLn6W02MGW2yP8JZMUihJlLTc2pzeee4HYyim9iolM7mkJKnR18Y8Ao58qz3i3wejYNGChvAv
fEpttMWIaayrFmsZnYjDXF+I1z/KLUz10wLdzrVGXgKD/MecxbS5bi1VtFUoYMfrPMbZa8rDZWau
puK/yygH99XgQcFNbyOwEeGVnZILxOd1l35wFJGX/fxGcpgJQJubwkgynJnSzuPj8nKCYyb7yVhU
dzNTt2gXXUBEtktpqrC9ybzuyJpS9I6w8zsXLLdMrMLIZWbHFETNedUllMFLCVHsXbhSVu0O07a1
Q435n949erKhoQZ977q5vZwo/9EUdZse0UG5sMm3AJCpWWFA8paNM8eKIlV7+HHB5QP8uQSp/KhG
MT4+6ibNXX20RCPhdniGCs6GndZmE4isSY3yeXjcYfP7Re6M2pRHhsw1Y/7V4KwcLJuqcXUK0e77
+mwaY4H8hVh2SLsVfwCDeVEe8/Ne1TwLUsoHaB0Ja4Nwo307n0YWA5R31umi9Kap4ZI/UYKcgQbJ
22+tQgJKa6UZNrLjJAIronVGhB0iZx75HcvyKcpaUO7TkpZlrML6zMjjmeGSS8c1zgSmwG3MzM1u
fSivdwenNXPh6p3GPMt9RVrVNiVHzcBCBT1AGdC2PT1NFYFgcF/LSGugYaAIJidFdNb75Ke0XsSp
OhERfHHdSgG5OGvQiEcosdEtduKnso10F1HN+MHwI22AhPYCbdKVwgi5NxTaydrMt1KdDrjB4dse
Bu9LHee/LbluRYdGGner6DewO9U79iJXa1lOYVgpV52skka5r9vsAu7YEul3B81YSnRLBAi3qyfg
AB5Aj+531hvxk4y4wx9MBQE/1ff36q8+gLqEgKZlaO166AbXTvyVgQ3i4/l5IWiDimoyD0tM11N2
HZphziie5wwbE3bdAKrZntnRj2WJevN6fj/bMOLim06QD5RreyBckGnySJa710ViXtvSb1keAiio
cEFrAERSY4WP+e8aWsed+Sb3uTlfw34dJFnXkZQ/9REhwx6B7Hb/HSiNW4yhBdJUX8GdeJak/uzq
KNkAfTICj7iF1f9yjwYLTiPdYrsaS321oY87oUhx4vnsHZF8tVDILkwe+wy2rP3O5VpRfVvPsZa4
xwcnodf/a+jyVD5b7RB1bIBaXngnRPfjnHxWXVMS9IismEYGvrvPce1TjxAjBIV/RLaRPmg539rB
14RgTke7fOdb5txf9PpUx9mjwIRASXZaNG+k8tJRg7P/RdoodylEOREdb/oiDIrDgYi8CxULyALL
XP2gwEm3OufaVoV2iRrrcxaZmBcDYyorbNrWYx1hZob3temWSmqgAk7lMUR4Mk6F9rHL2AzqFV7O
q+wxdGMCotHBtsoSpGLpJHtkrWDEcdSjvmPjJnOyH49YM343vLOO5HxKYZ3A38HmMLUe3mnPIoC5
kJd2yGojBF55Q24yCU0d6VfiF7B5bqa/aOM59FOuvIWaiBbP4Frav0QTRnfVscY0LLe9NHC53URq
jHy+k6011VRBNMud0J/QdoZeMsuJSBDCjJH1zZGGgJmQkROQYc+DWnXbPtYaeT1hgopwUcAHJnKf
jDii1bkBSWF5u5FamVUJveCJARa547pMB7HcS/MDsUkF6Y6vAQ6K/nPs44kUENBIw1ERBpsn/7yK
xgaROpHGi8SRSaxqcCjFaRYRiZ0bmUtN47lHd3KzTlYKHWzOhTjmSGuR9LWQnb/m9Ykx9QfXpZuU
Mq5og3EItlvNFKBlEGd1UG3azA4bz75SkyTXKzWjAHJSSaqhUFM8krFo4m5ZL0753Q9gWKPQGYBY
MDuSQO7E93wnYnU2KHCc0vlN9SKlIQNmjj3wpSDPAmmhVz4Pf8b1wTa973VabTYfKw89XopzjaJu
78j43lUGBgXa2AU1cWUC7qJsCR9MKBt5totRdoGzhtZV/i8VPj97zPqNHaVNKjaLZvuqjYFJppZ2
6wKXAqpyt1WQOjPEqIcVlpLChG1gV5cQWQ11t3JZOXNyVGLAjuiaaL0ru94ciPIGT1gnORD8wfRW
zyQR7OpswTx88YVn8dYutgDNyYUoqmKybTtTj6HvfJ2U7Ih7poHaTEwvYYhwk2b84GWJHVMHJNp6
Yp3RUcQwTsD5C2wiZ2HVWtE9tGTPqbs+HEZavEo0M7F+LoedPhMaw1/73LPSxRncj+R1mydHNHqN
VmgpbFeI0d4LxAE2MkocuWF4ecWrE1pSU66HiLGxOtLWHosD9sLreZoeky42cek7Jb8dYuTexSUy
6S+2QILlu4w2ULx0AJQsD3+MKawA2HzomxPkkmBeX3Jix4MOCB7nLK+xGfuEUp+b1V81ETrilQta
PNSFldJkRzxokI5/OoZCnP/o7eU8IpvRqFA6tfKEE5gnszuVm2kNj1pQJct9XpohCAFllRthmDdA
sNZ7B7I+I9juC8AfIkf/DaL8M6aeYjxKhgotX0Zp6WJHGeZzdRtGMZox56jYLTVU/yaab/HUpvvm
MngxK6Rt/SF+bBTZk1kG7OwKvUQ2KVm3mmorNQTWQ2wg/h4QT7Gle6ACQf01Y4+drniaMgoiu4U8
HlGF8WLOuFT8xCGCbXY28I0dglnkx0OLz5OostqX1FQOzCdw9QMBmflDWgUx+iUrnLho3IbntgT3
JGlWhsCJTvXIVTXzjY9jBRzbDCmdmSb+ejXjd5oQBuLDyiiwJ3NV4/BQWSDeJzpZUG6J0fyXy110
c4cQRA+OfEtpRa1qgXAQtWeFSbhKx43cbDPlwSa5Xgt71IMVpxBKd/+GNKuk1TJixos5zv/scM/V
3N7W0XNKdFnO6/CZeH5ZaAomGB8SAVnTuUYaL25e58LFNi+eIb7yeLdjbadsav4nnLHnvLCfiwdd
N07E12wjgSZcVoz+Mv3l0rEYE8CCdFKWrp8LEbip+wxR85PgCz2x8WKPGVbcJvtoOjD1rDNomyOi
EhCvoCD+Z9NU3fpuk98rZ4zOkX5q1nT747/EyivqFZpRgiQBCcQKlb1vtHWhQAa+2UcdEfH8Lv7a
axDzFFcfnuMP5Ax4yFdk5nb7I+jBsTfqM8lsIwGne2XfIlEL05joSJiWt7ejDeXm+HmBsLmFMrmj
9c3rzMrxdGlx1eW9BO2bHEla4M9CFU/30Ax6js8JNqBtInP7LFfBtj0q+vrcvK9s1Rz9Cn5XdDI8
pm7F86a0TzdsH4MwmJ9cv7kb0EK98jV3TIJUTpBkV1L00JlWtpRLoeYwMAQzoEATtvP8u3FgxUAH
rdFVSGgS+o+FdKT+Bj4hCKVxpqnySlrf8SlENOQLpfFmIo8kuF4/WcM/i3C+qKQnmvPuLhZ3uksq
/D19AZ5mvLFSkZnIyrpunBe5+HNEvE5l+kiFO1BGqG7b0ebqFCZgbc6tAlOfCHNbzS9pVVG0mrG5
bkpIoJU138WTcvVXMYFM1Nlsb1YkuaIIJSulbYaMO+BHupPCiF8uZKtHo/E6wWT3sMGsfcLJ9POb
wBMhMuKV8zahliMbmhCgJvZxNfoSMhRma/1boNC8kfyqQr2ljTtG/CMn7bdLYBqERmqh5D2SZ+ov
yCg89de+AUOo1+kgqoSAOB1BoiJvlYo3CbiBSzw9Y9v5XjhBww6gLX3g9jaETNR4Qnzd4kvJdKTT
EdgLR4XDqxzg57Q7jfZGKzt8AV91g5x3T44hMERHJo8GQ34sFP8wsdvVHctTd0KdPcO+WuIp5aPU
Gw2a4LMhdaJb8XRog0iJQu/85MgCIeBFoEkVCGxymELsVSriYp55L3VpYepIe0cBlUYspJ/wAI8P
N+Of7hwHoXeAi3h1iO9aTcTfUPt5EEQ6vnLgnRInlBVUttYzv8gjJ8N4LriFmkNOKc5342reV4kA
T+F7SGbRY+tn6UgpgAH4Q/m/BoXi9g8kBoJUJBDQ7V2Y9I2SXG0o9BZjQRbR7goKE3NOE12qHHGR
zyMj5SxZ0ERPr6z+YPSkvNWOvE7GVvkL87Ycqp5qHHWYDyEv/Ki07D8ymzoYvqiIAKhHn2VyANbU
Br9TNBSIFRgvaTRU+VWfO+tdrHQpwdzKXyfX44D4kuW8hN4RWDiDzRf5Pl6vrG5xY/OJQm0lbjW2
M7IwCk42EFis4ASISnSGSQ5lvkCEEY2OsG0bC0zz3HfdMick+WIo/gitrevbFrLlyTch1crw+H4O
+wxHrIctuj2F9ejMlL880azeFJ5t63huutOEkZxuPM8baGo3WwL3PMYLpY/Mj/FALgwEAEhUqW0b
J0BSJlUBNsnXS6iI+Y3Hdw0s84Afr0hybOAGezY0/IfSF/IClg2iRMSpb7NLoa9007YPbCDeCRSy
f/WdvgaEw7Jx5Wbh1ScmYMlrtc+t2LUUijYf75Gzmf1AvVmPMRd92esbAtcyiMWNXtxzsI3VmKA6
yC1pUqYV1vfVSxhjw6N9xHW/i8kskqDDy5SHB9mv8HUmx9ymPsycVz2TaAsnL9cGKcmJPeJt2bBq
2sJyo2VwBjUvSmC94hkOimzf8VgGgUQHUYuf4FlWMLQEinJvFwr2C1Z3FItPzjiIGFRwAyGY1oaG
uEkhkwUbsneSkiTeQrHnfDOyEuK8CLN9l2Li5td+0GWsFBktqYv62gPIrcQUvHZZTfz3RSDzqu94
PkelYt3flf9fGDLFGHI0+g8TvBCO4OVUdoehNyl79iGjZD1RPyw0GMUpDk+HdySiAsgy1KUdfVKE
2V3xwbSt/iuMLdkkIgYcvtKZWRLWRhuEJIdj2nu1nV+u7cohCDptssoa8rcgyMxz5SjlfTvXHoNa
03x6XR5+li9CyMSn6+yg7SJC9GIdHifEqIs9I2TaLzmLgRIfr9AYv7wLZXzm6srxS+dR2jNXezUM
hPzRmNop5ux1fQWJDZ9hxjI9QaKzCyyemIbQYaTG3veHOx4kP24DraSzJsCpj0nzdy3aVJ+pzRp+
v/CjjMKrrPSBoBBwsQ9DrQDOrIdmdjWDwcPibet0wdPkB0YozpD/7cYUJyo1jdVvmx9/4E3WIGCq
WphD22GjUYD9LbzkQDEnt4P3I0Jevy8pVCnl5xSYEdd0rjJNL9BcYV93UObrBSCf4SNLJ4L3eoUe
D0uDuuDohvAC7eoROTQmRZ5KGZjYodTZyaIpihOOrHqd01dhTbzI+d1Zw7VdOGjGZHGLlVhW4STz
CSBWFgbySCk1CCBwizZIHExBH1NbzYHW0Ux6R3fjRrhdhP8MtRJ5oh8KfYetQLqrwulM4iG311d3
16I82nr2aPu1dxxqHe6tP9/P0om+6H3Td2oEAbsqZ6wr1q/+5y0rFsn4YOrBgCnDbGByBZ8tl2BT
aII+ZnB6un2jxq8kAh/Dd8lTYl2z8tYbKWv917CZK/7MsY8X3u6kjsgn9iA1j0MOxb27oFVwexSp
+diXajUfnMATXtPH9k2rQwNS/tI+RjaRugbsN2tlP2JJnBRaQy3RI3nrMG+p4ctU0k7PlD4uphtm
2sf7VRxmh1X2ilS3G3hyybBWWpvrZXDb5uYvsRyIsilIr2KbkROjKjuxWXL/8QZhOVifqUkOxy9s
o6Fy0jit1gxeZM3BTiyndIhzySWK1g29K4qe72Ktf/1ZO2miA3jvYlHBTZKPEGgpE+c+9pFBxKgA
Thcducc1DIVgpIKpuGzvOOBQljl78tCPv3khhGVU+1CGoimctOIa5rZ0z1BZ+MkUGAwjqcLxUqFb
HlWLjlMw5W5VUPJADUt52iTfSPfGY/QwaH6jTjvWcizcfAbwxtfZLk9ab2bVeQ6NJUf3J1OLkpLd
YQ969YUuPRLWxesLtgMaEYZcME+Y/v9UEsRoZQ2XbMRFys8JM3Y67NQw7vRM7xuv7HIGX1as1RIh
MMjiINhfMJz1mDfOi/e9ZMFjQTcFUesgRAK1HIat5eLHTaEPHKZE5E+QeURfi7dMBudc556WVzP5
iNyfIW3+pSgCi++6NCju2FIZu3KWvxQdeiYe0YM1FhNmC20BdQvM2eH6Zhg29hr9CTlmJstJ8LRW
HWKbBl8JXGEHGtCi+usGpRL9lKEzrmLQ9Ro6+h1mSEFj99pk7jcmDrn+clBRxlC9tz3yh1bnJ3/T
70Y61fYUUbUsVuZk3YCa3Bl94n/w6j7ZocAlyiiNEwvDL/oePlsBKgmMuQ7cGNizUEDYJvDMBLWd
OX/C8S5N61SoTDrkvziw2efbZ3/YVr/U6JqSD6qEf1YQGNIHP+JdM2VnADGvbam2WIebLLZiuybv
zGG+NnHgC0k7MC8ea8Zugjt6oQOkt6SNivKmFR4Ry49icmxAF/EGa71qZXABtSmpi2VR/uBfFJuz
lhLHADq2rYNAV3oMFVhOWAfePF8pBBRoMuVcc15JCizq4MkPAKrSoCJ+atV4ZcnOSG39QopDej7J
KCjxaFyOns/Jne6l4iR432FKokI5HluxRb3lkWg59UFzE2Es40Rkacztfkkr3bznNXDahpyn4avw
sVWVeAWxbBk8aHrZCZgVT5hZb95bAwTrDKTi0OSXv+ib70UGWITdhd5/3ADcPpbFNjx9ZANvfIbC
SwiZvGyFnyg1TP43pw2yxJdFSqiY674UALgIhsywj8IeHc/Tl0MsvFbaUine3BwXd2+5+ea8xqn7
aW+XyflVgm2rXLUuaYrZ6UJfCpN1nbGeS+OdYaYuF2scKJaSkglnOn4AYCT8zPht5fqkKSbW6YKS
D+IMzj2Rlq+lP85DAiLXXkY8Mw6H8wkFlgY3g9Yh9XmaD6LHTNUBGwxiXXsk2aWM3F6r3ITAOhwx
YCRoM2VhzUGbReVX8qPCCxM9KF7hr3fPvsiNh5INaNcOFz65Txdp6L8TZGQXNYOibXuQjVIHE6tf
78cXzGZpcG3laR+E8VLVEvSowQiYHF+4OOoZYTeX9/AbYg7kElnd3ykgRV/mFhz7UZkMX0dyJdmB
TZL8eqLpfckD6X7gbXHkpTXKLJdRspkOM+KKMeHgRfyrtnTiRMKI+nq0qT/GT2eauDc9Ls8OLHBX
tCo3RN8iXVZM0pQJnxDAhhv7McUiLd2epwyFcOHLfQC+qWBIPUHat+SkR9iwP4H11Q9Gey4v/JMn
qwdrJ1rhSnTnTIpOrTbCZGsaUfvqjXvp38TZH522FD09vrx/u9nCUlsqxJAjxJQB548UTxelRFX6
1D2mzLNMRf/MunSplAuTjdmmVaKf7Xlpn9WrkTZnjVHQox2FYQjBHvMhmapsLEsNDjerFxxvEwSy
3T1vZIyzczkz/sbBj3+Xm9CW3mt1bKryIwjaVNhOyjLiD7gcSbMR/07txYmS75y0G2fGtMa3WVDG
7ff0FcHD8ivz7UfP/Uph3HLEDOvMTEtJ+DRpzVoCw2jFoEVxZjzO9TtV/CvH/YH4j3FTFjcbf+76
cXLpagUIvJxjr0vfz/9p1xgd5IAsSMCEsvrXr+YoG5CDcpQxbiLbnAh0L6BNTTzhiwyDZwK47G8C
VsHbJFKLiVRvaVfrjFQk9EEeGdGv/zbFssK+tG6JdCHWqj6OHmNUY5FUAbNbhOM/dWwsw2SnlfTw
O0eRuzcOBV9VTxq510grn4ch/C5jrXj7E0bKsg2ioP3fWJma16eeHIDUpYQaQwnyWsPEFKiR2aEt
UCg2xKEZXQLXnXUVuQZix9j85o/SHam5+aCdwy6uK/9HrkOsqcODshTz1hhASbpEyOXpe2okYFtE
pl3NdTO1gjl4o/AphbhdC+qr8IyQGVIfUsUXqmLCNRilfXWKjqpOZGyzwP7K8ZvZvsmgxQwebkSG
I3zOXDD4+j0XJH446toArL+Tq3OTUTxtRUaKChWUmrs0+7OfhyWnLnX6Vtp4AddE51C/ANao2LcU
tPqXIzng6wy5mZ5l5/zpTXWPa+42AjP6BNo4ZCu7GgBMGqheTDxo9ImYjvRZZuiAe3Xam2JZYnth
KdY1PImZZ+0tMv4aw9aw6ScZxNXPOJWQnTmJOevWn76uMr/05gpN8RfbH4PAv/xQYq9e4lRJFgPs
c+sfYckTHh03pc4JFjHLxhOwmL2Gom0PKOJpBWl87/XU4TG34FbUpnv4m+6IYLfQTRF2jaOpC7Ah
7SN5b4w6e29RjoyCmiDTF/cpee4Lw86UU7weKfvur4TURZ2DrYJ9af3lZKNm6AZX8z+5DdlFkn2r
w6UL+MwxfK3lS25E5soHM4Qa0xBefr9oSQxO+MD61OscgGzFk8D1HixSsddIL+W/s3yls22kNmdb
TKWjgkoizBgvZrDx71UkGPtQJE0hrrnNUOZhguQzQhZ4asDljYU6CnXdNAUUfQnmDhoBHPDAwmRF
W7ddBDQKXuMYv5IYrND85MgtH57DlWcVorB8XiMIj76yOQ6ig8o/1BvtlO9jWNmamkg8d2k7gy+Q
54p6He5Yf/trHz79hSx2cif6IlcHdnS7w4VSlbSjGQKvTD3vhpXkD00u2iJEhT2bLDN5/USllnVV
eEyfkVM2ZEhD9ysnS/PYUP3+/MFMoiY2MexVBNo4r8NRkPb5jJch8dk3S8M5ovWEPkBxPjAf/Gyx
3ZG53A2/6H40FNNe9QFmTwtPgCw8Za7tpQJkhbNQ6tWDMZuB827VH4yEYuCZ/1laUCbU5t7cP/v8
XxS9xSwYw84++r9fvw81wI1Lq53lOfu6ZJhGP4h8qrNkzL170NQAGQrgTrm6RgPBxKrFcWLbKKet
YJKirw/vqaxfFRzAlETnbYsK37zMdTlZo9oF0ugRpsHAoss8XbGThxlGs97X+RBVsXc8k9P4/DHW
nXe5e1MuzmnKxQaV/+hoHtVEmUy/uo286oUTrO0ElyQ+Eqm6cDxeQyoKYVG6zM8309K8Jt5zIGvu
z7KNUr1Psj04AABTSzqGX3qL12go39OrJ4sA3VpnnEa7zgz7QwnFk7nhdadV34lhCEt2V9I2pLO3
LwgATRm3uR95aYAN7ZdXhob2T70q0akEI18myixpxqYFZ66kRI89wLlA7Uc21QpWXv2t/6vuPek+
34jophUrsXjeEwI67w75AK4cdbbNMsSEmrRI/BDNiZxZBafL0cpwj3XsQc+po9uec+VyRwbef9zv
zaJ/UB2C4SDpAufRX4LO7eQG9wwnFW16Dd+4rJIEW2ZGaVmLruamYAXuppAbWHPucbo3V5Y3cC+z
BmnYC9Vn4CeNLmkN8ztxioaWx+SP9k6gRo/IYyumeGb5guMBj7ugoI2BVNmEA/ot+br4fZVseJMG
wSAMmihdiIg4ui8g9n0F4XPffAEQiYRGRx/dHxSK1fsJWimLEF9PaQS1isGXus2YUIPemV668tfg
n3FY7g4CSHHXS8igXpySC/+vUcPptGo7W76freaF0lLLWDoQgQRdQkg7VNfRanmBH4LqMwDtnzd5
rZ9nGEqXjA5BvF9BgzWTQtFlOHpQca7kTbXsXvFBf9fIxYw+/89gqLmnSrLCu5FOaw2+TA24oVfC
4jIT8s4ttsIeRXb6lKCE1RXZnlx93JjZpe/azkhv81Rotixl3hRjwUz4T8Ttw5L+6sMV9gbPJgR8
3rH0PgbZc55T2CiY22ZiiKJT5gE9yQQYxava4lD5ipQbpiJkEL7vVP4/IGXTZmHslEcJjb1slFQd
1yEKy7ZKXe+u4JCt3ldy0IpAm0x/Wzh2vpJPCtZjRpEivwa0YxIPeoIZquf0y6WRex33iIu8msoP
1MVNfDtnp4DrfGaQdExt2OABtYoTA62zd0hYBLst88tpwwpWzi0a07FAO3d4YqRKQNIVqDM/WjBC
gEWEGaPRa0kvqICtpHpcQIu9i1+4QeBpr5d+SUniIXRjrP9D6+Q9Y30IQ6alRZvA+YG3VFOeguvQ
pdZC47NTCeVK0udq3fAQP2bsSQEOBcU64LDteWSE70xIwMzmUCKu0M082cb6879rCvjwAHEHcGju
93FucUxyON49CA2607L8Lu6/YbZRtYJ27ZE+pUjQnVuWpII6QWN7XZScCVnw7JqlRspbTtf22sIf
mijPnPjZPZZCr+q6Ddrdbe0nkpZeEy+z4oDe2bEcXJyGW/6hfhGfITvGixZotHjmrW++pUl8wq5+
MV8IGJmN3MlgbawPV8h/3HsJ/DEQ07KlpW3NZB/MMuFhD+0ZG95zCEyDweCdGxn7tmN4iyYS2Khc
1ISx+r5QyljLH8vQcLA1zau4yCr3d5DiuinW/dvWVTktM3oZPSnhRo4jtmNqtH6NdowvjwxBt8Sl
+QjWfjDZXVTIC8nStE0ogCqiRhwOo8o3+NqSFUNkDChnh5ZNYeCGtHY14lcVkeljQ7sg2L0rseXT
1w5zXxnJUye4shSKiEHBh/29mUM5Bhsz5fYBKp4WKjRfuo1B0TeIcYIvprkM+Y+l7zT7Uy2L3Ggd
iuiSgIrA1EOOzHO7G6Z0+2nvlKhC8vBaopnJ7ToIhN87CSVbzgSB4lWiN+lJmRrqfh0nun1ke46d
rXOwORabo1uye7ARwzjMpl/AHdotL1w2+CddmtrZsQCEHP+tdJUInitCdzD86A1F2wY5Gk8lhNra
qpklVrUTjybxwMgFqp8WhonxCl9EQ8ZKMR2FDKz8crTntpeyzUwtWNe+fyYE6sNWSWZwf0zHHA0s
ikM5ysU8W7N86/oq+2Vmk1LYYu6VfZCwuSi3JZRNDgkK2N+th5Bqumdf02RZekq71I/46j2Fr4GV
0uq4bKNSDvyIwodS44Lhs+Z8YqK/atOE0PdsFvi8SfU2orpCcgamabUoCLWWqEyQ9kCRL/rwYoXz
8y4/3o5sMmBtJ+hj+erdkvyTAB4W6uTjUZe0bE8mICi+E0bBw1aChgG+xHv4WYx308MAIG9INfqG
74pZFbYukDFlm7UksOBcp0Egaxkryrx8skmtWGS6iDact+dId4hFQQx+q2cZkHGOc1zqeIvm4Kk6
Tbk/bJ/BpHYNSFTlsJQZB2btHTqy08/MxsWn8+quLOwv3nst6gTpXaFjoJNiyzyQ7nOgc6rPqdBo
JL9nyiVGqexLdoJn/vEgkxLFL/idHEJQ6RFEO8PSf5WXwgOx/G3f51vS4cQeyf2YYjsYLw0c906I
LWn7w/mFSP/Mi/pzul5blDDP4jl/n+yBr6Es+mxZmT4ffph6Dh5FQad0ScsnvZ0dC4HbDuImHW8+
6fJuOM1SeJiEeP/kKWw5RshpOam8jDd49PGEnX2wzrI4Wy9g2yu3zwCVOS6pQGAZ+YcP17aGXTcm
AlGIwrZsUPZdaJhcR20juvaYAZlX6yh6V4dytVCJynzxxXJTiQqyOpnIvsU8MlKfxKtYH9p2JHCB
wzI9MVpgUeZ5tlz8le6x3vqyD1TT5J0crEzr89dBr8wBYjDXGtRzFcGIEabd/LB6M/lbJoFd1pGg
0JorXfjHKlvaRd0xBJsmWyDcTPo5Df5RdT6LB6AkeloxoNYKrXkD5VAOHX2AuO/7JDSUDuyfL7ig
opSA3mIS9ffeR4T8C0FyLjmKU59YUwvh0L2z9vFDCDy/vAlXTxkeRDnxdpa5w31SGY2Td8I3mLSc
NQP4bduAJOcpMVqvGi7HQi1INzNiVmmwi9Pfpw2q+/jel5E/51sjPRuJEwma0jIzSLKyHGH7h7oN
ewcw97W71PHE1imolSsQdNdL32JjA7X0eRaLt2a7HCANdWZvILkZkG9FNqH78EAAzmSKhJpfaGy6
GEooRWTjmuldy8xLrvq7zDs7xvBCiMCp3PLEcvSxWiSaHCPL8AwTgw+gTQ61IBCTLqJk3QF9m3Wv
bP246FkJTv5S9mk/NAMo0ITuen2T+69eiBpRyl9EJDaVOaMF9Jj8npM/8eq4/Addps33Ec5mN1Mh
zsRNyZo5J0A5FhSptQ4X/g14uev5nd8ur2K/Ev7wf3ORFU3zIGlqsrTTh6iMLXVmHSMVq5a592IS
C2qbkLV6LRAVAgTRHpalNRnXkHx7nha/rU0cVry5wjM9Mb1BjtNoo7EB2gXrA9ffM535S1hC7JVJ
Ln/0vz/bZt79hY6AaAzQSMGPdx3vLqwdCprUvddgpnSfPTrwQ1taPItLz5Pr2YQQBVfSBdpZU/HX
v5cbgQg2itrzQWfC3vpFpZlncsjnvsna3o1uvAJ8TciMKCiTLISxfh4dDwbNkSDcDAy6wwGrVzmb
z7CbvZwH8KZNnmB4C2m/PBMquPo+s2VM07E6ZP2sjqxFcxAiI90EgFhhYQeyMX0F4hLQUolDBtS7
k+XT3T+8ca0gYrjcS+6IyayU6hq4xsgpysBiYD6nrYfKqP2vwpaKIn03Cd8FEFp3tWUtHDnWLkI/
wvcVY54qCVbe9/rZlepzdBxVrM9QiCXeDtL6zll6Dk7q494MhmyHTQTTuvqxGh/aQh/svjXaTC2E
TLoahtdfOTqTKdDE8RnrXbe3iUlWOkN2UtoZSeYRtFcY63xR9gm8TsmtYgUPKbmbUgG+/OmsFBBf
TtYaMUxs951C/X4DkV6K/eJkUSooiOm9YGyfHwRLjUI4C13C+mka68mxHsWYrUfsSTfRN+NS781+
eiyKZviCkE0cBiCND/cPnG4cinaEiipFUukJoobEvDol4wrhVuUDvoGLYNowog/PwGe+fiq97kJU
2nkXGTju4X4C/Rd8NKmfZhw4yU85J+Ql9qOKJOwahxbx0Tg2Am7Pxo/z4UZO7hjt7+ZEwD1srE90
CuZ2pgwJ3F2XU8v8mUbdnPsxJg1HkNC/iKRPO6kld9vQTH3PTdN6qW691qTVCt5Q77p20zza2L41
1azC/8y017uc9zhmm7tjNQuwksEwBrl6XO/spiWUMK/aXXToo3O/UbVsysFuxN4CmVu2+umOIsfJ
MxzjK2MpV4HubHc1sucdXN9CPSOshJJnXkP4eCbwuK191A7pNk8c7vMbvuJYYbsBkkJ1svUnxjRu
dzq39JcnKHfuP53Pcb7YPhYeV+szewom6CQ5Wb3nSDVKv9SpmiFpFLPpHkFJdcYB9F00zmlQLLar
SyaGQ3bt5UwSViUTDk2B6U19w8BY2hys9qFTqd0z9c3yvSrwXm9ueOjmoT2Wj+K9YtR/HIYjLvvq
gaV++eOSeuuFu52Wd3mB1os26nmUi2Ztyh/1KeW5PM9miWgfRDWFp5LtnJVfCrfxUp965MP6HYt2
DM9dqqpZ7p9pZmd1UGCRr0Twfn2fnuuFb84UqJZtP7z//MS8snLp4XgjvEE6WcmkzewRvDr/OuLi
JMCzoqJfM2e1XLr11oLEaKmHOl2BL+c4nva5wczGTf4xcg5/s5yKoP74hXcyK2FewNJH809dMIlU
AXXGAQ/L4ux9+dORhGqfiBXK6Hn7ytO1UQ0jMAlnr/oN5xOCZb2MQJVdirEXEOH2qp5sHvekWAyk
8iUJCFszH6+hKK8kHIlbs8qm1B310RF4FraYFjOC4ELXVCMMVyRNwsAxTyI75BCumxMist9JfXYy
9nlrGDo6Jqd0u6Otg12g4IDuBFPO9o1Z1sybWklDnZbOV5//ZAO9oSx+DGt3vxwFv24m2MBp2uRu
ca+XdFUGl2G/FOztNTdLqBbXdj7kZIGirg0N2vn9RssbDXW5lKXwg/bUQzkFBc3ExBfQV3blq+m3
C5oJMvHj0oi9SJoHFFc8GJ78vcswseW4M9xOSwJJEEbUfWASYhcF4bkam+TN6BdgQYqH8fbnbrkQ
yZFiMES2D6ACxMAFjhSDw+1OMreASHLzAwIjX0kJzgB9OBqZ4NlE20q7lrK3BjvHxXf/7oPDF/O9
JGQNOM2r6FbCrZJ9qZdXQ6VVOoFxwYHCUKYvUrO5RCfeUqHgmIkSbD1BETO+IYaKcjDJeDHMgby7
MLB58Amf7y+Fqhf4PlbdaMQEW4G6ZDE/lvn1guKRLdr9I3nhZmNSOejPkr9MgIk1CnEULwGaJS65
oHd7IkwNmqfwiurwyu0OeDq+ycLoGcpA1FL3yZJgit5phUNCwg7tEecJ79oDRE2e0V8K8VWPpQvJ
ISUbu7GpZGHPLLVT3M6MNSoWE2HCGmHKfVJENj4QTpuv1DrGKsEsNRMDvGa8cckYMejTa0UaRlBY
gO88YMxkjrPp+ukSwXquCgnVvDIGB1m6Uxg45dodqTg2tff9P+GzY77ECwpzY+qjfap9GcGP9Vzl
edgbG9tOOiAVApFZrO4hWV1foOotU9WxI38D5vdG2l7P1t6wTpErGhdsNT+fHjMdqo7rBM6DUze8
3xf6PorrHsdXzZcxNySaV/XBUwrNalDXrBHjSi65YKWIuuE/VvFf0yTxBHnMGDAeVHt1Fh+5VtHh
rIVTVzBUy0W9mAHyGGoZMWaXbvbKoK4azdkZy0ukrRayMp+ZCsUq5ebvZtXskssP2iQtKZDeS0wT
OqsN/9agr4/SGtshAObauiSv8nE5Z39yDKUQ8F70Fi+lYTXR0I8FnMAkrpnUvTdGT+w9QIFssK42
SjExR3QnsB91yGqkLCdRVXCzHb9Gp2qfE1MQOIsVTWA2x9dfi7TuRdOEf9VnVU4eFwr1DyLnxz3k
cTg6uwStGqrGIZMF3h82h7XbZDSisMSnQ3i2Ar+ylxS3LMIZtUuJ0OZbWO3Zd7fehiVWY0enfKqO
l6pbG0DO3+YArpgwKcAys6blZzDJ9hnP1YFuwu1mkM4O1W1p5dfmzek5LOnMhxdfuEnw3qLQZ4mB
XNDAmWde0pb1O8GDmkPXTQAr/n5Rw9gFpirUkbOWibIU6IrfwRONdPGZRt7VcO75dIivyXIoV8Am
rfNBGWwNi+O5+w0wi1TcZnZIys8mcHJJa/KVtblQ6mPxeArAQjntWUPA/OkE+w09Q31975Aqm7LM
Vpx+Dix0yTtBSB4iAf8RrRb7Qbz1rbY3skOGNC2b0o01wn/Oa0mCkr8p1A24J78UH+j5JQwjRdvs
aRllELzokFXDD/BeGM3U/S1inneJjz4+o9StJfYJyYXDC75ZGmVA+Uqb8o7sFUX30wXuBsHBtSKo
n0adZronNbeS7wYgQc+v2I4AsmzvQeLfEP597z8hx3KL1z6oot4Sc66lNGUoa/Cb9YSI4cVih6le
TwAchmWuZZbDVZoWBDYt9Q9yT7/kgOH/o3HMnojKdPg40Q5uso3pvNoP+jvLkXGXwG8OMxnbnTis
EF4u1uOFVe1swhI/NwXoazR5nR/gHKExw1Prz6/+Ig3uZC6h1FgAV9uoPZJX/+gSb4QkDMLVOsIu
4IPD1Rr6K0lfxCo0BP7fKIildPFtzr/XpxcttqYc3jwqBTU8rbZv1afdRL6lhbFDRvwj0CMk/nVE
ssv/kMHG7P/DqJ8K7aA5AfQsXbqD7CCi7FgwCszMMCICqbQM5wn+LJHEB+1AsuFhIX13IgcSRBQC
EqhtSBfoUUhWPjc1PWKsFU1l+hpWp24iG7KxEVrcKankyWN0XzO6xWYvXRqgfHlyC70fNGCL7wQw
A72zINnQ236csyu6fDVQaMvBoZaiwKDXMDyFKc2qIC6DTPXUjivtLWycBrt8taFmZ973dnTEhfnV
pWx6Iy/AAz+P6Au0Cvt1/jo8CJ/D0VH8g9o2ovjdH/mmi/c0l620byVISGJwVPh4Sl4pKScbDBoV
5VR2CM3BsSzWtSzu0W7iAn4nKijZWAVlhfhw/hkFAeLVNvRjUlLOLLTvg62NqjY15UoOZ94NK+3u
6GfB4NRawLpJfeM+Xdsy1fbDK4IKsPsz5SwL7tGhXI8MD1H5zTnM8/mW4yzeWPnwfCLV67Zk2KJC
VejekZRGfpiitAVVKA7RR0WvI4VLIaWFBT57R5lQw8KOkUXjOczyQPXQvmtO18Dvet3IWVYaWLCc
Z8yHjEHipjNehRRh2xBB2GOFXxbHeYtWQRqoMyupur4/zMRi0d3nLGORr/dgiu2nn34OTXzZfJHZ
/Swq0UQMoZdSi7XJy8KnjTuwTfd/NYeWNLW6uFZr7hgQ67oDpU4kf2S3hJ822FoUkBrbPgs9sFaK
E6regwHiE1BGrkdC5xr0/pbrpi5D1p4AzXM7IBqXen1729H3nrZ0HXm1Q52LJLkLfm4SEAIycUxc
3Sb3BGpJwCo3K4taKBGfj2FF3euY5cNgeTLNXhvxAGYWKo+N+q7OYqy1KUcixpZiatYBk6H2S0Iy
Qw74E7S495urUZHapFDKz3wEKLMnvRV4aZg88ljdo9aVgyl447JBvoIuzSdKA6Ec7S09tqa2ioxP
J1rrvN/URMnoO8cWIJEItO2CrErePQ9qoCh6OgZ1hqMT8Cq9Q/VVfK27J65JamepcF67dIFmeyKf
o9P/OrILxu8G8ddmTUmaMe00FvMv4TDS88i1ZrzhzOnaN72TqRxQ8/tFZTFYff5MyfE1KI/zjTqg
Nc11NsEdwTgeV0nv2RwFKIfPfhwRg+xQfgEZ3OSpcs5fKxyjKIQpHDtfKp+Flo9SQf4VsBoo7NEC
pcAEd+oXFpaAAvByOrLY0hqwbt4a3HpmQX1IE7SF/MW96q1jrjb3YbnArANJIJM/oPKesEQrAypL
bW4TUwNgZp4KHfhZuo4Cd9ujGyf06oRUjFBKPa2w8piBARrM+f/I00Y4yw+cXksXZMUwgsnqy9zZ
/SQ/lofs19E6yaBx9MIZfGbrF6GR4x310syawnQMYA0Jzqev60zghqzvHZKVhJ4b9fwRSyrdTr6B
0htct12pOQs3K7aXpqJCIMBx6wprU5HVqQ9ed878sWqzfj/Xb7aS3rOa2lPVEDl8McZ08CoKCh5b
9hrPCvYjts1lRRIarbCH0qE0R0E6r3zdhA2JpasnROBWHuM81FscX8GUUoyz97WuNuy9ZAVePCs6
EenTSsIKSwKJId81S20OsunxYSEwBX2sQKprcsPQ4bHSWp7rRRzQCawwt+R4tEHF4JNp2V6SF6TO
880+bq6vpJ2wqgiEOW2x4PNA8pMo7a8etSEeAWv2jzFruMwC7B7jh5EiY61+Tm0PAYsaCwQIZ7Dw
GDSlIMJMUmn+JSlFUGN/3MB/RsMsKN4O3/bqwflJV90L89W1NEHZSUhJWhmGvzKwJvCBGlARnOS0
xmqjT4dpe2SmARx0oeCZXrOv7fPQE6KAGHqckfEbzXikJMa1LFByL4KtvVxUwtncdu9l03kYJgS5
HyWc2oTxLEtjddQvJPE3RPrxgaRSOqPEIc5/xZW2OiZOWsL170WS/KHds2XwAvptUOY1Nkto0AEy
DIaYTm+YdUASQ5J/Hv5gejk7X5ZSf/4zq8Ry96TxeK9oxHZ684kfao+aUJ7OfqkTah8PdAe4kgne
wqLgoMvVaB9LBLoyQGnpECV0XPDhqEIPOdV4IfHroFx4mH4VTyyGf0uTklaHeXUWr96TZgU7LyDY
Qu+rZYSgEL8tI0qXVb8kk17Wc3vwl2aaUfgd44uJMGaL6z97F5qFphEHOb5FuEDgJTvWOfIQNFdK
5F7WCW2/xiTgUE2LVYR6USY0FuI+TKaQlfJhf4f6bnh9oRASJx59m2KyKiWkrZVdaU8NumQu7PLX
4kBpUwGzfW01dOye2zEaD52ssbsiEW7b6HwW2rhy2VVQ36fKJnRSOHH+IEybTjW1mVt64Hj9vCj/
Bj8X8f5j1k/fZrYbHziKX4+6dwIrKkkg/Uov7uYuO+vCdVvTNCAxsaOGVkUPP1VRGVUdcfQexiof
bZPxQpWJ/hbfye82KfPxIRKI2gR3Xm4H/sfdhvgDIdrYj0lE0HxR0JmbxuGlUUnf8hbgRDWFomkD
Er7Z+vPrksazGAoI5V75LiLmHIHFK2tNmAsJrgfdzr98suPU8/rwQChNe9vxWXqpvXrqAz5VpWqM
cq+lf5LVYokZwZNmsJr5OJvMPtrGIZsv0C79uSt01taY34Tc0gfVaF0TW1DtaJPmHMDC4NMwb20L
0MFBBBXnjJNFjwXlO0vw0sCw0xvqCylOGD/CRSAWKZXKa+gtyKj4YJeQ2PNapTMSimaAinp5IR2V
wlpBZ3B975nkVrkkRShyHTtd23mxonGEqZA4UTsvpTZkAnYl1fVHhGGJ/SYyfP5/H4czSn/PaxNG
k3JIJPZgtAamPjDB96dyOh0OGWpp2I9Rb8lcTpSfgRG1bVQ33tMlfTLbtLv3WhXA6UWBSfr9FnHm
lV3PI2BAscMKjpbI+w7GTWsn3agIGcXsBviecDVk5Xw8r81LeW8LWYbYtdhPoBQcITgwZ8AI9+0t
h/y1pQXh0/CkuLKHvjoRjwd6c8j8m6IzhipuQMr9fuO3DUPTV8eobsnLssgNvYEo0GNrdl6i6XlD
oJXwaaxnGdZPodN6uW98Ba8K/IdgN+1DdpbJi4Vl37wJulnZoP2MqcWSiVhKYQSJoz30d93gblHu
1ckUazuZvmWho7Nn8g1411/WzB0/hx24ZIE32fJiH66xdQWGlGDU4+00HWIqNHj4RXBimcQkD3XQ
lxeqWsUPelPaKb1aLcm9xDArMd7zO/unjPy1e3myU16ocNK31hj2liwS4bluyBZJEdty1zqR3EFs
XHDukarYPwsqK8ihI1cA1Y7BbxdoFxje4YUAA0LiW2WWhPt5RsKfcz8s89Vh15CA12QQUTpEBCdy
+gk85cWj/q7YgCcxlNfa6WsOy3p1a0oGy+mu3ZVSAx5FaLllRH4UGE/AHRp+fu1HptMgXkVGsjO5
mW0xC2QC9icHNQBl+ZCOAphj9NCxO+bitma9auTC1HOzX12WkIc8j5o/gBbJ0qE1JbitXPj5YeeK
acrtiW9bTp7n40OZmFrmqWCA/4ArsHJ3I8u4hviERdS86PzWW6bUMqbtfX4uxHkxAPujG2zxDEBs
rN8XCV51rHWWnFI8w/c1yDyYotFBQno5hpjl9BmlobyALbBb2K9pxZ4u8o0XZBKKh2dg9ewS9har
ufxLV5uqjygcpdCOsmkfUuUyL3AM16dqpSj2jwBu+1TR0hN4D/0EPy76A4UbHHfr+7PHVh+O6iR9
4Jo+g3SKvQEc1WH/WPayFh1XqZX6eKOaaD7XMf4ZQ4ml7B5zdm/JxiFZUJXm1AstM2UXhm2p56cw
/vz5TadpKijJVxKOk5frtvbLvZiJ/ebDT3hzmKfB5TlZ1U3ffRqUuExXNUSUe+7OtFkOmW+Sr6ka
xBMV2roIEDDkafbi78uD3VwLcgBNt4M8VsYGV3UJdQaZPW4FG57npxjDdBcjnFaSt5ygKQChAIv+
bczxq05DCt4EHnUnme/UriYTvpZRrsQjA65NQLdZmJmRYiv38sOoV6feSBZG7S572/7VN31Sln/h
RImz3edP2ZaQdm+81Y0t2gI+wLC/Reb/FquT2o+7iC4gDTHc6FxLdau4QFwiaklT6k9HMpESQRoW
09xZWKR08pnJfTd1cq8D5CbNdv9vcV6s3KhggMDS5i0dWEbOwj6vxj6biW+BEdTRq/ZqMzCmqP2J
wkI1CAoSqdW5s1AgOToPMxJdHd/+DboejsQDD5r6YcU6cXDaNDLHxzAvNNoRfpEvzpMmplmPHxFF
2vj5w1tBBb282PZtMFtKQTQuc8NMr622sTb6QnMUqL1cNHhaJs55+cMHY2Fx37v88dPm1r/OG67t
bqpWSk/i+6Ln39TUFMSPiKB7c9DUesgpQmG0DkQW72sPy/xAI9MUXCWvMYsxfTnTq/ttqMywqAoA
jxW4czbTWyGxHaTWrLDTkRHfe873H+77Zg/8XKiYFU/Tm92uJU8Ys3urv1fnXhL4nL0/dV+NfukC
D5A2xWRS4wsdxTGFfF9V7ut7ypKxGoyquadozdTGdPPvSVDfY5EgOxRQ78OYayW2SmDDbTPmM34/
d+Sfhx8SyeZNg7WSRMtzZ4SnD6Z6sGeqhnHCk8TpcnQ/ocGHBbA4mNTb2Y0MQzAjgR9OoLOJR6Ec
xXo6bGyZZ4DNv3JQV2cQHS5IOfhKxwIYt9LC8Jc83iJsPPQsKn27daySWXQOURewzlYsxlzGo2hZ
68Z/f9/IycV58uFrszhiDhYm07KCK8Ge+cMvqDXLGVXt1KD86Bwb4M5JpPL9Ajbcjs505AxgCdDC
ne/htbBIFfvA6hnstjtxKeVQyOHJ1MViGNTxbOtXPqkl+l+gGHzthmxMW+qbRoBhPEzU7awfPRR1
02Q7zXl08JTRi26bcSMsoXUjjXUXckdTdMoJywX70k33BjVZwFGNLHwBGrqHHPhLEoahf1lYXm1U
wTcfznDbcecBfVHb5kq//dHzNL2rfT4CyJHiAllzBIOwsAACFWxLW9OG9+CjZaJWVZwHiPLvOxFE
SXShurPMrid98TX41H2hZ7KpoTxgt5qeyFspd5UstJ0PUSw4klV8gB7kfcX4Hkjra0Q7R8/6hl8z
J0WbE6iZFJDwnWUq5VFEAwRSmmEAIUhGmTpckakvXdZbHseteBSL6cxh2p5y1flR623rz3KMQz0Q
uDKjJf+RHoMHBmBQBX6jvDy+g4mN9yPCsSLt+IgM6gB9/eCAxClcJe0/2uDy8y7MekPjpOOB2k39
FBLEzwomOF15XuH3375r9iX/XDMVINVp60bk6Rl8YP9sbSstcayv0FkS9MaiE6yYmAm7eGrDZ4od
4H0lIGDZfu02V2WXoDeAxXatI7ta8xCi5m8GgnOnXcfdvbj4GhXk9PBX/HEKPN1yO+79pQsnCPEq
+egy6QyieqAHbyP+cdjkxyKgLgnROfGfv4KftWzszzEPXUo4LnnESj63E8hnenYDnwlVXY1W9LFe
W8J5rhoMFTWgFFIHG6eR0EwlrppS0GDkfbuq5sTxN+zpdthACWZemJ4eK/CkXE2/vYGFlbHE/B/N
2BdsiOdSrQkuqqGIH3oVL5+wN8MEPnN+8fGMqu/bIGdO/hcr8Mpxs54ixkJtwNj97zUAY+z7Yspf
DWZ0tMqw3Fc8E9QvTQrb9weMG+sXvzNT36cq7/9AMd9RzSmqBsj6oPHoEnIxSkfR9F/GpeosjoUU
JrJVicOXaw+dW18/zrKAlGdlh4c9u6J8E8c3xCR4TP5rWRDZyF3qdceQHr1ZF5rXkutemP06dLPG
MjyPl1a5JkdSprBA8n3zjcxQBYVgC3FTWyuX7NZ2PYXYYhaWli5qohw2+L/D6Q49dCAaHi2814HX
cwTDeTZxWCTNVdQNbeHudaiS0UF1QnLloUtksRXmkDUw/RRSq88OmnnkrHmbI3k7TX8l50gRkmMq
LMzkp04U2mWgospTx8DKxRa1DN0rpWAVxbpvmCdNprek7g/uU7UIAbnoMao+2gmDPNg5SXRdCx7h
VMeraUnEyUrlBsiqNcYD3YvzMINe4Wyrl4URAfUkAofyXVVFuPdsq0OmtgjCPossUWT6bw12FFjT
7675p/y9N0tZEJYa9bG54cpsTsPfsKaUpzFRT6J9UN3G0YoJz8kIUs8SHL1HtazFNrgWlGpHLqoS
8fdeMwdnSCRt906E+D1cVYThdXNlMOJ9A51XXpFKqk7wcRVfRsr0cskhd/XZEKehMSRwkNi3Hw4+
fYn4l55WUlIyX6VxTiKbdZNX4LcAMWEjCREBeMDS6tXne4elZdlUNX9IARTqs60dLyVZM8giDzgp
HnUIBkUZ1DoUYrk1x6cBDtERtEAJLwfwcWHxqFXx4t53yQZua2IOBsEliUMDn/0srmj4Bs5+2xiX
qHPK227m3tSpInVwGIn6cbqEn98y31vIsHMbIId1+Xy7IkHRAsjjLZ7PI7/S7jrU3MK2q3T8LuCk
PLgy3bOpC2Dr3XQsh4SSNnwtasDPJXut+c26633pxfGTP/buMlXMjF4uvBMg/KNipaAXZiD9vHw7
2fq8GcWFwFgtj407EhbEYWfE1V4j9HdXraML1QB7Mskg4wztFz+I/2j9dhv+4y5gIEN/sPGREC/z
fUVjISLgXFB5LM6lTHwyJeGTKN/+Z+acxoBHZUoqx3/B0oLf3G45IX69lgoV9JQhPpv7+kHDJ0sa
tFC6g4lNbrsNJTNH+usDYkrpqeDjYQvMhqNV3YD6ZoHn3IIfl6JHTXTA3wnbl6fcaSOnDr8V+xJ6
cTLZA8UC9SvyTXBgRER/Ah5putmecXxXXi1w8MXuOB+4IryyPXQxO+gUOOX5vCqabaE6ljpjZW1M
C2owgtJWzqbfMU+GJyIO8INjIZc9z5vA73CK+1E8yiwu2RK797l0HviymN/ZQaIh9IZws0KT5TID
AOHFtuN2EcjsjZ2D3By/0EG5oPtL2DHR4FynBzsbuydD38DMCgQxftvLlRpQezxIcd0GeLACQ91H
S5T8h3r1PolKB0IPBUb+v2f/7tns4iJ7V4/NjNmsqb9z/if0DJOMmaNQg56uuQW91sQFQ9mvpTb7
zKU6iDLZ8qncrDCDaNnfeuKw3598VNvby6OqIavfa8ZL8pANTQFFOxG5d2sXG8waDeUL2ELNRXOk
l+e0zhYZqV2Unfod8zG/WEkP/GzaIJvsWDBJAAaZyzCnx6G031XdIL3zQIqiH9xOJOipTyRLOf7j
1OJ+DPmVX/988UCcn2+KZ00ffan05MsxsDNoJxDRRTQrXJGvquh455AgJsbdb6uLdQvNly1TzmV+
ymf7AjIbzqBFRZrEwcei0TfmnpQ28ChCXaFspMcL1B7HuGZvSF3x15e7tsO/jwaPJOmmKfmHZl6F
wvaxPzjQt2HnMCfbAYsNpv1CCwC1z0wWoyEstVghugSduLRqHEuL5tZLApT6WgVi25j30JJf+8W3
9O0FKdX7HVdq1dcFRgp5dExT8climtbb4yQPeJaY6mAC0+amd286FUGcfBRrQtmfUatFp0mU2G7m
gDa93cx/2ZFjDgHBeu2ujEMUMcP99Vn2DYtuMGfkvunDYr+NxL71WOjGhNtdWitN++xJCmKYQZUR
IkwW2JUR/6Qq4b2OxgqA+xqNdoIuwE7c+GC9Hq4rvIB7SUq0GFyyYL1x3JI2PeiOZIOBS2gBJhL9
tAT/lEKyZ1hQPt2R4nsnfIcAJQgt8TjYZGzpTHbj2HbfJfXbIHyBQx6bnV9N3k52RFSJNoneS24f
5OT+gIdD1p/POyriwif/HKlz8e5Lkhcj3YwbrHTxymln7oLS8XODIrdVZupKdyeQSxPKhlXANOyv
JRQSWOluwi+6sMvqg5IF/MvTb/qEFXjvgQ2hGFWJXaPYTOCcpSbCkY6OgpvCwaMgfKmUqreaeSx+
gh5r8LbXZ2s05ENDO3U4rb/bsDPe3976gyvBHElCufg+XagnRbQw/pZENbMOD2ABTml+euyerIPT
ytzX88V/GCv8jJbfvX+NdMfu1K2y5RT2wn4L4/DockX2ByR/9CEh+BMBwddyDL46BmHa48oi0ZcA
ER0lvtmGNEG7mvSU0727jfqYTBx+yha8TQOtwfUBLvVMCr28PyH/f81f94j20ZFLFCg4dwvgNj+V
JUKiMKbVdlAOoEE1+o1kG/6E6anEF97pAQ7Pq6xDnuRoSQ5t7BIVJb3zABTKZIJctmX0yc6Nkopj
EKbo5pFAzrWQ6qoekw9x+FxYAwPeMMkadlw6bP8hUT3/V0qjsAY60RSn/3gpl+tvIRDBOSKCaJzi
zSLDhXs2ci9/QXRhkwhK4pn4G0g4tit8NJeR9KTHuB6VeKf4dmjhOCSk2mCJlvcK4NpxN0NboYtL
oDMN0p5xydMC6dXA2win4NqvUQRSJDbpeL8gY9UUHES7z0El5aj9I3IWHN+WwjLS+iqjV6WjG3E2
aKSzS1LiVUBso/f9VOQW0D3wBFUz02KCw4kdLI4OsnXVnUP6YmXqvDSk2XPLevODranhntvPek6v
o8TwsikZ1mkQMvOJXmAbN5JB5YRfiYRrMym7cqdYhnGIE+A/j4q7eGCFfmARI/2OIFWUk9ZT4gm8
jyCEZJf7YZ5G/Bivf8q70+aWEUeQ5ugZevCFJWqOfEeXGMJ54BpyXrZ7EFbYN/76Pn1oXkZSaOgl
uD9BZitlV2Q6/Cc2susX2AwWhQfCaxFAdwPOHZoeEs95dU+EFz1Zm/0yZm+y2pBuQa4e4fOr3zWP
lpznlrfp1d6XpCIoTdOAxNG5XMWcManXket3RW/pe/FAhsD3nJEt9qCJHXg2hrNhfRw4pw/p3c+9
EFGMJzPk/JLDFp7O1FQ1/sL/OdYpOKglYr6SJQRjQCnXZpkzfg2dCaTex5xCAESZlXcWX+O05k6j
i//mqzYP2BNs2EySW/RsLKr0hDWpapsX+iQ2FuvT9lSUL4YfLKxkbQFwuAi2qPxIZ4d9GfvLFsAJ
EuKIMyC4re+INw4Pa+HswuBCVyUPI5f8JCqT4l2AUCa03rhyPayPMzWXUf51S4CAbz3Q5wIe+pfr
FLh2ee+LicMZhNY46lxBLvaohy1/R6+T2rmUD29MhJVx89hgE++GklSFPJaFmrTmUyvo4G3sde/y
WY342U7D1NDTtF+EVCyEDZB3xicijFdBryA6RwQGYkfwa1rnjGdifAKMIrv8wdM2vjk55BXxo74Y
JoINMK3xz3qxkED9KEqK5a3O3QRM5OtiYuhYd971lfFYLY0uizOfV9VJDApQbThr72ALHBJ0PbKQ
9Nq+RCiuoN1egmsXzm+wYXpeVjWj57wBs//b9ga9x9o8llWWBn1oyBf13+9NQHRs7MyRkgyydd5s
bPG4yZpi1tSqtSo509TLOO4zWn4pj9uBH0IR06FNA5CLySlAJcDmi8q6EI7uARmSmBlT1XrkwpiY
hp9sxXABr5iHkxTpXmSAz8IyZ5yUMAlgkKvOW1lDFH8dcQ9tFDKsdGva6n7SNPypiItk7ocWdcKh
zPdsmT4fMRehlxA99J3eDWDbKiiKOQxbjgEAdFVEdn1fhibErDfiIWHu52m6HzEGCe8JTfdXYDj1
leIugxlAGfqCHsfgSPLR1iy9GP4KJm1PiwsljGptIm3o0usqRFK/2BObOSnWVH9vuKE5S1PfItIS
M5jO8xbafHLXzg77KNafetNupKyR/WpZOs4plY5fWd3ZiPubQeAt6fn6mc7uk3lb6wqhq5MBgr2b
+0AxQ/uwnGksHe3IsAH2pjuUUcP5uvrFROEoiiUTbAy8AP1w4sPydmSO9Z6KCf83kc18QBgz3dqs
p4RaW7GX6dULIPi0FQQY6bhQrD85xZ6VZZRQ7bqmBrzFac5SUDUpNkkFTpsoK+GNOO9G5xjJNPc6
YZpESUpgs/IpJowz99Zlnl1WQMm2DHypajF7b95yb0RcrMP0b4U4FY6uoqSp1iv0YI+ri+tp3AaI
4NkkaFpXEn1QprldVnGNj0AU/LQ9rB+dmRMbQ+/3QHxj3KLTUqZ8lMa8YnlDBRTN2CM7oh346C8C
EBEN+OtSYYpZF7iLOt775jKmfai6XJMpGerF5nZAsB+L0D4foCaxjduoVkUNntnDPjcs27TusIYr
VIdZIoVnFlOO5Qvlp7SZo3ZJoR6T3YMUgaxEKbhoLAOMc/z7XX3A4HRAC2tGDbE0rlESjWmg19pQ
17HZE3gAAL3AfGDMmdCqHHkd6ldnHYtdFLl+QXvSiFD8mq3uArwCK3UoXX/0hn3xZTAqzEWKBBns
L1m6QSy547WcBve2/rulHHrkj2dzPDfqpMMqxNczh+bppwFh7A9j16WOScHbHKblWn2boPoPMQa+
epPkeK298HQHzy2Gj+Osht7o2fJJ5pnuZo6BG2UafisK2144zr2nnSroC1jSyx7Ho2epLVkyNFwS
gfy2LO4ljKgMN5yWvGaSrVNgF2JOHxxXiYhoFWOY57FHv6uOy/k8Exfm0bzcinUVLcYO0L1ITwN7
YW1tJUZXlq8U+eYZnqaFPRZ2Mu4pv3IDq5/ucMEZGyahnXp3+D5jpR16tLKWaSpWk1g1/YEtLPZg
0oEtmIuy+1xFUKu/hyRvCNnEeCBJmS/aeMFI8HgmcR0ltDzpXUV9rnpKCqliliGm/U2GFGUv4KaJ
r3LYYZ2YVwBQvT5FDTR/X0ws3P5Zj7Tzplydpmvn3cdkfzPm71DZ7eoEUSQ0cYCnMmZTo/5eXJEM
HQPjETvcyZ8m34tmRSK0C3SyUR2L2LTzpfSsBGURsvMoOMOHyM+dewNfsSvXOcLL6BuL+bUgHvzk
um2/zuXfoyoO6Gku3rr6c/aT2/gXmYCfffEtXenMh0V2+sHZdGHVua4chbAQthisK/Hxrkt7sp39
uDRuZdP6wCVJIY+De5Cf+NJJLxk3qqhdyPz7Il59K3EZj4HMK225DT5s61BMzSy3rHXnhICQe8IG
CZb17w9ipe7/EXsn8mgdKPdWJ3kPkWN4ZZav/K5DWtgt7orG2LL+81VLb0pXa+D+5/ZAQOeFHDIk
xJZEmKFrm1XHmL+5O3L5Lg7AERqc/0uEWfR6144ib5vk/vT9m3x6ZqOe5GXW5GRtajtj1LBnlvqk
4V30hyNIggzADPWm/mV1lEsGt7PtJs+v2sNZFI+BdBrPHHUm6RG3/Xb1kNEt6nm1K5h+9BKklRLZ
9qhSpr02OdefO0W4llZcWyCler0PrpgYm0JM3BmzhxVrc3B+2QZdUEfi/KNNZnBOgObPKf4zQ1He
7hD7j/4MWCjr7Yu2XWGAY3P2EKTEhwpqTcrpwakFKD7Vkab5PPcYCJqkRiEkDwXuewKvNtL8kZC4
zI3dzuk3ya5aCeiQ1P4j4Wzx97ORnGkXBQE322sm7Heng06q4QROeKR/rlUzx2OubtTP2jF+Q7po
1NqPQdB1oYHPPhUwW28s7TGkofVzcfMKBlAAyelL5cFBcBTsA2Q+v8i+SC5VI8iS46PTwgvIZgIY
aCqyEUTEkoVo8WKdcUWNxW63jRknP5k/zk+DJAPpdu98kM7173o8/G2xO2QP3xK8mjmKJOjT/qZh
wM/3YvLqP9bid5jJpHng47YWp22Aj4+xoXq6Fa4ANlyZ2mft4BDq3FgozoMZjDJJxOr/vdvCGgMa
vKMI3bnUDJ+gRDKznR7J1uZZnY50ZUVRGEi6S6DI9dHQ9dVcQdOl7+E2AC7mWVzjOYjyVGM6h9Ep
CInJabVkx/AkwcHdfWeFHPcgWQ8/NdGo/gS3aOqSyJ9FaFGl3rviZRQtCS++3rHNTIfypNI7pvFH
4zDGcjT5/+JaYlmhNa7NPpVfHLgahNi13Jt5nf/ycwN43tMNuZ1asrpfbiHmLLR4yX7lTnn5C44w
anmtrXzYi1OhMZbZ9Vdb/w9M1exECKclj5gyegMTTrc/YtQxxM0hsEAQDxSkJyPQg1EgQAoWKhw9
10i8bAIWno78lq7+vQjROEzkuayMoBFJbmKg32o3tq7KPqk5WRBVkq6g59dj5tsgAu/vSOY+XtUt
/QXILd/NA2L4BbHjgKaQgn2+MY6Ot6QKe0NPsos3Lfr1Zkb41WLjwjXJq3tTPLrT12S/Mnp3eZsD
7BYGfkNLttc1RqZ/qaeKP3CurxotyaMKHVqpDA1+xD8Dlx9XW3zEDX5/LfB3hQvm81tXWiME3bsZ
FaR1M3g4joOvwgNdMAvmSIjfosVyiz0X5M5u6OEYlSYk/z2EtnnXGszMAuHvS4NeHMgh6bveLp+z
z1pe9Vcc3VDizia4I957K/8FPpVKF1KRLtk14kQST6H2qua+Y46DkdWybCivrdFXJkHh3k7nFC9M
YpXLsGbnRF1EPLnl5+KPJCqgmbQntiLuAu+vHlTahp3U7EpwVY6nlTrgZ7Qpm/hZKsVu09QYNg5c
CleNBBPDs4vTB0+9ioG7EprzVCbj0yuKXpaZNzdd+KQSpOshdk+yQlWILX7sXJPukJPZkCbnus0B
Z4c+Mu7MeiCD1xA3iTpLGFllA0gJC6mvk52qOBjA7IxT349DASx50sWaY0m22ymLXfjYvoeTgmmw
CxKGDlWYwwtsNR/1zBxTgvnsvKQNqooAg/E5eiupsgvJVcpjpHfMv7Ri/sg9z6B5Xohl3Ia8K4vo
1w1+SRkOehSqCk4ErTOcO92ipKFsA3VvUpMwtLWl3HTDEsziR0LoAdaERbMqlgaaO6AGV0Y9Rr0Z
ENt4Pb/4kSl2oHZji4kMwuvKvWpKzPfMGDfQRbKY9Ymwo21MafQTIJZTeWJBiZ4GpC19RLAbZQg0
Xb4/dHBClTLYryWEN+e8CdCaD4xdLGLoX6ALw+YnSj23vhfds6ZyxEmmcFzP+wrlNGbgSfkI4P1O
9u71SUcWVJbvAvKmqUQERBDhlWhaJvlNK3sVlbww9NjwCLkRDaBV02mZboesV+nL6gd6MdGAOoFt
JABhiFOhQgEv3i6+4Ca5O5iZDf7GyFte6VPiJ2H0nTw3qyWP+NJjpk9coV3Oh4uDbyXqaKW0IRON
Iemv/ps+YDcInWoKu83eVlwrxkxYMt3rgkDwFWKtqudFNzLmEvnDY4uqJLPdA81cnrfAuu5OoXyw
1VE51SsxmefoDCLLp0QOrum9OJzBITVHr/JH8DCFElTLjVFeWf/I3f71D9a1Xpxjt/8xYxklbXMV
tuF9wzGeATxWXqHzO5jpeZiystU5tqT7UQQ1vvL/SdW+1Jc5LI8cXqOc4WMtmFWNzIdIFuJs/Udj
PBFCkx2I7mqsve7iHzevFAhhRARWKxvpTs71+zhoYP+Xd97Roe4AtZvpnTd8oBgz4NVIFIAu7/Pv
OpDyS11sOu/mUnAKfWI+tblSWKYJAG1qdZ08g1LW8Cz5g0ASJ9maPFIrmuDu5goggcf3JXpAMUFk
p7h3vhvKLjxcmT+kXkbuyUiWb+OaPordruWVWSLEW1DCLy3iyyj7dLE4PJhL8d5DvNliQzny+Lur
tMj+jPcWXgvriqt7ziTYBySs+pdBG+rxr9YUo9zJoWQSamozAQ/agwckKK6r7A6efVa7KEJVObZa
eb0zGneE2i4yHKQXJyoAfs65ll+QB7rD0KiK2Aft/N75OA3LPhlTVSsGftffpuO5KtdZAVB2YGna
j643lgtTrcN9A0neO+X7Mcwx0onScKrAd66i/oiqxpZfTNIIfqGZo26hrRuBISc2T3gFktnBRvHT
7UoH2XjCX5yhy78dozZg9s4F1u+d0OVcgGrtpz+oWbY+W3xod4dlh5M172uTiKAcy75+ZDtPjeQA
p7IBpXAo6NR9a2kpOYlA/xA6WPv0Dw+dgSXEi13dZTXSVAe9FSvj2AZx8d/K8Q7WffLUkprMdjOI
Y/g6fIZJHwBSR6uttfbzZmzQ5Y0/XxsR8mGRITYOIl36iBU0AbNEr+YIw1gHeaG6771ywdNwscut
Z27nj2WhATrgFHnRV1iRa0YO2KTDeYm7OFyiG8bz+wGrNruptCC0Se+/uoW7wV2MfiiVygTLhMfc
IBI4OV5GxNSuEQ+JMLD1XyfsH3h0ZXIVMWmnRG01QC0n5zQLi1iSiNXF2Vxwntl6NG3Om0j5d36f
ENI820mcZLnJnPDyjsqVhrjWjh0YJ4W57vc+aqDNH8Q6U+y8l1FP4EHs1xULF+5rFsTpOR9yUEvH
NlnQECyJJD2GhF4iPI67UwJVMZCuliTYoKRNIWIJVpNyrvBgGOs5Y8OZg+LEA1WwA94TM/WMs6Y1
BQ9j1Mcgl7RjhZInykOzh/ZyLoxV5t5LYnK31YMJ2LPRtLHhIGuOxSzEgRjWXP5xK55lPmCWw5WF
k+dTTWLB3d3w4trMZJLjS6TTFOgnHd7e60PAK5BSqtRHlG4NjPHdNydn6LKgtjA0bT32FSXGEsnt
ueKUHJGCNP/B7fI2QZQDKqtnrH+pu/q48XPtz6n8IrA3wh2egKdMjPt8TbiscvEOEE3FCK1JO1Uy
mjFkprA7metQf1m6Mra6XpnaiRPX99Ljn4M4fxUKEWKgwUarYwKzE5FXxfCnhzz+2FYg1ATOIBkJ
5dmK/AbD3Kz2Zpa4aI2iP8PfE+U+j4c3dAngY2M4If18su+y2lsVYTre+mjbJ9t+5S/1im97Z+AS
1cqCFzGKJcTNQp3TtB1UMkOM4TsFStJAuEZzGzoTVhPImtJwsI8pYXaJKUWouaATdJQT1iLfYdVV
S9IvPE6JD765rIHtjKWOSXAUG3fmqigVDvwjr/YVl+ZqgdytSd4dgy/i1aeM7dPGXslv5a/D6J/o
DarMKhb2uGKP4wTEKoWqZNviq2gIJE+qTk1N4dBB6CVBh2vcWKlABmKxTYQs7kGuCv/wlmKQv7cT
MsUSsXnpajnmS4KSDa6D7ZuhH0r1ISqKoxj4+EddkVfYZ3l64prfRviG38OOLLy5gZUNf+kjkPP0
fUZIBHMg9L/GKH3pT06WYShBhBrT2Kab46cWRgHsyA9mGNZAqUvFm2SaIlmWmqjWHWKKNUzTXJpc
K6dl+NAzrRecpBaRxYeNA+i2ryMyHbcC8Ub5a6+ymXAGyV72K8Ky4Krr52yxGyGEkI287Cty35YX
bqGh9MbKcIttiNF/cqpCrwhDtKjzaDzRdANvBDEKBfgdvWTFw7gyKvdvY2LLxo/si5eqr4svC9JK
j8vEmpZaSSDhyhZs8aLmF0vNj/Uubduv9X7nHwFTQYujZmma70QeMTTKF0Ed4zGV+D/zouhU+6TJ
eTu/8XJtRlktz6kFqIzQFn773DjJOSaOz3/h8J1kIi6XEWvx1mj6SXFBs7XoB394F2m+n10NY89J
QVdcCzRs0EPEOWS7Wcl6fLQJy8FE/bKSNxKbMOXPOdYJkRyLjM3Ma+43SJGJgrN5LWOjK/ZVs31U
S/NDRQC9uJxsTQhLCn+/hn6BIaSoXgRRMbvJX0mzSN3ktdhxOXjTUoKTA52qjP7xOkoTXYSM2dH3
DPwXIncGWaMBNtw8cZ9RMikz5AV8kNkA5UUJ7c8pPCVjzRHA10NGd8n3T26P1hpgSgDB4efwzzLd
TOcyGOXcnrLqw0Gm/4RFxbSy9VlCcNGwLQ3zn0OcfjDYkMQvqIj1EGCCaoRdbjfVUdYunwonl7nI
2iNrMn4Moo9FQ/QR1J2gwf6pPzfkx3c0z9DegOAb36B4YyiWzbWDWuBjaTQrb8smhxFLOLyfriSo
wYzyNVBg+c6zf6xxBvi93maDTs49cU7YUvNwwDcaVvz9kMn4fCy9WECgaD2C46BEN4xyL/USV2U6
T81jg9kCD3N9kjQ0ogNx/nXALVfMVN97AY0QxljX+MtH/26KSNYKMWDM0L3VRDylHZeUXtItW+rE
Ky1l/e4E+Uh6XHiJu5Koulc3PrECsr/X+j5rN9mZofZSKuOwK54MQzoYMEgnZt1Kz7ps0qqw2Kpk
BSmaa7qq8FHUTTnxdjx9Wsx52G4TXsHDGiK9CQiSX9WZGNmNgRJ2jDL1yBTD4cBWUVLYz+EwOye/
hi2p12MdhmWWLUTOKlPgl0qVN+dMngkxFtOpSQAEsJHP0R0tIUhlQmS/uOlnD1rtjPUVKXbUXHjc
MszcM0/DNl2GNUdWx19a/cyIefpQnkNoUIW1L/itHNyrGGlBx0rG05sOAIeFi2aciysoFRgft3Ke
Jm3YODD+VV+gTXokAem4z6+yS4Ut8OnbZhLMCPiWzNawPVUO83mlQhbOK9Di/u48DVRkSE6JcW24
4ppnLgp2wSyETFQYbuH8BI57rzZNiPXRfxnRVXyxLsU8mFhBXuQm9ft2jVVK1Je2jeS7j+mZJ4wT
qcGgn6f5bLI8/eWy+Kvc7TcQVTgP24HPPipvbtaW+rXnr7hwYlGk8mtRN/cMqiD0G2jzAX4mzoja
vy8+RaL3poHAZ2U+W+w7Jz711CdPuYMpyNIsOFY03r65wbmE8bcF+Eyaa4mKfIupKgD5/vMAuUTw
VozG47dcLtt0p1/BjvcswuEKxCswriwuRzP/Ma1yEVGyZnVrsFAoHvFrTO+5PpO6O5jB/RXaHXIk
n2dnDttvA7+aswisnM6Jp7KMappIq1jANAHNIXqSS0e2OLGs1Kw2CafLfFDYQQlScT/ZsFTgwEsx
aruOhaJB/bWX7ds2sSMyT7Hj0Oe4g1sU7iRwVz2D/IX2ZzTdmDiDzrOAoQzQBfjm7QjtS5Fw2PVT
NbpYCyeVR/KE2r8w6a9IVEojmLc/pTB1Zta3JCvc7y2KncBiSswvNm7GfHCXq2ft2lnFWNiFAgnW
8Dqke/Xr08wCyhkYBaOR/DRpwd8cmPjAcV20crm8CgMHuRjqN3d7sAAuaDkRPIJeVUm3yakgMTfR
Y+7+Fb5OKw1taec6v55DFXlYO5gA90nr3qoqhcOCttehrjI3uB8LKRgRcK9vS71crfVLZ+UCgvPn
V9G6SIocnyY7e28M0FijClbMl7rIlc80ojViV0sWDAoF/lSQ+Lu9Bn5Bh1LP7xRyRmU1681ll/lC
dzg7ujmYSXk+TY1ePlKsVXJyJVjy7wedGuuo2u+C0Kl/m3qJQzY9n/0lU+r2sT08yaDnoFKKGNTj
ON44WDiPeB+ag693NPN4g7bqPFrEk73VvWXfEbd82q/XpMpNfkZCvhngULNy4jH4EzrbFjY/rWuF
lYvxBPQSWduRbAVeJLfxv4XjCnxRkb4F2Fc8Mw2R+jvjXhc5qlqqWYPm6DbroYcZry7HJyWDyD3L
hTU1kUhge/1JgK3N7vQLKMKZPoZwvQpsKynUJ9eyphX44AmsFd8O74fCbCTpr1bbs5fqlUlIgvoj
pnziPckJEs4TDaGlSV6wW+pO6YkEIf9DGezRJshZNdpduh28bPcVwC4EXJSw0KzIabeR4c7e3XaL
cGPYP8F7Gz59ZHua2KiLfofbi8lRY7vb97+NKw0e3FUca7RnYWuuwSsAx0sMK5gTnJBXwjXJn65r
9Im38V16n8q2g1GH1emsB8uaqF91seQV8/BzoKqVEktST4/XhezlYExrt+rRZrNWXqsQ9jHqaTLi
7mdL/UZ/ixSvqbFXejnq5JWrss5Pu692gjyVDutNCdCFpoWIKR+HhIfiXlykVdPobBintoWmztut
WH1LKpjWVr15LUQWRwJ43rCem2iyoqTpgBErKTG1r9D88UFP9rrzqlBvO+4kuHLkZ290MJqyrW/d
d44HHugqcoRDcJZxUs8CPVwHg6Cco6uFjA8cSxc7dcH2hBjjuwQVUVwjLTv9ZWPBCj4802MCz044
ftHGSj30BdhZ4pIXXlgNJnu5iKdi3J3m2JdjUKg7gi1z51iz3e0ybf3BbaVx3fImH/so6/Afntab
v9yCypm2Z+OAtYskXlNQbKddTRMhgBoYWOOusUsB7tsoZCsuW5o6tadrP0wZ0/nQSSQCSRHBKn3y
oa2Hc59OP/Aes3VzFKsRehseSNDCgmyShqU8C8uEIgJ+VtQPBdCc8psIgAL5Qn3WguHVYWhfcNT/
wLgMoyXIe3sqiDvpYAxdbdCu3r8Avz0Y6R3ApzGtqCJxKYYZ5G9tCoYkrCMnCjFxPiVtRX+3OqT8
tQSCE9OQFDf1aNvZTifiTPeGd8Zpz4GITH2xRR4bXQFVxsjIS1LsbTep4EPsu80ugtVPREFjPCLE
fvLELM2Bbaj6u2YigdIXBlYdFCLEsWje4fwAzyRYxcIUnKl+MKgzWCvV3MjCkBDt/Ba0azjNJn8/
kWF3btsmJ6M0CaCnCw3wGFSZtWNLBGcCmeE123JPNR1hUjI8pGbEu8UaHRjGaL1HB0ep2M3jaCac
DxpE95vxFiMl9Z07sRJ+v/rInZQbf2fv3Wryi45zH17JmPCQO0D1zeh7ESW4cuBLTCLs2bSuH9ps
nN234z26Dc3pGX9qTJNJMgu3A1rd33kmC8nEtieIaAbHy5qt4jRHTyb+7hgGm+zrOe/7cpwmAvX5
ZIZfeeknwH3GFFoBkQhURF/KnZL3hDx5dMgnYS0keD2Pe9QCR2J7xFjWHPGf+IYWT+pDYGwYGN0Q
mkhx7iAFiTPIqTW/p0HuHMLCPK6raaT9NtMVHmBKQbyhKZ4ScK8CPg7Ci78XlrzFmypFRabVFIOd
1x1PaJdeFAuAWODEE6m0jlKGt/rulTBhZJPg1ruy9jLoSHwpRcymvkXTXHUczfZwpSZ3r1wyydad
x1m6Vn0H1dYxIb8hLMi7pyyP896VIqV7tRZW8q/18YSB1wh5qsZq+BxmSDnkE8NArG+5jU0kmihd
fGfqpZzyGqGOghLJVuotkYfD/GSJQJfL+kP1G426NQPrDTDFqgn/YxQHEn37c7lY4WteNA5vYBxb
hQ1Os+Mh6i0u1Frr291aHtkSHcbRLfQy3SjAJD/mgvL3N6a/iocDTF7c13MfsPR0Og7nV61JhcED
pd6WjTAcf94rsAJHCBav+sMcgTzoCn3M1LZffYw5ZNlK3zNT44PjDfQcKXEsF3HPn1LS5YXtyvaQ
V6n9mYOjDdm0TGJ6qxEq1gTdSy9nknTCHzibRXmO0UT0Q/hmKGXzyAdWfww5Jq5WY3IiX1iPqnES
+6kgj1zRnzy5v3PVHqAP1uIHpP06UFPHXg7Tyxiu4Vew4EC0ixc6JG5UmCKKSbI9waIb/uYIgNmr
AZqcFfyaXtQeiZYWplpHhHeoyjh/ATcRYoe+NYIVjj10U8R3pC2VwLr2NR1eCrUn4JnDybSP1DGr
D+pYup/+ww3rnhS3XCg2jPM13o3NaS6f+A3sVoCUq2qGvw4ThwhlrCLvKW4KZ2nKRlV58rHv3HOg
SaoULWRBoTQx3QipeZG9BMXaj0l9uPORxbgg6lTVuUWQYm6jF8LQUoIxLZ9n16QVeeb8xyVatjoT
ETDMjpqOtAKu4lM8aL3ANgL8vsLeZyfPoyUcKCUa2+Sww5eHDLnF86eqr+6SCbOje6PIlQVa/Fd2
IUEf6ACBkC0lXW+3X6UAktuDiIrsbjF5NS+wIaCPaNDwjN4DQ1piNWU10TvThUKBDC31dL5Qos2R
qY1bT1jDydOc1Ug9IAkNKYdgYIbZ+zb7W4s93oU2IN2Y5/tEMsn/1ZE8Y2X+48E70IoMYHf5dmZG
dkUyJnHHx/NVblwykL5Vk23wn90PbiCXASH2KeyXQq6g83J6g2aolRX4IFlJiE8anNPPR1cwwa/d
EH1G1rWwcTKCBdeHOvMc4BRa7VGp2clvjyGct8J2wn54v4Pz808U8Qbf6rU2qkNfT/jGI5cRenFN
+WT032/zuwo2dbHpEf1UX53pljnw7f7aSCDmWSshPSNMmbA2xsoA3dGU8odU6eEjjgBikb/RY3qB
dbGh1xmzBYWuw50W0+OvGWQaNFhem7EbKnibUQv4WIegfxBmOftoCZv1vvhK7C9pc4EFSFk5Fa4O
T0MmJfCfI5zMRLctEGqi/UHowS36pzughiQwmlcalipUUEDngqyGdbohHWgjjbIxylMjJ0e4bO5C
MQEuVL/123hLak/NNV6DgYkr/NYdIRWB6eRK0MZI3ABew4beQiBWxoXQ8qCMT87cWxm9rX9pJi6R
KJ/zM1Q4IExg6h7rCo3tMW/LcN4KMwgidQiJMdzy2AqbKLV/quueBh4p3UCSmWvugywiPsFMo9UB
nwzatrpgrhlagqtdZpthTTbclbGtozSr63lp+QhXjHihrK2BhUbwcoZfjdr4GAbloAozgfUnwDmT
jFoiBrXUF9qiprrbEWwQc6HIy0YWUMfGWdfMjQxaD6u4HnNHBVe0oee34QiJXGU3MQomX5Qb8RWy
MqT9pqJ/3k8kxUatRWQsJW+J0AODPVP/fSYlujwC04iq/0E18H/Lh/chdEYjz2Xyzn+2fJM3Zi4f
9B+rn8n7ulk5IbikliEHydpmFyI+OU7Hfpk1qrePae3qDoi2dPWA6cHbQP17eTURY3i+slIyMQnM
7VlMF8ZRr6tX7xTA1eHx5ma109+Mf7cgRbMAaj7R5cOSCL/SFz3vs7vOJk7WsFULp4yY3ez5YI++
hlLqccgzF+B8kAIs2yAuvx5U75X2ei5soH5SwzKl1mtDyooxMpPBBWhm7YX4yjX4fr/okgg9Jlkt
q9+oxdx9RhM/WT3vZ5s7BHvZaNs4vd6fRHxESrd54Z3M8Ck0zEh2W23GjbFjjt1cSPSTjva2HbKB
iCgPQSMtwocEO/YLHB4QjMATbagBwD3krM0DJc6uoL/71ySQfZQnOH7ngFyeCfWKgTT3+/SZVM1L
faHVIWd2R/8ZKmhQmBWaXe44JTWgPwsP+Bp87n/hbrfYfE8n38u7dC94TczM4femDI4vmRN6M1P8
Y0N+VQ8G2qR9jKC3ukg+BAOsp15a6qEBDZe0Kk8v19FKVCJwAN27jjvXWScZ9PodLZC0dynd8LT9
9HtLfE5SnvCaL126eNTNdcBzJ8jMe8DCCpea7CTuC6oK4q7u3QxfdMrFBQ093L6sCbghp2nXHlt8
h3LdqlJkXvNURdupdYr4nfUwg3KvlH+Y/Gt+rgBbi6DEdyMMwb+JsgaFClXw+GmQV834Oo4T2x5x
pW7/4+7ZcCzBh1bmm1znXu2YJuD9y8N+UhYTUrhB28Y+bLo5Km4LwpQkmIPX+ebZToCiGkCmbyWM
AoZd4PqFf17c26Xw51dhFAUUrmKIfF4AkcY3qGU0U26hhOjsukb1xlOOf5aA/2zzyzIgXC7rgafZ
gFQWtbuyHb5fhSoPgEOCP48pnLSR5BMxQiJhU+s4xixCZi4MP/ML4b4FhBCFzqtlkN8P1JekmoOO
2RgP20QYAR6xIQg8j3mW6/RuwQNMlhquoidEokI9zRbQjqRj4dqjTTnpOh19jBYMnRgpv1jxaGC7
eSuB3lxNm3Iwq6Zpe5zFcPdCXsKo2cM3zD8HGKtfvQlic+UfD7omxxLYtJEXgusAyTG8neT4HQxM
os+M/ANAaPv5Fckrrqq2bmp7dOh2QG4E67MYqluPhPtCpwr0j9kClt9cDc8J0KUGW9D7GwkojH8x
C7uAh2fMMe1RAmgXUkhzGzDKdp+9WoP0oDe4D9Pn/5QlNJMjK3GcB2TvgoeFyC09hWSfQ9bLvO+D
CFwcMDkQUQoCcnNNMx2ce7tD7IR8w5Q/W8h68uCC75QKGYsKTWmvtto4EBAQa0pXPPyeGix5rFUq
GYxGnSlM43ZZL2LnzTMFs/21kYk29HS5XD1mtiuOotiGm3Y+2Q7w78BpDoGEoi9PWCz3OfdtRPD8
pAhvpgV4QPNbdIFRwugSsB48YG1CsOFcL9d5qsbkuehI5BE/FNf/K6o7CI2SUSVdeBkDcpg1lMwB
NydK+OjZswgYjctYtZHMECiH/PGeT5VNqdxfDiXwn+5kwwQs3fzEuk6pOlO7UTfb4IXGSoxThWM6
qKKouK+5MekswJv8h1Scoc+WJuvfZ6chRMTO9goy8v2VeFWQbf/XXG8Y9lIItAbJiFIFFOP2vQid
LQHLyNsLmMT08X4DsHQrMhrRAIoxLIQJxTwW7ZDj+gY8mWnDg6a81C4Ui+ljSyYDjf8mbdlvznsm
WCYx/IajdU9PU0m4IuVRQ00zjLYXXBqMZs5RNJoQpdziMArc/dzmfg5AzwaSo/5kI270IBfn7L+u
L8jHCstqUjwPbsdtkYtrCsV5feHBZHNTet0iws7JDhiCD2yORAqVPy/dnCsDF3EfpLpDRbiUt62u
0axEG0qoByG93EQE9BWVxH1yiXiqh1tXhmssGlAHIf3KjMnltTVQjiLVID9qj9PeA3JGsULKW364
EAbzv4glgOB5whvVDy4C9FGKC2egMux+JvOV5+vyl6noWuOowWI2PK0v8Nct16OE53qyD5X2q0+c
AxlKCmdTgFLt3h4AITULCqg+L37MLrKLpOcwDqkl0z0icTAKcuu0iIaE6RW0gQFE66qVLd8v4Wty
+4r+NIsf7DHOkzRjg84K8NgJbbsDZipRQZT3Ca0Qn28r1TqKfWSdnUVot7ZiPMG/WnEbj4HGvtJF
Pj4MjzeJDzwBQmef0u7A5evn0uElVn99PEvsrsdmHLQdrQzd7aeLrssaTLMzpN2aM+xVH6yYdO4K
WgLYzu0A+vrRYP8qATg0NCyaEgeRT3BzJNThvjD4z67mheMAPoeSiUxKz5jgP1fkpscMnH2oGwBU
7OglUa2jHAHjMrvNATe3om3fKZt6RrooehXC//Qi4D2L+xuQiAwtyeE7aZxARwtegTCVkUx7MzfS
NFRiwTqCFSl7dDxc5AUZxo4cCO98VkJqu9Uc5tZbr+WWQxCjHB1xztGHkw3zGkRBKkhl+M5usAQ2
ZuPUMAkGKrhR1IILbptdQTq/gChRJgsHGFoQDrgpvapL50DvwwQ5Vw5MckXUNw/lO+kzDefoDCsg
bphMp0uvyBwWQNKp0NHrjLoS+WT8W2y3QcbvU08vrJpqP1LjPCQo80ZUlsqSIV2gt7GOTo3R9YDe
UXXcsPJOZnlApKcrNgHkO6b9e6t6lETeNXnLAQY5LWVISn+b+aK14gKBJnrVukxTIF30FNo2SXkZ
9JMmG1RBeEi4Gih50etcAoTQa6hUwGQ7XWs8v7awe5cWqR/wR2UM362FcAmrAcQGUZxRt+FNT2wO
0/t7di170zfMrzvQCNgR022hO7XiDDijhL8fmeVnLSqtTWFYxDIeX3PIrHy4SaQjr2p0AKacS/Bt
KkO7VigO0EGaogro3rJVOaj4fvKr8zQKcSUTDU2c0PEIW3h09ms7LUSBPNEqe+zHSgvOZLlFruUD
AygaueihDOE/OeBHA9eY1Vak/5HCOZBqzuKE+6Yl3fSo9UKV/XDqzxPBttAU1CPgasIIvsaOAThC
EakkRRYwHGFq5zCEvNRXhRhs8Clg0rvTzOTRuaJsfBOTCixKOsDWW92iafbQb/lnJqYcN5dSw7cc
cV/AGeryQqPriZnpvCKMesMCUnZDkfbxZl30ZCskJEStJ+2wNzNlOJ2934nT27Oq7SVa4rBhy/Qg
t/+4hw7cW2Dam3VH5cxZj2QSY/FHi0qpda6VmOFescfJbXacTAdUPyTQKIbUZqks+JXsTFZhGk6d
G3b1PErG4dISbmC+1Nf5cx140zHlPnvLiqJT3iSgjjvEYkp0JBrcyjaxy8aJaMA9gTqBE9uP2GuD
BRkG+OOZH0uVB0xTv9HX05XDtg7zMhtW4m5aq2+XTEEB+7MnDaOWKHhgRUoP8m2znrHZ/oxwW7Wn
tPVfH9X3jG5GdbvG7C/cbDwzrvgFvXNtacS0ahVl67YBm+f+kmj8YbdIb3F6MvgLUizCFy6DVfy8
+KRY7ADXW17uzjlIJkNxeADWmDenrWm2uYJO3+inLyI7OViHsLv/s9CLFehJ53Dz17T315piApqa
mXCXahzR2f61E/1w8sWy6HzX0aNozYIrNHezYkzggeM456rKQsgVExOWTUBslnREBE+HfetSXGcA
BkFLhsJz5ZyV6Dc7TfzSAAwGxYeY+WAZJ8NpPA6sWoiKFAf2LvC6uWu2V1eZujW9XftI3tHwPqbr
kuxrk35PRyQSJ9atNqtukRqgCwy9npFoLUmNJ594ctT5NmuSShS3XHcrtQc26FQ5PX5AfOYTdS2X
9pbp1TbZy5EkCZEE+Cdw/VDzfuqmwfhAB08n8Ew78ukDF9gI5WPVObKYp/iTQugEJLJeGsNDG5Dj
rL/+JpL2wQ9EGFGG58pQ0DC43QSu3k7IYrKXuOCmU1tZqkd82lliJVQnZx9XtHphVkwQC78RQN9V
jY4001Yo/vzSqZpyn3bQhLxC6hHiTKFIi3nH/jqTwgjwyHUJp3nR4lgz4azTJkhxoEiL0WfS1mkz
kVRdVlrrkdb4iHZmSSE6ib5VtkdV5IKayoPF9dp+AeTa4dpTwDkdx45kYUxdVEkf/vnhj0cphtAW
nCf9g5EOtjLhcs4STdmBnhRfxuZ0Hms2Ff1iyVhyBdDhaTI9ydNAxSeXXZwR0gr/3jmXts/aGg42
ZMh/cVyCxGaEdal+L7/0IxC3XpXrVctDVtRrT6QogLghluNc7C9xzUTIHATPhgVqGBk6iqhSxYJy
KXx0Jrr8rpvIU1PfIg/scUs2bRr5ublR7PwGwN+WJSvor679B/rV1eTjnV8WcLG6ZwudRMuCxEKG
6HTBhzTkKDw56aDe85MyIavLxpzkhFflTe25NZjEBJHAelqKvTjTsqI5Tp3A13jVZg4GPNLMLv0R
GCGI5Djn0y6hUE+l5it3Gl5SZ0jkCtp72fLV61NT1ExxhG1w53U4GrmcHC7ibIc0DG1gscxLAJaj
br/LMSb06nmdE9f4C6wa1KVGV7+YIpN9hvXlAo7ncUfaXJoptAoo2aG+phzHj8peZkbcHf0G0IIg
kgceDrWPalVYyaW18pSW11cvqnbVcMTWh9MCBdidUWKZ1rXpE5e0Ya/OHmrvPUE3ZwoJqLE7759W
e/Q6d+hp3Ry7mbLdDAkWyTRbwjNG6Gt/gsF+pnd1WEI+m4C8xe8Y4KFvRbeYrvucCHpaQpfpLfZE
uNmkVtP3hJb927gRb4dpx+nXtkhe0kxBjotagzq63y6Rot6T7NP7k4SQIev6T11++zQdiKg1VkrF
uQp17yIKzRqnnO9emHjdtxqMOGVrK9vZvp5x+7Lc+y47vJ31wxJeNX+c4pNMTvuv00k06DPWzmH6
X0/Zc5vOwTWtgz+/2G0+axS/22s2Rwp/ezA362HJu3KONihH2ZCBGJgNQgvDxijQ5UYDzmFDuJW/
RUpT6QeCtphVQNZnllJ0RdGISG4cqPbvNYfIH4SgxKF+uKYtCeemWOwNkrWahl13c0Cl4s2DlBPm
87kSeXSJeTngwsCwNiwHhzlVwubf9m2TJk+sV/DcNpGfjG3FBfoZ/TIGEq8QKAyCBwmorMbsC5c6
WWu8NlCvxwDueymFrG+pgm+2+K5a4yEA2DhP2WxJyJ/oorwFTPBazLMbTrFDV0MLCQdq+tPvgE8a
jlEUlj72fVUZ6SqYiF+3UlQJvtm4HVWf5wbF+5gno5a+l8oSNqIOJbJ1smFJakApGuaA+0KC0Bqu
ufbTgDZmweybZTMXqrkboC6z61T0JP1XUPBdcjW9ALdU/WlG1UOSfCz3Hnfr0fxTpaQycw2Pv9TQ
2gQU1I0bC90jp7NWyf29eZ7GknmdOG2WZNUtWVP7quuc9g2smKU/n/BPcYTDOmhGQMFvXhazvFlD
EwtBPHIYVjV9kE1RvcjC8dXKLLHDDKBcY7lzCHRs0pQIkaxHKdxJ1WG6ZxbyqLK9HmCPzAy9XlkX
rttDC/fvgarZySrzdlph2fNY2c2TyJaLubV6bUrzync33q30gYE/SDwzTH0EUqM91no/1ZaYuX3z
KmgI4iTtJ+02VzCOYH5tUNhrenNnjI0yYPnUZlHacxkVpAytwNDrvE3Y34o32K/w69zlFUZckMkD
lApBglAJRKmMFAHhIn5w/TzFM0sGNy8X8yktqkh9Jubvu4byBEgqiiQ7ZRT77q/mvZvnT1Ly/Hj0
poMOho1O4YqCVoGgPWyioby78IsJ7KpnqRLtXIyYVGpUKRXWYct0R6B3jZvW4tDYeV7yMdSi5QmW
3CHUZS6PUCdpOBYRBnZq2+/PnIp3dtOkW2ctzAHKP3Vc1fK4i76ZUilY4CjgyFKHfBP6BPZ0FVbC
jK148cY5JKsiieO4MmiO4uCN2s7ekxp8chEVVhkSVrMKVl/g2WbP2g6hbHOfFrP+gzIsjGkHVLle
w2/K8sn0z/otIr4QN0YCxGMZlePG7A+qg2uIiv8G2BNmnkAeqRZSAKqTrX1I93/cQsgJtS1aJ2Gw
rz28GS3EWihxTfrTmx2fvLh2EHzje6vIl7T7fFCkVH+WFnjwTi3I6go0EKdD7OybEN80XzIeikku
XguSiItz3e7AH2HwR9ryWOsLQYtpocD5yAACIpw2b1E6UURzuvX9pyHoXh3whNA55GrY4OgGpDgH
QLCbrf30ZZPQrpt8HRbRclLQRJzzS7HybahzY9opQViFPI1lwzlQCOXgeiOc1OuleYMAf0qS+OBd
ytxpv6rxXkcPQ0zqw7zN1Tm6VK1ul4mP99ikXYHzcLwCWZMh3mCc7+APfdiCzwPtIsGTQphg18kF
LbAajqUzFDWBpd21JNT2UQlbzXsk9zZ1/5FjQwheIvULvS83+6CqorLte0hs4hjBao2DiNAyk3iO
ET3F4e97XvcG+IAPKodTHU4/xDGWnYl+V/Dgu+RZJ0NYs2dGWh+5SY2ugVAeNWNcVEw74nd/25gV
dccTYJb3gxGTYgxuPdVWiLBsZTVSDexmPvvDdg44muExMacRGydqj/hg9zUFMxiKHhxVLZLVeewG
3h9wfs5/NYnAkCHhU1fOpBw5E1CsNaspEGN7KU+UghlCka3QXHQsxYhRSYvYacHMgXaYjnAbwhG8
XuSOmQaalBMSb+ECskyc1zYQX6WjxCry5iKhsZ21qxKsE8hl3jdreEnbVs/rKTV/hg5UGxxJaUBE
2fFhccM4vwE0gjCuaxBTRklN7N/huloDht4sWTP10Ds4XSEK1QdZBTiEi5yCmu3xKvpPzLkkaPI3
7jec8rl5mCbU+K1uzdVD/XvOhyKfFlJxU0lhK6LGZEvzRs6uM6wDUqmthSU3kGlFPRst4PeUEmPq
p+o1rNBPSqfBCscbUsDzMdBPacXFjGYFaE7RV0b7FO8b/6bs3Ndu6w5DziXSEtR0UlASIhNPDsh5
wVksMWihbYLstcpJ//axBVDfxzfM4qJOQHZpJAGSE1RR9tcuV1JUlmgCYpCmMua4Z1JuMDLvm5k8
xKHtKJCxraFSrCKfNb24D8zU4yhX8agqDlRtVk56Sk16OyKi6tgFtTNLvY90EhuwM8HVmZWR2VPO
sFZeRohGiBfLphgp3JNKXRT7ix/bmYxfrMisrTiAOMNXAnVP0kYUYZOIjsPTpj6WoDuHBjfmhpHS
KVQ8xJgDkjwWG5M+0R14w5Fi45OsuFTUA7W76alJLaSxuTKqy0UJMSHlt9zEY5uVpL+0uwRZ1GRB
ThlE3pPSGAKUVGMP7F7ctJ0OcSvsDSgbZUJjuX19ydped8C5S+nu+z0LvUP7ryMwn+3NyAYUAOCy
BDK+CsBgbUhyn+ZSzDcyZuSHfPtCv60PEbTHuiJ69hZ+OPxvxrfY04i+7YPhHLtm00D8A12nmbUz
N+O7yjnEboMFNhRyQq9mHljjhc6Rbkvgc3zSKy/P3GRebaXMTSr1l1FfV7Q5CiHo/nQAQNU4pa3s
BJFgQZc6enWT70Y1Cd02NtV0TprY1vPgdoU8dSALZ7C5n/j3PCZUqJ/0VOWbm9f9BilG2ihFAgUR
veQ/b+QhZe9Zd5ZSfpZmq2/aEjiDeHhwuI+xytLz24aqSh8kVGuhlrnGQvaQI6U+C/VTv4qLJuqX
rPvFzvlQS0dkcf4L7X41oyYD61GO4BsDFDxtECnlzFWD3LdE/3enZmIv/GPM49z5m3tavlIZYVN+
kIjjAGj+74ULvdaOTZoaL3zCTL3qRSrlNJchE5OeDIOBvcdZ3jLF4fG11hMoeVw+kMlRgyJoA2+e
vprjTo+zAtNAXqimICf0zlrAE2zw1rbKemKQADocmo4EVtSJnmqA+SAtk5fP3KmeCGdIN1tnLTbe
krc6WNKStGgnsRcD6Z51QE/8FFcL78eYTWudtGyVuUBl7v4wDk0bIG+z99VWNkfjbihINp35rEn+
pQJRjPhPMupv4lV7wLsuMdkY7eCHALlENYuoDENA5PPFJCKpdLsiuEaV9Ft+ChmNrLniXTebu7TU
94SfwFdcDQ9QOy0CAAGDYieu//PwoLHoT3DMnkcLxiwtRsCk2NUC5OV7KQixsiTk5eRbBtoCDTi/
P6yHrg/aBoo+UH7xkLfipW5C6W4+AFr2gcw6+/TJq/PnDPAqlu8Tz8SeX3wLM5J8SgtjV4apnGMi
AYEzUORQxStJGcjOvXDJjSJbrQ/Z8+NR/qRFMvlSjAn54Ac3MYNPqRigXAi09euM1vg1cs+Eb5ut
0x+zaR8CcUxNSBtbSOlNigEe/+UjaYhAiBhz7/pV9dbi/rAAd2izUzzmQIZJAT5aXDnsi2FOzEq1
WMReq0MmknryLxU23++ukp/LnlKf2PmMpuHCRlYkOSdfOLCWJxoWL1lKhYeeD1iTslJSMDxn5gwZ
aamLHYNQx2pxB3cpUZgZZ0kbi2+FN2+LxLo2nja/SNayMTQjx0/IkH0WmBq9eG++DdrBRFvBnFA9
ueL/afx36RaQ6NdIsu/4H/rex8dqkk2z11MZMhgCCElVAxmuNisHncCERDpNtQ4X1iull9WA7BlN
krTh/o0gr0Yh0ScUZfQFnMWuc4MSGAS2rDZfSf4P7G2L5HieOsO75ysAwfxAgpP5J5oGYBLaDvin
/mrR1NIfsRRrUqKxOqVwxdxzOpjEBU2y/K+7peVYthgJPnk23QMooJli+fYPfdRKRpUZO8y489pr
2EnwH924EQWePxm8P1icvwKC1wRrOBO47GnJDPbVcDuDph1WLC2Q+pNWel0FLkxqVbzpY99r762/
cauTeHmfD7t+LkhdH5gY3cqtmc1qJBqc15BsH2gP19RZgpzYLYXiQRZ24hlSIoJwduLQvyTOoIUs
OhGC+kdoMGDb4rF6xDhHTsyMbvmzaomAU1q4u4nxDR4NJTEaaLDtjBjJuDLBZLVKpiehe/ww4hOs
oqKGO5HWTj/XWro9Qw0PLi7lculvvPtB8DdYUjgreRMc6xkFqvzE9EvPSXZQK00JhvqFb2fpeo7m
SFIFmha+x0piiPEd8rK7ggUXO9xyWqanhaFOm2z1DDVY2WxhDDc5DE/pwTOKfAxCf3kWGtPCtFGe
U0d3gHZJGlR+zWFFpQCtj8jQ+bcGbCRxtGeVgtz57oMnotNkqC/6ZswvzjvUu9Kie0q7z1wT8JTF
dJAA9TAEM4LhBCbqK+jTeXzCMOCXTiJ20+Z7SC+kupv/9PpRXMJQv8jyr3FbfSS7+9RLpyIGEgpF
aIfcioxQrqM/LQdkrj6djcoXscd7ztLkBE6/jBG0fxjFp+9MxhN4wmgEApphCennPt0FbmlmoD9f
OoZJX+5uvRbLH6kkNRKqoiPHGkazPrO2GzgGLAoJUiBu+tLz7DOtR863NYEajkJ/hUBxy5UEAX7o
VAoqFX35xsPCnJXTjUpgppJvt03zw0y58MXT786OgvvpTO1ESFy2pJ8KAkXRhGW1lf6Yf72dRMqf
HrDhME6LFvZhGywxK8ajBdzPmjE9ifQHGQtqqtyRxYWFj5cW8l+QfWC1W9aXd8UaXB+Aaj3S5Ea/
qu6lFwvODUGmwomIv/mQxYrflA4GjUEP2FYuq2nXPeX4amRJzhQ+0x1tIwePL45Q+tQHPIxNwO1P
rB7kTYMZfKa9pmqOMe6hf4DO+YVDtv5aonQ5M+wpVXTYweARz3u7CVMYN2Vb+NQXxmkvkOMH2GoC
8MUfpZio41pSrNWB6ltdGaIKJAWal+S5iOBwgpHPFX+fCyjR+MMB2xorv+vXETMjIQKmTCxBsiyq
F8eS4Uy92oQHBCKc4nMDfoGmxcIjtOBOQb08raugwpdWJFnXoOJm/NbUoHcO66JXBeHIkLMYIPC2
h+CSGTb6s/3mf3u3ZoRIdzeokI5QiM0MrATp8a2332HD5R6X04NoJHHSgOu11O/fj6j0dUT/X5j3
HWKRbl5GctAGObaLEPgGDQOJoJ2CfD+EDywSLt4Wik9KI7dxgPPW9nHDp+opz5W6Zq6bCi/YRzP8
W26NK8gYuDokIoUiVUqPnYWQMqM9ucH0k7rYLhYtrUKfEV70X31djS1ozURFuhR3KL+3Bdm0cxD9
aCG0HXx9RkhJdOTmwKt59FIEr2a6IG7UTtSjMCPAkD7G2cvSWpXlV+hnyVW8rhnFBgoN3rc4S9aX
PLojdXLWJY7sguDJzVJyFC3o2C4lSo1h5ToKw8C+A1s6LuZpZAcBU9+wFa5Qlu+mINodem8ql2az
Kp9dnoUgBfr0G3dcL018UA+0L1FQACX+3i5CHQuZ/QMWs+Y5K0aMZcFqligZaFyesfXdXkxoG5j+
fA1U+P0MKjE3MswSgcDtB9TZqfA6qcauOetOFzgKTvLG3EWVALjL7TIfvwfY6f4zO3w2uB9njlBh
KrtS56/5c0DSV05RW+4NJULRjsDY8x4aWwbB6KHl+gAZZcRINGrTBDjMdNPJuweSNoHplbjWeBhY
u513KVQ+mWXWQOYp5LHlhGtxODxBlQDhRsPmNxhtkTIn301vn8WxcRr5F10SU+Jn214o3xvwIKxZ
NUrPOJHxVtBgwkIngFcu7HIUSE7l2TfAxhh10nRBIctA2ijOWYLCb5FEJxttQ1LBCEMjorK/Z7YP
n2J+yInWhxddUJ1KeEsX+OK4AS8m6E2GrMp0lN/7/HYeScyWIAt54Sef2Tu4W4IrPtllvKPeGYdw
EM3Ci2YEuvmCB3024haKjfLDxRfC9ZQZ4X324WTGGvn8x5lbesuQdrsuWDfgmnYjgjtN1Uoo6+qY
hmubRFCj2UqleUwiORU1Eg1hR5aBoHdyNP+H0RLaWqXspC1VRFjAkAfEycp/8DsfQ99L1CjPjorz
d+qZiLp8npPuYEsgE5jzs4RT04HR91zztWSsajiZ195Kr0XkthNHbJp5BktVPgxLg6t00kXcl22W
gduXdRSz1nqZL5LsZf0QM59HxSSStbxmM2O8hOlJbsYIpc4hYwX9NEpCAvGFw804KOSKPrFQaBN3
40hgb/pJfQ/rAM6xDFso7BLL/gIwbN9P5JLEUFkwsBgDmM/sWpj6QmLIXxwprGS7ewHlrEDeGrsX
SmItkmQlqpEqGRkegDShQWYy725buU2ZXMZUE9ZJ3TM/v5KD8G3y2FmY0F4qZK0Lsg8ObUsB1m1y
4rpRrCaVnP2YcbrupLhPttRTCJP2h3SlCkT5qiUqjHiRrlvXu01gUQLycNJlfMyQ0Z1pOqB8Qq4v
2/jgekmcydi0aVKQQf8XlNYx/8Ul8VPlWIHM5vhZrWUGU4h242YDf3Ggi7wiGqhjMjlL/wu35iYK
nDYdnpQ/83oO9OovbIoanEn6xN9NvUDfojAf1UMM3Gf58ZWrEKLGnuvfyECwK57QjdImZQIB30bC
3Zgt/WZ/N3+H4jMmB+R6pya13v+hBU4nLWerMZNX6ReZoNKQ76eGwYCgUF6gV0G1VekA3U8Qhrwr
NCF7Nc13FoLW+3AODMPuOgjZFvF03/j1dvLxJebM+flqxlpCEkcRRrtdlRL1AyKNXu7Ny3wkH8ij
TaTfHQ7OS5Qr3zfunvlVdvXhop1fO7P3RtbAQbzz9GssFVs0XBxMl6MS3YofYaAs1CkVrNqOb+Lm
3ksDTkCnLjhh8fBBwOBRTSrZsSI87oXwVI+XorCeKZ9mjCshjGA+sNmxTLYxbokHitPlRGBwFci4
8qU3+XAMBfEqQTGaKupD3wZdxofObVqAecIshK7e+g3MjnIVT9+W4C2kgBPkrhaoDaREQuY900zX
8JDnS8aiD3Wcw6EVFY0y+/cTaqISRiEFOqb2n+cc2peiNuLrgtdadvWvfLX2511iU7VzebLTRHsC
M6zaaLNGE0t643yN2hkX8hNIk6+P8v77QoN9LbJnyQfe+lIPiclsRWBY6btKEOK3oOC7rl0W7wWo
ncWlQd8mEPD57LBwRjKnr4Hwwu3TMQQ2LP/jggq1pWzxrvnL5hMhDzMJkMhKstFOBRMpDTVm6HuO
tNR+D8Asuww1kmVIcTesyMuV0mc/Kw/LyA16WvhSiGgVYwpiyWfotj42P0uNiv7vPWw+ol8/lnWr
1N+fvCAzljOO6QEk3uo0CaX+LViOJSfY8YnTjfMIE9RJREUFfMuKcZB+NEHHylS2g9O+xhx8pgkf
aMNVJGuuLRrMbOoPNn8jYh+j63G6U2B80E15l/TVg+9mJ1e/E/xTmVqyLsWq07zHqVtCC1blfjrs
FRxlq8PrxujpIJm9kdjY6J9IiV1vavW3KIerYT1PrDzskqgDAQ91GjO8RMDCVEW/dEAAIqzs04xd
bUlI0hxH/FCF9iTz11nNjhjQUOk5M15vo0a92uaFkqUx+U6JtwhslVG0wdW6kAj980T3/pS6gZiT
5M5i6wGB1LpDuorljSFlQYqIkr0RAjocHknQm1mrggjJ3zycxlLIYMpSArylqf0sIttZY0yfXJWX
SgfDTalSL0S2WOt5a7p+Eab9+5ZbkrdAT0yDzs1xjroXWpc2pNHcwDgWdycPXgmeVNkfzjbsFXEN
gyboD9lWoWtSaQlu4hO/HpU6c7lpJD4sM1m7aDHJbYircb4tTMWjId32LbWEoi+3Fafw7mkyRAVi
czdFUmz2Ueo0VsHCwX/snExO1Id5agV+q9sbWHbARYW4WsVoxU/lzhNt9MZYdhLowFV9yBv2X+4d
TRBMcXjpcZg8ZcKOLAOBzkrWRWvZYHyJBcvLM4tBgZO3dk5PkAMEi5aJ4T+0jUe6ZO5FnluiDwaf
FkeFn2Vxqqi9LKOeN5e/oyUYesAZXyRC5h46zVHot2X4+gxyCpTMHp+r44w8e8h89xjE1B5EBVLK
I+xc7NSVs7h/MN0CYRCDmKARh0Mqd2aES+cJ5BT3wNhUyCaWFcLSwwuJEMPwZXJM4nBSWvIt3+0L
+YNQT7pdlRyPcCrfKiIA8Rya0qk1yXrVGqQzm6rrdew7ZnU7VaohzV1n/4EpUPWJpdo3TMq4mLIm
fM1EW++H2uDk1GcjVmJVm0ggMD/D6VrEmra+gyDSnF+zr3ORihcl7YPRBqyRhebmQqptcw99A9tn
tbbJTN6cpUZ6aUuiLbigow62InPFMm8G+ssfBcFPKBkYRPK5idHz8AZbF5CiLxDJoCVh+SoR6+2Q
KYP8KW5jAptDh80yn5kx8d9LlggrqT2H8zUWaDTAP7S7FrACxTl/ndK+X60Aw9IiYLC8pUl3tfD2
KfdpJ0ibGNRVcpriImhNo2gJOyr+dDsmoAEubQutyQCmD93yyYNpjau3NZILNKNe51juHejPdxWm
twvauT/QXuWqijD/MJhbJg5ow15WAXlrkcYC3u7DNFXBg9sDyXzfp2qgi9UWcwhsTpzR70S26VMG
Z6dl+giovMrb7MEgJLCFVNmpBMshIdE+DiKLdg66s/LgpDxFcUOubvBy7knYXpCu4MWRJGNLMjFt
TIGD2WqHhsWOxubLDubyFHMWAjYPFHaBC0IolWCYaSyMBplzuxtVU/Ef6rVxuPavprQHxmpHkQTq
5ZsjW+s8gNvvNwbDyYJIWzGhLDPhSeIv/GhWg1cNnxI/dx/6FcqClw4KriZ7S3Ouvyx4eiGVOlH2
K0ViJocA9uRZ7A5nZR4wFrMwfnIKxJpO6ac7Ey/03mkxA2LZkbREWTZtPyW1t8m9+n6Pmr1vh3Li
TulnWq2ujFamtfbStbkWuoGvHyecWMUsT7KBerw/nVMH9fOqDgkiRa+iyLkK5kgEBPlP6vko1dfp
FAThHPm+KMIbp0Y1qRInQk6kYCNj7BJRPYd1S83jsxQ4u8p5ZK5CBx4Jdu/zfj2MRUyH/IlBRDwc
lgxWsgx0oPE9iha2Vat2ofSPVTJaWi+wYGhTLfqRn0Y8Uoit3NZWS10fZKGMXpGxM6rrPWqqTpqp
v1r3sDs9ORFH08cwlGR/ERtwWvj90K4IhHKauz8cuohyuFjOhs12JDni3VSNE+0FCgZOr8xC0oov
zw23c+FMBJCLS418pIsS2MXeaZspQCNObFR49RE9JC7W+2RIMMcMM9GyueBLdwx1n9eMpR3s9qtI
VqhahTJZpSOdwfuWX1V0pBc+NMDIH/aDEJXtIyCEiOJoriozkt1yKx8ccupd5I5swnmRGSxcfy7l
Tfbm+1PRQ2cLHL3tkUInOw24h/3la+64bjijbJnii16okI/LgjsCL4JYnzZGo+GV2j9FcwqKSQp6
MnXTdD9Zy/YjGq+R9uWkhqybIFXoJBUSJuxquH1kMrlK8P0EyRPxGNlBqZnhBezO2jCYlVtNQuKI
8wTNXQFmnzwFDlMzSEgp78ztprxn/eRseC+RnJf03z8bSo57fed9UmTJkzaJiXTg9Cw/fGymCIHf
uRd3qphLHD86L/AbvD3zinPNbG3yJGJL2JievSAyFNLwT6CPDoxG7aKCL+PERNWNJuAt/ywjGAui
AsIuQRDSqeucWAfGPfig4sIcFYIIsqfvAC2q1UNnhLSABSBq1NMy5f4c1v46K6afXk4m36S6YeMd
To7PkRzqMVKOGjbKNH2xsqS9KN5dbjoPMyaExoIj+Yxt9u8vc5WXLRurcWEjxlhuWtcl3+gANX3P
jHi4i/tpM1XbTAh65RQoZ3BA30EzPR6BmtTYxzt95ERYVBTTOvl5xvOMIJH24LQ/RqCAxi50PVNx
ZZnunU2po2IzjEjliu/W3FspOeyZ4Y2/jz+//UhLE2wfDbBk8mRdvLu0ORip6acYrLlj5dHhdimo
2DByQokJ+yEUmFyO/p1Skdskw9aK/WJptLupZsrnagTHVSDLBhfSTOhHZcXN6cClMqrpDMWN23SU
yPFnAPtmPIZmdSBydN572kWpOx6Rth40fDxpHsXPp9TrVEfut2DEgGFFb7ZjEfkaaZneeLYYJL3B
jDnNQL6+HsumV0EDMOECr6M6ed67/nTaSzRsxQ2w0cWzwomU1mavpsodj0AUhspKR4tVENteaNCs
VjTwvWVwsFezuImLbh3keOpeRelzUd1MeBL0LWizu5e4zM3yVtTI4MwVmrvc+r5Z3NDv/t5O3qeg
wcgCa3ZQ6DGtzIie+CKCi8wo+TCZFmccftS6W68PBDSWsLxTPv6Lld77pVPXbU9PUoI1SzZowleS
UiGdjC8s8ufhmNtld1LFNgeKHrOkFjj5x7V7okHZQW5pwxVeVYTId3HslUHccRThQJnm/4HE87PR
Kuzj22vLo4K6gDm0p3yeY+Dj4ZU/k2I6o6z+khLcxGyzMTrqen7wgJUoUhf8nkCubXHa81R0pXpE
yY+n8fJ8Ubw7QoqK77euEfgCRl4D4aJwBg9aLZu3NhtlenaaHCaSgVTiLPM8ZamiBLy2gE8lOzvY
/ZgdIO0NYBz7lumTay8QDxvWuE4Of14CiQ/VulQ8FTp83qjrve/RK5ZfZtM30CywlrzV+H9lFG4c
fan3cAY56bwCQNVYbWhb98nGRd8j79xo+7iFG+sNU73Sk6E83npGqK4EYyRYfndQvXVN9JkBnn9E
GhnJP//IFVfDIFZWWzliOybUYSAXSaPFwizVY6PT4dF4nKPr4VukqczBVGzNmdE0I4271CNlqykE
91zUoadQx5lEgwmkJJeiwMoE47RtxtloNw0IjErlJMn2RXWW+6zYM1OmixqlkFHI1ElqXXz9QM6t
FAhoObnRGAZcEDdKuVv6XFDLgMLNnurGQ7pGMCtvsCu3twsnUmVRJOdou7CdS58IXn/8M9f/iRP1
vbyxf32/uWE6NeAXa7cCbteK2Qpqn/wij5CcXysL4fPQ0CfXpmwWQQ2v3HEEWEvzY+LtN/86khQ/
x2ChE/txonyT6uOVw7VJzo3cCc4JlVayDi3iQbkF/kBUUSaFTAqkTHH+lGeLs6+YSeunOjSjOEQ6
rvoAeZTyMBcK73rU8Z+iHk0kfhm3dJrX8p2KQuWEkb7AUbkeGdWvErz4p+LDYxxTHGYZPaBbuKRf
4Xvo6amEZQoWX7deCDTXZI5jUN5hB6CEGlq95TEr6W3SQMWZC6af3zNTf9/rjJsVAccoRwQ6+LPE
DKJUgnxH3Gwg0KYeO2xa7wV49hlfeiu20ufUc6mc2S86bjOAUK1YWWI+zzXgIMM6UDK8PVUO5lQF
eeapoNoCXk58i8iZcEZB96ilacaKQcjyBAyfA3XgC4fjVrvQCJc4y7sKFu0lIay8Yg0Y/LWBXNH/
HPZ+4gMoiDT1mrxyor9nkcq9R65K0ro4FkAM219scAP/NnERQ03UO+IYhm+Z2iQdeLKhfdrlAAR6
CVYZ1IbBzMiSiOaE1IQNE7qa/USoS/GVtd4LdGNrEwZceg6KC5PR9Pu5cHgy2TiQ7QOmufMTli8i
0Jm1OxelzoPqF8vfV/ZHHVn16uXpMshH0pD9sEwJOR04nnVF1WzLSpIJ7BLOgar3uHnKVLRdOv4W
HDJEmfiGIk93pyIo9Sd/KUwDHJtyXoVytt/vpGgiCJZVccQShuVVpipfqxFy7vkHrBNueMBDndY8
f2Afi2qh+kSh6jE7Kxl+Q1FVHW6mS1RtAMlKIQbPI9RbDqjn13RYrLL5QWDG2UoEpSnqus3E16Va
qtIwlJ4sjxOqAVQ3caRC+USjM4bYd2ZtZaAIu+psr/7mMygu/oV+JSso7d5RvPV/Sc9e0tE9V2ab
bYCuDNC0XoMD5FpOLIe1BjmOBM/wp+Dz7wMLk+4FruPnRxeXmJFY+7HBl5bKB8WO/xWXGxIBGse7
RZxA42bgc4xnq9ZRkqkzQsOIltrIW1ijhRxKrdYBN8xyUn1Zr6UqrO5BKDJUgdFHOUy4c82m94ja
Pns/YHNOcJE6yR77usWQPO6fac+eSuUT0aAm/PiVZNAGwcVFs+NsbnRkzwVol6MmkzIknAhNHClF
jIoGLxaLSjH4epyZHq5R/0s+eVDZAz9trTBEvX3ZRQd1wmavdoqx0eDlWbTZEeP4eunupE8BLKEC
xPT9Gp8e2MI/5pgqs+K+de1nv9M0gy3SpqEMnB+tJNELfAS7oN1v+mORkLskZRnP+sTbTtXzrQ1j
baWtlzJddEmvPqxppR46DNjawjZSSWCTvRU/joR8Bi21Etdbj36xd90bpx6HEZFuwojoj7zRzEUL
9UBDT6QKjupI8AAzxmUFW4WCV+Y3FPPpgwVkv6sa3ovgCmEmOBUBSeaaye2rK1uLnEch6YWuZ1+4
eW1Ls+YEkvWhVtIE9sMIE8oyNmxciV85yinQqknvWrYB8T+ZxcvATy4ArtPKT1QuDxZH8TvPtQVk
bH8DZwGbEEepkzZ0VgI3b6J+Uem5r2xSARRg7YQpJLDK4KjY8LbPTO93jAgNHqDVJhTJFTAZWaFN
hSVAYZ7mrBQqbJz2lr5OTHFHMDqdIdAaRcv5PYP/lqn/zSvPIxrMbtEOdaufwUWHsWKUfSKw5IvK
KZ5Sihg7KyrLUzBk7PJjXobhvIELt5mJ0vvoWe5FJZWGUiQzNB/ZLv7e6OC+zJzdQatJhaneaiJK
wS+wi2K4pWB8Rt7aDwaZjPErpXhYE2a8kUmNo8jxadOgvWWTi0rqEkL3Llb7Xh0JrCCwr2xGp/sp
FS37Io2u8+FZ84ISawXxuytMy5UIRnHa08Gg2c/+HsaPwksl8X0SuqWtDIh0FmH09vsKre2x7iXh
H4VuJm7MVLPdU9IYg2rI3bnOYfJbDGp0S68UN/QSbxfF6MUtA5TeZF2gFFiokatHfU5NBFA0YrKb
ec7TbqnNMLHdqrmcNn7vARiq7jp3Ei/mXAmab16a26P+WVr/e6IXvvn5plZXC3phqjpo4yrblIeJ
i7uiPKwMCXB3meLIuyFXOwc8Oys+fhkDRuk+8iF+eab9YZjjNYQHcRSd4KZYUIS3ibsFHHjF/4bt
91qECxIqWmh2tjYvgMXJIzmTocJtGpuyP4xJkkkaO25HJdUjIivsM2KpAylP9BZtcufLq6rGfpie
6UNo9urod4oyn26CsabWjOlM4uvIqpaT4otrMp8Ta5vU7O2WJqGfGoZt/5CBqsMleoVTiDuLxgQ8
NY6bC9VUDY+XEqaY6M6jSYZSksLUPLdQTA3KtfwL42gYJVhOMmOZComXNQnUSkGE3nzSuBIVXj0H
u+6o3ynskHBfHmggC+Uve8xZ53n8TiCnBi132zfH16aNof4QdM/4z8ItQdaOgb8wJDixWqaTeEUL
d986bLbHzI59SY8MIo95qfF8ocPFqmkMcloAngJNXy6+u5WOzs8IbLn6RqZT7DrgwJCYV1BbClyy
PwAEffulM+BLZEh32AzF4IMdstY8qy0DkS3O3TWrpNQNOOjYVwPnR+kt7vO6jAzLIUg0QseVYQW6
8wZvsnHcLtwwaHvD//0USM6J1aLBnnOekHCu4JurGFh+0A6kLWCbumaGM3/Wmty3R+snZSgM+mMc
0cfGaS+wjr8nIMOpR6CmmWsqIymKfTHK8FCsrviAZxGk4HLxl6Od9GpPkwDDgUkq3wU7eKG2XZTO
ZVdb+v+YXM2syYmYdOCWEcmM10xNJJNfn1Y+W+Vbe1BRaMFyrZO+HwJivcn9JdW8mWTBs76ve0Bh
odL5enES4mlCD6Ta62YwmJf6E1JygCYHYdg7DQisGjEg+vQjrfd+ASDOGIVa3OFszu3dXDMdXhWx
a3qaPciksngkcdsVTD587zJkb3VvVghNwxtfShLfGUVuC+AfMljFO1EkzwGS5CwnZ75d4Gbyq/Qu
JzHghGJvAAZRWp9RVc5hoiZD2nA93OfcedEMTGJ1BTGHaQC2Lt1RzYaHZ8CCRZrYZMgU6ZJERIdh
GMBYh8k4xAL54vAFR/7e9LXMjuoTv0Xpop4AfRigtgIlZWUS0yiScRDxOSVL+h3+5Rp4WUFUkDQT
DNJ1AAWLKOsyQqrf3gTe8UKgz9sXKDxHjgWM0kImrqwxlv45Klyc+UsDU62y/mqgdO+rsim7761a
d5g6f951URWXFWjYcTFBzLMwpGujvKMYL9MtVHo4j/AaubihnLGKAIy8Ddsr9k3AeH5DNW1AR+iF
S0OMPCl9dTS66GxiG9pOGFLsbPte6Y+ca5AaPAb6eM4jrP78LJr6e2+p7ZlATKBonrU3TCmoVLsi
OgMPaJInwud2l8ECKL5oSKkzTwtjxZ8HWCt4fkOxV/oM3TXx/jhRD5YP9HY3TzDF5M3BYpjbAQyA
juhkzi8bv51JcTkfttqzpjPT7X3+rE+hF7PtKVBMRyf9cSIDM+49GQdwrlmDz7V4unnOqrPeNgYg
/YO+vm5JGLRPr+fNLt2NGqqJSy8frL15Pf6unqiA7/WJwmiN/AhGq9mt3IGu25QBe0iEt1115q8W
SQoa8nDmTbS3LpFRPIJQB3Lrnfa/nxDRCBdu6rc4pGaPh7pif2RGbxWkoPN6EkFQa/R2ialFFYQN
X+tIsGqDQQEEl5qnRFe7ySH8tQkWMKol8JFdXxajD9JPtCZGCKZCEe53ZyMEfAsKIPmibaMrSRlH
17+7Rn3AsmyfNywTrbXtlbHZf4ymeXWrN+HEGbjL84EIX93fhOeNkeSnkAEq1CTa0Rwcs6D3i79z
A6kyGvJE99vLGlodBIBdmhTKIaQAqFUe/RqmaPDE4d8ieMXLHHXWPXk1EIIwzcTk5fQ9Hi9UAo/d
a1UQh1yfEW4KI5QrIhptPykzvepiNyHoBJio2YmLDZcy6m+CQNOTsSZUmHhIRqkvRcKS2PZZfRWx
HESIyUmNXgG3blSFSYki2myXWBCx790ZpbJtAqf9YHgV1Qhjujr1rX7LtuoRtFZKWeZb69dKI0y7
sQrhAg0/FpCVAbl6W1cWC08MYinCBWj+dNMnZUFE1/H+SKD8mF3ZAgHsusnMeg/UM2uWy/Juc7Es
YuRz/9zIBb2iomhHXmC+8jbv/IAnNUAc/9WUESqQMUC8ON5OG5vdUZROsxnlolc+U6EgIRcvF4vw
0c6F7/Kx13vCF5e27dDXqrTJo7OYaINjt5wQcYh3tBrulOgLE21rvGURkjXR9JXFVpFFbH5wX3/S
d/Kmi4n9BlvULJkCvC3pon/+0EIeHOAX/HHcYyG4cVnECO4qTaNfVknVVTkLjIXIoPJs8Kwuwfkg
aDIyhdJvPjXUh+KJ5WuCE+ikHeYybGTSeB0kuf6qhUDv2BdLeR297dVC9dv8uqXumfsg3+ueGBti
D+vXhmJoczn1abyjsHlBzH1Y+m2/0vSMVvjDij7m7NkjNTjtDfvb9BbYyAimHHlmJ42v9V5I+lyE
Cetx/ed6Fw7odaeqDJE7gaHEpBGsGbvoNgxA7MePwsxosHuRi0i0h+MHhVMHtY3/JUZUx/4xY7sJ
/aZZL/iOr6NtHNO4K07S5wl2ny0w01/48JPazLySSfYk8lJAaac1GtJgvMY3Ryz6BZ0vuujeg4kU
UuLFFQXMgr6gMuEQEnRWIT54WIASsSZQA1a8Z3Fv7DxE+2+8C1k1mSBJuaB1t8lrbVzkrsYv4M+c
ct1gn4VP0+2lF7hd4JtGHQxoD63ZuXxAYW9u3kG93fcbq7LYS0i/85mQojp9pxHgunjTIn7BruUn
uKZa2YsS03Hu7nfI4/lqBKpCXorvJrvQuTOcM9df0JfN8lrEHSNX46uctd7H76qdFvZkanXWv4LJ
NdhnfJS6QlM2ec/VBOFKDmT4raUovHX9r59O1TPnzKuqorQIdwLmh3SwQdSG8qY5byAexc0A8zns
HnFQRXrwxOUUrOPdcBjuTaU9BBTORwty6994r84ufeSPm4VH+SWO9h6GWIyJk1gR3l+8eFLd6lHH
5En88evnZysdOhY5V0Hn4RVF2HogUmjTIPFaI08pAZhcOjxbrK7X9vVv7FZJ5SeEjXgyc1gxi3Qk
taNAg2AvIccUb9I7ZVUa3ckNMbC5/hhdfgEnntObJxziE/mvRTGyHeOlv4nyB+Kfba6lRZ0DZdxL
yMj4AQGZenufaD2E77ffxZYHHh7EvQSryLuSQRRRG6mnk98b5RLxbqLOGaGr0VAei4uOgGl0ebrS
C/Yhg/ITH7UpdLwNcqQfohiuIHsAupV4pGgmkCH3kAg96dh1Ltf0jn1TyoAAAC2Q8puSRcRjVWsH
faziPWfTxM/wFvOvyae7CuhI6BtTIlrIbfmfaPjIzvHTb3sD/0qfXdbKTh5tBbJ6KnDMwe0lUx1M
pCM4L99PH0FzVWQblWioTdar4ii1cK0G5+HrduVmtnmsR+CZjkx6a7UfZtmQfOF+24b5IYtk0lLJ
eQO4y9G8KymwxH9kAKg+0TO22PXEaKnaycxwi+bsu75+b8JC2/u3zC+mVA2O2ImEln2UHJaS7SxC
wr3mPf45nJaO0U7w+GTSmHDpg57pOHFH7rsrs7l2RrgpKpPiouy/XedyzNE1nvbylTFyHIx6qFRX
AHX7nsB47qBXg+AyPuFlohZZZxHpdVkM8M/DaBEHx58NDUvpEt/ww7P3io/g3y/GZe9S0WQ7Rwto
Xtx3PWjwqalLHc/UGiJTi7lm4HZPKe2RoumumFkVXcfQvgfWlSKoYH4Qc2tkSuR/1TPbkWPycEaN
TyPXmUQ+9Tc5lg/zfhXOmGCLIAz/lnpG75V/z8cOUS/yuNskHjNVU58+Kiq09qfVpJy6wzSyTAhg
dniPSlMzSMSvzKXA/nXxRt+icWtPUhS26qLIgPA6PyvXhVIiChfLrUCLme17rL86//1397odK1qJ
VOL3TmCeiSx8ou9ne4k8jx9pcO4cKAAyvIziUliFhASNnpu8k0N65CES9UloatW6TlwuCrAUoLn2
CU1mJPjF0sWU8Gtr802/MJW3etCFSEjv7oHXrAnXuQMeW6B7ulO4m6/uDhPRAxVkPBhbxzNQX41Q
INBSqKaOcANQ0UKMWmgzb9bm8m+yuqUib8/WFjfD3wTrb5vcb4VCP/sexJgl5Zv5nVjLQYrEBCBU
tGXaBZRJQI1OLwDnuV1PFsyz03tycva50FXvDL5Dqod1XFX6V+4+o5v8s84+WWdpE7efs3qNZOnJ
7AH2FKXB8IAiQC+uudd+FGJN26KDR8Kk929QNsemOPaDnNDbFL8idj0hblYhC1TYoE6WXKatnAXZ
zH2kw47Et5rklHoLct/33IAKarDhwJ9Kglx7LRlIMu7f9/lwLp8t38RPnsKaODPk4P2U27NuQ+s+
R3sHrzgvJNLRs5tisEkeb/F+ticDRjHoXZOtDIkgcWcc/j8odjAqVz+bhuxS/225FY5cTAppgr6S
KzGAGjV/UiDaQpy4B+9Fb2jlr7BKRBuD21/9JxgFqCKLK1nVfQ4jh+go84B1DJeD/sZoCU27cRGE
fAkIf01CZg8gEQ0oFyFhvLyDEJPGlWdgD+eNJv3dsLD9kWmcNkWqPX4q1ZsHesViVPN4f8mXYeXs
c7RCvaxKr4DQ5f5rPZ6JF1YtYI5vZ+eEMLgS5zbcT0N4Y33vU270ewA3tJ6rI9iks/HPxeyLRHqU
kLHAOgsAqs9yORzL42u1GeC3yl/rEvZaxbNIw3jp9Uv2WppK0/H1CjGmXpnw6s8dSr26UD+estXC
Lz54yJS0E75txrQ2sjWmoJvK4uw/TMINuFhDRwcBbr5nVrpZaYtj7PdA569Y5EpTh229ehrC0/QZ
pkLhgE5Xb0lf4Crbt+hIy0Xk+SGVYMbo6KzDBmez5i5HAbBDkxvYqCOMGZ1BIPBA1imftbEwPcvy
a3ntTs3yo4soqm9zERW+e4kaoWogggT5EyhaSzbQBlG0ohy5Sy0f7cKSw7ioubW6leVQ4ASZyKF9
tfdA2rWBewyCDJb2bDMjnHQ6eoh0rOpLYCI/D30Cf4nsOWDfTJHWOKOyvmbX+1LqyOPlWyrzv+mI
Oe2w4vsfBvl7A1PwVMjzLjg+9+yC+7IeEjSvKAefHUe7MqxwVMfTYKYf+6wvQ46tAyyFeW57bJDj
KwBm+ov9WLeXXuFj2nWTGKYYGEQXyBGpUoBgtBhqfU2WIMYH5QT/zvWj40AmuAqVIohw4ASHSkOl
lKLPDdWbn2A0LeEHedecPEKInCv5256eHzNKwF012+OhWYPDPWS3WksNZgat4mCAIe3CxqaIuDbd
7TaD2j7D8CNS26Cx9UindDutHhiiEwenSPD50xJmr2EX4aDMe++nmaKXSuo2iBkXTtIxh+jupMw+
hSxx97VlzKZ/MfMZPeozGGK8L7Rl0UGI1OAtFx3xfwaj7LdcGP+uVjVMPQ7Q6OyPV0hpPQW4fc4V
o0AQxh6mTUDcGHDlvtT7M5y/GSrF9MV4yDC/6SBxBQvbUjRYIV70Lp7lQ0HTsOI5lCWrB/lLMm8O
kAqBqlmnBjPTs+vSaAqzWR+meYgxO9eQDiV5Rf1Bjz4rmmEroP0RjoKG5h53kvbUX2DcWOP5fRlv
xvpwnFgWVsZ1UyPPLSQRjc8w0XH6X1TWuRBJQYAZeV4D7EDYhfYExMDTk3lOKO2QQg720zn44oSp
0l3Ts7VDTPcIKUtbqrSqO/Xbxca8xvdqty+UJvUc0+ZVOqyW6gTkOEf/WG924Qf0QPsNttgP73Yc
edS0bj0ulqbQAuw+591viq8FqvBjLb+aAaD//XXpDxMxGdLYdj6WXWRw/7tPZPEN6O8gQxDlfiP7
yfIqRFdlnPp14ZL8h1OzcmbykpXHQkqYDCjdRfQ0zqmcoDOlsEKy9DJt9U+jb8dn3WITxn2FCPTA
18TrdxCSGKs6riA02HX7Als9/A7oHL3qcRsy0ADXb5tXnHJcpynzkvKU6flg8dH7y1BwtSKLIm3H
kBhC/Y3tFQsiCIKWyxIjtiQy4WZIrnPFtdgsmEXgHayZP2fKjcwwymbXF9oYB9FPuFUwFFulnJZB
hlBhmmwJpDXeQITdVTcnccSLseKzzCMNgRBEn3+8gP+o9xm9gIxJ36e5uQ326uirqYw2DeqyXpVo
99kzZgsyzFF3jyMVFHiO3PelPV5RehanrcwQfj0auIWaXyi7+Vej8jqn6SO4zCfGzdahcsGT8lc7
dg4pZ11iG5OpRvRkZV0pRh0vAeAwAv+HRMnG4amp2K2RxwM/xMh78KC1wsa7HCQjTrC+PI+oGJF/
2OqaNeYgft08RlZEVbe6e4OujXqh7oj894GHnwOFCj3kuerF8Ucr9fnAj9BWIK5NL1qDzx7lgg6C
kabFz2e/bshfjzUPztHfFdKzxyH2j/st2UjIuog+E1lXV5hgxH7oPayD3Iu2SNlW3rnppD6NVGjU
Y1KaGcon2NpFRIFol3o0sbTgTiWUOoXozwB2ke4Kobve1Q/CfLhML56gZJRi9c/5aFTMfNd/i6IE
szD8XW/DSjgpOXrVUwBl0+zMN2giGPjD9LujlP4S0RddjniVeAEM1xZKPlUcouJuiAyCsq7xQQWe
Dl+ww701jmPN0xkcCZrPpmfS6w/DQOGj3ruch+G4BUfz1wH4AKUY08byjZEHdvx4vqYOd7ZODQYw
SdYPgI2RbVOGUgGz1X6Tctj5ob0rYDhn0E9qeAjKOItr5oqs4DIHo3gGFTBKxcHY6w1x0CAj43e1
cCVQI4rSw6n9bk6MA4CxJ81aeR2Vsko31tuugVh49vpIaNGWsqDqQduBXb6YugqEv8MEQZWzF5wh
JB1cju/blzbX70UbPLMapPudFIgWBKLnO+21udToT/s4XOijuQ9gXjAYQVJlNJ+S1npMrXUXuRk7
8b6prTQyV7Vf3yQMhQIJVSyNaXhkZS4jy4PgjGJD3w/WEvCv3lc0rN1FOrQHwGWnqZylxRC76ER+
6VpXWtoCUmLPbFCPALxO1l11s3ulAjS93ZQMN6FuW5RDjglChLDUlURfpW9EcUgFj3MaOo7lKRv3
7MCbqL/nFHiS94YeQyrsTeIGdMvzN/7tO1eDn9c+quaPhsEvx6YB/vBKvZU10KUBw3SDgEU5490u
gn7QCRB9/yHxkMQYid/ezd8StB4n86lyLi7ZyQgZDD6FvqrRvf3NTbqOzk2QQWgA9bcC4XjdoalA
dLPwV3OOhdqvl2BmCMrNtojzoV3PHbtrQV1ebOCfyh2hhMr8XaXMOleXE+CGVMw7bso95DMKgx5M
0Y9VZUhHysyA0vh/GvJKnhQusaf12F9pU7f39Ho+UXU0gu7wqPuUJaetoMFrgBZDovFCNTjWNBMV
xrTV1v8wfLqJrdv0MdFFYT0iD5hsiD2wXfKIgcJpJu6ZYTutciB1hNdy8SrEtHXyK4oodBoZmalE
6AFaBOzkExL/yVMoS4TVIPeN8U28KdBR8Y2rhjnSQUSp/VNYZqVPYQpPzCSpO1XtRztbDLSMcjuw
iNkVNEvKWe38iOpOKN+GRmacdioFkeDE7KgaqnNBh4JaaZkblnPaNnzRRUkjUZs4+c8UMIEy8/+R
fILTIz29ubrMZ/aArCnDTUuKNhZ0qe56T/ai+p1/8ksWopJaJidpuT2aaWq/cl2k0mD7V4bhaXIp
W4HQubDB5uYu5PTqfR6y7dhQCB6yzB5MDl4iNug95vF2AXGkU+bxBohfCAubTDcTYEdi4Ms3uF9h
FHcsMoGB7ivyjg9jXxerzW9oIoNb44yt4GM2Dws2x0AVH/MqiLsFfB+97e30rt+fSAsi/BEjT+aZ
NT40kXIb4GS6RgVG9lBU9OELahgPa/UUGVi/BiF9XqXf8DKCVnXPN6HDcJQuBqC5MzLsn5LLeURP
PrNbrdOMiR8Pbzq8zsqc1cMuPr7q6CAtZBMev+iUeXO/OoH3k+5kPm9o9yVCF5wr2ihel1gWg+XJ
/Ezv52X7mqSLEcX8NiZn45MUrESlNCYoYCumWAfB7HhhUfPgXXhQoUuwsKsXJbFN5FZSvtpOu2lK
R5xnOkOoHsrPdzdr7q4TXSLU28XajjivWVCFk+pLzB+EyqQpKstrKEuKoBr6I9oSvPeEdMaL5S1q
H3IXkdVvHL73fk8IEmw5QmsAUcwUV4stlSTXgh9Wa5VjWO/MAQEUHudj9j5Yy8vhKmKolMcvnVJ9
AV3epEwsTloNGIFLb7l6z3HIgOyuG4IJZg5blC6f3jOOpP2k7N5lHCf4s5P90sXpF62eUhdmHKF6
ldlm0qIH4rwlgRWnICKAQ8oFCYFcJj1uh5yCxhg8DOIhtb7R5dZ7JAKCiqYSihmkvMC0uJFlG+WN
OYiZmvWX5F2J1OxLSeukL80t5C3rDiKphxVuHH2n7hk57oHwCgmvjfixfULbbpthjOHach6pPbcs
FjhpW9vlYBMQlCRPQIOGEF19+OohBINbVPPt9zs0FJAvcV1f5n/cbF+JYioEw9QkuCYuQpKU/bnE
ZIRd3wuMyou2pboSz9SxLH9cAQktS0Q00MnplpZNBZJjf74P6mn3AgKLnmapPW4U8xCYmtbk7Fkl
SZiaJDaWAFxGLFs5NnAgtrbuUvhsR8461SAtltKJ+ZyNGNr0WwcMDsfJREO4Te1Y+t4H3sOHBPuH
JAXQ0neMUaF4J1JnKQCeb3MH1tma1nAhibhl6o7osxezdrpzU9AvRUTtW324USrXxlipndgexVwp
UPE2AEbop1R3sz5GxhvF6t+I+P8EjlMr7qGMNqD5CUwEm/h/l7izzWekFVQh9J8GXKS6F9SYqwP6
+TJ3ReDA3vbiEyHpaH33kkR7FS5kcD4tEC8baCGGMC7cOqNMT6e5osrOF2aSEf+8V4njgml/MthC
SiyeAZNG9bPIQl7Y2gEqnwJSlX/5NXbENSUGlE4iQycHz/ZSvpAGFDe78jUZDrI7Krjja4CuJxMi
PHpuPeXlSbemQBUdvFmybSnIajkJPmna8d0m7z9cOEPO6zwaNskJY+5sdjKam/zktLSxyDwoKp2Y
UQlCKLrV31iJwbsM9BvYWEXqAsvNmLzTV8RG/Kt3TKz23oa4C5fKI4z8rw8Wbr8yy3jmpwowiOPQ
q5anlOdnKDAH6hBmos5hw2lrWGgWgQJ/i2rFupmyZ/4MLrFD5v8hs6OMr1WvjzMP0AJAdpUum0Gq
9uXODnZURXzJJsDrJ2KAWhwB78vxMGnpn8fPMosDV4TvutC9X/cP+1vaAWRrMgZjEJxg3D0CbsTk
71EgIzsx+v3qgspGcg6Cv1uxILdKQTQeKjbz6SwckjCoQJf3BPauioDtbDt4HmLpjbQ2K5aBOhO3
pzIz8DHDLDaX2bRNKcpv6Hq+E83nsLwKBqCQBO3rc6VIhNyF3BUdsvYVkPp+EzQYpxSnrP9iJAOK
rGzdauKB8u+/rGITMJ7Vk/CztuR96FWnRY7hRMCCLDJugz1MKkoJVcwGvAekm2A3cyOAtWGwZSvi
Sg52x/oUCEX89jc4OS2VP5uLg6w4qsXi8rfy9S13jdrDtK4FKdSiUHdydeRLsSUVno5eL0SWe0xo
8igGKj8pTQVhaqqGJ1XmozjV3DS2DuzQdvVi3jLzs9+Tkbmn9TlQsGgbs5b+Zh/neqZdwLW/vb7W
vVHQYXL6tYlX6eLnUB8Xb28IVw4F/WoawhbgQOArbHyZPGKQ3fJPDlCuCommC2gO9RlG7EqKCbnY
D+og0+G+niAED3KvqrqHUTE49f3RpycQLTuuLv6eY9JvRzApjruzdQPiBJCxx/IcJC1HKhPPTkYj
YjvBLtaH23mPHSSka2Cq2GS2nLeCKUclfp7CtRK9k2HWlUQp8X5XumtYGYesDOwxVuK+ht2tCM5v
YgKRfVXRKluHb2lJi9UMPgtmuaKlggZ+UsaGt3ygz86+LB3C74n7MlC1+QdqwdLxyIItkFHSwU0Q
CJ+jMn2qTWJGNjERMlpjzwdQ8I+OT9jKfdWq1yx6xY3guR698Kpajt6SkWGlTE20lkLWgzloNThb
0fiVopY35p4jPkT091GMI1lLsYSVUijxwSiHHHXYA+Po08PUiR32jTrSExO3An+udlgVs/VnbiY1
3RIr/fhueFQB874kLfVEOMB0RSLsHsa4sOyWXpwaZbJR8OZ6pd6kr2qD0z7I6MflnWz77D4HhFA3
Dr2bGQUjEmvc9Skz0r5AiQBAaXWire7vS391GK/q0FnOcgdQrZZNJpJ9nrZxP+OpTgFAi8j095TM
fI+D++U1Wm+H1ZfSYB7WufoaAaF/Q/HKbg7+H7JKXcefZ4Xa/62O/4aSzVNVOLHOTIuNihR8egV2
mrULNoBoymOWdqM2pFz0QjfzGHVEa4saQGrak5pBjh7yiFLh5aKf2lHazeFUOqQNEHKfPa3kjpM9
fvdALPGzY4n0dn6pALUwt3dm8NwNDQtFhBkWbj7XbMS+97p0tfkaX8ts9w8xAHOoqcshCM1r/Vm5
4VTSBpGjQRoYD1eqqMgn7T8nlY/+3Cnr9LBFBm554HCA1DyqKCCMDUlHgrXP6BLvYa4TTy/UlEUR
bKYz2pX0Y8JvbiGoBhApP1nI9krvKis0wqW07Vg+N8gHeyrTEvZjtIRlbG25DlxdysU0u9zrlxg1
GoP8AgbIMcEenOyba7OklS7jiucUC7cRhhBBP2/KX6m1BMtkOiTuhZHJLfeF2/pPJZFJZ9w2ZV4g
dl4g16BV6kxUL34hVphWERznNZzE7i2YYlGOeSmR0lPlry47Mh3whtmEhGYh2b9FS/WSrDzFZCwH
PsrkYv7LSryLp+29SolLbpryEVdOl9jzVZX/eP4aBqkfINBJhXwQncokGm7+a6nT/gOk6zGmlgMt
S8AI0pnN+n9n1tk5q16Xxb1i1mLTpgqKBYj5ssyKHjL15gr7MvcbFeLUMDIuXS77XFSlpgyuTxd+
dHWGVB5bPXLuDWxn41Az/ftJosHn5Ms+wBEMTy2mxYo2EFeyW6niG45+weoTrgXcMQkivcthUBL9
EkqdBaDKks2bh5oAB9mxiysfi5XigBuJzrKCxXIV943Q7NIh+vKREdSrFek079+vDT1/THEFxqbt
Se/V2kMgjInv6DSJZJopVmaFJuzEXMXw5DuMHc6NcnSwJRKh92CpWoT3dmZLTZGpFr1EQG005bJH
iIdJndmzEfAry9Qm5Fcmz/ks9+Cuo+EybhZR0KL4fHHHcqGORTapmEeUKnboaYweGxuzRVRZoPmD
ZcDQ/0KiSNkVD5R62Ml4NzULDISPMzG/BdfZ4r7assBIIi1Iz3DJ0f5IlzsykmGU0J7azak28xQx
0/CEJMQhEhk2Uqz+kgjZqVAtiqakYO0LowcAFvJDRl0MywdXchW+xbl7PY/jmjjH42gHI0MofrB7
fgpvCG+BRq01B7G/lik35FlMEGnGCaNdaMLoFTnivxxdQKvYk9Vytm7QDWwNS5MIeXz6R2nNp+lX
Z3eIQkHJE+y1/7dI4GzpHsEr0UmjBG9w57K2J774Spx8G0rYwsjAh1bcbiHNU1+93zxBiaLvbwR6
qXT4MxdmMjtIhxHfoL4d84nDX0ZOZJ5PaOw/gUNm1Bo/0Svi6TD+L+eztmu1qw29pFiJZ73NAOIT
cs+vu8OziWwHBz3t/OYlf6Mf/34clltQuf3w9lIK9pJKDPDJ/vw4Wr9buS9i3RzUTfpYAfmfDuC/
m7bKD8VdRoPTn9+Mgl3XxWQpZIZSlRP4mpIIVjuL6Hi0kf4X2tixz3jD8v+n48Jr9MVLE6HGFIkl
/lCYY6FooTXs6+4dZwhNGPxcgsf97KIBy/vw5wtXAIvKeXpi/E0nyKTQ5pltvxCfaifpMpwWkdIN
3HaIIdtitxGFemnVmJRf4zoWmt/aQnU2WvPP29XiWUpazRmGsByJs4aHBw46oJgFYlM8I0/3nhwt
ktbmwXb1s66h6wmmP1BfxlsffJdplfG8j9TTa68vK1k7cI17oNBvWspSA2ajM/2HGeWEw1zdvwdz
2z59/dKiGYUh8RiKcxxB54op3DRi07bjNwSV/fwvPZrNBNqvfh2B2q63j4qFUhdugiDhzg/0bJlt
K9jYJydaeLWZPgHOqbcGCwzA8Y/Iudk10eP0gfIqIOYx+EZ97/rnia3+gsyTRZqFSNG26+O7EgFm
ouHvchRe/Bs8RnsnMo16Yv7P8/ayhP/84qncqRzbk+ZLleKjXz2dwLpfbWQcYIF6TlmOKcTqQyAs
mmJDN9998pY1gWbvpCAg5h1pVPWxk2jvfEAYEDlFAFgwQsuKY56a6ojlQnJFeduCu1LKLwwfMnu6
t7vpzpFHRhB3bh0S18btojAUbui2f2nZMzW6elXyaMgbYlMDcZ2JkTiJ52G9PUzqsVeDk9FSI8Xw
h6oKVsqrD+0p2wyh/aW58TsQaGK8tSmT1P4fmCPohTp4YOZYCUqJZtwLGAHXzJM5We7YDjnvU2ou
LG7jtqvbf/RgkTJju6eoHz1uR5Kq1Ufms5Sn5L5h5RJ2b1972yoCR9ksRL0Qp6i2ZhiyBJtb+2VF
ey0C4fG0PqLzipiV35PrL0KA2L2VM/tXNP/h2nIFIY1YshN81Fh3RP4jPENRie/sCq8iw6Wjceev
klwjvYDkXaXKImqdQw3tWTYHSVwj3HKEwk7G74TlydSI6PQDaLXYEuWVnElw21pxlthjMrQxU+d6
ktZac5plkuBoC5pzixoimPGtFipBMQSE5L2uwqeRYN0ty/RTHYViug/TFuHnrOdI1NmW+eryfZm+
lr6/izifr1yf/daxJAKmabTepf/pYcaxbhw+YCkDUAWBAJS3yk7D5MhLrW3ssrI1JhP23hQnGHW4
CLlJURtIvReAl3x7CI1Tf5uYr4iplb+nJCigbUfH6RBQvFg/riT7fetzq91si8+EJMCix8b7fvzT
Hnwny1mgWI7E60Fh9QUV/V0DyLpCIHFLArffalXg+s6IefUd6sbg8X0VkZseEvdAM3ibMXj0Dnv8
g7VFYCBdXUzHUs9LLWf+E3vEC0k9YOIbSXcBTY8sQwUN6v63O3Zy5tQPJRTH3DZUwfl8Opl1UmYh
0mVzrww0LJ9qg1sbYkx9y1jXjsdEmB8lDLzkafPqHfRX3gZ4u7UQxnY+NtAGmedNYLezqd0UjOuH
x3L6SwKZL2aIV584t2x495HIQoW6txL7zkW6q5k+S7RheF+vDRVyiP3Xr7CI3FaJMbj2nE4v3Ch3
wkLjaAqsomuT30IzU1LP50pFYXprh+DsHxr5WvRCHzd713/AyuQuXzA3VxNrDSS227Wq8LI2eVjv
rbLISsgYwjHFppGjEEcruWyf//FyMEfmUKd2YQfLEFNhzhMS1seArsL2r05W+IMJXgIf+OMTTrVD
CXHk0IzFpAiPXRNolFWWk1mwQZE4qxvsJk8TLmNXK9Y85NBjNhoj7RujonytO5d6iyldNHNpz8nh
GEiWXGso9GC1rSoxu1QKC64ZuggDm1vwjRMHotSVnVwY4edhDCC2IAaop0XDz6stYOiA+k/EInCW
gpIQCPj/yqK6pKrTgOimALuVip8v59WwRe4kxxN5QYr88VDb/rD50GwUoR3MynSKrVmnFHzmqf4H
u/XeyZ3YsL+VDmwNBoWHFD3MRIoue1BrNJVrFRqO5wsfjN0VkSw+MLuE8d9fpn3u0fjv5WfFx4sZ
zUAbjbXp/1XzvbCqc7Z1Bze89majYT8VOqBjvwow0S2evtfJywDuYJWoyd9gFxwDvTx9MU7GV+xJ
bgy1S4660RK5bX5+2idhTI3QdxrsQhtGbvuVhscUhA3aE9aG278rFILRmbTJoUn3yqwRrFLSE9yj
zdo7G85suyc/D2z7Fykvey6ADqYRP7gEaRoqP8Y0TbFqK/LMJ2nIZ4eXzc/sD/LZCH9Cf70QfFac
dwWDt/VoybDlP8W4uVD/sbACQ8lnGU0hqewxWaNAQkrU9hewm0NZC9dh+rVa9i3LnUGvJ8tzx6QF
Tccj8vDjXv/KTExOCAIe6oOwCJAEI6uLWWBf8Z5SUwcV9UxWVjC0M/Aho3uH33JfmZX15pgaBiJH
yaMuJdQz88WGIEbfk1o/shM8y7e/UcYel+PWNrymL2NvPxLd1erlpkfaSrffwsNwnrdG8AwNiT0j
hC0elJO3uK3hueB7a1W+SqvfUfWMc3p2kRV/2Z+sKUG31U5a8ipE8UBWeFWzVZT0cFAsCg0PEpF8
sSAVEAI6hg9NzssXg6n/XKlCOnnmZ7Hex1+9dlhWYJKXPT0JJeNNQIBhxlsnCxjThpF+nMd2XKvu
hX4NN0J3CNhcaWiEhGAj2LGlJJhKUH0mie8krveYd/SEGF/NcQHp2l8r8pNhRqGy2wWltOhMuL5k
qE8HG0BgegE1XgJ67+bLZ2CIp9aGwYDFQWPDbgvPCL8B/TgXl6m98MQQbmhzkT48Kdt2B7/3fbgf
wtIYexKIc/z1epBJ2VUwaG6SZ4vRi6Hb+bN+ovdXVOYSrk8cc25REM3Wv1u4QMkHwGL4QwDsgHmy
Mn3d15uhoM1I0gMxpfQP+GCZhEx3wJIrZe6/ks2TamVhuZYXm5bMFHGL4bRr34SY0sZBPP08yAil
9hpcyq3/l32OR7p9M0RhwvpgMDoiecuKzsRhvue0Z2DHV31WWW/zKcwNy3rL5Ryp7OYeZqSTD7PE
n+cbecuhKJ+g8oSaS2AskJoBY9BxOy91hnriEV7jP6YxsuThZf0xDb0yjFM+WAr8AeALOTgpKC3Q
pfGM9yekJ17XIyCArGnV2kbYUe3SOO59E9nP9hPJHxgdIyj8k6RewruLWVPkfhYjzC7hpfpiUoe7
jyWKBZCvZvzVmzWaqnJyjqheloeqDeUjkPz9RL1vm1u9GIspwRPlHPGWZulTI6v4BRKZyW/mZkzk
u2v7O1SvrL/YLfi4LqXpmYGC07HWjFMgOedVXc4TGmcNBvU2CB0HHLaiwq4zI+/kr3ILUVhE+41m
iKShtAHpRU1egFHnC11r963u8TZBMxWSIZR6KMjdbdlkctEUmq/5qDZy3IqeTQ17tqx2iymwtmGo
RO0wJSzd31BHtPElGTMyaX4j+XmQJhM6pzsUPfGGzEDwW0tiQJ7NXFfr9mEN7kjhfPzB9/pb+MKg
9wmtZpzsI/TnIL0dm9wmCR6puC2rFakwUG39DdRuNlEle13I/HRxydgpnLmbpx1tQ5ahTvb4Ks2z
gVjERrxabe3EbfP+AZflsnAZbSMhmWq8pPUYt69pk3NX8cqK+RGhN7pky+/+5VtbGHb6OUK1ruCb
o0NiMdyLGWXPPfPrYn/hjJQISBMLbrAKOruukZuTU7GtriZYxiu/JhO6p8JxCaXJ9qZMDRdjpNkm
5wJzE+1LDHIm8N/Pff58hoXSX8ogaB80/N3xl8GrQgXic9vrORMlVIxZLByzrxpDprpN1eSlePxP
pToZNqAkb5d1Y1WQAGNZ1PdAJ1iMkft78Nje9WxwdgvC/46QNsToRXwcOrohqFLGdvdNTRLc7PKT
iYVJALSk3D6ZOHKgb9DgFvBZ4EV+ZPVSBWXWne0KnvKZVGDbsuCvaYI3rySutiPmxr4IAwJXWznG
8Rnh8+pjym+GGGY6GIC6wm9Hw2OGJs8hZwEvLcHYhD9+9ExYEu1Oh1mzl2zDtfoMICvgm0L99ppQ
9QpeP7dybRjBHbELDPVfy0DNtbl6ZtRpqL1BtrhPjP+AJ0vnQa+n7g0YZleKmsCOm4jDMmTXWqsu
LvAm+qYQpWBVGN2SvqPicxOw+FuJm2/szpQVVpeNSxiq9hyrqfyZH2217JzcCaUiZhHdpk6USEoq
NDOI61J8Y71hIbyYBzMqLFDCGCjNurnEbH5GJCIxeFnYaXk0ZPrdJsVTqGh8/wRfGWXkJDNiCsAF
XSEaXhelLh/oMXsZx/k3llw5KLQNqIi1Dw/D71pwcbwgmfJgOOeWUIIarVpIYmnyYve9a/VcbCZ/
g0IogNstHXgxEzQ3B/NrRUbYydr8Dv78J//QCzufQvfT2P8UAvyDH7r3CnslyA2r3OLc9JpaHCQg
jpwZZvps2gxf672ftVGi4BdV4vUNX5BnlhZqVXv658RT5yg8zP/rGEm9nR1jBPT4tvJcD+0roKO9
tcBjKxqfyhlTsEz1MCBtiahCQBMrqdn2xotVPdvDWVtxnEzEVxKf2nihpuS1yHCFhsRwu1bJ/NAl
W3nV3bvc7kCN3QaDfypMc/SCSYVptViO/7VWnSXm0XoWIIbBvSbobeY9JJQaJ9AERNXHuBYIvKmV
aT50Ek6mh4chRnpRqqTEDIi8wUUa5fTBw6VZA7vIQI2kDwusC6Tj6Hl/olqmYa0kakdSq/E9GGUh
ydHadIQvSs7q6Z6lRpmI5BGMgf70R9fc+56e9A31lKc83tV2JT2/AT0iRYjQ2Fn7q3Av0nZq6J1G
t6ohhyDwGweHOE5Ab9y++es/pVaA/O9mFNipdYhvS/HwrwVyize1+lEwgO91fUJaGHKRwQ3hxGli
etMyuJG40bBHYk8Wj1FQt7djcZQ3se4QmQBasOTXapgSCFc7YfRs87H6hjw9CKnvknqRCF9fj5Zv
RsG+8PNDTHv8Q5wHdvVwqZWQuLq1OSiwOB5nLS9AX/M/YheKy6y4FOwIYCLlFVC9L2Mp2UO7Pq+Y
2NHNv7hhzyTFWcbbksI0EnGPLwWC8G3qQmuIiVqZYzdOXt2lW0FZP4ZiOwk3KD9dRtr+yCjeWLM+
ueU7TnhOIMJ16kYQ3O/trDbUFT4X89pcoHRYrF2bl4FxMcQbs2PisU+pFYVyd40FEU3nBmCvH1dg
s3ENXweg+Arj/3wFDx014bpdK2XHllax2bKODmo+eL1xrc45RYaEIwPOToy/n8c1P4Ksk0Be1I3L
KkH2BKcJVksgPLoZfJ9zaGQvjb7GkwhrabiMl3uifqcWF4GROFtqo9LjJB6k5x6RU/khP0rF2Zyq
UPb3T9KYg98RnFh3s2W6b2IiAmmmV/RY5NwiJYczd5lGIzdiDbqcx/BGK/OtDHDjMIXXQqX9ZyDv
loIYJ9deKfiIy5fdl4sBkPqXm3BEsSen5J4uViveiLgfakdR2CANiWH5itRbG21H9aEPLkK6vTtI
yMcGd63awCGdQEnfrAmV1/lJiQ/C3IMse/T49Yz4l8hklGKgCVBbEEjLtfp2EHGzRKbLDEIqJaaa
ttmNk1+BuWSgNsM8EUVUiFtSwbhe9NdruyKpoZQdEiUnI9G7QAGCxrZV2FbMRwrcFm2aPKT8JwS8
Z3V9x74ME3NsH/nkCh1Ga866EB/VKqz37vW6J9cktWolpD6iQY+K2bXEYOgL5T/Rb+fN6Pg4mdO2
V+Bty0oLiWoIy0Gn83x25C0freHcHkDIrdS/beFoBHIRCqgXvtx2j8Uewki6f9sNhdS5oNj4Ub+U
c4/Q5gCdpx9a1kULHZWq8DBQJ9eNJbXKDHpKuIdUok1DeNceXCCa4YfdOLoidOHaOsK+NVv2Ab1W
UpuhtumIBZR50/+0hV3tI5wKH7b0/etsP9jLM4ePvzkxl7mMrPAkNddSS1stxioDRNu1dM9Scmv5
+jl88E2XOL/EL1yGRBW93FgEk+yl9zX7E3fyiptHPrtVltrDjlUWLD1wy175EfPnyVcYnwvb6NOK
BXEXOUEnpIjnq1KIuN8AVXbFmbGrDO2XNy5FY24oqluHQ0RdTV+tTR8ERHNs+mFdLVuCiCGUFaFp
CzTLHhXFqUDziC0FgztZUkSwHfc4G6BUF1tbI4ZpjeeTVeOHZUOkWpb98vWm7TNbs7sTsywRx7D9
Qc9gRc0Ic0JgeMecyo09MQN1wiQVNyftj/+nDNE35anylM6DXj/lLNKGxpMLXyFUTkg1Y50e6qg6
QWwW3RYyW54g9m2JxnmCWRVcLUSeWinklGeSkzjB6JmpnX+xaBO6volSzXzp8Ppo3dP6f5kJOgvm
tIcvNhmMQt2BEAlqLqIoUAsllltJWKSulqGXyOdvA7Sg+Bwz2IS1ygqKxtHDa+H+UHHmVmuR1fpZ
NlauS/dKqs9IA9qTzOuUjS5OGaI3KWbh6e6f0LeNhsA2CWvsW35M7JYV0K9Bm+1Pli2221ZbkQ40
F3HzTAhjAZ+eviFo9fQ63jFAVf/YvsK893s5XeIiyctaTX7Qk29rU0WgYfqOlLGp27kwynYkgwjj
uHwP7lKLQjJBJcWOFVS+qQIRBCpqQVjA7VW3N2RByoSso+Z3PLe0RWz4V0su/leyRpyprbCj9HpC
4caLm5+5Zk6Ejs7MImHjt9AfktfpaKhgV4WhiYPr3RTVRVEbh04vvraFWT4dHwdeHrk7vHcpdvWa
zAuJW9xazPrVJ4MP/1gAUjBAiT9N6OqSFpu/yAOHgObtCA1HvfKGrgz035CtnX9mHyIHCgSu8TUS
pSwtyjTT7lUh4kew4Bt1qQ9bxnP2aEtHeaXT858Pmr73zjpU/9Zt//0Tit9x03NCG2J4CfgqwE33
H10r+jYI+wH3nNswe7k8nwOjfLvMPnxFdYatxZHEDnegWaEnbIPMy9lg1fwZrcXM/CoiwNGTVXyW
Qei0blblg+0XON4NBFHyizpK+SLbn3zeNhBc/MJauoMe6F/pjYrf/w2mfZAhnFhMWerWGRDiB4fn
gXNPEGHyewxoupASSvNOSvCAR4bTlZbhU8f0J+sAKWQmLWKto/xuic4ftqsWLZTnDeFelaaxJvVw
szi4gGW8njh8zKl1oxnJ4BIDkJ5durEDk5z9aKHIYit8Qr0563PlXwO+BfWtM2ZaGQrl08xkr+Lu
oIUMlW9shR/eDxLkvZDyDLQQatbnB4dGQKVeh0Px12gcDIzMXQb2B1lO5UnPFlevAMLFLxoof/s4
escCYqZYMoPf5c3NqZcBl9rfbQ1EEjnNraMH/RQSQIzbj0bcQkaj0adKR2Dq6Hkw9Kyx+c/UDCgH
U2huKk+IX+EoXQrst7D7kzE3jKzwk3sVTg0NyroB1sClsM1mjNg+JcLNUqcV4vmCl1n5ylbMGUP1
oq5u7EtvJBF2JPGYFkZvAJ75ae70ANHUA8MfvHutlkYqhDcVkj/QhzVWR3wv3GW9WDMtdk5son0V
v5LlyLZx41ToO805p/AkRya9iKsmOC4l+RN0gTqVYCTp4ioOiq82up7CSkWVejLgMlRxQIkxPE+L
a0vlHQvfI3IJeP4grX30fGDZ0NbwslIMap+E/bF4jVbe74NKA243C6xOtIr+cj0g/zehqNVTqQR4
T9zBc1RDWXYJszyWgEgtturECcf+t6mQhFrBKNXH/MtL+VMiseQC7FFTrs1oHLpBTKcHdDxEQQH4
KCQolEwYEIks/D41P6PLUD+XaKrTxkN+pFadQvBUuRrDjuHDLXl1bUtHr4novA4X6AHCSdCYOeNc
y4Uz9qb4oPaQXD6x62tc7qRu7MhTIws2mKooCrxm48x50i7XtTuMNoQsBFt4dfH8pIdLSnj0EzcC
Tmfn/KjYCtRRWtJ2LPjmtS4NGuOpQU09H6OvSsAzjxmfGF66PzTWE2JYxRAtUjv3KEut88UvzBK1
53EfOjK7r2ue+06NqscJKRAdLStY1cXvxWmGSSfMxz02mVMLNROMgS5jCtk9Zkl1v8MtDczzKoQb
aSP3CRkTo1zWSEpOltOXt1tB8iuBvNjkam+RFxxMF5q3ulZ59lI2MXtqBBdnujogHW8EFKrkGIBa
rwrOIeWeucO9pY1dhMGKS2hnV80iu0YTFEqGJxeSqu/5gyiwQW4IgJj/xI4mR6YM4yvHOmxJivH/
/GrKM/SHwDM1ZJvxtli08ZUTG1j2PS4I2a7Jtagj28JQrMqScRDT7nmQIFIUZmq35TpH5s7Hfyc/
fSGPRek+fKQCXgFlXH4osjhQv6Zrl6KdXyRmumHAMKwm/Zw419X6veBsDdbBSjTjXcJbb6eLrbnh
RD13x53OAloHenS7GFwPOIv+zcrZ/Qd6MWPAajce4bPPl3AkRYZi1wZ1FIS6TgmHjhdAj2aNxG8o
7I0A9fJ4/Qmr6I1G/vymvNypw92GyUfki8MABFBpsMQqbypssFtg4/hHSwOoT9BX5PDyD1YbHK6f
KnfTSiaKRBJfUt2pWePhIScRugrpJy14TDxkXmJnVIAAE4rYIq4paST4BvLADTy6IZTY1mxdPIbB
t9g95poxJjPeaCTvNPBlIAxjW9Ad9GR6QSADjJjR7QwDUfHQC288LV02ektYSdK2XGHJ0kibR1ja
HkeV0vYkOORZQZIM9CD2TWTKK68RHcwPQOu9rHIh7x3mcgzEpwfrzI5y7GVH1grhw7vjE+10+Ctq
LQjIqkYMid3ahXvC4Y+0GxcqkL0dxeb2k/kz+CB9oVFuVHvCRHZw8+7+eHsJK6ftn1IXy73HxecV
T6/GVsOYvQEc++Z/d1z6Iwt1n5Be7zfwYAYCsYTxA3wsKq14asQTJWT3ylaZryO4BUByhjrncb9T
dfGliEGCwmKH5TLDIV+zTEwZ1Z+MH292dxYEim5Oc8D91okwp2dD4tEY745qsO6tk1ZRjbk5qT4z
kBrqjeYujedhjghrh+1aUInyPzw7jTbe1EqBvrFL4QMyndPJQzFSu8azrGL9Or3lH8GV1x13pLUG
x4f12o+LQ8c6nZWoWoyyaoitLMdD99ziHQp2APmTLFNEX0RS/U1xpyTLE+TQuhxYZ7ipI21DmgPp
X0oRO7zXEC5AP3xgyL6hABKEDEJar1EnMPpHf5NV1suwZcECes6NRKBof5jd0sNJAc3Wp1VeY7EK
sESKtpOm8wwq2s/Qod1XOKnXe75BDAB4pltO5AqvgxJeSfYeg/q6THdqTYLcSxM3Mj71xF1ijPGl
X1WyI2G2z6pq4+aWgF1y2Q6ixuuAz/YbJGE+Fg1jcGxgvJR8/HdfPaFNTp5jiM2sWoltQKFzTNHt
fVgN5/M6XPPnwkX4bCe+7vKDefpwJgzr5bPrO2l07uYMRpaCnFC4thqcNiuythgz7rKwHlnwSd/J
0R/wQXPaR75jaKYLRKdryHdlwv3Q61O+m/R4bZN5T7EdO6iMocxKEfpDIkG/SGmwjI6C2CgSJrqD
bAre5V7H8jqRwFDeHJdR7heCqh4dTPTcIgRy/bsARxNwV4pazKcM5EGsJovdQZffMQgozuHDjL1J
dcb4aLDI/Y8qsVCzzjPMxfxUMfJe7EXXh/RNtzcYFBDfda9DK5Hrn5Yi/LgapqsvgiwFWwHP5yB2
1NUdriv9OtHEGJWdF3EYS+/hGj2/g/dLSIn9uiEgQ4OwAOjTswJcDlznscY53kl+6Ql2MeY5sfxu
6qjw/BfVn7U1UTBFOxojAx+/HD7yCUii/Ak6Wkw+iWGxEb0OXt4IPsYs09x/lcM4WJjNQhZhkQ2Y
iOVtiqA0uTwXrCdmZrhw5h/VvEP6H8YbCbnrd2ZcyC96XTEBuikNB/i4dVI7npNV9wgfFmZ1s65g
LZEuwWizOqAh+PcHeFOgQnCxxnH+2GK9rpMKAt+wE8PKmcRWCpm+q4ITCc6JBKHDH2wpAlIMmxnC
G5w/h6NNceV4ZwPidOx8c9Il0+/kCNNCABcRRqdknP4M8XiNSFZWC9fzFjADRHTiuaRRrAsjIOB6
iSRclu7LokDFEPSaCt/jZw+HaVGBir7fN97dku/mq1egi1ODs7puT5UX7z0yut7aHpcHLns3U2Bi
NOvTZH1oZRhQ1++oSHd9Z5RyklAdswGyeNKVBD8hiqsAUyY5kWrbzHVzHUW4BWec5MfOpvvCT6ay
5GhwijzTCZY/MfvV4hm3gDVTwkSml6qNPi4PIoGLAF3XRkkQIFlkO6xRF4BNNMpvbubTOJkmHhcx
b3rAuTNEKStZZKGHSff4BVU2vMUr5731FRRv90fXDs7A1ag9RKtY6zS1lKhCTSGeCmI8T62+0i/R
RqCnsJqvBlijARv0jRv6VuYAz8pf6uvEHAVrKZpsgZBFM102zDD2BEGhueEKwc9qNwpC0KTRqgA+
CCyUZbfm6Dw/RqsBVUCgpWQwseF8lLbwQpBK7inBl6ZUxMQz5zw0ph+rmZsyjpMVgd6YVLUbGVq8
2U8hhLJPrsEJuDsxO48Z7xEcDJj5Xiq8mTvV5Gi9d+9lL/dbAYh/nrViB62pwNvCn0QBjhz5ExVN
f7RZCpTMXPlXwyeQTUO/N5kZ30lQUl2OfB45rNU2Gds1V7QG+F9xmgI1MPV3hhnKjRWMeZb2ucVH
syaV0fXSvy66euzCeej3i+s0i6yb4qSdX9XlS4QF06gpPHV2gA+ldi2SsLUOFaiud5+TauRJAn+7
zM5tdO47GlqkS2qK61rq2n4aM1/P4ZocGUmdHlEDoo5/jMFiJvEmT8HAOfbkWIX/ScTf9wdi0kNP
lTvggoa8+9WXhuPMKKrwqDcS8Q92xaxZK2J8mCXu4UtY2t45DBIHFSRfFM/KMo5dOgQfs8wTuFTE
3St76s5jwlpJtjnMPDvZur66I5BizWMmpXOGnWpLmQevM7xqDOZcp05nuzum0Obtq6bspxdL5HK+
LIvgQUD4ZP/ekSIm0nMDAz2ux5d9CvlJ5koIkiofCxovJaBHXqazUtzM+Zbn8EzB7VhRwg0sCVXb
F8RqcNvR5Z0/ujtd5uzL4b7ejas+8+fycd7g0ctqc4KM/S5YCme3UKdFjIR/WSmTTy/oyBy1INud
06L5gmQg74ejDca1shifCFSgA8ZYsf6aM0wQfk3Yoa3LgtN+FAIjU+cHd/01L6sqefI25eFHAqvD
E1mMpAuP5rsZg+AEKOuws9BkAEA2eu+6LortD3wXx6ZQEQ35zSxvYSZpBP12ptpJrU3exlC5vJzD
M0p/slVgZnhOCVYFhhE+3tyNHQF/HPJDZnug74uSkYVZnGRgPhZHJPRKeVI9WfxTLTTiEPKspLkM
HIvhWxRUWHBtuKfLH81UMVAxgjPk79MGvsvJ6W2WwMxMEX7EkFl6oQ3GyUggKIOYpRscLa46em57
zHTmm412mbgZmyRwuEPT2umiRqUJirEkboPJsxGpqU3KKcW2tzFR7MXr3te0IWO1vdB48Fxrekg/
AzhWAaZ1mAg9731GBKRo8qyWTAcwKXMShX/He8rF/kIKu844J4acvzYtr36SX40IvFczdRzzO9sC
fq85anrc0Iw6D/rE2W2T9ZU6eK9eEG1jFLVxocyc/OOchjk8XewvPy3zYCqKpyLIKyyhXfHYNcQm
spwHHiKbi2J3L1Kq8CQMMA6zQ4KzzVIUmU71UOIhw4W040aTmuSttTHkjo1XCqb17b+F8mKc57Hv
1Pb9L7+sTg1g0Fz25U/ymXk2Tqr0M0h7jEFM/H/kB6FvLB7l6hkj0lz0lRzVDlU+GW99zb93KBbs
735csELBeS46T9AmDqbFFQKOQROZEpRkhSogLBlr5IA8JU4HK5yh24dmLe6yQ6muegXq1i6MN3Vm
aEdfG4E74fjK+3FdUfQz2Llj+UQ+P0IpUDUhMcYjmIy5QKONGaUrT24sv02HiozZbakFqn+ZiJJD
0MbRSxGUQ0983KtD1UWdHg8ybP/6DpmOhIjeKSXqN3/I0/jLBOMywa1dsEONu0P4FlSPX8RcKYJE
ctS1uPFfAULcBwSoqIiz04t9sZ1b+dHpLzVaYwQF1ePuwLYbU0wGWSziEKs4yMiCvNHF5RJUHd4P
mJcVfh57Nyi3UNk4BUuwTxVFCVgnBz8HQJMHuZpFJW6pUUGfa+qOG+5gWUl4b0250CafvAPmv3RP
7pkyfSw36wKSpWCQ98MQFNQW1CU9/P+8FPni83ZzsJESwl+L6O90Ou0Thocts/vH8wU6xQb6XrrB
mGH+k9HXbvmW8CWxNu0n8wPV/A0tS06cIhqD3kYyp5DvPuaeaAjRfOzuRVqeZV1FGgSe9+xGkCoq
ZOi+p7Ye62Riwrv0vFB68ZmOehUs3/dlD4XCkAM6+ZwYRneWISfYdVQUPVnuPOoPGu2c7B7Slpgv
/KLTkJM3/h7sZQ7eJTDfLjhO/1JtccK06VE2+bz/AmSBq9TXxQF10dksSzuMtZRwkdqE/+AFA3H5
OAiPo/NOvvTPKteuDx9FNAGNf5Vjm5rrNhjd/DpveeJPAOkwff2bBaCcLFXamJ0++KbF9L5660kx
IadwJL+3uil8YzrGaKmj626aOVGJhIP7MMoLiIduUz/q6ct6jukZgd8pmVkH12V05LEwrGfjgIze
/nQN3Ov+/2fzpMJl+FcO+v0T56UvFUIWDpK8G7OPlHn+t0Jpbat/ASzGOihFIXcPvjiedFkU9Yme
nAA06LezAxid9r00I7jG8BGO3BxsaeOeAKHpmOa2eDvs1EVTSHlkg6t6Hq9bC4UzU8kK2EuAJxCy
+Ti650scoxAO113OqGpKCo7MZ98bR5f+JOERqCeU8lsEQa52PeuG2Tr542IBZzpMo5uHhCe5gVqV
JHYpB+Co77CO7oxD1KyVrQh1WtVMTx/4vuOWVC5eaIerAdl99N7/B5jtFPLGS6MarnzSFXLxOHuV
fiqVhNRKw4erZyfrYaKH8KeqIHb/bAjuzVJLM/hsVGs0KuFoXl40Dssxrfu93GB6vVk6Ch8poIgh
q926D81ELbB6eNwxw7v+uTkFjLO+PFINgYiAKtTw8Bz/HgZmvGFsSdoMqvotMiXnwmvZxSv7FghS
fgj2oNaZLfOA71hBgXAqRTntucFs9Vx/5WJHwnbhdGwGJFKQQtWy7buN21M6urPukT0T+cxTpKvi
pScR4vCQQS/7Rg1n5PyxHANlFD/zFuJEuPw365l2DvWWwx5aVYrv3hDjoxE+4qpNWYooVowEVKZV
aLyu3RK0NTEtR+k76/w/UQTfX4NHE75LC+Nhn/lGJlgx0uSJ5Y7GZV7PsMVNDO7NbCULCVbO+B+9
aRrDRllB7eU1kSw6QngaEvO7IDXBSSaobpf7DA6cnc9X2bn2CAKCIJCr6LfNvmp5NZtKJ4U8qQVq
hD8Mjsw0kya0NeeHSH1wKdXJlKWEzqRBPXv9xEoUxZhTM2+mBuMRlFK3DbWljcNAldokk6mD6ybl
IvYYs+UoZGod9sfmjk0yGyNmObu9/k0v0s+bzw6Llpqj60QRnYmqlnOa014plPocUiXFECniVkSs
hTqeaX2oNJdZBfALZyHU254af8g71wXtXgApjmPyrtQqOzck1+q3xKf0A3C/vigL4lx+3lej4sAK
+MBvVML2SDt0J79yPyYqbiU65Oc4fkGNH3siVEcYXyYv4XrKwsIdBlRHsQRBx+DzgFq1CUu5gr4i
lIbHBxiMyqCyuw9PP3mgl6hsjgj558TSst8agzxrxTLQpqwop7xzGY46h+2Dmr7fg6eGp3+6i/Jj
JhfMIg75M3XrLG1wyppXjOD5cvlS9QOojg0sBvF8rTtXKW4+Dd+HY58SUHHq1xFENrU+cZ0Ji5yA
p2Y14/7ZSACGZ0IEt+pu3rmvck/l4WWuxSLm8WeTL5c+VZ2hYi+8JX81YIj81TagfMv8iZ1PeYfE
beL8/6k8sp+LWzHIf2H3L4vZ+3pSnrreLYVADimocHfB8/pC5JyL1uLlhoGy4RaZAewj89mmvRbO
mR9h6nJce6Wf/ahmC3wC7SWa3vyCTS3YH7wrbnnkaa3sqDWP35CFKS3uauqTMD/viEa/jA1KFNCE
p0vi4glA3kalun8LmX7KQfOWjgflI/yuicaTe2xQW45iB3Y6WW+QYC3oHfAVptfLJLuAPhr/LjgS
b8qQtX7xXl9GkpCaPiRY6Awo5bFM4vGwprRWZu6IeEqhdXj1sGXjr65h8B7kIi/Fy+Y7H7A7zlmt
odlYtx7yMKdclTL1TPuLz8YuD8CWWsocG2VLZ6CknXLLcm7QCQwVZpieag+lj2jLcQSY1yXQ45sH
EGl5mE94++3IWf585nDQhXGcFnXF6pTdObeXCygUbz9zI8MQQ46uPFkM9/3kRzuEiYf2hGUyXx+y
HAJUImhyFiHmcgNsHvi9R1siG5GTtays1of/wtapG8hr/OYl0SvNxzlQqegV1E2uwayH8lG4HF1A
0ikiIP2sn9ec9tMzQSgwwbQWuQtIelxu6GIyBlZsFY3UwVSzj7/CcNnjrfzog+wvGFU+OlUNXOPF
3uJBeKCrhyZkmeM/TM8tfh6zbE/6KQe7E5mGrahy9h94t8RRtNxdxRTdNMHd0SbIaGy+hJs5OwSd
L4XIHHbFUfq3kKsAFJyWKrS/+4cCTUfuKzyfBR5JJoG4ztlRgXamX/gxb1cqlGaGFkAWMLsvpZLr
SSe5I72Q2dgFQQCzT8DnPql1/V+oMIcaLtPOEAe9TVcv3wcA0oXIsCTn5q2CurL+GI1gQpg+M7AT
0Hr/+yyAjv11ZZhOxct5Haz+BnzZlfW7XxO6IhohGeI1kzLh468oZJbUuzND8wGkRZFrm+0BnuWN
MgF2mlYFMh7Gns1Oxj7qmqh+1KGZdCKdVX+6rJxzV45FxSXZwQi7hCoMv7Qpg5voUqZfajaMlPQ8
jO2Ll8lFQx1SNq3bemCqm3TB9TsIXfljqQqmyZa9gZSFCq3/0Fuwryu3uMRdHZzG7ujOmuA/nG9N
oVk0tYJzDB+HRzHFcSOYGHbYW+cdFDspngeFll/l4K+DV0qKnPIFOrfb+V5hwJjKsle6hbF3U4Gp
XkX5ESOn35OWbNWEI2eZbNMu028BxcCZhLSefewsfJISl9f+Y9tfFkMysuhi0HxoqaXs0/jg1GND
9/Nfv1VA63pOUyS+Ac2isFw7Q83DfBT35V3NPDI9BgdhVjdaUQKmHlD0CJa8TqadRM5Mcu8ZI5fz
r5jMZuBm3ryfHI26/gzhb0CqJp/AsOnR+2sPm0/eAkVy/ih8g/wm8xWadyfWW/SiIXqIn4QxMYzN
8/xJNa0OMJRo2aTgYSisxiqk2f7EiPkCy3QhWrpsCET8SlvA4PjtFoCHd8DbDRvuJ7dcKtbnKErW
E0ezwcOTloBf+XCHHMuHWHcvrzZtrhZ3s5gY2SiYL7NiPsX44f3Hma9DZ9PijjEJXCcGfuq1bcCw
9n5t97aUQWY7p/IfUpYa5m5YpLDlbjKcFoI0GHa5PF2oZwJ56cvdNYVf00xZ99qePeehP5RTesd6
uS8Ezq/ACjiVA8LT4AbIBp45cw7uo+7ETw/fpe6RoR9Py63DoGA5tcQGdPT7GeBz8BZEOSqjLdQZ
BPhO6b0J1cmHIRN628AAMiIlKRPzAKTk6GeRRLvEcJMg6fipVUd7Z7AxfkD0sLW+H3g83Suy6kCq
c0KrKEkYttRKO79DxQiWHNUPwHXSJ1WyMqQ4U3yoYAjBhO19YDnjJQ/ol+cGSZhboG0uBC/EbrqI
hsA4zYhnSaNANhZH068vspigEoS2ifH8KKucuZ1tHZ9Q+S5heyaRRX4xiEW1iZ1ZfQ/frc/6oHZI
YDmmuGyiw4dlXlCrqO68TKsxftEfR1PtYli+bd70POkRVfXW6glWjcbphPhHg79MzYWBlwWYQHS6
sS1KNnOfhq0TW3VvBrcGvctujsXu560RK9V9kkT2+ceY/t1NJal2XLJvOLXMWv/UgWKUJeyIJlFN
k3jyBI+RuvVyPp9fv3yPPMYtbH8rUxLgo4R7llOtNsx+VgfdXpKKrD615f86Q9YntlmOYU2o+8+B
QqApIM9PMvg1vmb6MWYKb+Zb0bBORZtn6sRgWmTjgRLxzD98zIv+Iq6YUUM/dNRte6LKdv3lqng0
LvnRRD5skOpgwryvaX+iqKqnu9wUpnEbMVdzFAFI0gCCCL4vL40/VGP0ifkdExp0CojZMo7cyrRc
rxsgX+2BZxw7PLwZyHbJ57PmYq9IgOiTrFSePmGXCUTt0i0NpfNLv2E8AJMkVeG5Ube39nERn8pv
RHNILBSSdnHPAAFgaaiv78Zc5hrwulcWtWQTQeLzZ3hS/i1go+nPyKWiYfwVVzjAUyJOgCzsuf4Q
z+D1sl7Tsri0H0mGDk9GhFPx34WZ1CGtjb6yfNAPISJuS3oR+kH0twVzTPYwvjGX+W8XpO3vEF+a
DkLEJ9lKkFcRRByABL0YpYlof0B2UJSyBXS8FyLiAylG0izafrqQZD4B7wqLqVpRQJxmtSeJCKT+
rltESL+ndPE4QZhPQoTmg7FIrxM0JWrcOoA8bmB5O9ND6EnGDOIrOtveJFwbQsuqb6ZN7M2Lt8af
rqJqJGxPiiHhZjSuvwDA0uzjeCh/PeBttdC+mWJTdPgsezsZ+PPPD1NvehYmO+VFbwP1Quogft3V
cfGkSNS3VuCEdMI9O2Are+folL9HoeBLyjkctmmRe7jzYeJWsRz4S1cpE/D8a3lkVjPVzYfVWUxS
WBG8F+Hk4YsIKxnyIJzQ0DKo16JFpDwgI82a+GN79GYDtXsuUGpps9YgJl6JwqidI4+l7RT2r6U6
xd9spVtdEMaNTEgc64valdhSyq2z6Yoa9uahabSNOS9CH0UfF8g7GB1vTcy754kjiv9iHPkh0PaS
630SFipHSCVHI0uhD6vZQbXaxceJNoxhybSKw63TmPP9Mycoh1mrHUdtB7Oo6jb2i+jfZ/4WBsxj
r4BlxdF+WEbmQiFeK4vkbDG2viJ0it4OxlE6VjkPtwOvZvA6og+4hEdgGDDj7Z3lPqqTyAuaVhSg
QSerwKNv9buZJJt4nVErm9CoV+xHsmrIAZn/x/BuloTWMmdFLeZWS1UVrA5QMaV1/0l9JXCyK2Rz
KYRXYOz00mTMx8/YfKtgRaIB3v+y7w3irXGdyYuOlq++6BGomgonJN1OxxSei5L9W8qLt+Rvpuwz
K9cxBZK/unFVvXq5XzfIdypRT55yPT3yXcAMuzgXkeNzp42Gcc1M++a8ZMU8eWBFQrEk7LpoYwml
Lq9FvqiL6VKi21Brmr9uats/h+p9Y9qPoOq5awEmDnApNibl/+nka4hjRWNm5tdRoGgH937os3mU
1s+xUVpaqle+/xovApCCLhXB/W+Vf/+4AUAHXmyzDAGFNAqslVcxf11htP42ONkPkZJOSCfxsxoX
Ovbm7PU2yNjbuAVxf31T2+I5YBZvnJBiAk4v3YQCaqkgVufW7/uPZbWww0E+nukvKplbwYj33FAJ
UYze+hW2Xc+LNS2heBL4zNAiJcD+/99kqs20t/hWsirzNxCk4raElQIEOB9K6VAJHI1gB3yX7soJ
hjsMAmR3lqO+sigwwFQTXhQPbwruUqxlkUdQ5DeJx5t7QfvrzYWVMLRHSU5SAHb8MaYOe5Ar1/dp
6t70G0WL+veDMYoWeZkPXsjTLRx0U95FRaCLPYOR3W0Jz6qLb4ygsNXylCxGTS6z88Wgz/uNBEF6
DU1n2xKj31l4w+iN6+pmaoPFK+MBjtygYNsjY7gOzLTLfNymxUVMGKXS+wt1GTu7gutoS0S2EIRr
TqXvb0dIpKkaHqLz9qD+uTmrSMX/9BvOJH+Y7MrxHvHQjh9cCdXtBeh2mmcV5KPVKlRU1wf4WIix
URR64mk8IgX5C5ArWXj0MR6u6xOdDCZgwurG7f9Vr8Ev0IqcIP5oBVoCGHbRDrGjAmryKmR50ahg
NKhFaCoWXZde5HlFJs2FEcV1S/JNo6CkCi5KiOXxHfubb30tJURQb5PNrGQlOILH83ZGGQdbBH8F
PizIS9xF4Mt6V4ybdLv6UP+aqcZj2VUYl6JVmeCEeJhFDvsaocKl+NjUZftWlyJ39/PeWB29HDMn
4a3SE0wlWTGkuft/op6Dl93IabkZWEl1bl1OKj38XR9tRYAqmoHiCdUdedcNqnnLr6jfY5hWkpYj
9SeiTXuWQ2y8A5+w41E8GgYQ1HGfU2FDMcO0X0KKrNBL7MxgA60fhjHf22NsIYbZHjh2SG4CBepZ
JKZuz1J2NuUdWm9eCdoVGZjNSLYRMYMlyUHuB8B6S+t6WgRnwri0qM7KHQzjzuMj9LWsli5QyaRW
bF/64rBq5P0/L0F0IJkUwQ81lQeECpL+XbcQpcJLeyM8DeTkalto90SkjPf+xZqHQduaTw+qU695
3kLJxfGcO+NpUt4G6GbhLMinIfdiuX5VSlY2Ztk/w2q71Uc41zJOpWNh2svW1ySGqD9wgS00kaE8
0BhNjO7OPb+83ToezY0b754pVFNuf8Wg080E2Rbi2l6ho9OkiDZoABrbFogSziRxkWSMCqkY8lEx
XwTLo+YDzipvnB5dUsas7fy1yshEcLe+awQiMewMTY16CfydIsS65xZ3fmp+UrS2/phgFKXEsgw5
vmh2V/esPg/oslm51KJDZu312RnX9y6v2tRwCyjiIUf3COFUo/ryJQjWJPVy7Bj7/lY23qK9e9ox
Fy2wyO9w4o2PFGi+77fkSitJbsHDDFF6QkV6n0NK5VN/RqnURVw+wEROp1OU9w7Z6c9Ghig7zlqc
zXN4H0k7Nhm57Ti+7PykBrA87WsqqQP14uMIDUbEqCecke1wRD2S6aP8ZFwUqNhugq+68YFoffrb
fX9DsEiZpu4ZLaYgrnOMWageiYt2Czmr8QY9G6pdbr63XAwLwlmZV7E7iTtchAwiExoDhNR1mHiA
5QLJ5R1byqmbhfO9d9ejKw8KJ6j7eZv3F/6wW+vFIulOWzgbyM0Wry3xFQJDHsHu4/qPewqPw1sy
5V6kDzIyhY69mp0f8IyTD1jh8QN9/9MhOaIDwRO1fFxOOAsXIMRziAmXnEOYoETzqHehtNqBzrxI
LoTF3XD+0jHen4FOl10M/MCekhSceLkjHIh7LEBp7eb+c7SpcSBtjjxPXZL+Zn6i62fdJrEuflCY
FfM3B64NwT2ltLOtZJbUmjgTOfY+d1qO8sEYrdHQt2X2+dXqjXDqGKyb1l79ykNnpAIjbg/PgKmW
HHMbJlkSWC4q8/lTh5tySDrnNjSk4ZYUSZHTiGU40YQeIkqEb8GWEr49+rNYBEKeEMJiupsuJq0i
s6YxdUzjVRv/5UR4+6HUqozMrq4PI9WU4M7OpFYwBMV1WJ/cE84nboA+BBqSiZWidDXAhRdZBRP+
8a2I7GH0VQcRvD40GcbXiuU3EpYpRZaD04oi+JzawU2+0w2kq9QxKZzyNkiqM/rloBzJmkQeBlm4
HATCfLEAesB+c+33qLOaXt1THIZOywdRQhqCiOUGUnPRofxM2hnAL95SKXJJTwQGHFecaq/KOoRj
T5sDdcgdLfL6SMOJlpRn/UOSm3WONk4e1UASfkloWy5lTdGXa7HbM4d6EvYmBj0VBU7wz6gOcIaE
cMhhxb30TAn/9fvLqHfGwkkt0dw0bcX0lazGd4cZdFofoqhYHSjzW478vpSPNA34n47k7XVq9hr4
N8pbC+GzFCSJybqNiJivPAuoXuDeckihlUtJtqFjRgxlPxKfr8O/5CKNVa8ybVuyL3S1+BXZfmxx
RZ2NvmYVvTXr0ipcQhgSumezENpvRcew2heSvAIA3ClMHW2CsEv/kI6o9p5WBTHmy6Z8coG5nJ9D
TIhp/xCvDqu+YRczWP7weJz8qmtO5CaShB4YSybHXcDPp1OqHHACwNy+S/v/e4vpjpwQ4ca6vcjL
RAWvqZ282xDcZkhUJWSjWr0uvhPlgfFN4lQwV+uheBIUHvGcfPLCiCviRQyPb0xv+M1YMINpJnSn
+ubIxATlm+BNJI5vSudHwOY3jyp4AXe5Mt0ob5cRQMpcJ27OwFXPpHIkKrQGADmi0xSjOq1XcFEA
n4tNEg1p/jfOZ6ASEY3dhIdkjlWnTRKqaGKK+uZ/cF2CQ2ymadmzsUEjQBCs6s/NSAvJUgUsSlC1
MQwqdxJZ4O5jOvKqY1vPh+PVuQeiprsYCK116D457ZYL2ZJjBKTt0O1zroOVd4GXYKdJi3xSDoEz
kfz2hIPNzsk3SjtpAIdcmd8tw6UYEHADutZjlvOfiM5DRbW3AaV6jhIFaTMiJe6lYbVdsceLMoFW
sQKJypaxQ/AkzADkbTPPMHAdyX5DmTjGDQ0e60c4W48hxJtto5WiI1AihCIrG2C5Fouiwkqfp7Jn
PDOVjFAqd4H5TAj6zYFFo0LdRJ6Jc7AxO/IHuydNU42G7eGmU6VwMvH6n4r7+2cxglHdPpVo6M0R
EcX1s/97QVw1Ao162T51oQotnJ/lFg+4eFr6hV6SbORGR3MHwqj1WP5ajNVaOe16zi1lUMBV+DN7
39qeFMqh2IF6J3R1LCJ9U/zAtpPJoS4qN4e1zxIvsHXCsVVoIptdy0E5W23St8YY9rN9a11hapc6
k/muo8WFJ11N+2y5sSfa79rsL/8tM7oTftzHIPO8LUFRIsPEYMLtvKKvOWENt+uRBH1pncKJh6h1
DSSI8KUU8l/G0jJWoWIxpGvT4q2x863rpqODLLNSebxrIbCmM8Txg+jlSOsjLGGbjaXlZVHly1wv
ku5I6438gT3hTY3kldegKNPYZ49e7qrJihqeb22mH7+0DcgJCUkJ+Cb6cjql0tKNz7EoqZQfwXyU
1WLFn/65/pkspDnF0/R2/jnDZ9cSCRZuWbQP41mca/mRWLC630aa5S5hqrJMkEWxjKlH3c/ruF4d
6U8oiXzKYVDFP55jR2bT2BzrFRAZmJO/6engjXhBp6BbtoLaIj27SAEv3g/CvJ1ULFovjfUdxOXM
Xo6zXXYGcpb7PQ9Mxr4566S+bdA1fK1J6P5yikU+TsCGWGprrtsH/oO7aPD8atvWdFNZYyueGxM6
0j/B8jDHQHJeov6MDEYnUjw2NzFkFUVM14yMPq3zw4OCotBnnLax3+B8mL0c4hgWBIVoYFQR01S9
1BwPYbc+D0Z0Vp+outrm7MUn5rDBBnL9An+MenbTU6Ud+VjImNChWtvrZYIUdBeQzNO1axJtnQjW
8YO9Xb2NMuyafk1lF5CQkoXy284pM+GmlJwS6EJlLwmU3WOnHFMy0j7hguc6hscQHBSnc8nfmmx+
fSTbur6A1K48ZfBOIDZ3BhaxgXMphpVUn1PDMXGD/jw7gFCeyHYryoEzPK6z6E3mkh3lGEHyq/9I
sEVwgqxLCNuuYz76bjVCUQ51Up/Ks2u0iVQiWgXXNmmTmKADkwvS5Z4LyOsSDaQW+t651pC4j6TJ
5fo82tll9SPOfBwCLech/DqG2d4hGXeb+yzHkpY17Elbtimw3JRSmqmdvaky8qCYiKX+TZYHJjdO
VbzWa2rlHrz9Bm5MUYcBv2i0CexexTYM5cfoGZQ1UT1Uoz4/4dV96L7BiDkJUORkF2Tko0TbIn5G
PrIU7Andn+EkJP9bfb13TnYqACPGEW75+mos09Dp2vLWGfMeIY65wICExW/E26eEFNPc3PsaAuir
BWoH540FHi46JZAFQfRlHvgRundXwlrvp+X6j2TnK54TWKxCD/A/oOnXpSpIxpJ5B0CL5y4nEUEH
v17eaAAwRaN78Z9ZWyGWOvyA0SiEySJvqBI5bon70Sb/Th379m8/dv5uH8Ryt5Y0b01F5jzloxJN
F/In6hL5++Jl9xWDH7e8u14kZOmAgvb4cn2aZxQdkonJH124ZJX3SZ3V4GU5opn/MdFSDPRSd1LJ
ciuNZX8OPP4QGrqt+HRmdWW1PqMRApLVeuFcts0dUS9jz9hZ1Vcyngkcf4h8vMy7uBxOG+s41F2k
AdnwomZwyV087Xff6rPuTDNOtkfayfPfRE8cKDgjXyN9VBX+Tncu11c2JPJhIZ5cVDLWeJ/pWh0Z
Ws/dDrtV//i4EXNjOHfy4khR4Adyka/EfVgnb4R3m5v16qitPG7i4zA/wg8O/tAnY7fQZ2tozExZ
jJs0dCohx5J6jEKMX4/70fmefB3egRyuJPE/1VgWiPosBd19eTXYDJ0llzmB2dScxeWTXM1iwrn7
w8cXbwnMhFHwRWaphxUPSeXUo31zaMmpxY9aXbvTAICHLCiqv3H6DmYP+J/gQNHo6Zx5+YNmsg4/
w6crKoeDTda/k4QizYXqVn41SitXp9PoGx6luFHem+CZdsGNWKN7NjrMT8YW3sNw6uMtMMkPJ+fh
7BOE+PpdX0cZ4EmTquDX/UPNGyEPVLkG8VV9XtK9KlkWs+rOX7wjTFBMcqhkJt59hpMUj+zGpRxn
U2lQiy9Rx2RFR5HvHUpumBUjF5TwpZmi+2GwHV6JaQLKqfRv65YxsHC6Ut1w8IyI7HgjaecbxPEG
jhEH3I0h8YA6f/SQuYYw6ibET0ORSiiyD0gkfTfs/rRHSUtEhr79gb0EcpKkEU1bGjQaZhRJfsiQ
s/m6IXOnBXKAyxfVzL+VidkTFph9uVNOSm4DBSs1g/uoFf/iALhWuJ5dHVxRdgAGMZcdC6QO0Zd1
fKL31dlQufkt8rObL/Imz1Fl5MBXGY3IseWaamm1OQlR9Butr93KbbPCOFrYIGazWTrbsYbojDsK
LGGRTX5qGUNMa22P/oIBBPZNlYCQm49fXVUl/sJmiwvDXn0QYlST06pA9c2QBrBZVPn9h066xd6y
PPX/lH2DaNC0QnY1Frre5vGt87NaSJs9DVyi3GopBcNYFhh6iK/p0qTzJgGRTVrcijD5PickdJi5
IkVdc9B0YmsBHRvyJVhWqSsUBVGttIv7ejD/cuRDxuSTpKNF5yxyH9MwA80sI+Nu62GbVB9kuEN2
5PQG9ROgeb9xmXGkV2v14P03BcP5+izBzOtyTMl4f8Y+ClnJkT/yWbun2wFOZebuVTt1n8ENDt5f
HyPiWuZWoAncyGN0tnRjOwJ/6cMI1VYA1yllQYzqOB4xoBm20lZ6KPn0kxsPEjZLt+H+wU9V0N7h
g9b1NkZ4Bb1IXlbDQoqxmMPMaDFCp2EkcgKBAOapOhUJnhadf+DAyHgTg2uEaNjjivdj89KfTu3C
JGe6CvB0S+5AxwUMFRdRPE+jZm1ybjRZD7UNglv8noKZWPDSxozrMMZCkfbI9bBnaq4QW1ylOiA/
QOjxQ1iXpW3z+lXAnn0C2BqAG8tfE+BwVEORCCSx9VBYUnMquOb9HCw6ZJdG8eh6rMHLRwKuVHvM
qtQyoRqsYtQz77Lw9w95nDpOsCzPWovzeRYvMu97lgM1tiUpefDxjQy1E3Q0F1Wzb9IwVUxcF5iP
oFAPNuRNXcS72rWviKUguL3cqyG3lytEPQ6X8AKQSrbxypZv6AUEluCa1/ZC2TNepqNB1jVZgP+/
X4NTfO1qfC2ujtpLwJlcbMbhg9wnE2G7AA4MvSawNB+2Mlw+yJmRiibQLKcjmEfGLbsFQb2D2y9Z
jrT5sJqniwOhlqyEqs7OzPNttvduOONwhHmYbAySRoqnZJsBqfhIsQr7BvYRZNqWha4Xan8ggGgD
9swWCM07NJHmOwd8K/qeHqSCDFgkZlnZBxXfz9lwf/dGcHw63SMbspGk587gcm46awLYX6DENo3f
Tp4EpYSpp73A59zmcj8MyFBZ/Z7CfiPmrqpcMQN4MIzxGME/f+HCb9MIBKN2S9fdITmJYyjA8mCR
fh+zoDC8RVsfAd+c5AhEQ7PaFfnX3lwhf9JNhLnjD0wkMjFccf1ET/D9UkIPdbt2kiDagsKNu6uw
JzHBzFP/3ZBJ1GgZwnFbp2+/5fGGLmiTU0Jk5U3Hy2kXJkqXzyu6GsDBhGz7tl+2EEqVAvUvlikD
rga3NEXlznhsHVRbLlx4llDEosXZ2QjqsGVh5LW2oqmk3qfVKw91f+HiBLypjFuwi0kvUzyyW8/G
F7l9e6mqRmQH127y4buWNW22vt4/8faXf+i5ZKwSMZhr5lHrEsJ8RTUQksjB/fy+CPEfwz4oy4mw
z9IsTyyAtcHl+HwrhmVO2My9TIiT843AoQ1v9hnj3gOvp2CP4Ef6iYPFxTRYDu6N8S3yPyVqwe6I
OSIiqcSHBmZ7R5mpXJPcFTPD9/w6gMY1Uc03mbdSz5K5pzvr/NjzTn85SFhiI28rez1a5/KAFZlN
IY1DxfFVHlS6ltbN0E+m8thH7fZIAh1GMbsQck4vw/52Qk/YcvpwwtIv+gausVbEWj0YBRC/pVL3
o9JI1BAkbHctfcs9txcNaF11QmxtVNwMKCxNu36Nf8n9RyHI62OhZA6Uz0PBsDOWXaD4FVEaFJsa
gJtGFIbcycBVG5rfAJctHTCz0/m0Qs+1AhhAq3ksq5Jkr1xwjin5AOW1UTbAx54EuiU1wPJLlXcr
fDsD3mO+/r419cCugf3+E0IknxzIWEWbP0WdEuOc243TNYdz+iYquSzTKWEmDJoaFeL0AALmIOwF
7YJ6zxhNGO3Z18FETAFNFwfxLaB9PQWRgAK50VrogfUJWHrX1xwY7qxIq/AOoKpgOUKM5bsmouAd
EPId3PujWSQ3xHWpSMh0ngJ9eg9V6wHh+reiYj4OTwwaOtSxrC1I0E0w0JMhDkUmKzvCRuI+saGG
vrODHwSnDRQS8YbpI8/LVcY1qlqd3BACruYK3eJvqpg+pffSaZ2ACyeuPsJfXFJMQpWJtvzWS/+G
aRqWy8DLK2AAxVM/9v+gmG3Lvt8OBZe/po0XxjCjS43byOdI+FZsP990tD47hg+K6uPmPmSuqKRb
S5/fv75ycV0fMoP7S5yxNSl5wNXwv0TqFEnRwL4M7s+WdCvcSbr7YwX+iVUtZ0ogyKjSsVCRAD/1
bEkZHh0waGP1WGO1LadxOC52ZEwyawpxUSAtir8lVS/ubwUWsQLDSuQHDNj9BePJjCrxbD39lIt2
KtacKyBZN795xxhVr0Bi6RoVIsCLCmCWzhpBAZtGZJ7/DDUDH+TQ37rDE47VpzNqZrgfd1rmekWe
ahy6E1qvADnRJB+l1tc6sHVJmUyS8UIiczQr/GodoJvVUdsaqmswd+Idy9Ry3B7xD40OsmHUjGzi
0t0TBRnBBstOpigIlNgHeLDianqXwnrTqh06vrSWrL6iDHu3OaYeQa1DkFiDGOToBCfxMqPD7TNO
8cZtcAWsgpFcu4kXe0uapo3fIUE6guROd7LV9bkug+svYuNKp/Dq7wlOXA+7gVBCXxIroutPVyRP
/d4rQH28KSLXu5433RF16o56kGfRZsA3u4cgGIb8ZaXpuRSrMm5bqDsnlPruC2/KoN4HblMEnFGF
6qnHuhLw75CHyARP3vRSJAwUn0CmsNE3kiNLRSGMQ8vPD6BNL661qUL8Z1ndjXerI6UIW21/ADeb
DOINTRUh7ycSJZUYUl19u0/HApIWwruT3tKlbYu7oCB6bUaf2ybqfNxpjShUHMpuBjEeujEw7vI2
ZkMlWUnqsbb6Ch0Kdeol71qWsSQ9eHmylWCOF3ZgN90Jekg3lwFlhZhuBAxNwwO6kZEnC9bCbvfr
TfCs+djibNP8vxSYcKZy6Q/TpDrmybtrnCYkvBj+ONoBow4Rb+pwoetl+wDQmAOQNp1GtN2hEIk+
PuSPBnpfxxw3AQzROfM2oR7KzV6WyXiy8TPE4M+R+vWRftJmt1TJlcX+7EBupXz4dU2W1p60nEMH
lfqe1BjZDD8aDQCoIscwsNYWZwUOXVEZmv0gLIKEXlYcMB6bBkjqOylHn8LnOTKDynn0xQmNe9Cf
NtlQ91bqIbFiEdXpkFNLPQ03KlPSxVDycadFmeW/sOH5XkJVSA5/amsSm2anTJ5kiHX3294pyRZC
QaWWGeLTZegUxijqtdgBJcLej1BcDdYZot8WiDMB5QL2GKYXrr4FG6fML310KDJzLTRfUtWaFEo0
lSto1/LU1sdncbekF2JYUbB7NkUm4a+5C2G0KRpuiJoIHvEhCXJ6eTw7XHR0xwqK+GwePuCi9NyI
dVQ2JTpgEnskHQGe7DuHqrwTUSss44u66NQL3OKxhvHgZgR3snagTX8q3jF6TIdh2BwJ5CRG8uNz
EnOqgTzCxN/MApy9FBW+P11Y3+RDP2gqeGNPGNVBqwwwCjxbhHEs3VrohHRWKMNyvT52HK+V0gBB
5ftUBT+QyBOzA+/lYLIruCNL8Fz4077/CqEG7SbNB34JGFNNiwjquUply4Wp4ghZSRMQcLOp1AL9
/QPS0oMpMES1fGooGggl9meKMWCZj+diCfLjETVMmfVkmo6pbVLp4Un9djL9S2A0S9kwdA2lXfyu
6kqg/+Ce0W0oEZMDwQzm6EY99JkhGC6ujLRndqzly5yBB3q4+9tSQTio1U53r/f3bWMGsNWk8NVx
5kqLi9phuk0CbiifZt8oR+nPfcwLLnOvhd3USl9Ds93hnCfArUBVZG5VijJqP8oaz0bph9yCZlmD
SMrYxXwMehJGbs+HLmLNLkAnZS8xxlwZxL9BuPsX7KMbxjmFAs1LrJF6KXUNFEsmk13qSYoxrPcW
PSb/QQUzYgFbEGkYXsMuAEPYvH+JI12Z0QT5eX6h+1iKHpELqHcE4YERCu+ZdaZpPbjruLVBpo4H
Q1aGL5VENXzler1Y9Bc3pSVQHL8uUi5QjO21P2hdU7JbAuzIvzlwnBLP3sp1YYpgtZz4Rl6zyjkR
E08YMh1C4e9zqKpaToHoeCz2qt/ehfFfxvRBj2RhALdn+L8qEqxYSQBz10p4FMOG/+6HO21uXnbr
yh6K2PK/faFihMHbn7GXyNUdB9Tlg2c9DaIPr0v5Efq9WPaYfZOmIMdPVgsNQoW6855WuHwnqkmw
Klzhn4Ezyoa6+j5E7CHgHo4r4PbIt8EP4rCBytnNpkNoscyzEjUqEqa1KgkVkxdboGC5KtNfZlHY
OEbLTOzRLsyDOViq0l6P2VA9ZoSRilkyRlszIEm4hLZxq/LB8eYlQOiph9VohdSzuStoCZAEVvyj
p6YGAehi10sY83DWNJsK4ldmMJdcAcLjotgKkDClY599hFFK8j4sNK+um1otZHzonQTsTNQuVhsB
uoB5lVSYWRYIbLwCud0muGrX0TM4LcXPLs/oH6wYY0EBNoSwZ5ou27ttnOmWcS/5zugmYx18LdUl
sxpfVay3yZfrkjdHBlBrktf74EFp4ydcCnK+huarUzOtjUn5/OkrBRY/OUQMOb6XuWOzAeZBfKIy
WmpwnbLt0sLvIU4BuCcpnetaokqwBRKm6WY8t6baNUQCNP6G2S9DAbvuqvUToYkmE/11ZVVb/XvH
Sg0ZAsz7G34C4sDWKHFtvMPl41yg5pUv5W7rYN4olMpJdfrQ9QKA5AwSyKB8G80yqbkRTPwwoOci
yEt5FEhpX0NzyEG6Tu+Omh0KtcxKGhAU6QM8/2ZZoTfLXYz+66XtXnmEA9WGGFz53pxL2R0bvEM9
i3XsXkUt9QPXiVO4RHiIT77vZhlM5LPRfsceCAXrb2qgDfP27aprwyb+fjoi76xIf0TWfvoic51o
FZ5lHHY5K5D5Zex1btAJu0IQEpVZR6s778wWxJd8ZOXyc0wmr5jCrxeB5gPErEuKFPhLNgzkmtWj
dZlsJLUeLWBgJ56TBRocY1x7COCjzfFYQWZr3y/wNI8oJQDnHVus4/OYZBb6Wl8aUOqvBZdhjUYW
i3YG0RMHcvYPxK82PxTYQdsHg5wI0cVzrFcWoTseXn4An9e8LY3SkgXdzVf8REjivfofJ8rn+xOj
zcOzwlvK8ISdA0QmMXOwyJaxeASi++SpffH8qXOpE8cAEzqk3kaFdhOwQ26Xmqpamy5gygJoxHEY
1HjyyjFtrPE0qjvl1hf1BoeUXeSrIrkWi71q8C7h8UcBrdci4Mx60VKDmsGG+6cQ02+Q/PU9w6Mx
sP1oap4cwbsar8K83zNl5ymLGnoO2NXEOZ4R+poisZZXveEN6nflHAGeEYX+6Zx/PdZ5X4KP3hD2
g2qkZeRm06lr22bIHBB5xXc9m6rCm0JmIE9CZZUaQ9fX2tNRIfyuuq/uM04S1IlKmYgvsN8udy2a
Wm5oxi0gMAyddfGf2KBCuTVIFMvxCMYlLyg3IyRd4GjHzh0i+7SLKqGGO8ASpDjL7mA+tfut8dJ+
DP5mSDjYY5ctmNVX7S+Bo3ePNNC0UipvTjublG8KZMLUSYkRmFPg11p3Zqeo9XP8MBAv0FvZUuhb
tLtXfGaHB5zzlrevTH415TlUjQoFGSuMUHMsMyMDNlPjRgiJErk1R8uf6XBEpFD2gMTggw5xJxzQ
PYKK+NaAU+uqj06Lyn/Va91bBgnoSu8G1li+uCEmYS2gAw+iGc5LBj9tv+wBNXnIfhBFLru5cbG9
X+bYIja9YIiUMnP5ig2XG+86/nMHqZwNCxK+h9YkF4HNI1wxkWmu3vCdVX4V66YA5JBbyDAMGzkB
XBr7VpXPSfkEZjAzMkH3VtRtCsI72m9VRxvov6m32Z72Eu4gSZs+cF4bEJ/6c8p+lpf+SmhuaEPV
l+aXPP+7lIsZeAqqqdrkmp3Mz+vWA5GXh73qxLM5A52kYC3P3dXmaAOe4u1WmH3N92oMO1lqGd0a
5jdW7a/l32dy7UFiaxcR68MGX8ffawbmuIPE58r3cWTPy0kUCplnrpSaPM+bkwvGRuYQRbQcdUmi
E6oiv43uWUwfBsY/+OimW3p0SI5MHv1XmWoY+HXOnOZbBdct5VVY6S5UXcmXamCUkMOnMA+p4Xja
Exc5JQqUxxAD6Z6BBfl2t9D2oDoZznorLaaMu2F96z6LU4Jj3WJm9ifLwrbYkka4IQG46kWLlwbB
k4WyiYsYFDNONB+UTFXGXGDsXH9o6OYcZakIhmOqIEM7A2kioYYmKQ0XGKGL4JkNbgIwqffjAdFc
hac5EzDuhVZa9pzq/mYTEje9VSMbYwLyuUN7XtrwIUxwo7j7JwtrFz2CY8meRQqZ3IiqzSnTbHyP
AQSpjTpx/9r4fq/Tv50PpACKMrTX+vHQzjDyZAXL8B1pkM0qrFSGThY8NEKA6tgAMSi4ZDjxaWcU
ixVlSCuH7hOMizQomuYm7Uj3AU8F8kbpjUzh7tO1RKH+e6FsPzv1PRcjnqF74tYoC/w1cOB7wRpF
sUvOS9ChTnuOqnL5AoZ1LOPJKDOnLLvYoCl0PK1vfRz6TtKWu74ihupZ7vCu8Kr+UeuE50w/hG9y
NqTxIbIBLlD61491xFmrVXSqerPkjcaOh1X+f5e+GIqT3pnx6FkHDZPgaDFqHbw72MO5pIO/3K8H
f3ini+pKv5TNo6G8V2DyMfPry7jkW6UwsgeAJcaRE2BXePGeWhZkVevcecOyfHmT/lP6+P82lDvC
WTgxwfUpj8+Sec6E1Q3rs8ZZN0oPErRs+MAeQtw6ooOp/hcsZ04LaF/ZqL2JVB3GFWITmHs3c34A
k4tFNraUj6YqOrREND3/hte2Y9urYStbF2WtCTPCD3lXSY4X9cewixdZPp1aQyTPpIZ0JJVwA5hV
8vxL0SvXMxgO8XB1/U8yWjvFIo+v8J8rsy6DmAkEUlyf5jLiDmtkKktJMY7Qf1UbI2ZDPMoWIh1p
bv8aO29HjHtz0Qok6SvQJ38uo9cNQEEa3h4DcQf2lE6WtMCrLSYVpSR/1Gutrg3Fd9hM3t616dpA
vw8d42Htnw1lWvDp25XC9096OHoXy1bhdi+W0tHaYCL/YaY7X+B6DUW+yuxPsBUZvzvKfy7DvVKR
xGg1UbDkfVwdNsXT4vf18qLBR1PFRr3lRJ78ICJW/W9iNUB8g/BU2WFUSAxoTYl0ILiyBoxvFYhg
SsdZP4YszLJlAG4X+piWYaosMH8+nEVkTfkC6n7+7KXxtiSvKTvQ0TmjiaFiSrVlM38ihoZqdk/Z
m3Z0w+9HREiLSYQgfZB0FefmYNmAIVAanwIts14DtnIrnAOZlB6xKyZ3aK0zbk20R5nDKsR7cvk5
eHb7mz9gq8u04XW8ENG4G8ekO9JcnNP9JJu5Pe/5lSaZvmDSxObU05lmeSodgUfkNbvgBt6kQBhy
iXUgZxmX+0w0cUZKSf7rmjcJTDSdXWYwe0zJ52nQ8VKTcyWzPBEDtv/tFl4PmFOLLzNvaBrvwN5D
fvEYk0ZKdlBBwIrtmAUCmr0KpvSR57FuxZEeuSZkivCA62qjG5b5Wd6ap1CjqmhYaa5kVLhR+MJK
K+Ak/QaYHeZMya4qd6TBn2To76NGVilYieBOhRoB4mLJCtjPImCkYAiyx6NnpGl1nC1u4ma8Ds0H
xrk/oPl15Z1cJuCMODsDQKV7Qu9/coefJMgNp6hfwntM+2EvCtTGwYILHVscC4tt+IWlUvQno2i3
EiQVExVDBWogjdrtgJJ31pgYbZO6V3V67UMsukMLGJftNx7JctmwjHJ1M9TAqM8F6dva2Y+Q5ogf
2tbEus/G4CjmhmY4gJiNwb2jUQXuz8gH1CxutzbeVQbp+yw3BDP9afFMoJ9mKt6gW75/3eg/yMjg
6Yi7ThgR9jf3giYB2BoIHiIcIqTjNoo7U8o45iW7iKp/VT6iyflxdRLoewlz4fwgH2HLF4KLwW6X
+lJJFNO3RFWF/5fiaNgtwLUcSRZR684UkKnGyDYRmTkbDTK9mkmeljbSkYLM/wLrCXJsGaMl8qwX
KTNQykjCgRN1Bkda0aapv0YnW/xFfSsQBde6wpfVF0GAjHMRRkD9rek73Woz1XfofY+dAGNaBvcs
SZsIi1/6klWwM8/wU+PoinzQZY1eSF965n/TwxU+8ZXxQc/kDfhlsOKT/zUWT7V96OtXDn4ecoZo
2UCgsYJgVEkv/0fuUt8lu1ZuHlcMYfkjrLxF8XqO/JL9e/q6/hrtgArOf+sqMf5snsDep/M9LpNM
oXA8vGkXGks1TfqbBl4F2Iv5eH73+XLZ5p4HOYneRA3ZtxC/L84dS1IzkuV7s56UwNpYCWjAjSCg
knrhehbRC3iRFW+DsXO+x0VHX4EX2dErU1sugqekt7BZChQmyUly66k1r287WWGkq+tIEmXIEeCL
BErraddP8ymNiYtSJDwjDsxPcLrL+Ed1046GuH8clJ9McqVE3Dxb0BSSbu4pHn8lLk5v+m1FWJx1
+LQm+oqB81w86r6NVEgnHQxh67w81+auAGR3wnYNYlho7SudC0iK0uKAz2E/jHa1FvABXzAOJvTX
8EGQ/h39J/CcJAhCkUfYCno+pU5gmWgxOviIk7cGXEyND+I7F+fW9LeEn5Ax+fdIVU+b4hTa7+O1
n7OIEtGoi6cZ51oJRXaOhhq0AfMgF6l3K3MQ1NLWd1sQ9AErm3LKTWYpcN8b8h3UwaWmNkBcQxBd
bbbZotuCuaLBkUvbo+uGHFKKwvRAdEjnE3LsHl9MX4j/Bmcz44Da0bvlZnoPE6nZi1G0FV1SIR+C
8/xAoVQwbcA7ExFTA8ANmzLLREpZqm1MspT4yA6mt6QoS5aBwcAT3gokAx8qZeDpylDfUIhk7Vwm
WKMtTPi5XlsDdoWBJqu7rWaYeGMDC6m2iUM4iQ0m/uxSaTnBsEcg03Sa99XufKXbe/H+8rIs+v7c
n0+irwryK3dxAGFJJf0olunRLuApI3jfJxrW1Q21RdczphhxmcDjnHFxvkoRjbq8O2nppVLRtbWV
msHaRkUlEFi6xXKBN0PHMmb4peD817ObpIEL2YUZ9K6yKqe2GyG++FXxorSo5rTbb/g9fO3Ycghi
+cnBPLLh4L1RqBzkcNCtToN4EqvkA57GDydfCwCiPfJUJefLeRVXDEIgsSSGjI/++m0CVCqCsKO1
ZTVYT2EPviS3aAI4+vtFBVIk+1s7ZE6ohUWhQdCJHJNHmVA0TQ3o/JEn5Ne68nxS1I7MUtfj8tOI
B+s+kvL1NqxQRpcedbTfxvCYhd69JBwSfG94jtVf9teJ1TIYXi6NzZLx+SVpPNqpvP7Gpels0aty
+JfFpg==
`protect end_protected

