

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cJ9uuvmph1jKHnJ51H06eO5xJLD2E2GBNiSQaG7P/dwfiZIp74ayKWYuQyHobWTwaGEZCCkf7Q+4
q588LXVT+Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SUnVLMGAdU88ORnhH8PZWn/lqGOLeslgmsYuWOVpHKCRRN70Lc0BXNIARhkcUAM7LFX7aOpOF6Cv
QEEu9O4c74tBOhvgd/y1NdC10Qd3kR6DzylhRTOzg5GywHRI9pgEEctM+Mh22QkLK3G+meUwu3Yj
CBzrxnPuRSTET+W+gOk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
13eaU6Sg+4WJ5OITHwP72Y5oXTC2HP4iu+eCE3pdfpGRUOrflhDSmziW1ytsADKAZq1iZ00Lg5T1
StgWKNr/a4r9TU96+L0eAbjBW3X1W6OUEZa0rK/R4dNdVca32144igusHNiM5n04r+zV6pgW1g7w
xazh8ZMHCpKS/j1lDv85PKjJV6NsnbrBgCFnWbcakBlxjAYvc64TFCD77HZ9bEPBXC1k5rMpf2ku
VUVq7PSqlkERhtk58TffRueEMw55EcT+qwtoIGCm8QylPc0huI3LmbpHoW7NlmowRyUrJ7nWa+Ld
hcyH2kOpGSrBPYjWUmR0J1qkGM35R2+6Xmj26A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YCquRRMSVDoS3CiUYGVLeD+9mPjt9AW7TW2bB8angCB99ZxpnrrDAN8SOlJhyn8B5tX+NpMQ9yGj
ZSWgOZSleb2ih0WefXQ8OltF28ZfzaEsf8mUexR/W+Ku7nphq6XTJL0qtIfxxCn1kfj/eEkXECB1
CuxU414Ebx0X6R/ywaDEI8gIG/0AAHzENrPkvjaXH8bn2bq3wsHQrLkPRQh4Ngnw1rvmnoFhm4jk
cmrWWvg83RPMwFIcHxZ9M3g2yUX6d+77OnDqG34YXH1fMJgBDRCAVHCw3TYsLKHJ6+UOsbnnMuuf
47/MB2//Zy7jHFoEzeS75x4ZbXhICqqA81C3Fg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FCb0M/ZbiRMj3Hk+SVNddysGGZJEYiCxC37EHMDYeuN2fLgvgMwZcuMHlU1rU2E4XRbFp+ZBFgzb
Ey2m12dInVtlCUQWcdvEd8puN+XTqHQJMXiDjWroc2i/US8wffBry729CZ01iLefyubFoaVkITWK
f+KdFwXGVXLWEJ9fsKc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GVfMjRsrrSS+qdjeL6E5Gdj4t/CSIURBhcR6ZHRRU1eeJX3riaNrm1KT19BkNPmRRSh5TWyPNjkc
ZiGR5UAO/Okgco1e70zIYF6bMh203Q/EMmijte0IMz3b3lNZXR9OobLMgYKyyOlCoWAFJpzejvu5
ZZD+euimAc+4FLmXuWghTw7pZ4Zz3nur9efQuCvnePlQjaAD/gbDAKn4wg/yLLkOgbBkUgcAtp9N
OdE+OE1ipoC5j+7q1fF4+DnxJAZjqCA/MKNFjwzxPLqVmqBo11g3adVKlDYpSvGBOxlSqUHxDenE
qcOIa1Fs/8fEtY2mw1BeSlNFLZPLrD7ILWi4Fg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NAKZG/SvNL5wedDqxYscfqOuv7tomMRRCUtZkyBWw63teU+XDZnpZwUECIamvdTXmPBMZvATYzNs
trxURnffffe6I4mqEKJVQU2GeAzD2Nt3RGgok4XiLTADAelNoxYBxlBRc63Puz5GUoUETvEnxGHw
XMp1SMrjg4ZjdIS7KKX1wByNHKPG9lsaFhoBKhDLHxKwOpJYQKhUh9Xvr+d1G0N/2lxH80swtERc
9xussNkogu42JVVlLGT/VfARso1lQ9XIaVgbnjU/OerfYXxoCZR4xNTKoLen3zmd5k1wI8UKmuPO
+So1iOjwUlqCUs2ANcAogb2FhPaqhFmbWHQegg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qiziz32uC62c0pwLnvnWs6dnzkvXMNyLh68w5CY+k3Ogl11V+WBbHaQ18kXtPFIdy++3a4vw1Cbt
2Isifrkzj5xOGK4sC4hDSLLoZU5j/JJJQFmiqfZEd28Vk6hCSZPQbiCOIMxkwbpGDXyx5i11ayuf
SIKS9htw9T5KlTxU0J5iAZ1pPpfN0eEV1DzNggu9rDZAHOf+kYsV3j/xyyvz8EmNBMgJMv/oIOLh
xChyCm/0N6YjI1AW/51mSazU+z5GMgYBbX17sTpN1QQpE4WULtCGgbEYLd5NpofmfNRcTWjYOFG8
XlkmEM9Q6ldYtI+TYWmxqQ7pssOcWyXrAFOF8A==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mdyUk2rJsGbOkHOgSxG9f2rMtNhvZ91qZGcfP5EjZlnsBtu3w5GUbUmoUXqbCFXctEIxk9mwrZnx
6xgA+E4ZAhO0Ca9q+rX5vwFUvfJ2zmmsY9MUi717nJ6+2gX5XMK1IA/uzZLkucnGnqcf2ye6ivsK
6OkxGvpAWL5omj9eqfPAbg3ProcRadxNQSiI+/zdinNIaTPCadaDw3B6UgKniTvjOc/SDXshek59
53yoGMWpFBH79n8ctjIoixaiprGTBIX8HLetCKm9H8pUeJEsT2lYT9P9tU7BTzNL4I7gi9AXuwuG
m6UAPhz3ywthY55L3q05ZuZp2I/P19XyyOH4dg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 121872)
`protect data_block
w5ospHtErDZ6tDAj6HY6T2J7nyBXiBrkbaC5ACcCwwsX0Z0cW6TZNHjvuw178C8oFhTzlXmQyI9Y
uH10tIcCcw5BtVxSsMwm9J/cMf0IPBEsnyHaIIrJJpe9p/EMCI3EaRDXbNwjdzCQiV/BUPt2j+3L
dQAkGx9pvGu4bxw7lOf5ujAkVDXRvrYAXtqu35ViCKdUHCRIaNmOXgKJJlSLBbtoyYV2UtuY5E+o
GTdKjD5hPUeEdPuPA0w0HUkwESylycmH/u03H1iPSY8VhH6n4g5YsySJrk3ciXQPrwKyhgEtVBXj
1ofLvO37k8RWFAnS1f5RWhuJC+ihuA1h25woxwCB/MEzgWdfPzwci3V1CGtGJrKmYYIvSqyMHAkW
GRamkxYpAow71geB4kkoKSgh/JV3QBvMkP04jHQRHW9RK7b5wSo6jLCzrJeUgNHlRrrle6P1X5Xj
mGT5Ufn6ifbftFZTyNfvUM/OTsMhaIYL0bNkbcndfLxxhXx1PvrMPPgLhr4rvRQUCgHCJMr+tKSJ
FiiTidiMPWQ3dwuwqyF/ZaHEmC3GXoiCPaM22s2903aOS20aE2985v4rsv/QVVjbFOcggiQsrszv
fAVArdgRpx0jWUL+DkE2pkzEfth+z3TdTncbj3MCF63v4xlEH4M6YLn6XGGwcDXoneVI8WSjizSI
3w2ytfxk5K2pS8YSscZrJ+cfDV7S7ay1lAg6Iz/KW7ak8C800AIYjiSchamOH3r4piVqpTLpNLi9
+pznAuL1RL50PIYbi7oRQP3x2oTulx8xf22vipds6FXKj2mWf48i9mrwhMRnqtYgUGQm4pvFR9qh
pG58u2pNQNg9O/UasMP8ALkhRde85zo8tuzjHPAqEusRPFqdAZ2g3y8vWbmq5dApf8Q6dI90R2wh
wp2DyN5hDNK4q83awygqiHMrEE1UuaiFJOmzQLjnVAf7GBBIbx/HyB3tn0sNeP9WNS9tqhbzwEc6
se2uGWQtijauLPN7OY/RKmzn0mZGkBhUlq8MEoVufPZdTwKnx8sri94/YeLoX9dNUqpNcQDlkhlt
1lgOe0xm1zQPJ6Vork2yw+3zYWrK4ri6wr6lZNy+tm2XuBL3ZJ9RoeJBYSzQKcdYnb7bxf+7CNv/
MHGqKrfg5iA7loY46clnc28Eooq/K70mZmCElmd/OjHP50/Gx3nbDEXn0pTf4IipjP+BpCQJNli2
qswqjsSU3BlHYVLdQwDPVigflMazUPV1jaRbEEvRk24pDA62DBC73PHR/VbHXk54D0xOl6vft2Xh
QI7XUPtZyWb10Enr8dWIlOZEfz9l69jDRenLfP0uAskcvZZOSlV5rDLyWa1fJsVUpIgSg32IGkpX
CxTWX0dLVT1MQaUpOFLVx87ZaMtK9wEvU+2rZlkurpTsvGCDKTNX3PpaOenxvmr6A/2rcneZ7XxT
Nzf/iiQZgqftF20pawJcGxa3ZNz+SBhx/e042HRS7D7hRTShTS4FBygcEd3mBEfLPSHNk2aKxe7y
K/ZLBZUBg33xSWMVcswdmvLkkMRe1Azn2F/I/VWszRmSrPh359mZmfN4ssm6Kw74gloYCVsJIdE4
rZXlA9n34Zib4Mw44FJmwjMcJzi3XY+WJrqIiUH6jHnGtteBKchlJR3ND5CwfbsJ/1SslG5oGl9k
9+9fNJcG/v3k7JooxH/FPRYt28373R003jz0J8cxOz/edOtx3P1yu0dY3gRGo6mNj6Js0XAgtWln
Rwu1hmhLua+sKrD1IBXbzC4pxEepVntpdrV68J1JSv14omhHyOVXN31bO2XprJ4As0vI86QLRUCU
1pwdoLih5ruwOhYTtGyqM4dLhpPs0bggGb669UUB1qa8WD28IMFBo9qN/6RrlaAZenTtQgNgy/rP
ZBX02xvFXjz+mA5eHa8VCspaMrDpRBV5pXtd4FlTuapfbnC5E0jDcdIjYhOG64DtPqAIhL71Hu8I
/xBNHy1dX5p9b2MGBSWkesYdVZg1TZq/AdJew6JftODHqqXjpX4fwn9tEmujqtJiKykyjZ3MXHAQ
mwnamvMahsN0QuYyx8AwDmcdt6JzAPUOY246iSkcToPbFuP7dkloc2rgBJQ3WSOeUJpFnwuhoTcf
FKgTJAe6Xv1rm6VGIL3utmq//kJQpFxF/jJnDEinuiaZC8I2ei5H2LvWG7vIFv7G88WBicTkdxWT
VjqlA0FTiTEdO3K321NW0taaU9xHuzSM1Xk6RyEiKUrtcPbhZsAWm+h+oU9cFuDEF/sO48z9fH/d
P0M555VIbooL2xGK9DS5wdEoH+7ysx0rwzcxIWZuCf1fYlwqg0z5KKCPtRwGfnWPjXtHL+dZ46y9
YF0ZMT1H74HHcbnCqY/mLoEgo/zaAX+kg/y0hwlzAdaAInKmuTphrF/XWbqC4eptNz8SxmdgPphb
IXuopi/LnLZXdWUcWQImsunJyhopzxER/kZem9REv6i7YUwqt7shT6OuAYAoRcOfb5tZh4+w1zxU
tnDlK27uPV7/KCHX+a2CB0wiZaWVa/dTlYOSP9Nkqgr5sbn4t77DrrrRB8z7o+cJNPjhja6H8rke
wfWDYQEPAx2FARMjI5rkVfoBIYlT1vPBU3kqDKhoI0QAY8zdLoKfUN8l5kADuQEBItxmt/1vqz7M
7OstRsCcamFbgqRFit3scISQvm5YRFpAybqPDFKIERF374JTuvlFAAuFJwHXDT/mEHnzCRungBFp
/jWEiMNKwZfnPEFbkEXXSFWq3MewRFeOr2CSdHA14dizsjFrazG4EvyJaAsWmvdyzHWvo1O+K99z
EE1lsqU8Z11JEGAvlJFzz752yIDtjKhzw6nD9vrFGtE3qiyHdMhGR9H0RArankdBREKEMcCej80O
r89LSlFxE7J8zgaYtRbPYjDRAYTqPGS5P8zsGy6OfB29b+YBBGdCKlamtG/dteBA9fqrHC5kVcyv
e9w9e5wuho4+IcV69YXVFHyp60HfH1SP0luf3M+TxOtkuqmJ/+vbwLdzfQQhanRT0Ixs28qYtnp5
szaFJp7Dg+su1+4c07HIQAVlrJtt195LzSBdDDh3vhji3bxrV2pp293nZom2OzuKtC5YL6xBivf8
HVeaORsVhx/sgrZqbjd+rTd9FuTaEaVrZKELeG47c4MXOpD6OzQfGyKhLLCu3iZ2OCNhpLjiqUSm
Ptqi0QASYIOnZ12SZ6MdFmcE5jkuoIXegb6J5InKBt27JYDpTng5s57ezSLrSgLL3POHvc2J0oYq
tuRBOgzZguKdR6/7AxqwA2rC7tPFP7FAGfjv4ZvMnRruSwwBqe6qPnBnad6QShyH8PoNQm7OSv+l
i+WeD3mSUqhl8D/9QJeiMbtqPinKp/5sEssyQGAe+9o3cGsOiyTb7XILRwZWfqHbzwG4ZT2p2UHX
L6/Kpo/rYH5lFgAZ3kH/w4SxFKOSdy8oD3Igl2RmSE6mhdPt/vif6ndGCMhOEFrQm9yYK9jQAWf+
oeNZmeBQbBL07g95JlRfjjD6xB8UBBCZ4G5512J0qwDrAuMQqeuD6XHDhnrG0NqqmnVOHsmovLo+
Dqyh6M5j+0oUAgoh557Nl65huSjGAY/wCtcDOg2IGp9IpSnIwQXQ+TfDbLbBnkxoJLlfHHmX7bah
1+F5LdP8xa4ieiDWPHJvGRAs2HYtoSfVMFjglRB6/NpRCp1CCCgkeHZl6ndSkWF942GK0a5w4Tap
f5j0bvVkYFdniez3i96FReOkjFpcYAWPxpVdjJ4KuIGO8yxJxUkrHePFxN1eFnWYAAMBuh7/jNnK
dxKt0GEFiGqEgZkc9S4ONoBPzpnYHFzDcglXrlFPno4dlWaLWmd7ANOF4V2fLJC0WpvIWUr1fpLw
bdFFHkA0c1oHMMAF5f/bVAO6b76CakmGUEXy2GUembVY2hJi/HB41B2YzXQT/eKKwDDtZVyHe3tz
URE/yJA/OMg0onrOJGpOOVZ61S6vxcXGxYS5K6VPQbsOWhxTtKqP9gzkIyBNBYYWxHKw4i9xzEwD
ZRC4y8tMYlCUxGuCKwR//mpxPDL8Ev9Q7+qYdRd45eQquofjllFBYjZVWJWdrQwi+r0MNjQDbXAK
QQ6kz7SOhA7ym35MzzmHmaufIuQWLE0wWf2O5yllGpvJPP2szVlR2o7osSAGCb4TG86ejdCi95A/
PR0Zk1gvHAtj1p4fJ8HxVWC2O0MddukNv6o2dMeCeYkVY08jEcOiJUYTIaNDvXSuynFjnBaJqKSX
Dw6oOAdkVtp86UseAGEOnZ3uBA+nJlRvRkxFpcduHcBrC/9lxIdxT8eIBNmSa1eGtXiKJXo4xMiP
CuxacDPCJrX+uT1VgYLyFOzkceYm1edt9i+pd828GmWHGaHK9VFe7KoPCd9zwhXVVIf0bSxBdD2z
jBQdT7qdSas4FcKVPUtzG584V7r8u8DeBWJddj+HBwY2wY0v3eEWF0gU7ZLVrM/EZ7shDmjZ9IUv
l3cMYtsGO0wfgRF0Qn2hp1HLLUmIRKiFVo3MvGu4pUgmdDgc5lgB/Ae+X9ljMbjgNQNjVnh3QB3p
F9ApItWK7TBnSXc2Q9vCugUb6cOJVAo//yZY3g8+1y0+4XhaXhf+SYaRzm6f6fQwPIzJF+Ao2CJo
7ersli6cWHZHyJlx1vWPcaBp6Pr3wG8KPm75cbpEXoEEjWqcMkITJS3/ICtuF9ff6bp5LorlOHbe
Ofwfgx192CClRnMZ9WRHyPIokKdUpED4D1ItOIj947f/Ye1/0tIj9cs4ujCe9WnGEiSB48TMhhJm
Uo95l7+Nk2XCX8nYJXxAD8c63DAHyM08MnEmukHIdVlycOcse0fOtFjsD7MgzxOQMEq3bRwT7ZaM
YMb3lyrYXOJv9ak9nX4nNv+GC632M/UwI/v9/u3eRrzFAGPAFy7Mwgzn2Qqu+pGLlFCvpys6O3Qo
1f6AZPYA97i5LxhmML9HBveEm0D9h430EUullJYoOqOx2kPudpXM+3xIy+GO4Pe8GX33MrYrEDGl
2n6Fl/0GU+bm9SvPgCA+xTICypMgugYKpVFPG3Uip69BYzTxvbssBHtHZ+7EqXSf5j9CZHJ3ZSim
ZHOSx5qw3yNr8bNb8p6PgPaErLjUS+7ro6v2KmH7iRoNU4c+kuweLJCEgN3/bIFwB75Dnf2mB+2V
qyxx7kjKA+Ppeu85PJTpl8cFBMay8Bv+vlCd+T9a1/KXskyYb9z8CPzOmlzGIDJf5k6hdf2qxiJo
5v8K08yhAHHsWyEnvAM8zSIw1+wKazAAeZAuwPcRwB2Vf7IeAiNM7R6y0LRTLBRGfkmCg8coaWHh
aJSKX5qc4pqAZ0n9G9ci3CxE6ZJ8izkHN0bjubozHiXIczklMY/wv0YDT11L1goh/5ygWxfjAQkg
7/RIHdUAcP38RlqlPwXpuxFgs2bUV8nIKyVwgwDfCmxES35nHw3oeemsANDYHvlY0pHeoGS+Ljjn
bw8pcwXP0nttDyC9PZEV8oxPRR4dFBLSBBDnYSt2s6Kbqy07W58YaU5oP2ToqgXHVuyADdXWVq0L
M3R1fXChNYvT8oQRghya8gVlWliQT+vufYOSeiNR0H7U/vQb0xISWHz4MALbLrLJBlffpOwAo/8C
XsrCuz/7qAU74cD4RKbRt61Xpdzxx70za1tkYd3c9O3ilZ8zGRLWTs10HXxrud8nFEkRcPzwjDyz
VVyma+GzKiirJXCZtAiZwUSAOtDU4THHBEmC/NGSmz7ZEaixMz5HbF/VUDZCLl8z/1S6dSjnINDC
i0WQfvtFnDwalBJsyF0yavwrJSwID5J3U9T57O8KyRMrCrhkUS63r0hVHWzuCOvzwRzhcylbM+MI
LTFzu8n7uArk0GbWh4w1fa6BWmkJy7fT68I2kbGUDeCgq/OavY0Zwcsb4dasS92wWQsnzzCY+zVR
6eJRXc0DvSBpMc2OG9EkmoNaVG9kbGt5y7GbY8EIBE2yQ+c8Ui4GmydNTrOOFLP98wDh8NagfC4K
uKVAM6mH3nqmuRjDujRPi6MiErNVeNUSan5Y3rRo759/f3m4O+fz5KjeZExm3pQ0vqrLLibNoe8x
gtJ3Xl3P1KMdiJrCnctGNo2fIldvXO1DB+Fgej8VIMJX9/cCO/o+W4uMDbSQ3HZ8W9xxgWbO1Qwx
NgDXvCOY+lijYr5zxWQBOM6vbu/MZA3PTMcxE3PmJwctnxMGJBsSNLNbfaymjWgCBJ+7P/Ocz3N6
gnl5SE4z4YyW/vbwvCQdjKyutoONMc3K0b4SAIOsqNYilNi32f5NCEBpmGjUcqpEgUv1WQI4QOD3
ybK4IUvnISjtGXgpdw/WzAg4kKQBhBpcaW50pSITJXlbMEZfL4As/FXi+JkOkXMeKUQK3pKYdP9d
uQ6MR1L4n+Ftu7+ojtkkDyobUCP0YViN4JAek0Df8p+6oqrF1HO/ctR3JTPVn9xQvniA/6LVnh4s
alVVRnxEHgedhU65bBKkBts/ucKPP0bTguWVoLSUNfrSyKA4uM8M98fTsx87ni+lFx4KuqG6axgG
MOhvVh0pbgENhKglIfuEDHHvxljVFvXBZdvDEYooe1NP8C+eEqtRv5LTOOq/eP06j512bbZZP49P
ajf1Jw7ibjHRQ+6Ev/GQYA+AZm4GQxa3wUiV4SJLkc32t7XNAcgeWDYyhxgr4xf3WTwD5Qj0Tw7G
1k3nenuf82YwSgJd5H24ods8A7zjp6TH8nt84xp8xQnowHThSze3GsLWQ8wypN25caVNQUSKdxVv
eVtbK3jZISftqUgEWXg+pA7Y4lPlpmwJgSiJefKxQLv6mm4G2MkQ/wz/HtlZQwg8+yMN7n/TMuex
Y0YhKclrfa2pA8/t4XrXG+MjXacwQUgcWlvBeRnC2iU56Ns69o4HRNuKz3i3agftzOWXvC+OvM9J
YQw/S3eJGx7ihMXeQFrlZ814hPz57iIe1U8eXihmPxAQnXro4014m8AMjpq1y9PkjG/VLpQzxjIV
nJkHUN0at2r1f44tTqnQ532oQaFHCpCtDZRo0LLDdaA6a+yoAMvM0iUCX9AED/AsR8Fg5lfLDuhT
eck9ElgJINozuXEuUM97sUKTtUb5J2JiLQv2dteVndscqkwiVNbLzpzniaEMzusga3+nIG0npdRJ
g9P8KGb6UN7CbVrMSbB+i8uAU9PvyuuP3oDPuswLjOfKqa5I+ei+RbeGV9Kqu4mzfYLNc5GzGPQV
tzoSWOFfM7WUJBTMP52X20xqGcaQsgdUZIh2zok2IriA/WJ73Sj0UhenqxX0OtbdavErfz8y+QvU
ma8wcEElbeKqkOBw2kvUOmrxxKiMge4FWzDbLti6L2maAnpIaWqHGl7qkXg5XMaVjtlt9ksbJBSC
xwd8acZ/C+BLguKwVa7cT3DJNceT/b2hvwuzREsX4VKlbfKLLBrRBfuH4l9njW0e4Ksyl8J7jQyr
Pccqm9dL1JJwuhb/RsgQQguvx6Np9Ls+yz/s3VaQcAfl4VcQaw6JOaudNqYwX5HwUwkis5O4Bs3+
v2wc6mxiJtvx9h9Vb2gdh3AT6UDk9mLlTJP4QNy2l0cM87cPG2BJsFY+QwtUeMQhMitKzpD+73sb
0VIhDwnP+tnxp3zJ8vGQo55tUuUiohPO9KRfqQnb0aDxrO1OOPkQYZSbhReZLykbDLmtH85JnJ4J
si/NxHD8ltXf88V1bVWRqBGfDl0Ey3WwlyZRLux5E8wFR2uVaGh5AifMcPYHEgMLZ4HpnEDPaKSl
XAfaVWZSyu2LmEJPXsLvCpvlbuKa4qQekeAU7N3KnlJvIFnutY5hNNSJ/P2X5fUaFpFI6RsbnexL
U2byaPaURdp/jr675PfCIggDwjLZkQqCH4iZhTMbtndo4R4b/aDRatXNJ7E7yYARpYL+PeJ3kXNW
85hbx0AZx1TDuYjJ2NyTlwJ73VFve9vYU0AETmbqOmKVbBtRMR6eaBrDzOnIoXzoH9ZIbuhTTEi3
3A2kVtwfe62w0oQgPPeB87zqzniZgo0tkbIXwg0iYUsWiPthQGNbc/yHFIfJMeInkBZhjCTCVXdy
AX8NXE3yKhZGW8xzjJFknh8rWHroQ3KyS9RyGNDW20a+Eq10EHLx4wOnPp6z5Pk3CEdbnr4sPsQQ
ONfRrxnFMcAfOmuyrT0rwpXownFy7HIot9Ph6V2eWEu2G706Kt04vmzMdrwKPsr+1FHh51zE8fw6
eVpALkrG0nUelvnsGfdWtpTZ+/OwfYtq+AsmoF0A4I13HYfkQ9v3iKlBfvs9Fr4ISTl9zOWEf1sf
E2pp0Gk/jUzmeCGH0Hgcm2p5ZMx7BENRCwgBeqQ/HveaVoufQ1RR644UQJCyypSzBGbESgcfXtW0
Z3CJg4bEhLx1zLddpNJYeRur+RklzjU5FU0U3nvp3/DH/pkEBMZLbBXMaBx/IH+WWzJfMFW4zuYt
Wq+AwI2Feg0qOPjSdmT/4D6lFc/oQu5BpJPBP3b/Sw1dZVQ4VVA2UtIKnv0xfwG/pKZ/qbgN9r/o
udhc3E3q4QgenypIbeQ8oWplsmki577B8xshBk3pdp58+yG/WH9aH7kSiE/Re4L4X/tTuUXWZbgN
Eu1q3o0AV72Dij55f0H1grZqtFuVDggrN4zPpyz1dwv4FLaC0pSvhLHKqxWnup+qd+cGuzu+nhXa
ywtHcg8cwiug2v9++TgcEzYarM16sgKTcdlYshgTtSXm9NXc1rv8Nb8iQPRjP9BtbkiuJ7RLdmqj
d/ClmY+1di4ons9c7eAdDgQxEAru5VAPvExgjisqY2fb9jY2dRJ0ysQs4MOgCO4MSwsdefcYrt80
TxJGtpZwpSwdhnJFgirVqLnEn8m3S63FXM+5AYlo1YwGC2QXbW3+ZaVNh9c1WD5fFaGSRNL+H/xA
xagk9M2Mw5orfqil1vPJO9swFUtA8kLjthRWDnn3hiiuSzcf5iCQNRIVf7Bo71APAVtkzxdHjZh3
hHxXz+SHba/aY/izBegdcrOHuKQT5FISwLbU1OSwtD1Kvz/dml+3wPvlat/wRIdizkPIi5SSnkiU
OmKAHZt9WgbgaAbf44PzOpgBdAgAa3A9BB/1MhpHrt+5z+oNEzM+iqaWFWbdf5GHLpkhf6XSgt22
IyEWsDvFSnTWXIe9J8CdwnkP9EhdWNMMXffc+dQ0e5wToL/qTDXkb9XPZaxFILXw9+K0Sx5VFRHU
Lc35eEfvM/TOsKNTdvI34uNxfeO5mlzdQ83DgY3wLA4h0DlHBDMYofKvyXZEfWcP9Mag7lR613gR
SnFHPdXFhWHu9eiu3JopURFmpan2qviKEh41fJyHv9DNPWoY+stk0HuK6mNYN/ou23lLn4mnL1rq
jxp54smnH3rGGmILfPAY0K7ds0nZ4JGf8znJVDfSzBOGzCwj9Cw9N/SiGRL967Bpc/AsUxAzUR39
XB+5haWNxYHW+AmMyfs9NMjqZoA0+iTrOzsvPcOxtwGTHJ8dJ4v/iyXxQbls7b7Ier8CO+CW/WTP
2iYWZ3LuYdkKweI/QpNoLSa9+56r+fVSXYFBXaS2DWeSNCdEgEZ4CAhsVBzy7Bz5/r2wdJy4lCfm
52fwcYCK6Lfz8bbIEuvaSRPua09wf0ZjJqJwEMbdSPfpaRLyndu4LpQm0i3gci/mk0prhFmPDlbb
Qykl2W/dvANZpYIjDukSofiiWFmWyzhKSzgXC6p4OaAEq0Co+RM4mMpHLwlClEPzdH9SLe93F1LZ
7mlNrakzQh/ZWqnJaJ79FBdSnRSbPKDEcZvYa1w15HAFS8+4wkjPVQkXTFer4L0+oz/lrDe9CJBP
tWq6YOPoq7/EIs04OMBQukznMojExdRS48SwbZ7of78THyOoUx0erFNGZZor9NatVKBXzo6r2bL+
eEMkwQddbABWW0pQGaMrGKGusaCuLtgh1vDu6sEarfH2Ni46f3xvmsAhH2fPlFyO1cokscCpBbfc
vQ/5Dcm17WHrn0XSVByGPzTlxdiD0xcXGi/VGO8sidvZyiXI/dc6uJIfJVLqRATvDpB0UakjlrVT
7XyTidfL1zxPSJpPMQvr1jJljWNjm4jVVMf+yKZ8NnuqXA1JiA5E5ejHbGSYvmrfaBl9D+r/4Rj8
OIm+dw/YoZrD/sTanxFIfxbtemHeQnCmLQZyM0Qnw7c1uzvz6xfeHiEbV4A33pUXgdYDnPh2ElI7
pVT7jLhxwBFFAM+c4NDL9O+GlTjKmjsD7qywasz3D+RzSMCeqexjwSZr7u4hkPfRm5yRIp2fmBjm
jxN+2gvKzo/cHn4vuAWWcRL74wcqfryq/tTAk1pQRmvY2zyPA953rWf+5gyu+5CE9rYiR8Kbe/oh
jhGcn5kKr0DtFgt4CsERB6z8deT1putiLNAufeRPSPFvsyaH4jxd3uzoVdze6Y6LPBgX+g1OV4ng
p3i+huO8E0QE8jC3sQeTUpAyGE7p4916lEvv+8Pi++JLiwTz2jtZGHjZOSQqAq7pJb06fIBJOdID
jMvwqV+BFSlkofVc1JPz8QU+cdhMd013RS6yzKT5Dc5DCwem5IxEJnPtRAvQOrGPkvXdVPBEjF8O
QiCbVcSYHm4ThL05IQ7cX0xh7+K+jKS3uWHCB9zXj7vbA8z5pp84WsH006lknqSyNEttT5tWm40U
0/VA7VIiZg/1obv5PCZlEDic3pT1tjlfZzPdL5nCAG7Z9UK9/mU4UVjpySzflAjdW3NOyrMNJsl8
GW7/uPoFaZKMRWxhU9KtM3ds3GaA2UxhyQbIGb9sOanwdfI+5keiQSvL44O6RCg68tLNX39881Ux
cKIAaOIjTPBER8t4bnY/CPQ6I0TSl7dw014E1hk6gILmpBvL6F2PV0h6KjuytQj42QEXvGPaB1Yq
C2dSRnFkdB9/w4nL3p3ATcL7mVRNLUQTDquIgkzZxOowvttLluugJbQ8UeqqVAuzMqrnp5rLk1LN
QKsYoRzt+bEqMwtiaFwaNvucfszx9QhQVp3Z0agjrQ73aSDbXoPiuKD8vwCi6Q1pAMji4R+pBhWe
xSZEzR/qRHGxify4PqMpRXC850cSUWgx3r4GUL+T6I9/tP8wmF0KH9hZVnVYd4UWTEL5Tss7cXpM
RoMiVzKN9usw/aV4SmzSc7qfGncvYNi0pVMol/RV8AAJu/dZ83reVC91+r7SodDuhANyl/DEgtON
oK3S+qAffbv8UjwKKtbDPPT9SSCAOZiH6vA53xsNrFV6dUnvH+p5oVZQ3Y2LsGaS9zoDiZvnt5gz
77emxteqcshpHzCtDm4jfkltVIMF5hckfQkESazARFWzfIybG/OwOogVdiFxoINKfO+/ka1/3SVR
00F8nidarAykUzjzRDc7ktTePKF/r1xUuhkEkPLM932UduFWNtmuSS6Z4wvWUq0vf046y7G2X6My
9H5vIiXcQximD5lbUliDqKy8pTZDiXLwI0rkzQozMWEY4memWMrkoopuYsaE2gVbCYpJAb7KTVq5
sLD2I7gErssOkKaMUdX+syaP/mH3NOaXtJQgw8B14ZqUM/6t0G7wf3B8TtuwLX0itVoSJW2SRcT4
36WQkE4oKIs2ObVaJ95bHwrUfB08vg8U4g3p1EXwPVwhmolSfVyPjtF2c8oW3x2iAIIul3Aw9aIC
6QFnw2gUN08G3oV+FzEpfVAyCzRWnP5bIhhEWrr7oIN2DEp7NacOcPKBh0O3REw311KzmOJa2GQd
spqMsMKTI9IZscUWOFA0MMlJmPLOd6sCuoUKocoC+OvzQHaNZmxHzmOlM2esR73LhreQzXfixahc
BnSplcY9qEAzP1ztaXaU8+PjvxDovyGOhaxyK16tp6zVRa2J+jPR9QejoPRYc2uNv0iONtidTJf7
js9jzxUwNHq3JvWWIOkb/Ug2JNs/j17751D/VugymOIcw+45U8coRIqDUKsKzv24fDoG0xIoP5Hl
jn+avDAqR9v5QbBTiuRkkS5xOn/iISoIYiDa+mJAuKOBabdHarvXSbfGu5ZglTSUmjendYwdeXSu
vnlgjXFZM8qqXPWM+FK+rHOD1FQ9/hx9//PZFBtIIerumuZQFTjtHgh8IQAyQqRG9zR8IgZr1VcL
YPpt2Yc1P8+IN1HvxI5K4vK24nR6wBD+zgfUQ8AotFmjjRfzX480aDRcZAHl3kEtCuOqU2Rz/f+r
D9tNAQEacU1SN3qP9O/q1jRVj+u28C4Qq20K1ae3+QYr+lTKxb+8WGLFtMA0itfwi36vgF/n+wFH
1lz/siW3w/KLvicEn1uxWCq8tdh9OCuu6cC+ZNi1F0gnyyfTaZ7yrW9oVQ2M34H4A7up+pw9DOjM
MwU0yYB95DALfEgzT8XDr+BP4jQuugMO3ONrmP84dSkcVnZEXB2hmTAeqIdHxeFOZ/p0vGYDO3xq
CLqJKeagOlIHFh2gqLVvstCyh0UrbvD8hROwJNXG/1/UOYFsZMs4u7CjL32Lnt3KwNmG4YavHPtE
4Xso4ZDGTDaVJUNAxYLOwnHBjMJjNs9BlqAhYZ2mjFXfWWS74uooOYeMDem+9mwL20ASqu8nUtnU
UfDSd14G8KQRJzwFlWArvC23UohAvvW0GBqq1jlJXrr+LzxBDBS17H2jvdO2k+Ya0liPYUsUOiDF
4P4r2KLAxBX1EiTzmdLRrBCRBOcKMpsHFt/3yb8Evjf2aAubPriLxUD9YfGvd9fbaIOl7teHlvNU
ZFmdaL+CiFmqjIhPkbv7VnClvGIMrqHrAPT6t7MMjLE89SxcfivhSEk2Lww8KeoVlsgk4n8bjXri
3pb5PW5zhTqvkwjPljDAzQTKHtpqxB+cjMDXkMAu2P9VJnAy7A7jsPvesKx+s5XZdY+9FZGNw7Cn
F1sCx+jHz/RfnsGVvrQFTkI1VJF9/pTqQVN0/rO5P9IDond+dMi4eh1hdb2sXV+T3Dmwt87cd2Rj
kRm0TvRR5zNEXd+CgE6Atfit2DDMOVg2Tkynjz5ceC10bNlX4yRn9Cpd32kHHQhL4xQb0kEdCYyF
n+JvUS2B3Hmx6SiYXbETwSJryoW3kZ5Clqrj8U0CroggmU+kD1m5r6UCyN0yyomFKQsP7TqUqQ50
Kv5gDaE/rtWmYL2ATJ60We8v0EAkAP31jinaPooMjlk48+jsu0E7xZi78ewg1lbq3cdW0M+ziUy4
85sz40Qt91Cxul2n9VD1rbsD2MVSZJ/NkK7SLbqgEG8Y+hP5q4OgTPojruhZuTbsM3nFz9PknD2f
9K/hKE36MRe7kvbb7NsPPaDNk4Jk7c8ZYQg34NEWOnxRqIzj+kQYwVoXlC7PPXjStM5AL5Tb31n8
86YA9EMOPWORsb/Nz6trzeERNvpEp6EokUIXCbLXrwfsry97j9Na1zmkearLLPlER4/EHPjTjpv7
jHX/mkKqlnkLxSrkc3BE3hb8MrJbxu/7PvM5yMqfK+C3zD3or1xSKROlbymBjA2HA36tKukJwCt/
hXVJYCf239bUHlLkhAJw2emtzPb0Faiaw+OhArThLMKEQWK0h8CDn758/1kkWh3ssL8vHfynxnvo
kzi67Gmo52SmQqNQgM4tA2PtMpEK8JXXT6R5CBsWc3J02oyElPrly7oPm3C+ujz58GiWu8zXNyQc
/lJJihKqZhN+zKuWmPH4oT3hdKDONm4uLpFYsS4QUKzQtE0U/GkCXFcLe1jRxsKUoWBoj2mskCKE
xSX24AiJf5HTZJlUiQPKCOpuRROL2Gz/idiaicong7xU37H5O0i6nuHxlazgsFdxAAsqPyaB5B+g
oAm+oxZarGYLYUKb9ScG7NVB6xv07DB5edEiQeW9UwpKcig1k6i7wjL5qc8PY7HE1PnocVr66Njp
YRq8K/cNtuD+FrZDRBNMm29Q2lXaLPed76rC1kecYXpnG61/7zW0yTNEpeLSLQI3tfyH9s5qUIqL
Bn4Qs8m68q/F7GKk5AEoQf/Nquu3KWH3V52EBzfwZVLCmDlC/p4/WttbtqHSQEAdM6v8ZSLnvwBn
14kVKFzq5A2wa5jEGMKxiRe6mKwIdkKKz6qXcfuVohbC0Zz84pNH6GmAlJ+WJGOD+dbKg+Rox0LV
MmnXKjEQQwoG2T8xDRPPChoo55yLsGsESFt0IkLnl6lMvuFY5oD01blhn0RnQOrO9jjfdFy+o6gA
g1QtuQwqz6ce6svkgIaA3nDP3NPcs1QMmXXfE6i1BHIdNCcX+glBMdxYAyoV0CN+ZQW40L/iUnRu
Z21yEddhitJ8RcLQWzOGo1Gbt7MMd5xZCJhsXogCVpggxlU0K9HdEjj+jKPwwzUfPhgZD/e/yKSB
8XvyiY/Qc9x9AdhLm+SYeYHQvEsXfIJCoZDj3A9w6dRAL/HkDEq1Tu09TkqOMBmTEitQ4CDJG/Sd
uStMtadfYZJ3vAGxYEX/ShivB002tv1wWxtVSARF0GyrPJ9C4Tqa0Jz5uEa/wJGWMjxD2KEjoPf9
fQOPoD64CL0avX39F3alB8F7+0Z9sd7t2D46FIqnGCfdwl2egKCOwTQP1msj6cEa10tPPxrVMQgZ
OP5G/ZpzMAJnOkWghhPkKqAUv1+2k+cVefRG2eSD4C5d1/ObDgiyVorV+8J7/uU0GzTwp+62s72m
8XGt/CZB8wKP0W3sMoe9ViQTUL0RdFNlE5W+07DftiaBvxFm40W2QAf2TTBxsjLbPbbBI5wVkpjE
BiMeEWOwBIndykPhlsIcopIRMNu+6KCeAmxstr7ja09JXdEn1jL5C7Afdax2PQvuR3DdoC6vnCV2
ZDUqfso/kV2JvaINeFvCDYhwSnLtFLrsLN2FFr5k3oo4pee8HPfQI+WtkJkxVYMxgb5JrYHD5Mds
+vgMk6mgSlvel8Hd/gLBTFDIAgUdw4+RXHtYoanpJcKO9qxu+nQ/VxpHCMyMNEXOPimod3Atj8gL
fODUfFwj6RI/gc2fftUfWFCzGlpPmOSEgwgLWmHzylUagyyweWm11+yhwncNIB9pg87xGoU4zg9I
nrIy7TADryZqxv96R9taAa/lieRD8Qm/sr06JcYDKbkcbELaF9GGhVcyZhtxKEuybONqU2feCrV0
Q1NdgAJdUKxJHSEaEAgtVpPi8cKGjSmWMgKotOoC8JSRnOksekZfIKUMRjAi8m070if0PnEWt/gY
djay7QrD52sScwNO0sfz584y54CJlxQWbWFiTwWL+M31vhC4VQsBbU5lxDsjb6utyW2faEQIUS7e
leUbl4M3DxuapNPU800agxnhAz1DcG/coPt/iWw8Q/jwIpqSy46pAz8c32674MLKBLDzkqLJnUYa
z0xR8EbQTQVabt4dKr0YjWrt6EACE/NuuAOWEoo7sFPHinegzjC9xCvjnYnwMPYm0cDxHThkhzFg
8+P/EN/lwj26rDx/OO8VSXCnMH7KIDrbJxCms6NuGoIKjWxUU0h1vdI9NKznhoZXNzEUBEUA7Iqo
P35GN45bto7DiGs4DCX+3udvFyvlZvLoGGYx+7qgP54ckStIMP/Ev1lSuov4mWndOTLcaJgAhKN6
zqjf9b3SUrnug8lCj/teeSFutcqvRTM/aevtKBDdwEKDjZzZCW0Y6YhiqROKk4hqBaWMEDcumg/B
eVp22DVa3pyMTO5j9kYtwK3tjEjz14cRJD0w7bFJz4tSL6QPrDEP8ME3RsYhG+Ght1wNcrZjec+l
J8a2Vs+rYuD6SgWtxtzlYrGvRg8sRcZmnUQolxBGdCNImUH8zwUn8GROQ4afCrv1UFkJ+PNIvfbf
ZP8EfYF7KpR+nKNawC7BBuEm2UDYOJPjVpTO/TDYLtswbx5Mv30h01qhbBmTn2jSAgRHIvdz9KBg
CcexhI1dbWdpZSMVyrn2H49TMiJvzGzzImV2rS6kJQpIVM3xeVPij3q6lshMWNgA7gJ38bUgLzaE
GmYTsO8orUbD3U0hGXWpeIsQpHe1NRY1MkWnYYtAVmy9CtCoPl/K85tHY/0kqVZZk6ZWd5oJG5oj
l2fMT9XRJ/7gXQvYtYdc5SQ9dkwcMg/P4A4A+7jKWWkdmSSiPqRooTBBUMFwwoLPZFIhBWrMYgm9
Y2XX7CzSkbf6shIFpUlQiI83tY4qhll0oesSrmYiJab5Hsr07g0HKuDvTRs/JHt9B7lTgMVxj6v0
MLjEi6T7pNXbETQ/SRFECno1WW81BXSZMhiQDD54Mkyt4GqHHIsHGQy3wMokY2TM0+YWkVl07Kcm
JpfIpveWjNjgDhXrTA7RNA6dac82t0oG6alBWTA83ykB/ufbDjnpMJ+scsW97dfbqIKTwTIMhS5S
+n1nYo+vlxb56j5RwrYmJCJc5Jvf0yAS7jtxz2OcPpLhj6hDAhJkc3SiMJnQDLoug+34oH8Lb12C
h0TES/do3axRpFm7KDJD2I+/4yw+xb6/P5RqXbirDbLWS8mjN0Y9EUcbxkkMHu5sjgjMhnVMFVgx
tC6p/rN5IGSH8p9t6GqgCmnGTu+58GcjiHSQGpAB57mKoknCc/Iv9Ev4pfakeSRiwq6vPQ9rvkz4
bDg/8J4V6Xcj+2xkSPpOYiAvp//tVcKUx674I6/KP4OCqQQKVc5SsIkZsvM9nPARVG2HevHevRiY
Gd2k8AiCENdH1zzkwmEE509C3Ec6CGVaBOJtwDJFnhWVcVxZ1ZWPegTFiHRSfJBJOIoEqO7CQo06
Gf39wpTds+LMgX4HUeGYNxiox1mDILWsDuhpriD9c0DRydn1YJzvrldrSB4ORC6Z0bKkacj1HIpT
08YTROeu2tjCT/OflCn3G//jqbw5BWfyXOCG9cv/ogDy2ER+BZyPpYfBlGPr2n9WTM5lQ49HbDbI
g4Tjg7DBN+U/ABiSBw5TYekuL/whdDZXZUgBNVSd/KpEPLPFFKCB3TzJOXc1BDY9Y5oJeHbWlQ7p
Lv5nvnL68qqlL2yrwoETRlBhodjKdvIEmAkOm0UVfTcxY9IqALVyZ4kPAlSOXuymCOeccm9oHE4p
hVXYwe0lq06MNn8yluGcmfGyuuNxBk1yhqYkaz/SYBQyfP/5IePrinwjDnyBC3UJBMnpu6XY3lwM
AvDThV0Np/bUEw8s9Qf2kvvt9z3RqdBcRNQ67rQoGqsk7aP2U5Nh6zobHCK/SgTiNYCZtQL8znNb
iraLrT8JKVjPt7cFn/XPOWgdOSyYcXmnHnHxIk4pj716Spg1zPIPpgwqjP0qPxZnGgx7FCDAAmw5
1oXObgxgHizPdEcm1l71xdC3Q/tsDf8U03HQ116OlzxEGqTviHJi/qtIHYAHG8I/d+Q5My6IAQTe
sdGwfMFs8+Sx+8EtEJxDlA3gxqSfoci3EqBSJRWf7+bpHqvcKi/ecwmhMeJdOjSvXYkNffsjSNi0
gr310Y1SvNNcHiki9c8EoOdvBADCQoqijwOfz7GnKCA0H/H4vO+9CI6piqiBYA5b+snCA7r9fGE6
6JhWzPRDzPiM1e/KvgWbyhXMSdeFXV07MHtMVghhkTCEteXDd53jYgZlZJlorf2fE1bJ8xQcpLrQ
Fdn6Cwx/RI6lR8hHwEN2h1sDGVJYsTfsNVpJ2Hij3Hk5Yt+d4OPa1SWV5xhbElhDyeDUQdM0RFwm
BkfyIm15JzMzL5sqA/9FJDkBFNKCTOxn22wfpy4Of5wvzqgplXnqxuWWJlN3Jf6EAsParC+ebO++
JWDim9vFEGd0wDZYdLxT9ja7se5ns3xPgc8IngF/1m6PFvLZtARz6f4uR0IsY60vJ9ehkdt1Ybgq
5Y21+GYwe/zWtwfUx6AO9vV3M+mwhPxkWi/MfNmANzj0/mFxrhgFob5J8BK4nCucZ8ofwMwUFoqd
KKkKw//YZA/tcuWh/AmtiPkEPL2k4l52K2Nt1Az17WsE3hVqPX9kljZ38cFgQY+CnEqFHsQK8+hU
EKdVs0wTlkUDigxT7arbNbEQyGUSWLetC6Q9NML74vzIOJgmkKla3eTMgKjIBfHKxNLBrhGRQEuT
4R+LUe/cdtTDSvkJyNKPsLNnxSXFdcjPG1KB88J4GsuufWK6nvrWRPue2+NBT4LzeGZq1rD9Hoh6
8OG6aKKsYRmnI5/7fGG3fnnnGP/CZiz35ch0mETjRTysVmH+W6WOWCVdRncME8/Ia0yEZ1Mv015+
GGByz9VlK5EJ4clbXFAzk6EDkLpOOsm93TKrMI8CKx4RZyY5FGax2+Y46upDWQyEqjSsYLLxnftb
bxWTSxIgPUTR/grGmVdDZt+6GIj8z59hXpkQ4PUvcgEaaTtI9wNGqcZ+vTdFrkFcdP/eK6hv1M59
2xEGVv3JMi10gyMr/2kSNvXhSbzTnKi3WV65ZVdjZhXAHmVStElYWFCW2ZCmnu3f7betFen5lOym
fSR5MtUQXaRTBG7rWA822ChpeDsHQs8UfrahjAATxO63WwHnYppRHPERreeGrhGNfSSzbGAsxp5m
4Zo0CjtWF1yHINUavDmtnAHZVDimJHtWw12lyxiiTGP6FD84JB/fs2LXkqwnnRcDkG83GBIMwmdC
SV5h1kwc3xaVFNdwzlpnFk296gOLnMpscMz15H9wMg2egHdhy0eXiapemlfENmN4Vj03zaUaAsYr
O0xcSm5CgYu91IoYiBBrbTfccPUBJ0mfsXd6mFysIcUqk4Y9ItS6QSeDhbLewxNG+Fl/HqGMCzA+
Sdeqo7pkALgajBRb3cqq3BtV29uB4K4ev9k3dV8fov5WLluYJXW0xXdA+QzcP7J1Up/nybvJ4lB9
Zue3Ugoqkj4qPEwPLSNvS9fJphlMOUVXT33VHXaT+/dQTMyiCMEc2yD2BF/bI1jMXgWusv2r9reV
h7AQDzilrHvZwO6hsS+8azWCroBJIT77IIQNVrw026kerinbF3PCLsYOZrBDmWbT6AKrrJINi1r4
jygAFm6yDSVnDyGccTcs3akAXjThiW8cbAyJCD5SBNV5HkQoF2RS71tX48voJWZgnFoWxAmp0619
6NBLeaMZQeA2jYaJkQx7enmoX13eU6WiV1LnUOXlal9GsHoa1sTxHuDriNrj/OR55Kr3p7RWJQKy
/MGIcJvxYz3vOS5XfV8oqa2th2gjcg3iQ2iOh30IZHOpaAJnXracZNhYw2ebnybDYbYcPRMEsAZ1
8jaQC2tOUkJC7kqECSibABXTLrsNsstoFuTmhgqVygC2L/EamP2wvfta4Lk1jy103Ut3FGvKv7d+
CIF57cprRAFl0gC6yFygm5nl8V4xAT/hedwSK69vQOsk4GWnIv7h9zKdnV1rB2dgxe2IyT80biHA
5J7mVLrZ6DI8w3MAKiIUe/eyEYmbCU+tKJ8CQig+ddIOtvb/V9b462j96/tGsPO6s6qcNKiJdfdv
FEaHY6tsw2PAAZnrtISQr1YiVRuob/qgUR+nC5AmloUlXLrcko7OMrpTdTFyxtS931D926SbpESq
GIU3Wvl7ujVBfX3vcVSwnCF1vb/8dEqq/+q3W7+muO8l5k28JLzEaj5f/MzA45247OrJuxxeo79/
QtE26N5HBGWxZvVU1JBbhr5iWwM029mm59Z/GdnjYKE3hl7uC/zClFqPcJv6FLOkcJtkjqq8CyBv
y9ocUAnBdb6o4IHfvktp4W296TZ5D91xbnVbPQzde0E0LTnJ6qmdGkrMjfTpNPaCnvrAIWRRE+gt
aZlokkvuDkh6CjdZG77vqIxfH+ut2LkIx6ZPA877YjMEfNe0h3jmYZlGWVq4li71xZwCeGWdG4LG
iqA71QTmUVmpcOHY89NUpBriCdycKDxqDA3cimx6nuF2RUDjOb8I8V1lx0Rl4loF7My+pAsd33Yy
NFgTniO3YDmcX1zBRjvgcFVE4GAKod0hvQFESj+XNd16+M8QKqPNz9ua30m2No40eJa5/q5PJGBk
4Hef0bwf6vV9fUEvsABssNmqx9U5MYq1cUSwNuJpgtiFOKp1aW1iUEDx4S8YaOJElyUX3NAHHsix
U+c7nDfoirQ+ZnyxpP0f+B5atgizFwB9thw00VZrpVqzUBgciXztHW9NVOx8jtA466ElYs5H/qKN
m9InYZZC2lxdcaEieDcX64V2k/blkdUcY4hw1ABdtxiwYZNuxCDf5zJw+0RCdVZCzSO0Xt9aqlg3
BNFpaz1IvCVzIIKNt4eiRadHzgrNU1ZgC1RWtDGmtyCV+XqDN/XQLLZ9t7NScKK64eSnkw0qhO0H
6+N5/MMrhO98V/ms0EEB74R9Nso1d8JKlVSgHcQLN2r56M6fl61yvNSMhHbjgy/IUXdQ1CdaMLcO
CVglRbg0u6aaA2A9GUyJc4i2EAawI3DuwaThD90KT8MTntFm7TakINAUocj2LkZLvn6HQOfmR3AZ
lmvfAMHh9NR4KiHWZ8rjp1NagyFDmIbzVxdKIp8hTqmdLYHRcFC+w3SPCdTp4FQryI1wnNvl+f1s
objG9JEVicG59jKpE+hXSv4X9T6HE1gA3kHVQmmLXOot/SwZudi1N/QWXiZtMRjK1LuircF63CHg
uNMu7tnTlB3BIZ+kN+pvqN8KkHcm73UP6vVd9BdSPC1hsL92KQX8UBKVZargiWjrHi4koDJc4Z5n
sU59KBsIDtFp/nkWzZMExyp78w3TxEd+FmhmwazCgOY3K4oRLxOKdzyvBR3BD0UdcKWPZekHJs1t
tj/H/dQLdwpz9qJnXNFQKWzfu68asC9bAQxZU3tjIqA7cUsQfgQX7uamEH3n/d/U1gk+GnN6vYHj
NFn4FiV4xIxe8wonWryO0pz4j6DpkTsN5BVq6Wo0ymLLfNkN1QoY0gGOrBbB/zlMfJpqZIVFW2Fy
c1lATAL/GVP1VeBr5Ed9Dn5Vi2sF4373QXBCACGVdk6QBRG6emsxD69eKKIsiA1pg9Ay6vb6hxBq
TPv6Q/pdlOGgjok24RZRZjCJ7jQiIKi38/32x6tuBw7xswQeqX3Fk52vRuV8KsF7p4g9SifTuXcz
31MZdiChGfiq/9/EwqISSKP3K/rl1hP0xEOygF+59jO+h4tmGKSwRnvdhN7Qr37qyc0KqC9QNCZI
nFH7JzRTzsqZ+dyPhA6wbDjeDjJpERg7eBb8QwgTkRd90DJ6Iy+u3FOUSnKd0BUAQn86wNJyGBO7
vCPLjtn4jauraGSPSkOMpY/Z6SemP1uDZ5CJeoWPo43IVYpmogQqwMiW2KXjewEvh7v3jPnyB2Nw
4uTFjiJZcIT7cloM9AZKCXDkBG4N/UdXZljsA7UPDHBsBc7D8Flq/A69v9cAW1f5upOu61TIw99k
x09vcbglBe0EtUF7zl+Gsgnba32qK1sW08/OnP681DNZam4bbuhmhnn+OiBrFTuAi6G26dCRGjnW
cQQ3YOd7xjJCkIwGuPO2cgnK+ucNKDgsVgkHa5ZYXu18kxffyq08KnSKzhyYUlN+YYjThONGn3RL
kXbhRppdCccGVccg4f+gDMRpEhXDoAMC+ZfwGuyMRBMuIL2fg7hZjahALVPyi3AIZvseCKfP51Tl
J7/NyelU6CJuJOf38Urk9efjLTGDux8TfcmX0sXdaKi15Ec522rJLtWZif8Qb5Z3LvIiRYdwW+ZX
oHXAfUBKmjcXijuI9mgt4v1a8TwtORBdWnk/JjhWZWXIAydWihIj6jngBm9iE6yYxWA3UohWs51j
9xWh0TizutF3m3qEE0GjvMFcUbhQAOfphwcoSNW5kqWB4Cwlw0lfnaK+sKyi6Jd5wS8btWTdoCIi
wPPG6T35Ijt4MV3QcPV8zVKckDXQjKHmP7iaIAM4SOfQhC/TRaU5403hNHhFZeJ0MqqNEMz/L/Vu
Z9tKclT+MHepf6R/99u2HRsigBX93fekMBAyvlZUT76O3C1wcVtjnPWw/Sz6eBXzMZc6CiMw8T8x
AwnFp9zmjc/zysc1h0LnztH50QmzXvBZXVPm+pOyHhXSzU4G6wB2OUTCr/mXLTxSP5xeSrzwODiW
a9vydPyDqZf+1dQP3BlHcW+IiMssRGdhAxUMiW3pGR6a+OuJVJXgYf2Zq1U9axzCncpDGYPVbD0x
0KiliGQnH88K1T5I1FlatuL7P/yOXvPw82R7xpMeMeizgTbqxmmcs+vZU2fS3jOxEtAKHAqtMGah
XBDQSxqflig7A/KEPFBZATU9z+viL5xH0pbi7AIx+Bg8Zd3kMR9TQhavtjPaGM+eQklDEhivVeSN
WNoDdrVnCn8yEfAr1u+YLEC7RhyLbNTKbYdGwGrwIhCvw7KXtAtF2idU3G5sfPcj9jf2egvvLol0
I9g6So6dt3uEL0Emct3cnBxDiNCml4D/MjZKM6at8LgSZ1vBTF5RhOE0KZbYqyVA2aYKnCkLb/1u
c3xchbkUUsRSjMIR4/ekCoyiYh9OFLB19tIxRgNc3L3WEWdih7wlrtLlEimOlZDqdqkewe8fL2C2
Jo9BUTMNjpb0S90J/YADSHNSGG3ea8LAQWX3dw6OvXTU0vwHQn6J7i88KZL6Fjo0j6j2CzfL+tXB
8VHzJmfENzJxFTFJrxs30v/+cxleJGYsHWHS/XsnEc/73q/Q6l+hYJjowYY3cXtur5fKmmGw/IzZ
k/T+ZCeA+fj7Cs5O2ELREPgpf3AQErZUgqMGd56lnM16ue0WGFNQJXQBIeGUGGUlS0POkgKPyUJA
a+dWkI6hrnptM851TD88vIG3qKpR7ZtjiKgtgSL/gHsvM5jzaaCX0PTswYdFbKD1u7Rcu1AFXjTd
tPrGdG7mzFpgNFBLaKqKrWuLYQj/GPG36ZzM+jrkc00iD0LQrbfi+c4PlOeX5e3+OC+fD2qnXxwi
ugaaxs1vplwo6w+MxSuK0UCie1MTWrNlYhstgmqgOn1YoX7AbuG6jGfz2ne04iwr1RqTMG37EgFm
VY2rY4WY1ROkuS6LDFvdSgX5QvdypNTHjDxnh3UPj2PzgeRvUk+mBEISVnwnJ7wla3t4w5DKUEhp
uDyW+SPEjZqpnEIYSPVY3UPm5hMhhrFWMT8HtvfHq2ruJsyGSxSLItiQFayOkbs/w4S/LQf+8f6y
EH4yAe4mSlP6zq8BkFBIlGVH1LgsyJAeYspXThkThJJVWbhggjGfmCfmGqedzVDoDFhRNOT2Usui
OP3O6HE8U0nj/x9xeKABAfsrnz0nlfPk9qT6RMoadRU27yaNQ0WnLUkAbb25PKVHDLUdRW13shjH
rxTQbMCkVffSRlYn+S5PV+zxkEutPVPB50Lj6vwAvzEb9UKqgfREkKjMLhS+S4RhhyfJqmEEH5HT
XYEUqrkGUMA3SRP1/nosYGYldQ6BEStBuc+tywoE1big+zIQpzLmbGZ6ZQ4FkdQWDuZrOh9wnk7Y
R2cX4hy/HSeRGyduQydCnP0uLbxRm+Of46G/xoLOainaNLz+iNVMcJhp2ZFsy/aObUqBNXPWDcJY
lG2/1MYwwIaz7c0MO3C7YYD4Z/xJmJyPE6O7p9R5KOaLD6uXsOssr3m7fvXgAosAAi81s027sWC8
Ky3VKeWhoM0hg0JOftLSL1obHMtjLGn2FpGN9LfAWwqT7liix7+MW/j1+FiSIHALOFRxxOHYooPp
M8YkCW2ld893+rGl65i26x6HSoPcswimkCrONw4ieL4QAPR1i+LHXT0wowAlawUMFDT7/rJJiHWp
iLvDdVGYXRMkdsDtmG5VVCfMhH8LYiRvacaHBdo0pl24pVE6CF193WeEBL+ws/Bg54gbpKp4eyGN
m6BWlT2165ilkABvGf1vq2/ipJMSEcEMGP3lbOIv1UChN3TuFzRHrG6bV0NDwYJItWNagikGWKw0
0Y7t44YP3/xMGBzHO8lTVTF6Mh2p7imeApPN+d7a4i+0Q3NV6tyWHHHkZspY9uqGlEk3XIlTAKYk
RyWRRKNMHAH/QB2ZNw9F8iUnLRMeXa6ZRz2RxzY90LZKqm9fFvKVnvRoBvll30m4fz6EXzP2u/XR
3dO/2+XgDTLZN/uqF/DcA1dEFMX84BQCsbQoRjOBx/dhW6kj/tLwUpMnUoA5KXwKp16Pa+La7JIM
0m5MDzrXsg6KESU9ThtVFHJtS8uQyFdOOA0NbW+Jk9Zlt2xxdq4OPQcce76EO8kq2yi0Z8kpLsGe
ZwOLfXlqyGP2zpJrRihNUdsoBjIpntygFa4ZouqS2hhsYPi4O3b5c3RswEfXeoZpUdaY9NrJvV1U
VIz3eoRAfhfMn3PDNPfw4HEJH3gF4iQdaOjsioElJhS+mFVPk1SN7cSo1WNnoLb7Cxw/U1Q+CN8A
nF74llqpQ7FZcltRvc9XuZ3r34wXdUHhnf5BvualrOMvkGMNJs5jgc8Nl7guHbRGuCB7ktxDS2JE
4ISP9h4TXtfXhtX+urCvMdnv0DmOHF7qvIJr7Lyt69qMRTg0c7MRxbzC7/ojQnRDSedMadL53Slf
G+qNkPfkx2vDy3lI62JddbhC1kCnEv9yP6eUqJ5OXKY7JVpY4AMcFOLFicjkWnYM3w2onXUQhXjP
R6t7KclUZstfWgCYdNp44FD+DiJraCndVgLKui4tMf0Pi8CekiM4crkVAH24p7TPGfhx2+aonHW7
qHFw/POPLCXHEw6UhpPCTEPV52X0Vl82gwcpNxLQX5Cg0LXlQ3L6SLiAzFLfBt/ERHRJOWBwXmCm
FYqa2s4jhs8dHawYZqTMacZpLG9Gqk6lu+RZriCnhqCfHdUZqbb9FQFctg0DbfrN7Q781UDHuSQS
hntkuyx1MmLOl9R3TeMvu4nE54Vt9QcslsxVy6NGKIKV+VN/yd7d42ONCUt/Zh0+PygA32EbnHDz
2YyW64SawVMU1ADCQ6fMAHVoMsNE9bM6YGhdih09R9OziAS8TLH1J0HK0uU90+CftbYM92y8lLIL
yt/7MOLarBIOG7QR+rzjogygaiv9PiomNwuQCLCrdSbMB70GNG57BCIGywsa37EC10MQuWsA+mUo
/Ea2KFN6/KV5GafL/+xbHZyyXdbdt44SeCpoanWWWw1SL6TkAUNBJL3gQJD+qo6B0ztSXiH9mCHV
HqyY0l5msRpU32oLqDvktUD8SNSJgpVA80WSSsqpdRDC3OfUigx01KKEwsILpGDnUj8KuwxEzS88
Pa0yaUuQ4yqHLgYVEApYI0yFiD7xBFm0cwCgSkPIJcLRDU0FgMsTOPsL0zk2eUHpZUgqzjyl+KE6
0q2wYPIqwEgyebU+r2MBAxkHi5eeWWtSRxttkSGICb+m0v336QHtVHxmf9CzTfpm0pjIt+IUIujv
zBKOPUC2oHzJXHsIe3I0cXvNfOiaRpLTsdheUNj379Cpt/VImIdTKh6lCAmsI/uVLc+Zzlor+Yon
iSjml6SU9QkDb5J6S/U/znR3POUSAuVVXFeY5tqkBEvUdVZPL8KBofATxRTqgJthIbyD6Oq+cceE
Zqfvxv1HkOFHqSf0cn/JJAp13gx3OEIBZgaw6HSNjQuNH7X2FL7UFqhGDRc1YibtKAQoF2rSrRzL
nNwvxxoDXIThQ+wOgbI5GnETHq80ckUQgWOG9MhPi9TMxXQDzRlh3vq7J0MhFS1t6FWc6zce6fTI
0WBP+7wlyemCqOVKUnvNtsDENbd+f4DvEfqV2O1Y0r8kmILUxZh1JHUr+KYhnsn6bAaizaU/g+yC
8IV2Hmx3K/VZ8z/fuiFxV6gB+eh2++q5ie8M0slt5QYMDO2ZiaRP1sKcbV9zLL1O94RBSYhkfJeR
x7eO/K4y+4eiWdWOGL0SN8qpXBhf/4gFZzF334gB3gr4yC/bUbQJVyNBeQ7wTxwzSo1nJnzAg1Wt
7Ta3Q8Uqr2i8QZQFOndGV5ZFtsga7pFkW8cTvHKEarXkJ0gfYByIWJ4p/ZmTYGMW5C/waY4X+XSR
od4OflDBegb0oN59g3p18bH1fan1xQjcWo2k9CBNEAQW2qEAc3PvYmJhV2/oIFtMJYSeJoX/gyO4
fzGNwGU2asQjVCTWRmi9p7HHK/wbRMFZGVNd1clE1sXgk6LwQ8u1/8Yt84r7RDW1Rhps6MTec3Ak
9a2t0V2jE8iKkJUCwbzzQUbpwWDSSJfscxsbRAqlVTG7m49gPIvslTMauNW3Gd8VGZQyEzFKc8OC
D2zcLOtcsBhoXWNGsLhH3zUkaDkYG5rVQZvAghCwuQUmjFcaGOBJi5DEBUolEEMeMhifsQfzVayU
9Sq0q6EH7hkMWDIIL7cIPSoAprlxbdKzAWfMXn3wDplgAxhip2HOgDl32QCki7A1Kk538YHpViJk
Ssl03EE+Q4OibxoBrzOn3ZZlGhZ3t5xMwtCuHP+03iXvYqBae9ffm5/vNxU8eSNFBbmjR/292BG6
j8ongF5egna2I+C7KAbKqE8QOWPoFwjOaKPwOLSmlS5smJLIIBx1m+KQPGhRepgaD2Vif6Fm1GMK
QdglcZLm/FUzijdoba4VDkwoWjBimOblJ05+BGHd5Om6DVDSKQeWdD+VvtHa3kr6z1cjerOsQ5rt
hCloGLxJKKpYUQP9d/vsQLxnqioi7Rp2HTOlibGu3p1SanjxKJDfkV8dyyh0kAEsnXswhvxRWvr+
AQSWHeKBqMjDgkupOR/RWvf0KyfBA1oGYMQkYVyJO/YntseLEGaoBSwRxi+AiHem/ilMMdnQ8L1Y
TTT5ycVq8A5jcO1arlvKKoh2gdjoDS6+XOAywHnj2+oh9hkzArEzX+ZqTTeRgswwV1V/40ZRB5Qk
zj/6R4zi5pLBzrV5d4hGOvrkaVPugwMTYHkuur0BooijRi1l/5ZHVQKZfXu6RlV8H4jIXyp4iJ1p
SYE3HmW7viViiJX5Z8xdH+hv7ZJ3ZxIcSr5tntEy3aL5AYbwEPE4GhJGA4MbykoQYgbpMEDIbSrS
05xSV8z3DmoYrelAua2cD1PL4nzAJoyutxzFlxNnEaO4clcx8SNUfORTQwl9zoZ9ZfP4C4ixeOox
OrW9QoXcSR4Az1dM2HvN0by8JZjoGcuK3XcTWfwVgaCS6MFL7Ri+fXrj/Q9IQXWd8pMXRawtWZWQ
7ErSzkOAzqjzKMTlp0owX8AG0qmu0az2iHymKJTIEKQmeMut21pQHINpfW3Ih4osnDEAXjm0WreB
jkeLgF1r9oX0uYDhTqFrZrYwJ+MNAWp38DsgWIqVAYZDwpkADzg7dOeQZgY0C3mbmgz0UL30tmXr
RDo9kSQ2PQ4KX/F/7Iahxs6Zg1RGQgDQmB3OZlMPV3GFBPzemP5zWVieANb0mZFQCJo+hp9+XXow
0Os6qZkhgTH0FeN2l9D6DsJf820f2A0jkWhiNBH0sugNVINWgseJiydogjO2AHk44oI2hLd0rZN1
TvUuUejY4X2TihdQPkKbeF/Vjpe7qxrlv0XJA3eQ/VkyDKQNzDQUDDjDKcmQnBzh7zrLjUEBVy/R
hV8wQ3DDGYkOeV0hYaJWQcqVKei7rfHXHSxsJafAqm9oTD4lCZb5qhh+QE46tYTHt+GzPa7ldIrC
4lUzNKXlnrhUQ6YQHdveQt23Kk+j7h3NiYsGbtrPG7Pp0tX2zYhY6fS5WpaWMpIN08cdKS7uqVB3
bIWhMt2jwqdduTYAspGXZo70nUt1hpYrQYgfdcVrprrZUz616DAnR10S0YjX6eq8wRoVCeJLNLv7
0E9XK02R+rl4kYNCM+OAGC6UtPXIIWsErmryryoFK+UInjJGwz64B2X2Af9vCq8Hx+YJZeZvpJJg
BQxbuvKUzNQZnnuxwerYNKdRNuzs5qRqgb8ntta/lUo8OegeWR9ch3wfVzW3NgzVDzthQCfr2EUE
XNzUGLk7gE/pm8SziORSJGd/Ic9TyOUw7B3sdJRjkQ8hfqJtK9Jn8Nim6nFUmXqVd/y2ENGMIqRn
MQQO+kJJ1n86KwWu4vS8z27nSrjGGF6p+A/y69YUl69Pp08T4kOfpMPZdtIvYaObu96j0meTvz1D
d07XIc/HDrMCRyoxPzVxz8NUG844oUr7btLF2l31X3N2p5t/5VVvuUZgCi0vo6CgxXqVbLviOL9x
eyIOiG8CZpMPP0dDJL5ztUiiMLXyG5NBZeXBEUuoEEB4hkKWzxAuHB6vcLodXsRQiLwJqO3O23cc
0rIyDEKG3wNhwb6DsFZMbpDyA2ltyhxNiIFAWBlvlN/6hrwfIZBzLzoygv1HDMt8xsrEYUCfNsRe
ybUr2mLgfhqak+kJTQUO2/38ykNlOqdSuQH624lAzycW++5SCNXe8AhQFazYx0aXQct6ck3NFNHf
L/dQoy68LecbOuicold4DpePmMYCHwanfCUB8cP9q50HfOC35QDyiyuOMiMK6pIx0FVGTB4ba6Jz
9i2IBt1hPxJCatnc8ByOxBMXghbvyYXBImML9UktISY+eAxeKdsXxQiFYWtOeacak993+ZkNiESR
UEnGldrRJCG0hV54wg24GEHSgPMlWbFFTHvvAC/Dr/fQJhl7VfIVkoxL538XV1RBJs/nUCZN69v8
cQll3Cc62Z84P0cV8KKKvk07Dtui4nVlqlfN8vgRKpaZJHkwzYN89n8ZO3t8zodnRTkqHCVqhakk
xzfcPgI3fot8Zw6Wu32+6VUDFFswYy3Xm7CNN3HopZSbeG/Ideql/T2dpdmBxtdE24cyhLuWBKVF
FlgNTTv8tb4o549JnlJXZjlVF7PJAAdSOK5fk1w8CkHVoJ9UeNFNKO1v1duJAYZtWfmqsSyDeAXD
nnoML+S0TlN2LPFG5qnnPxTgLaBqiuypPFIe9YWbskSPnAZJw3LwI2JZNfNUpZR8lqcuc7mA8y6/
PLLxPvSBQeG8BOXu6b0YVaaIP4x+3XlQyDx3418pyot9j15Gysw65ACWibtGN9VGl8+/u7d4ysIx
2YxZvG57flbh0LIZ4rW27mfl3jI9IbaKC3Uwfp/AyHCpeHZHJzi+a5m32kR4gZ/RoMgtaumaPyxd
4IN4hYJetf/0xPckLroTCeHLQCLecKcUZxhmpSZAjdRe0oskYjELUlzS6mX4qzC0dqPNEg2K/k9T
7ZxkEI5wMM3xnHnu3bXkoMzgsM/ynTAhSnP09n1NJuE7xRHqtyLvoYOUKvH7t+Gk/KlzyxhLbntJ
LyLGwwMs4XFW9RGlEy4Ki0Wo0VQghFJN14Xl+7/sOLmgLfNTHeCv+0z/1KaEFFwSt7InSdXAM1UJ
DcsBXlEAV6Yqhm77ff2mf24dSBKzkztgo+YEafNbw0N5B2FrdBh6y6fkMGXOkXOf5B92f5OIQKKy
0LhB2dEl2tKVNvbKRivl7y7kg6a3fXSZnaORKtn9NX4Sd7x1AiSDJy4ZuKHSfi6C0wp5F17PYaSg
Rpevt2Ebg7W+PSNXY5zpvF6x+QiSudAzzxcUz06p/rACQTugWbv3Zj0RIxklWBaz7z1KMcWa+AV9
YdqLyYkdqIUt8pbL+Ltv+s1BoFFquY+xV29f8ZH19hkt2UJkBNz41LOFjcAX2xppBMeu6Z/IxyFG
MfE5HPl0QGwh/8/uggHsSrPRTLi+20RsxlBxkUacGjM6Lv52dW79AdhXCUSq0OVJdNu/NSmO0VKR
KI5OYej0vE0MTF2s85btkgepq5kQ5OYMLkHVw4rQ1xlNmKVYzWsVHDq1Argcy7aril8cIzmEFIyY
0VgpnywXMMrF7vvP4pNFyfq59a/11sXNFAkuuPeN/G6M53B3Gw9alQ+hEyqBezH4iOEilHwOW3zU
O5DXUmUPhzaFuf4Y4ePG1IobkNfA4RO/ZoqhwHPAGg+2dnIQtuQ7KuYBZcTxsv5inUH/a4Zv92uw
apKJKY3PRA8uZjSVx5WfwBzAWQ1ItzorLj6qzUMF0nCtMgdlt0q0NVdYU89ITtne+b5rCeUs45cD
tLzmVwubUvZp2WPm7GAZQDTF7JhmLTf04KplmLF5xMUm3NuJ2Woz2+5aZoBWmOknVHAzo5PWLwzv
v7nfbRBqNmB+iYwTk7o6jgAooQzGww+n/s4WkPnJhv/ne+h41a3/OSeJeg2Ld2zUj2OKxUmkuNZa
I1WKAyxcwkZg0NFBsmvb50HqW7A6rWwVr910ailyM4EduB7b8uwBAGAJwxNHi/6yYICXNpo4f7AY
MbqFMg1KTkgzbh+clLYSz0uDqOqr+esnN2yEtLLBPzSvhh5FZeu8ijQoKy+IemseHGe9YwRjBo3k
AHHNDqD5HrG/SGSoHQeqhu9h8eRCCu8lrjVPnr182liizqxtnlAvAf3c0zPNsmAge+3K0553q23m
c0a08w21wXUQYHP7Jooj95bJ0DySwJeMQzCA8WALUeJCmTuMLHKzaKr6j4Y0Sb3VQlhA8z4vT8WA
gCo38Gp+iqg80Hor9XSibYsJweH34Bt6/VcApFONKrJnt1rsbjLIZn21JKOK5Y9ArNHU8FK56GP7
1osrr/Lf3RlAcMJzPzI+gPy7yKCz5Nmo6QT6H/qZ5i71qfXVjktgPQxxNPzqqNj+X7B8Uqv40kxJ
K8yZiTDtX5hCGtKNdBtU+VdbUXQK7s33/rQ7VFP965gQ89CibVOUaHdhMnK4l7F/5+aU3aHB4oS9
XLGgE3pNxrhxRMq1m1CCqLQdBXT9kbxdFOPkMJ0QnA0TWCvRbrW1sMqwVVjbMuuk8KuOlzpHocfF
9MHpxYPFE8D2VeZRXMQOJZHwFEpIDFjCvhSFora4k+2P0305vuh90Lt/RKsZbSRYBBboQqBmv9ya
yNW624eh6KnkxVN5GtZ9yer+n698MN3pk1BV6bGEp+GmO0A8zZw+T2IKqvlvqLlWdbsERCalnCDM
7yAzVOJ5519IU2Maow/qli0I5bxFzopBSrV5BzE0j6Qcdgsm5qtUB08ECp+HtjL73xAbcMdO65TN
R0WP27dLAeiIek1q3gFxOnsorszot2K31JevO7162Vxg/jR43rI9lJQSUopC+h/lXaHWFILQekMz
dxsXlk+IEfOGNDZXOdu5wHVEFPWjMmW8tgNRSO50hHYpW1sqw8tS2P84q+pEWgXDuH4baxtrc0B/
ISXCoP2tGYK+zZfenH7ARq3KGPJdVYKuKW6jSLph2QnOpT90a/Y9Mxw5MZufyCmDoqkij/1kkcso
CbOXzVNQ8VfQto59g+Ad2JkVbZ2Ayimfu2KjHUW8BF1lxTWj+W5E4NsrLwbLuNBa11+aLRznWSia
uifH5xXsAdx/dtxMHMaNZN1wxh50scjn0UkGe8Pa/T1pAnwHi9Q57POUQfZbo41uZM+TkoVPUIVQ
KwjTKlNMoYLkw2IVG7ourcaJsbqsNYVkkpRgkIjdsVdz1xiT1H3zLLWeSeGFncd0pyJclEB+w7aT
c6op4j2vJ/I7hKIWOxGBTwwX/xMB3VJrKE6G6qN2EtrpB70p7N+l9/ugRhibL5P3iNiCiXWQxXbK
EAjZ/MmouWMZSeboDnCYCbS79YNBu7OQgFRMLSaQZQFneXwqwhMGKxiPrTzWsutrmPbKsOQeNBBe
A8xYHSgsXgUAt+i2VCYXLPHOaMWnxzxc8i+9yImhmhuHMHRsOoGxVKXwVFm+ePkRP3TcTIW7HhQy
YEaox0Xn9VsmMtwpa1b2pLlVS0vj0plIz/YfT2ya6WHKf3yf99ZO3RPpmIqr4ZlMaO3o5PZaBkm6
NEO8AwEpdAxAuFiuKUebeo9mw64LMX5jNVN2SFaWv6fvGNzFgUE0WCmqklWemZA+HwdY+dnukwD4
65+r4DJ87psWg4c901pmmnik49qpxIiMLkk+G48x7NHzMmeT/ZQeHRLiMuZNZcvMiXHeoSpHMVyv
yOOE9uynvrrwXsFusMcCgDU1QFfWz2EhiXmRvU5ovx1izAD3UDKs0CWdMlW2BN949DMiW61MdiAp
GCwdiraD2fwMYSekdrifn3pmE8D9BekRFb6481HNEdTWavZhBSkJtGG5RgIrIZDFH/7zGY8bGrnH
aVEy7JQz9BUjoD0JOU325YwlDZJWsVmXzerB4NKDKcbMSEvWkf/DMqm0Duaa3+mMcyUPcp/LO1iq
+8Io0Tl5tAkhTM4j5wswrpzYTqUFQqS8lUjaGtna+G7EB0lLpXEZhw9lnMm/8iuqLmn63qHeuFh7
cnBuoErdtz1pm2cdbx9KgrdcyoxJ4KAN03/WG9bNrl9jPB0JnSNZvN5tsD+FP6aOhkDDPAK9gcXf
rfASC6Av4WIer1PD+lw4j83mF7mWOiCLEJe7xJCRaCfzx77PhbQBDy+lGF2/lV+U+S4n+TPafAQX
mB09QxXiF1J1PaFAbNXLC7eW40V6elwYaFDq7T4g7R6dRCeCnoPj/OYA2B1iQjdp0rLXo27SSZTV
1/0aMh+FZsdQmOSbO1n/1+k20H93245NvTtu2IC5gPK+AcfRPLTspX3hSBD8dS7YQTfWxJCIx1ah
k1fYTmNhx/uWtiG4yyuN6K0n83GJTazUoEz0RykgSlUUXyesisUAuoawkMR1FCQA5A94YxmJSvM6
UXq7dPZ+gb+w26xuQZ5tc4434cM+uAAbYDqK3zsv5/IdslpBgk8tM/TG8Ccngd01XAeQywUbcI+W
ROuvihr6w6GDonTgsGepLnTsF06LveFo1u10DpkDQMoFqCS1bebQ2zmBjCDSRDDtyPsimUth8a4n
OrimYMwjZMEC2dhUYoHNpfDq/+4kv6JwAZ/H8iTSFiDjeIGZLccXxluHdGZioCzNozF/LbExrAU1
ruNgkPN2ZgoerDqHTn33eS8vsKwewADYEVg8svMlQ4muP/AoQ0AIIRyQ/phGujNdhoXof2jhxTXi
Ik5/VBOIemZ6Aze5O21VaDkyJ3IHokpku81K9UoAdYEduLeUw+1oldEI6x6pD4XyPu43mK21T3q4
2Iz+gm19q59pO6y3V0sempqmRP629ELv3doprSc0j5Ym74e5yMBZe6fu9BJ14ECg9UBZzkdbe2A2
CZROSLA/fb+IChYdJ9fquazJm/hJwl1pK2KkU7+N8N0drhsTnm+BwdZNOmTK6cic7hrwPB0odODJ
I/yWmdjbtjcKbV4I6YxdrleskMryD4AorgmhdyrnVmrxNt0DgGrAugV56WFpYk2YWR7JB89bKOT8
GqtgCMgYLCWgqqqrv+ahfcztcdKmLBs33C4UQHyJbN0c+k/JzcTzy8Dmp7rGMTsoZuPmsPac/30w
2IWwYuPBXTdZKRiH+LUTHM4EW3GC8Z8PEXkYTEmkwCxCQurqS0tbFimfKm8WuOXFQkQEcGYhvLoB
/hOZ+0XTcHktuj6pDLwRPazr8xVNpHgic8+iFMGMr38HdUj5OlfmNvtMjECXoyDBEhhkpYG+0Q4E
Epp5PYBXlG+GgqTM6hCYHTz4qhcqrgfdtFT8UUyevkssCRotGjwK2SRBkDGaNi0e4BFxThXNOMr5
smPf4KlklCAmvWvHP7qQ8L0lzZxmlTKPtI/J/Lg3vdw7ZVDRBt7rO5T41mJ0dDcKH/9gibvJ8OJt
zVrXlyaEj33S7L5251X0ietWNr9rFrPTxJNffFQW5OKd/oR7+95omNOx+Thj+ZoWKkcrU5U+w4mP
mxelSoOS+A5YwLaf6UUbvq3ma2VG6X81PaQSKlD230XDfbmM5Rq8FzP3KvEKKbwFs9nCCY5EnOz+
mfvMcdrUjSQIrGFGU12chY9obtk/0EWqPMMc2Rq4GZQi7xdydCWHK2JidXqLccr6v545YFeFkOvD
zjdHPFLiP53E2tBkIGZZ8qv+pASiPMHiCdRDuKtOcckWIllFMB8doHamK0bG+6AA3k/29mFUiB4N
aJZ6ZYBu0/EonLwOgNEL1SOR/+Hqa9Ia7VEQnw8UyNbJdwDm8D0dSFmugTxWq1zgyxK0AJX72mtR
IDxmBKnXOPHfxMpRg2pMwEuo2Fk3rr88cetR0XzNnZq6pgsJGR5nl//nX5siWgv39ROmTckcg+Mm
Uaj4iXwSqSoxdSNkH7SUk52E2Y4OADsGVu0OHJru7oYCiS3FbckiDTjgXWLR6KmMNYhq44u6Hr7Y
FFpRCPItjifOmnGgs7d9fYLUEJxu99tgd8tpB9aRU3D9ntJsIvWhSfPPmkBbIVfK975RzE6mhaBq
qx7g6434QVYHfXHoWkoIQOXlZcX3N0I6zFo45X0CVL1kG2zzri0iq0PyX6GHe8Xf/ueU96s/PPnQ
UjzNkFvTsptNkacUarU7drutb1ykJs58HV4UIVf26pZxnK55la+DpAI4GouXKxuQNkP+l3rLzjkj
avxMAIjvtP6lxS/MJk0qBaxe/pk9Av8FqkhHuxbKhxN17/7+aftkQ5qQRUJp/RSo21v1cNMbZEnU
rJPJFwHcceZEZj5/S8XBOeGN6UNjojKnfjfLFPIuVzWzs5RtHzpO67kzbzksSqAi1HmRxSJt/FUU
XDIUUNpmKOGzKcwZ0Uc5ytQdUxTS9rSSX0sBuI8L2/eD7GNyZDjzzC2Y0LjlHbHptWPxU5L9S+mk
c5xq2qMQIGlHniqAoUZZa6pOunf0l3aIr5OX5srssjUQfHEC8WySWYRTcH4r7XRNS390JJ9Wsq5n
5GzWuI0w3qdaDgWBEqsW9RUtGIu6DA017ehoxmKWThHEOrmWMDcJqzNaWUNte7uxOfUjPO4hg9w1
7wW76mS3tciL3S+JpK9oiblszRo0I3uhJF0jyIM0Pod6D5z8x5JXbLZzcyfh6AHLtTerY/JX78WJ
gV86f1+qk/HUKcTJxwr1nC07oRs3gVbWvW2VWKv/8iT+qQHu/EJJiLV08ybjHT7U08B51brMroZR
Wg6iSj3tqg2W3b49M/Z7pTqYjJfTXF6J6o8KHqol6QXc0/dKjXbVlSP55zZ6VawoLI4AR/98RTf1
0i01cZh4W+L+T3mpkeJOHWVl/QLDhzwS1Y1DZtzNtJd2q5AUDP/U4O4R/A1nqPnGbsDw0QZv7mx2
bQ5jnrYIG9V6Z1u3sn6drahIg9JJOIjHEzoT9te2T7tn2UqhzFtg0jBvWK9DvHENmARFltUX2ka3
7S87IpqYWdgcFFf4oDfRCeKkfN5+QFu9vjar0USJfWhjXiPbLcbJas7yKdahW554HNAZMCg1jLso
EO1lL2A64qZYcnrGrhwaYcv3A2tJ1dk3AC+/OY1EaR6BlNfb0P+fVVfewXQWPRsxSkxE4SELMeAR
lU2FPdnBiNsDjFBVHmdLJm/3PZCLGzyEgNJkMQpcr2EULUMVfO9OKtwmL0eDhH42G1AaWOgSF/70
AdlvJHzuYQ8wKGbNC/Kfa2BrwmLOR9gIPEHtPWvvSo2GW+SiGnfn6zx1WrZ1mhYde4Wir8ag7RcE
ItejV53JQNoYdKckDQTTtkdSthc1Lk9VWzFN2u6rd1jLGP0c5ofr6UvNNrvRDPYn3WZDBkTiCQRG
wyc7NfVoN1iklI+dyx0QAiEzbCeGeJs6bPwQZBt4X5RJ2sSbc/fcEdSAuboQt9UBd6QToPPhoeqQ
EukA+Chzl7dCLCXv3AXmObc/9iS+LaBuw1EiOBjsu/cABTkarmOeCAIJEx9IodPoc+6Zttqv866/
eVcRlu8a9pqsVcOSD9CzV6tsi87mGmyeZxMdoAB6NsgRGWp/JgAA92aCEvoTlMUZa0Br0QELi98I
4C3a1q4c9FwqkcBnioE1tknp8jjxFqDm+3iK8YFrRSCiuQ1a4aBlnJKs30Ml9kS1aHULc5dCp67C
MLt8UtmBIXYqT9/qKn31NuXyTrH9EVgjz8Kb+0thgRbOU9NhKccJ2jnL0Hf0RxzYyEuEZEqFi0nF
w2tgAQNsnGOQtTS4gSTWsyETuZ8tH42CLyq2vqQ2OTzilrCi8cHW2JRQxm2Ph1hoYP+VTWMHYeO7
n83RIcKzesLr74QR+mtVwRlhCCYxMRW516+wsPEqutJFocqEB2/pR8DAHpJuBowNdlIEpR+mNKZ3
SsmB30j/68W2ut1fTQB+bX3OsjPDt/DErguaGEznMHi4lvqHAxy8crgM47Ueg51H3WkDCa8/Z02f
ZK6ANpffPxPkxPIjOPOPT70B05bVSSAuAOE37SNVRfZhy+vlzkmeD+3cprMChepA+i/AngwzZeKA
mobE1opXlRrMz3G7UtXStqNJrQlIfMohwvmgCiXS4MgM8pMEggMHcifZxXcRAm29kIQmahysrYEN
08LJxgkQYM+1IL78inEtfgTOyjqo6i4TixwimXT4PEZ3aAHFbVj1x5Qy269vnbvnp1HBbWGn7PjO
tQBPXGbHWv3b1tb0glTlUhNtorHY6F9/lMeokvljewcEPV6BGtfoDGEZq1QaDpq9BEnfLdkyQ+c2
BqZ55eoepqtNHotMix4BlAF/X/V51xdt7FowzMWqEXT4n5boUF6oB3a/1tlIqZGjfY941LgFUeZD
UsvuHVI5gsIEgvvsc1h07Yrvgkg8j/ejL+/WB10ed80WWiJAqmKA67FFc8nPVxmIlV71L8eaQHjV
8Db5TQ7PXD2wfM4dty+9Q1wnocFefNwIWFkG8DxjvVHwpMzQ+gpIXaspNvgkRHRXTtSAVxEa8Ifw
odq87ei/HLSD7c11evfXJYQe52g8JZdBpaSGAc39ZFqZ+akGXrTQzOMgj+hYswrY6L878kCLT4zz
hG7XmQuyyKr+juNebr/33Ee8UrqFLeSHWuvALFxjrRL5SdKXWN1tlEOswCrTi80ZMkoUJc8F/8+6
9AK/jVXHVONssyzzcpcY0OkbN/qntrkbaPxNyCcgNRdGQ2LmwmmMFMLe2bzpyc0NZnUVc4yFOTN3
VhQIOC8ahr6sqsIOlCMxpb/4olh/Yu5MLLyfn4nsA6kULnmwuYlTqD39pq+xv2BKMdCvg+jyKNsm
rUzDiWMxYG0XfNGKTj/jDiKlP1SNU4Aphr0Tkr9dgivTLkrpXCp5rIj9NzuY0bfcxr2nds3lz1lR
TwNSOpR2YX6GbV+NsF63S0JPd3VtLmSn6AjJvcImD4ZDs4u0RyRq6X1vauB6+5+M5kWW6vSOYx3J
qxtnjTdHinK/xtXMaCgCB2fuioWGk9PYyzRuspB+uynMrtv9Z4X5Fs3eAjpKS22/jYvHZwwj3fDt
3slB22BnnSXYok48OWStv98fVhR/XP9VJEZVVty2pf+eXcOn5MVEVWp1i5JMQcUMdnqTo1PhD7Q+
DZkPlSsMHTujpaWXOuugFK+HysQFuSNjxZ6M/Lv/H2eNFAQsj8/Mw/1txRXg4+OwjNQzFk3oR0Ca
eDqEn3TNyxcYJAnL9sA95C2p8T6GkITiH3NDVW9e/0vfcUcLhFL/LKJYpO3iEZmsxXSrn+1ItqTJ
dm2x+C61+S9Zyoyljpl/gcf7gLURhnLPFsePnvWDmhNqHkwBQ9181W7/6dIeyz9t7BadMZMTshvA
x5+HOJ7GkYJhGvjiVA+jYrv6i8TNa4H35bOR3xmmWPYchP9dQPe4mjj9Scngezl7UVwkJsK9LiBr
fI/U6D/JsEXAeuiiVzCAnTPIDJHaCDSNi6LlxfAfzdkHvfSiZ1rb9RtPT9QGFzmC4gsLp+PRwtdc
LhZM6zstRNgmNIqyxFtYmQ64rQejKRArG0WhSjhLtIUumsYoDIGrF2bvbA1zbvB/CWi7Qsf3CRck
MxJoCSwWVGW/uvu6ePSSueHAfokhg7HwxBcmiv7Sf1LIUs07zMCuGCF9T11stHHN/61O85LiJ1da
yaR6R0Ak2Lqez5VSW70+g1mvJ6QYcSFk/FABsaiGi35lNT/y+TysjyR2PRRSS9eptTRGRWXH7ArC
aPL9faXyG/EV3738gwaKr1jiM8+i/eGKP97i/5h1M1sfkdttR4OnpqWRmQS8VenCteNYLKcIZz5F
myWeZB6D9k7hCx3Fz071ZKqoKNtlmUMcZnsNicbUgNS+5RwSjwP026pyGOXoLNfeJpUPiptxMIl+
isxxKncKGDJH0uGjJvAvxls5dg7Na6aREqYFsg6NlCwjg2j0t+JHtmLvJ32rbtKFpvezCIc9mnZ9
C3LWyX9ZFZBu+QS/+CBcL19SN7M9ejbmjTCjWQPhPMjjS1HTPQ4WaJjaBkgbsN0FLud/zAoHLjUq
Pj3iyfjDbGQp1JS/rgaWUR5K9gWNDMuo06/H7MjhebEgCY7PXa5sWzfWnrtl5hdG657RRt7hvPAH
59XYVMpmhkjlwn4EPalMjtm1Af+z5wqKCn9xUEMRf+5MbxaVdFb7nFHpSfhNwi9nGZts3a2nJEGi
zzfZgiWV9UdNhvnDEWCZEN2KM8+ALQ2kPGhFyT0vCPOabdt5Q9Lhf6TZ3wJeXVt/8Sv3zWSR40Dh
+WLleTQsLYdHisLbcHi2DJ1pJCWHNkMP8QfNEelnghGdLImzBBnrlYtGSQ8AWEnAy/fS/u/R/1C2
bnvV1+ril7UaIgHe+P1ZGkpfCn5IQmbO/gF4pbPH0k8+EZ5rCeN9WNy5giVTNEVHKuNknHnOCEgk
4b+HaCxrv6EV8fOmsAEV6K1C3jFJyA0gGNKHSscq6pNhDC4C47/ubE3noXHbAIbudZsMMU/+qdIk
8uPm04f/suM8setsm6DATgL0+e8Hao+KwMwvR1ba9j8Lbu5AjtCjDQd88zHi+QU7TwEL2wONPpmd
f59onz/xWQJcTxshbVdaolIuvNRotfWfaMXtpGkC/5K0nu/yJMw01T44m9I9PSy6PHHU2aPUpgxG
oDGB5KSWi+4z1Ina8q7CdwXkEMpsIvF1kPWkBC3OOOK0mH63elegWVO4cA1mhDF+vMpS024g1311
hXvWs4NioSbVd5ejFi+JF1gWoH0aziHzfT3Y2fZJgr8kciLJH3/rdpRK+PMlXcH8gWoq6i7pC4LU
20cwaEjajNUL90jF8iaozdzqehlM2Tvnrbxv2qXzHt0V42LLDyObqs5/knHUlS2LG/EtfS7Ds6tQ
8QChT7j9mnrOLCfxB1Rahu0C0AQOh935aXQt//0MIKqvhCQzmZi2aiWaVGvHPsuwy3XGl00g4Zdj
3vztDx54S0hpxgHGw0G6ItO232cd/Um3dqGvFiPOOqW9eLGTMYFXduwGjFQrPA3sYATIQpdiWp0Q
YUYR1Smd584+AsI7+iYc5ndl+jvVCiH7kgUqfsZ10h29FUPVVgct2P++YKKBCR+U0eTnv+6wiH2d
g40kU4VTX5n587fZk6Fq9gDOaEzzX/sbOs+84YNP93O/8EsPXzbJKozUhfD99L2Oc2I1RDxxA5B7
/qapLa2VhJ8K70XaBZemfJvfKQGqwth2pdOe6vb79fQLvJvPeJv1Ese3x8gv+a4HEu+MXY1nQRWX
o8SKenfVPLJcf3dHfIV2Haqv5qVZheeAnUC2SOw2E3+JGzemcCRvVBenLDRyD47fiYtTu73q3+IL
X8c6K3XWnDYfckW7LFOnM9Es1B6HA4EdSGIchET2XfoCGedHvIYLt1PGiQdRjnYPMLyArT42YP8n
/SRsY8Z5hyamvsEDp+IB/MjqlhsOA6okNQMxLH+NjlNms+wkgP/3HUheiIwDqW7ejdbZTQW7Fs5Y
eTuvXei+zgBGjrvRMjRILO7LNQPTehNXvZESIw1jrdARaQCnrXIkpZtrpP30+WAZ1x21tPAhcA4T
mUaLvSy72GG+GHUo76IaoYCujn10xtZ+TUv0y32S3q99MDopGabKO5J3GVsg8q9HAPCXHxY2cHGd
UA+7G8NJDSN/Pg9PfTeFUGOCOachel8K1Ij3eJo/Z9E1iAcADvwWbEigKivdNgGU0foyywLcFoTg
tpF1wZVLlwAZFZsmZyfGFS26zFV8Y2Ln1T+/uUYdsEAO0bynDEu1sWMH8R5W/COGc5GV8U6y9tep
ts5eekO8n+krd8TX+rC2hr08EbJO1Xdq0pDoXsQGA9ZCvd5k2/sTIzylt2vJ8NA6WSWAS0/Hlicz
SYie3tQivY5664OaMKQ/gUO1zocD6kKmJ6OIvo9p6UN8ZvQhBZ1SX3d4YXjXgJjnBx6U6eyDj7A7
p3LLah70OsCnQP+VJ1tGi5R7XfvXGzQq8pXiMC4tEfGux9xAKM9Sxtehwm0yuEIhWKGvRgWPF2Ps
VpknEvz+E/jaQf6QY7I263KptFgd9LBb4QVC9L+4vHZhSbbbPoNRqeNJpbFUU0YRY/13PsS5CwOM
8ukv7/VWuKKxwt9uWKPoTveXMkYqzeAH95sWOyod/hrr86XI1f8MiDgypkh84jLmbzdGLXk0OAdX
ukkHXaiEhOeGMeBDisKJLJ9bTFC2DhHOk0e57BMwsfH95Aqz6uBVXaFST+F6cjAAu4sljXxAVQ20
z4/BOlG1pYfk3sdQgMwMItvcpvSWyTdQM7NwSAiGEtZJSZpe/E59iBrrO3W1DRJBT/+pe7JY/Lwx
UW7uifG1L9Ly2R2MxrsbNjSwPTr8JJjuFo7500XUHGEZt+3Zhym9QwqGNmcJwExmXdfidoRAJShp
DuPreJzsKMqGBMb5KCkPri/G3bZimRIjxxgfMxxpCgar0J5YC8Qew2FLArMNiMlDUMDMlfgk14eH
sHo5/cVg4fInF5OS7izbXF4nvq/ysKoOS2/PYLxMYkAHaxKhGS3pFiujBhUQT+IXHOy19batvYyb
KKVTYiNLykmLwhQBZK/cS3sPhmd0olIDz+hCxe2JILbUjtdjXJUcRSh69bR3PCSQjJzbYQYQmP5b
9p8MCiHmb3ro3rKRMJZZh7ShnXUL7eKZgaLLtRwTlNyAKZi8CApDT9Ajdz0lwd9imea+KoVOK7TH
Flq+BG0vRXaAcYe3zab4XzxiDvkQyAG1D4VKxaVy7dW40lBfrastpv6/z3PnxoMs35zYLuq89QhD
3kdiVFKBtWT1AooFTn8usXiiWe8iK/kQCQq/HGZ3A/24mg9tYhvI/+2R5rU+l2a1wwvEn9vh7H6F
3+hE5CrbBjYW23Zl8ZJMDQasXl46LInSh4JIrL8rHteO5iaf/SaeHAoWKcr1MNyM/euWEB0P/lj+
SeeQSTYv215ARdOGVoHqkCnrzcJZIadG2gdDcVpm2590rcJtb+7dOWxPQUt5iNNglt8yzrTy9YGQ
F49F68ge12JPENXeF8nDTYSM+F7UQf8OvfXqf8PlfG4oRD8FON0AXfMQh5851AY/Cp08SX/MeW9F
KoV2V9iO6aBrP/+VkvhhU2grzg+rtRqveQyexOEr8SWahpJ/RKtsCTAaSCVrQrfsgkOAex9A7zCk
2Riv/Fo5INGEGiBBVL9wWcuLD0Ff/Er80yq83RWCU7rdRKXEfPJyfym2OXJpRTAfzhwOmu04SGLK
RI+Z1y28vcWWI3BeqEUu/EsNRDS8fHYuq6U8vyM7WimwByW6pkue3BblzbO55J/sqSHKYHmqPoRN
40pekllc5JP7MDs3pblqMd1HiydvWFRzJsV6U6RRr34E9FfDexZeBYAKV5QeKaMzhU0WSfgIvSul
zhKjRxm2nMPdtyvTLbvWGTjBLj173Aqj6sif/kKi0aXxMzy7jSqy/yusvoo/lV+zObBjEj+igOjk
4qI0moU5x5hxD7ysDki4uklNT1rulAU50VknFwGan6n8UCYF9OIFbwbBGWKindKdf3W6SMp8oF5s
pVoZ0fMc3k1YI0zu9Bjm8WKnco3c2zrkoKVAjhNO562NZ7AMt4Be0RAHv0/Xw5uJrze7ACkQ1t/n
2yqX3EizDtj6YNKXklt567UA7uQYH7e0iVFaAuziTtVzthhh6DY1+6TQGBvW3qnR/JXCr0wucVbH
ZVGO3pPYuGFJ66ZUMkPuVlpuTdNe0UPVZ+2MLq9oGmm0OWYADaKDwAAyqJxCDEBsfYAofObz+k5t
LYmbwRjSM57/yNEWguhdvKRKtDoehP+oktgOOkFy/jjp81v4kf0fytCBVK4tfZKbhfXLVG0Mwk5H
CysXZhBTLA7BA03YBR/ziEspKR70OWBRikDEYGqBZ9lkFUmHfyNjSq/hCMr1wCprFKjkpcSWJ/PD
AB/X6bFHjYvwMrsMuVDn/iIfNPa3ZLGN/gVrRfZ2SHl7SbXr537FFCKkvI/NaIIAx4M0l0eQ+s/8
l3thOW0nYLUrnbr+9MzvO/kg1W+HzSkUvUKk9JgTRC687kWDoq7g0PJ8dc8bjx6j5iIiUkCLiVPl
4J+FkvNkeugv9RbYbqSSBjPDIA6saJ61D1Amb0KOvoDqR6usVqoSEnmiHuWHkIPLGqf+RxqeNLgs
18mEKS6m2gK6Od5QNApoXJQBjDV3jLrqVqdfqtC+W5yGGUen6IWWzL2ZBJ3oMi3G2HiOBEWV2DQ7
tnc+DHy0lHQe6bSkXJwKc0EwmLVTuiSvGmU1QAT7D5VYwCz9Dsz8uNkx+w9n9hhLuwyGYnns6326
d5HinUUJxS7FI1aZdUXR8+RNR9RwHh1C3F8u1DvZabgnyee40giIE7tM98yXeSxh62oWm/TbJulP
H1flWNcAlkFM4risd5ge+v+CkbXSfFdMKl1qKIhQX2hC6ZMqzrRCI4j+bud6KvsHovxmXxYO9r8H
xRYBthV116Px15fvIzo0wEhChecmtBKmOhZtcZPs/8YEbFV6ty7Dcd6l5LjzSnMpgjZgufMDRNIg
5qrOpny+a/KC63HKvz4dZdBQOV9m9FtMepkACwqlrfWc14dXwvr5V0mx9q9mLGROK4Fw0gOZC+wI
X//Hjyr5Mex4VpWi3dVCs6q3XrPayc6QRFmgABSV/gTIEzGGK0ijPtdQTY27uLUwfwhBmK2TzDO3
LvWIBEMzS2BwQ9uc7W3xGnkYj7ot/NV6H6TBu2ET8ADb0/K9OuZ8L1bM901XL/Yi03eW8wNNnMlX
peUnRFNWnQkiN08DhDt5xRsVEji513Hwi6FvzKvNVo3dowIl8ksJSSyq+T7WvcIjsBBn5BFDK99s
2Ffvfr1w0YNnJg8KfuUyd43vJBRLkgUm0ZNnzPS7X6PU4+gPvvAqYtGalMyLYJ7UMqX7Jg25Ndy+
85lC7IeaGVxVSg5+s0lZvVVF3AOL4FFPbRsLDCk+OCYCW/KiWSjOfu5tSuxdxOGYTghb9U4EF+MP
Fbd3xIFCehw25zD98MfbxURuuhY7boNVt7xvcE3SUvX9B7Q6AeS93yZondDJdzJx9OZQB0xUraRa
m7L78ZF3BErONyMrwSILiyK687WiZbePIvY9xbaLdbmejW/ymOOlnEuKuXLPV3ec27oYUiWnGZvN
szu3Nx8yYqxdgD84sJrgLLBg0wMXya/73f9ir5IPkA+rlSiqfpLy2+vr9pXmyeWTvx7sl1FBjx99
L3U2xko2/wU//04lfr3UDmPu2uM81y6fuOiZ3ogHoDynmjmkbj5mc72s1eSCb5v4v1wET4Q3opsx
Em+Ur6dtRgHpEibWl6GDlH4ppWtyKvj3I6g4jAicbzWBqp2a/TnqRlCN9vGPsvGyPiykpzkVNUkk
MkVMru71FxHLBXzQwR5bljILjxgWznlAFA4VQoaG4/RQTyHEjjAgQvEWcpU7PqRrjiOjgq3Mo9Ui
6nGgNZauLoYxfW0Pd+Hx+Qd/7ZIN/VDsVQ0WWNZKe3XT/3V31mT/YvKfLEXDBNPsR1641tFbFq47
nsRRIGq2VMCVu0DkOragq8yM8MFO8JdqCNJyPFuBeXpMFQZKU/KWprMcShLGYmhLlDbDQF8483Dg
/7zkqftxpwynkiGWkihQuXXRJXato/3Qq/z1mTa3xO8SnqjW2kqTxvarDHrtxQvXdSPJGQIk1q7j
kDvyb5U/FN1DGzIWtvMCpdBVSB1U0gjY59AiC3+0byMiL90jBJ+q6M9IsFdgfGPTC760x93B2pxp
mkrtSbgwC22mGaYhq2gMja64+UKkSNKCXTv3rlQD5RJRl5CU240AHOXT56t7qxPicJAICw7wDt+U
HLpULHOU3cm7BCRB8Lz0BaDk6NtTL1Kp/M16UxQe45J7pt0xejqUq5t6umAnWNV6x8H5PYCfIQpR
ik9dGDiLf4v1ASTKH0y4jsXD5nTIZuzP3edG6eLjScoTCQPpSpCXlENR89mYn3/ul7J3uXKqin4J
bwEHEwXdlZCgXx+fUaarVNJuibXI5cpMYv5aytaJVCS9k1kq88r1BmkUjOmbvi/1snV5nUMYFIfI
3MVlERDso8ARFboodbfmF0xpwIkWA1/82LVnJ7D5lEIljFjqBdCeNy/CfxJ/IB9I7vFh9lP5YMim
hTdIbVQSXiRd58I4YLwm+hBUkRzMtVJdXL4t7II+EPn7jwKBKPROeEfVQMv+XjzCr9AglL7mgdWC
M/k6XplF3JWlfkiRazQhX0xX3QWWf4r6Uo+5d/iUlqs7RMJPCfeAiE2GUSCT/gSpkOx158ESYqdM
fo7YEqFW8uXgAyVhYfaNYKrTNB0i53PfrgmUZ1nQB86yI7teDC8ZCP8FYvISwVl9lDZGQAQO//Hd
IN3gOqxUco7px0+Du4Hb5AANwmmoM318CkfkuxkMAnAKz6vqlR7RVNvof7eM624MYeoP6JWnJYoR
YwtjgA+pjdIaIvOWeWrcquM2shh5D5BfYzLpcyyio5epE1+iuY2Pxq7kJPFTHUvZ9iG8Or+MEqXm
vS2RoY2bpNKLmKCwEZRxMY1uhV9M8auEE0Lp0mYyyL4XeO6OH/GTGXfsq/Tx7LwZ4/HF1LDPCnCc
OJN58cKSn0xdqHKtuO1yvesyHWe8vvIpf93FhUAG0c/c05GEydNt8zFv5Rcrh/L/HqhZwoY4SkVk
DL9lMiHy7Gw2UnoGal4JlalaXej7+gFKs13/q17wAmQfrByMi1BN5JRqPHr4oNQwqil3ehlCmsaA
muIzlEzlijpzm0dbrE7XBzh2t4ZchKrGN8y4hvXKNZZUjVbz1p/KPtZJDzbzIhVDLTd90puRLUVN
tv3Pg7FgVbgWlf2GRsR7vyAxryD5l4NG9lwO2EOZ/mLIfR0VTYT93xoWD/pAVKC0rzKsYhPZ+TKV
v8yG4U2JO5Jg4aWEcwyTWnT36/pJ43KAhMYYatHTif15pzV4SDiV+ZZroyDCSBtlAi+jjTiTI6Tl
IZs1oNKcV6ORIfUJUJTyNhf+51+Qo8ymudh9D7Bohn0k+f2nSgET+YEHmpGXl7gTO5HM9/yHL8Hb
0M8uBSIG6ToWraXj+i0LNZHXDXKA+l21lh7n5fLq7jTb4yFVanIx1nvxljLYroOyNv7U0/4AipjB
1g7GmH2MpfflAL/4IfW8vHUa+RflRt8PQEFCKIsnGWvZxDfbX2aILBJpJHvqyMuBhMMRd6Aw6bEj
CUXhGvDw6C+bSETJ53RBHZurXXTKjpZKUDoSIC9bImFxtQpVs6E0Kw5miX/dv3wRaP82zI7BOCvQ
m6CNVWpUp1H/2R0nq3+H+9OBhOOP5MjqAISPr9FMClrnuA1gk9hP2v6GKWjp+dovsUfxf0fRwkBG
5u0bk7n2XVDfQZ5WIpqXhjdKdtPc5M/LsDAOX/hwk9TValXeuxmDbEtlCbbd1cYP/8QRF3OfBS73
IZry6bHq61kwJHX1vWy/Hv2fqHlCGPWukdmDSgqOTmvn9PNieSfvB0OFH/6hu4Dzp2WAwyqWNdXT
HtNBzVguCMh1Nq1zZ0s66o7ZvFzhdiV5P3758e5u5GfmFFn65hsLfDm7aPmXOYyfsxfqxD08ggr4
Jh2VDAiwWj5LX9z6UFIXfm4jouAlFV82KqzvLaXpo64lRg5P0HGR+hucR0e9H5gqJkIAyCTXt4uo
QTVQSVdf/5eX9iCXssbQ+fOhz1P7Qbo38O7NX35nspPBJNOAtZjFlIkPkjuGLvuGHFRblq/Kdwz/
CYZZG1fXxyOkiVNPAQIY/wID/x507RMZFsVZ0b98YMHyXBvrZHpLkEDsrHBRUC9+3Li7CcsZJ5NF
5FxzGILkVrnRuQoL8dPsNW2MXLORxveVmgKYrrIvE/nvdWtBvM5VCtcw08i7+qlBYjVWw0+o31M5
ojrZb8s4Hx79XQiK2QNZAJ89r5yawxI3WwAZgBOLh2cSiNk64meHDwuA1lMCYvbA9TMDGlJO8YR6
9JbVHzba1R3AH3FW5JXZiC83DrzZuPAohBh5lY6coiOgR0KiC2HFa+PfLwX+sIntv87FC2w3iCjV
VJmJrF3D7s2wGoyREBk0/HXdAI6P7yZL+lnSAPXl5xJmmMHMjWJBxxp65ivlOeg9qIdSTCXnwz4k
pUzwrl3i7qzjPy5iuJcbqd/OhmANaOEWg+DtDIIDPDev+PPn0Q+NdbDqmMzxFkcQJmQto08Tqzc6
zxOLX3gFB7eM6gxp6rxM8s3eoH8FzYrldQF1eFwL97E8CNAUBoyMzAs6VXUf2M67LJC+Q4V4kZwx
0+j6oIvMoe9eqmCJmTjfSz2RPL9lYzGUCdfNr46OJk9ZJIG4evaEZMnlHQpzm3me3FOpkpKiKMRy
TBAEyhM6XXspv8ck1fJtqhWppfVShOxUTmJTAtoqlIrUgGs68N3wzLvEGUsAKdC712iQejeuBZkA
IO7/alkmORtKzJpsawxVnB5UBxgq/XJ/OrUwaULu58jqQEUWCuB3sXRszFVC9h/8yF2nw/+pYR5L
aJSvWlrD6dFrKIR2iBxl8FAL8+3VO4Cru2qQCq8K+3HNcm4OwLiAhWKrYvqo7AyA3LsCzZorDf6o
Dvv7PvpkeGN02AlrqtVm5nLCdzMhTPP7qvjxQ8Sa9ls9wI8PVOlVZ0EwUR2QRLwJZRJKu8a7UgDi
HDxep2QT5n4iTwJ/qBBpLVoJhyW2rB1L1R4TAHdHRpBxFdeEeGbL53eG6Z0y60gyvsPUW71UQz4t
lnbL49MS/j673lMEB3XP0HfhlsROOP3D0NjsBD/dJbVfB0IMyYCwdnw2XJfy6QzP4wADGDBtatNm
6kcXTghaKhRhHd30EXjOCxAMpiYJEpHZEUV857qob3w+xsbwDsFmdKES3FFr8yDMz4/6lt70pXKn
lSN+T+AufRuvAhDLFFDlRFHQitK4EHD6Dd7+cDZeUcUJ9YlvJgsR1kcurBS12j//fu4niok5jf6F
I+iS6wP0UkHQOkvaA2SfsZ1bB6D/u4vZ6gPQMyBGn11PrxTJEF+KGx9CEpJxElbhFSoT641wK8jn
qBc0u+TsNjYRDwWY2zmyynkY+grVaO0uh/byZuwP+uC8od3t9So/HxsiYsRiJ0a1ZRUHNfMRAQfm
urABlJtNmpn9bVnoBXooCzQVc3nCPawz98fr70fiuOslFlz7eY2FZo9zkOjfQqFEUBiK32m+UCyS
zIr/ljJtI8BBWRCYers6YV8kqyvRJ+5nrOWy07RHI1hgevNS69vogTXDTRdF/hRxUrLGx9c5xKUt
jGkQXzctaFwesCW356nbvYrFcSIM7ohEZgM7XGJmQSGvTShvNr+2Jm3+O/B0eTB0RGVM1vg1sVBQ
cKONbTbzxCZRmw2W37qke7w1uqwszXOPpnnDpuxjO695HzASwcKtLo0EsT43RLfdzS7zd5oBfZxn
F+S6fhoIDsvjXE/CzBEFw1pHMKQaIwSl5YxMeo4SgpI+rvSeqwQW+uVUDVTv+nRQ7SzcE+ekR9B8
fRoe30HYz5OFbChFNNCQLh+X5RMUfYjhrxGYMqe4Mw8qfcUs1dcOGRSLehj4Li1KYu1f6J65Js1H
P6Mu/0g1CwMp90pJPhzWajyirMjJUddpOX63M2gn4robBi+WDIfUlgLnY2lvg45grpegl7GYQJC0
TFb3JFewj5/vQAJ+cDtxB7R3uukOsnzDlAsgx6TeqowejD/l9A8HKp0ge6g8lK27IlRUpnqoytqW
KQa+qEhSI9tTfLhuR3DqARYLUOzZr5P+Qjy51tAe6CPXCNyhMETQdmRsHtV2sioVOCVFqnE2wabM
C4WhJrEi/uI7mfGThE17G7X+uQaHyX+6pfBjoJZb39eDad2ZSmfI/QNydtZApTnjSoNbbPpBrclf
iPxKVHee4pj8qhJsKM39FKoEH5Xr1kjNdNPWneuLzhejPMyJdGeQpeyHF3OE0tsvAxyNBeZdPrqk
Ge3UrHtWOT4zlNzAnwVHwPSx/tqTaKNkNFV73c/3UB7fB9WzlQ3BK/gzhx0QsrYD3E35sB9tM5rR
mhGlM/O8WmuRB+Lg3hk1UxC6vwyvzmfLc86S7RToX4QQPKIbBz/i35bKnaaxBmitoPZfWvJXDzaw
PvZzUQKE2JEvUooIbCXfJbsyeVTYkdhLp078Hi5HzvJm2rW4+i4bTCWFUHq0pFj4pvCW+CYy5w+3
83gis6/GwVYPh6DBMGBzB5M80Dqx3xesMV3FK/dVEvj1tvGTXf7vf3TjRf+7187pGgMTucNwfOWC
JzcSuDSIyNvHsApxu99ElOr7Uy++rSktFvWGk/ue0D40/2i/hTZZjqjlL+WeGHn+HYO+tKnhcIV8
pC/G3f5VDn9WE+PSlIopqtTH0xF766aLSlk7imSLxCtHMIrMZwapQGQH0cKPbodINBrg0nUQyM7F
U/ANxbfl13Fc/1ldli8ZVbHCA8Og2Z9XXzPszGdDiMP4ll4gaxIRbGlUOVgdHuBXwDMh5v5r9m4I
PPDzhd16J6gUOPtPsXWEHRUF6eqqCUPg2ugHoJOL6cWCHWw11qGrfTcoIH/R4+Om3glDz6/a70si
yj8u+BRdnlvjz5VwqnHzteHHXV7KjUBLNfx9MJNcpBy3dfwfxyzOxe6AS+P/VKRO7vxPF1G0AIts
2SnDYn2iPGGXG/LHV5M1NhtPX4JuS80R1wP2rf4v0ByH1BiyC1rtP/b/mexkd4RQhMKabyubmmq6
2ZOMx6tS3OVAguaTbocXMBzpp3ElE/Q7Fny8NcPyII+qGMwf/lOCNlOQ2twXWnfgw1kPZCRdX7FB
TG/Hd8JYMpuW23T2dxow1u5cEVWTnRw8K6wusuydM2uQ1YTVC9wmiDiuAdfEKlzsMzXG6MCD7Tqn
N552TtSerlR72doimpuCwLLWvJYzF1iXsDT369dDMgL25ZJ8J2XYXWzCjOpJJzjXqw+svNwmHY8z
gmfPNAajtZntdZmh7o6La02O9+GW2zQO3DdwTkSwr7FGJPgFjFzGn1alN+qan8ixHRiyhJOAe4jF
oZnb+xpiZAahUTM7nJ7yMAvRqtG+KNn/qL7/zi/yF6V/JezE+coBz/h8V06zTXLjHuC9G929pXsx
XFRXdHsrUu8W5iiG1zKGMQzl03tz7KjfENRiCKhwq2R3rP9WS7LqvzbxvjpAS2hDOklHXNVsKqYU
opeISu1ZJKzTM9vrTL02ABO424qEOo3GtL4vWAhyBT7UE94KGQgwkMKBujTMwuHKLMbEtP5Idm38
mg2Op5cZtWaBENRBR7GtodS+7LgWfpUxP0A8kNRFBaQXdb4jyGsItGCAfXcT3P7QBEcfFogFmACm
P1PpgZFtv0gZnYL8j/tdB13RRE7ddy7Wb6eJOyqXmhy2LdVEN34brFmJDeIc16Gze3uF613G0vY2
T+PUPY5VU2wHQgJbKrOKYpnDHxGcYDOf+xkLev3U7ilhZCIVkO1Oaga1Vk9osYvlzKHiIBezHIHb
Dg98lFEl8gKmyLACHpu3GNH2WnJLUT0bIKN7Ue5BhiBF0MIFceGuVhIzeErbgquiQvM420q0mg2u
aTvfRuBZQ5WMYKqhXeyJS1QMpDuPFtZjLTO0i+RaCYGORIkAdoERVMxIAJ4Y1ZZ520E0+ueZpc6R
GaXsXxQ+QsD1LGsUvYmOYcQyEb82A3qJ2wwcUbzKt0raKm1g+q/zQd7M5cNV/w3SSPXtWrOk05iY
n4hI3ZEmeg63sZF5BtTUaoKvxH7zI12E5s6IKwc21Q86Nt0GNg/nGMcFn2QwvQtBZ/cKxsoRC2yz
Ng4sGfzAn3lhNa3aJsoRkeqLUbRexypl/hTZ5TGFFG3epguw0I01U+GxnhQfbeJ00FoWWU5iZm3X
uVoCG6P0mmyJXRRHhllXwEihfWtqpGIsSvynzwanbSlXyS6ZoqUTDiG53p/5ttMG01TsvQZGFdrr
W3w2vO7b7tnRFiiJc/q4vR3BNCDKBN9DAnLqW+NFNFl9a1eJOSrbaRk66iVLiJOaA0g+OIBg3xaW
8NjLNZslhIE3k54+o9OBu7nG2gfr3i30tWcsosRTOUHEWo4Vy5kVlZvAJBqNY1vlxRvkVBk1cgLx
1pEuziNrfDsLMQalUG1aj0DgVUuFegJnNqOKmlY79bsNdYBTr7ITZJuqL2YP3f7+GS1aCONjwlwC
NcnWT+UEEEfRIaM9JPxKfJ63LS52LMEBB61oRFP2MF+Wt41Zvg7ZWJA0tBlRR8kKSOy6ZfK9HWqQ
TjYVGeoUBr/ak8dWFlIAfZnCSZ6+UpajLc/wetW2P+QGiP3TygDJ/2oY67p4lOJfaskmcpftjNk/
UogZQj6rKBuw+V8U4Ou9SRRAM+cw26aP/+FWASJ0oAh480qeuQ0Fi+da33D4dIDpDnvXlbYWAnD3
/2bQ9MTui6dTV+HXgboCDuipSIQJCob16Oaf8mfXfpAZiznInfZF3G44h89fh38C84vYmiK1rSoo
H3CCMrsDQNfem3JL9RaBP5s/EfP/LSJqMJM2ePpo1WYymo/OCyJTMbV50w5rEoQMM8HiugGUpfar
AicE5u4P6iAvFo6IQujNDFfz0fpb096xx00MDcZWab8ymBxfvctE/FEaricCnl3pb83l6J+b0eDQ
qht5V6+dHsmp5aBbY/lzL+Ugv5Jh6YqspNaKHccRL3HOkCDSQwGxqM8qaPT98Y4sOG+td+3ds9Ih
16VcPGqZm0fnIY2DiNrEH70XmiYIJT0qZH2Zpmb7ed/+hC8+/71OCoxmW/FSE8id2X6UKoluXNQU
Dlm7UltZQjR+gyIiEJW592dJVFF8fDQkcerDYgKNhRK6ARcocF/fY6xRWqkJLVdVD2QVJ2Z3WqtZ
W2V81wXGdu6D2pVw4lVqtB6gtrfmMXgo+M1ru17l8XsVFxWWOwi0JS5b8nB3npOy+0mrZXg7Th38
NeTQFgcaSF51Jfa2LgV0V9p7iPBKHHJWBtXcnMKA5ovhkOrizji6eDnmjMBYykwUSyXLW7h5OKBC
EOWYR4agy2zrTtii3q9pO6upzDa7b8uj1QByGjKpAH/zXioQtC4QfhLR21AaAKGXv1Z3oxq5Qu9K
nls9r2etZlDLwa2JnhXd7SYmyy1WiHuxl6NP/KAbwPRk/DcC2iKU8epKiXIF8emuWL2wfjoVPp7h
AKwBJb0jyA4oXKuCMFjwN/YoKpASoPf2RwzH7jGyo3GfcD2k6hwhKy48SgL45NR5jwZCFG+AHa8R
l13l5LNIvrCfC9xQhbF1tN6cyCSvJWq6i1CoBtEK4LAruv3plyHiqXPXs7qxzoyLC7SxF5u+qrVE
nxSww/ott7hwf4TaYmwLb/RDlRM9xWAAv/oo2lFcXcI8DCW2/XsTaH3Uu3ylXYN0cEtWZqzqrFer
MXVbbF6IfPMC0+AM3stqVz8gQKx+D+kIq5+C5y1K6KUIPfqdY+8H+e6JJV2PwN6YLk89tZE06eY+
9Q5lRto3b4bxblM1huafPEQJHDmve7fxZ6n/2Bof8RBKIx+7KsrpeP9YMx9eAVLC7Ua2u5srpc4V
h/aaeglJ6I/kY3Pgy+YdJ94L6+atN7Tu2U7EMlIIxFtlRGKIKVezHtpEhbR7eAZ23STWxbQ4HeEZ
QuTS5BsCPUeH3+PDGVYK+WbOw7JJLk0KLvFdwbcn7nYi6oxF7ijcr3nY4lmqRt+BBhJWVCYOdvwZ
wRDJcX7nsELfWIWgLnuzCKEPFDUiZgbExWyoRiSXXWk+BjtDzSdljF2bTgJUeDE573MEsXb/07Zd
cBalajpZdQfVQhA+dvgBBioQVLa86KJ8tI9SIAXEtAv+jeelYcX1o6bkPcErbNEyaoT5ZJCukwR2
BCvAeMD8QKp+t1VDrUsuJbjvf+C31y3HidKqFW8PAR3eoXFonOX8IioBGpj9LO0QK7Dzlne6VlGn
iSC1/Y0chrMcq3CBV4F67p7guLixq+TGVvsvSK1nhnAOQDcySLp2esqPvq6PuTzjmzQ3K3jJHs3i
azTrCKwcnVVUm8ntZPYG2uXm8W8ZOGjw5kn3KalGWcQ3poOYV4Px7cINr50HW+Ro4IH5nuIYViPA
gN6ejf/CStjQJ1Q+7T/8+Xywop/Qwkssta5KMeLTDHB2rntMFaZpIokpc/2sULyFGqgWNt0erof0
Eoms5FGYBvdyCW8AsV5ESF6dmNU8I8IiRXbfcnPDoEh9Yo7Y4lW43AUosfT6WsC/5WEtXcJtSis4
gxp1ULk6AUuDYxQbj4PKlAuoDI2PnlIHwD62JMbO23TW/HTuxQFw4Oxtt7aoN7m3CAt3cAAV479B
PTsdRIKRMUspY1YoBjyvizfYXBgprnbyfNdeUF78PClKTUCMpo5BAF+hmBCoI9SCO6rSR3likoWt
0zkjf5QE9VGn1zH0txaBYjBUuwUv8QNOOBrc99KVHg+Dte9lIREuL0ywWS12AiTliC187rzNS7eU
JACMd6CDcxd9F/8hveiKqPFtLRfsqsuJTyPZoyqjh/k6rwZ5WGrmV0xnBqBsocvdRgLibIIqcyj+
Pdwd+Ji2Rn9Lh5MYn+6evWL6QnTIB3z8pWQX6s02ungnCc8dicfKW/X4Yi8NzgFx5fHBFgoqcT+3
vi/F1GFk6Aq28eDjaDumquQKagVtEXvDg0KfxcYJEJeseB+bC2SVflD2z/PoOYm/T4h5re4f20EG
tsRhjgE+l0jfI9dV87K9A1MVCyvS9cyjw1LoyJZMfvzkDl3a75QfgmaDjvdA6asd15PzGJwm7KPL
YhL84Aqezhq5nejZcAHGiMleGmIjnVYqnqBopYi+Yir5ymoOqRvbrwq+5OrmICJgVs5aUetwt39m
4voSceoEDMstTuQqK3EtZKGjvJJrTT4c3MLx61ltLYdRr0oD1JgXV7PADHGkVmYmOeIynVn7VZqR
H6w58+nYYHfzDYJJRHB+irEeea6l6uAkyuSJssJVPJQgosf41Dm/OKPkdPviRm9crPYjj9/1N7Hh
X9YZHNzxgs5Qm7RAXG1GWOnYyP4aZrJ+iiw1ralhCFZ42/rZIaUhYKZ/uG8qFVzafFgsorVXL8/r
FF8GVRpzCyMhxnUy2k/QyOAsvFUfSi9D5hekeFB7dI+lh30qBxSUtoV5GD2ZEAGhBtrxUUMfzLM0
nl+m+Jy55Yq9ElVVPlQElr95v2q6w459Hvg0DzF6Ci0YrAHWjvbGwBZjsr3zXEoSOfHXn3/NsdAh
Cl6lHes9gros20pOZjTeDBcLHOlSgBZ64wWq4846jwRuatNKV/G4ejNXEzVJO7j0I79JeIJInIh4
liYBcsHdSSpnBkaImsMjU2xGUcowZ3PvTXu8hSFQWHvVk3LlH6l/pQnaj9fLhO62xF8fd0NLkdOY
24vFiCFwZGaIv6cs2Y8qbXv5I+pf2wLKPTN6jQFZv8Sy/K+JaQUSa7Z0Tx0WACg/F3sNU7KDcRCH
/m080VH2JyM5MXSEO45COl8qjslBqtvUOOVlHCJclMfq98L5oZ+ws0ZLBwz7C2WXnMCya9l3Em6S
ezZLLMscClrb3cFZ2hfze13IBEpROYpkQUjoBlmbI6aBpVYgkAJlbnHahvh18AGdWQUGjzApOlnL
cDWpHXmpJj+CZcsOPO/vkb5HAYufMq+NtluJ7mX+E/rLLqKUmSGWlzNyAKjzV2rS+xI+21KLEHbu
4UJXq7TPik88GRXduEJa5QodQCKbNCkaDkBOkDyeAVcJYhTMbzrF9el/WT5a8aC+lqKno85GGKdD
SDWpBAHqZ5HaQsQERGbvmcac70JjNrkWJ0nnwARUkOJ1wBbGgDpVsz+SgQQRFyxRwjr15WRkBY9Y
SzSHyEz3CnYv4kqBLBQZkUnQ7PqeOskBaS1tIJCaRXHLd6tavlkS8TI9gCiswcMpK4XW0uYaCP9j
8ch8X6CYCd0Q656/HqMjBsGJwl+G8AfadLXQ9zkbx8AziIbDqV2AeJQPFaG4mPfsa9sVznu7t66Q
lfTWmldyhzEV92lSFXmDe78aCFUfK3o+eqp6Hv880e90IcIosRM/ELUY3FX9ZIOpFn0ODTf6bz3Q
t4vzFXH17Tn4AXTtxj2vPiO8muaIrX7DH08kJEsxv+vgH4LJnn3xtOrWzzto/ccCz4svfEylYV+u
quPLDdA1bLfsUW/0fIdFXdL5oA+JU5ptIBxDxQ3cYrwTTiD3oEGLo0kVVTcte1G+GqHRu37wNTBs
r+4lEK+Wo4McAjhvAtC9H5MiF7YANIaJvmZH0CrA2aEJh+1PploNpRaA4IrCHK+C5HVW+176D2cy
xR7YqU/+JwUCClIIpHIvQd2gl49QO8msvkNxxA85ca46GLgyFfK0ahr2JmKDRJf1RRuKGXeL3XQk
baG4qDVxL+ko6uKeIhxpACUJfCvAFbJIFu8xeM3ZpyQbpeuR2yvKLw5hxSgYF6Kml2t5A/5TkRZq
CKYcM8n31mjNLufT6ZEdmC4duH1dA+RFkYeBujlckOBAjKjFGotDEY6lFwBRgNbxe6ky6raURhwJ
+KHIAAMAgszB8XpuT1M2TMvRyRCXMje0LrzwHIbVR5EG6fyXNAe1atQC3q0q+KRPeCvzprNOIS75
/s+wj5yHhpo+3Voxo5fY0LfWJgQt489ZaaCl6fCfBgv743G9FQkaPljMdFzAm8+h10lVMjZdxrZ8
NMdY31WNkhsBehkDZml+NFPO2J+EdjA9pYldd+HaHf5HK1G52YAlI8wn3/jZyPLyJzQQTJNZSSto
qHgW3Nks/mluiAb40G2eQqkFc0UL+bQovxE9gV/7hPBxnzZnLcGwT2E5b3Z7WGGxAR6ibyN7AmGF
o54ZzQ+KXoH2O73wS/17sXiEhvNEXImu1lgyhXLiArc7Wqy+MHMwoO65dswCz7MT+M/2cicGwXoi
bsFR7uDmRW2K6zbc2L9UYlCI+QWXg5f0rF+5dv+7TDShEt/8/XSOblgqCu+iJD4h4V6m+0OyNyqG
+O9bMkQFnONxwjCy2XKohPC6aIFfl9STpuy3GsLrcVOQqAS3psQwCy8NtXMEOab2IwakZISSnLiU
/8SkMUk2wadreFYM/SuRdzuTbSSJqUT247tscndE/QbczPDV9kop7qDRAvbHhZk/yPBl+31P9O1g
AijW7x0IlP3Ap2FNO99pAduRgWrBIKHzFQ8EqwSlUjY0EYYzq29XF9SEkYqFkc7XAI9WPqta7E4U
DEWUL8SgXj3fbobEhMTp+A7+E3k3x9smjJ1MidRvzcJnwssb9a1YYwq09Xt58ON0KGYXzTdpgpP5
/ho9tXsEDCK9Cb2XrP2E/ke17XwbzLuJZPk7UVPVoDT95TOGNBakAbxe4F7l4RsH64X1jiOqgbYE
bDwyC3ufpaTDPaUithDHyOATml9ZHg8d1I0QmFpTHVpjFBw4q72iNWwXA37jpq1wpKOzS4XJTt1T
DKenhMjkPZ/gDVhGkm2GFRoOl1tX8DawHw7LLdg2HYndjEfiIqDpnlYfEIUYZIY8B5xqZj+PS2qc
O7Q0DLspbmshE6EVJKL7ug9H6z9TvlhAlVanxfwFfZRxRvZKRTVoDivJZXYN19ExHVhgFVANEfmJ
MxDLhcdkbg1jzmU6vWfqiNxXB9aOyJWkAIYE/IpKxFkPX5+G4VmcOyApbggbrEEFOZYllH6tkOSH
xbYISq+Ygty1qvHe7/sFQlqXoERUSclg2vyRAt90kGS9okcXquwunhHgyJSQ4v/9t1f0ep69uV/a
0GlDxD461Qqp0K+3yFcu0H253VK+CqoDYea0Dc14EYIeVQHeglbaLrxyJXWm4JoNANnJVPvIZheI
jWzjRKcTneAsAph7duQsZxpWL534DBYel21RJR9odwnYEZDkyHNyT1fRYjc63UXKABvwB5slpmjI
g3JUH6c8UjAqqYZ6exszHxXFAUBfTOWEOPB7ivn5zpklJMkrTH/RxUuQB7QJXA/f7epqnMinAmR0
YafkNT2EEkKXz9T9W/QPPb0VIGXt7QsovTvMy5EBKKEHat6G7xsr1aoUjNRyUbN6ySBrfWZphWbr
5oKwmTfCHku4BJtDeP0yDf1mVaBhY4tX2jn6HkrCf8AK5AUEkDJH6Q0iHeAoc+J3c+10x8hLutsq
Lqp+7+TEB8/CfDMO/VpckOF3Oqj78sq1Suz2Vyv3znF5Pe2Qr9GXOFOHfOf1PrBpsMeEMjcJbOz1
IczBr26olzh012h3MYhUtR01EhTWRJZ35yS3xBux3V5Rv++ws8L8LkvJMeURXVVH7DHZsUsFbv/V
jUDW6G8PcEVLlmNGs3ZDb7YBcsRzA2fD92nYDJmH24srpT9Ht9ilef1N5ReJtozypfxOuTVAAKas
C0YzRFEpw3MjQENzJIqVSZH2EvaJo2w33sfLBnKwj4ZGb6cHzGh5rpoq97S64NBZIEMKD4KAv6Gn
n3v1cDscdxHKoX6XJ/2yvZ5QmKjGy2ojHQ23WZD2X9vzUNw9IXWjELKblVn9wZmEf510xQNdl1V5
oxMbnZ2DgNWJunxbhvv/C2z/D4mekU9aiOWJXcLOPnQss3Frnts0xtt9VZ12hrBwhRPexJhjccMY
DlllUlS9yiPdqWpe1n8UJjY+ZKfMnGVgho8b35jWgRPmnOczVbhPVNefnAeOITHYAZTZ2k6luyed
ROHcoJRb964hzY1oGM5DYjbrqDZrHfdLBcKXAsMXp1teIymzDdR/EcOwmniMofNC6924w+hVsTag
sHkwskOkLrru8wm/FAdtKikSGnkX4H6nnpJmKFZiWOZmWgNO+GB8Vy/g92B6qN2Sp1t1gCPtKH7w
DRxM2O6ZBV6GoNZhHIkoiSdacEfntIOjk+Lbt3l/LDwBQgMA37jpEJ4dkMBwNHHfMUHn9yt6vbSc
X0KG5tB179kTxV6ElISdxkhVmIlqdZvABZPzWPh/q7O2J5xaTTcokHVXcp53rLRhufbgshlDuB5/
7LFD4UeT5tutLI44Pdd4BYCqugPQlZILQQQY9ILeXDvuPk3JglFBejodBofR+JU2qNig+1Nt3rlU
OadLM5Hfs2rehb5aUVGjkxfHx5PCXS2mO4UD1r5ht6/2S4tqlQ4NKWwiu1c7RMJdr694OAeFBMZ8
o3XsNCRRd6grPwMrZEw9HWSRHZclIS3GjzAfPc6FAJasvIRVF/6zJYddzH9a7hFiK35VT8nuvWOT
o9stNv9BgmxRbG9VEWRPid8IKKRTAqR/qHEwroL/bC+kcc0zk3zRTFZLE6iq00ETctUfVbT7GzyZ
SbKMDEs6i0200STAl1brMS69HKeHTy6gFhIoOHH8Ttd/RRKSapR8n6k2r1/AsDujPhbP18LUpTkR
vLOfKILf121LOQ9ZzkzjUsjs0mttm6hohuewG9dSNmv3kXcxqTsPXV7DeTSGbKoGnvw4xhJZ1ebP
jCkNqDs4yWxBQEVsUqXjfuxztUgrWlq0nK68sxhb7npWJ2bexzCE2f6AFle88Vgd9m6UAMk2FusA
cADWcKWzoFjBWDJ7tWcTAAKRqn2MlGUO70Z2E9JlboSCINFmhuJqbyQpdz1SXvK8XlqR6cmIPfU/
icwgjNoF+VG/E1+IVWBFS/r8T9q92Q7/JeHSuNn+gURS6Sg8inhvgfhr0oWZQfVwjdX7V6/aQRaY
NVIqBCkUwd1GSNueQqnld53ZzGk+fSrobdmxM4OQx3fTFApOL0CMMtY/4drct6LaEfA4D0mYKWQd
vWWglRr4Ao/wtuFV1O9Gey2ero+M+WGMiCAmsA4b3vP8ISgE3/dlWqGxETBXtg+YWs+TjR3Nh1Lf
ENK0rnvMMh7yKmrHm0GqpqrJm1ZiiGSUiD0HkL6n6mru/Xq/KG3UblQVbsF0ieLkJ2fAdGARj153
hnhzk9dlvASeNDurywjBU41fVgMWOGuGxw1NUGTLQPTZ3HhETPEUjcKnMW9zD0jYKgyRiUqFoyGO
vw3Hd3AI2m+yv01j3VGB5UAAEJkGUPOLfSir5YfZTK8XO9lSHNHyV4myrcKtn6AJsrL8YZlhj6Ve
eMbPpYGXs666f+BH4V0KuaU7LquJU4vOOd7uclHYJ69Pvpfp8vfP2OMRwKb/UE/qgGVOVppaFKUp
xh5NNJJWXNj0LhjGScm7nPP1V2ACkqikEUYUMrKI2o5kIwra3eS8mEkulWLfQ6TliB3oOSCTnDfy
xvcPZxuN+wxAC93VRhiwPEFmjLnNW0gmzkWJpl0DJBomfdqKHEVMWd7iHXKRwRCZYPVtmcKttNqB
rz26lt9MKSsNMB3z7kJSd7tcE7aggZc1trDkZxRn6oBbL/CnGgMb3LhsJY2oX7xv5l+ochjS8tUO
RHJ39AMbm7SIVqqvT03I8ucoU/4pjUjf4I8volANBLrJkAFXoQ5J0YoimHPgw/vGVUc9ctp8teht
HlDOl7hjqsd1ND86D9AEAUxkCM96RfY4w/WdOGyWZX3c1vKUPiX4dXLUITTvpGJSHM+bxHEiEUGy
5W+4k0Yk2o9pBCJ6GcKpLOK6uuRHMbUzHVzAmjVsKstiRfN7tbFS72pxEsWFaAxU9y17EMLQF5u9
XgsI+Vcp0+wTwT5LCi7Ssq0KiuQYfbPfPpw2tl3f2Otls1nzUQI7G+/aD7C1IzZM8KsMHSEBEQtj
KB8/YwRzt4zVIHH/gfYriIvhwKmYWdznLbCY38z6/lK7RALbceosLba6jcbhL5M/hDqoiPoWF/3V
f0/w/Yce2eZVF3s7E44apLwJszVfFzCZeNktAPxlBQBZkStbotchzZ3bp3tgoBzU9iVhoZxO5Sab
aIFZuXCfcGF9A8C1zdZV14doltXG+/XVPo32Rt66KooTlV2f+4/5mi0cAFAA9u5mZ4BiToS7AezJ
QRldXyoGLjHM9Yybl9yAIc1miCsptAC5MgQQtaa19cQsxYWlqmCyTsq5Bxl12k1+NNRqnbTKhoFu
nEGQ0h7WZPX618iCacBaIh6BrqOfziYiVvKDLfvkwQkOWcXu+8gk2ugKHJdkpD9hZy+Hq2cxJtHS
R48GMz3RqB92WJcQwkZmQ9IsgK3vIo5ogWCaZfGFH6fweudWTSI6VC6OLb5lgjSzQA4/HY/IngNv
i1T+8BNKhEBVZJ+V8v4HHnY2iybiHuUPzMrNX6/FN7ZlIHIEC9tXs1Xr03DaO9eoU8xWz+7G2vCq
+jwcPhF24NWs0IXTf/oHC6LEFpFYNTvU1VL1HVsUpY2ss1TW+NL3NyHnAB2TvCsBP5+qn/S6SPxu
l7QAmNbiys9VG2HayQfxgnePREZMWHBn4BJgKH3s7tp4TciT4Dmw5DfirhSneOAGJuheBNqc68Dn
hQ/1xdnns+SXLgj/RFcpoTOErl4swlydmSSiH1UN+q+7dLJFwHC52uC1Q6uyi4Zf8giPqVWMTc4t
qIjSNdfLHu3LSgnDzYJk5RI6GEpDM7NEAMm65MHt4r+ufVBJv43xzUevM5J/7T9swPYH8QW5tkEi
untegy3oAFJwQ517Oo6xF7ENhftoM/D8De1IgM4VYkY0NSqQNGwWfXhU9i9769tQJK3e8TxpPMZ6
v144eXgU0/ZDAGIN6a7lQLrNdifNnSjdD5nna64LGzJs0O6M3FUWWPObr0CRpXqyBsMGuKciF4ZB
1v4rTXU3Xwu2vgaAGG5Tov0VP4ERHhrnxy93sihYHJtlK4kTb+S3uWfFXaRyawx1lfryHVSXesnF
UcT9Y5/7gOa2UGUNbX0FK1rYqU0V7b36Edi8rSXB1d1HAvKLWFO82xJ7SHjL+1A6eSQma9Q6Tejf
IYGoBXpCUPw2OQZ7a41Gwu+gohdzXJ91h3B4ssWaqpw9Ke6EeE1Kdk4YPvBkxmLStEZzaWzFwsyh
Ax1MsOl9BAbxfVpPo2nHHAcn6w1i1Ppqx6AGku8kVGHjjYdk9NpRNtZPiDTHpOj1hKcjbvZUz982
1tBIrU1phL7nQ92XelW/MYrUQ0ibqVM7091v67NbPCFydXDN42v12d+3mwZVq374XbahXXndinEI
nhEvu83UuZa1pj/adyn9p3e8xuwGd+Sqw4IF/1nF1FD0M7sQ254nnVgcYXx5kGvgZSLniwE4VRXZ
QLXO/ZORXE3O/zEO8sGcFr9CR4wHHckfOm6ebYiU6DN4ewUxeyaakl2VUzOkqwI2VN71NPOa10rB
2ScmuqPAEHgH/6Y0hWgmp6AdPgG8Er6yUUkrzYJfRWEZcKibsAP8LYLfhnEXttHMgBecKum6L0Cz
OvLmovbhW8jMiia5RtKdnyT1MtuDi/j4Q63OXuh+qziWkjTs5+A6SHad4ysEnbxM/LTs6vwjLaWt
VW6XBjdd/TiDxmPAW8ySOJEamQQbyRK1eLHx59WguX4yHRJ+tN6fSuggO6EGbupp8uaILddHWLuk
gtpo/B1oyjCEaDAmn3OhOSKHgCAGvgXEgE9IsvJfdvRlsye/jPs6KerxdxWIvZV0oBUYOPuGvrzq
e/FeBUxNRv2gHZpqOMB/dSUw2JaHKh2wWaB7Lk6bL3/nhaVnF3aZCdOI+59ov24B4Go7pr4iaTRv
gG7BE3N/umIW4ofnqYD9JejEVle19ffPWZYZUzYBYoaRomtu3ZTRo3Ym68Sfy7yVkwlzfTpLI+CP
c9jkRbh3BhpsgFcWvRy2nm8Fnvecea7tVY9xklE45srs9JNCyWKJ/s6r9i1CFgifrZxzqVmCcXsY
P3S3A7No2fN1UCYMvGj7iIekimE3BffWoIEcmPICFgvxjRHgYS9RCaLmQddcdz5kbsz6HgVrBu18
IPuEe+rSRTKXXIu2ex1EBx4z15F+FQcSQWthWt4H2wWujr2eK0d6/rGWxPWYUk5ci2tUs92FqwtA
VT09H3opIgTGmwUq3CHPUs9X8qJTdR8ggvRcLSyZe1vFdHfRf97WxE0xY58YRPb7du9YtQH2ZVM4
wLY42qX66+K4Cr6ttEcpLzVsQa1vF1A+VjNWXaIbtuh1yDo21gkezpvD8PfqjfAk7YxIZh5ben+V
ZJzERXIIGvuUj9aJrjrwXigxdHk9JeGS8/lcMFVEzAhJUgkZafnJNw/4dosoS+cuJcZu1+q28WS1
58sy+G6hL3sLaI6u2mEK8rRHu3lV9Qr4XBgYHR51XgPH8GVarWSWvtAq0z71Nav0jlALwhqC8JhR
mWKSmTALG1NhlpbErJtigoJN2kUjmWB1oFHNqS6VTw86i2z9BBrmtUnTIXrni26jwl5eVwBLf0F8
C1VZM+G9CJ94wJQ18C1JlJ7hIyOJXDTFHaM//w3NsuaRC0sGkvmiBd20o9iNl5ijxKBB/nRkWrVU
9xPtVjI8pC/6Q8zHglQ21GH2EONLVFovDKgJ5TDSRkUNFoD732CJhUTaXA0s+2/WUJ6JKL2X0XOi
GKFNYotx/aY5MtFldH6Ztz2znvQawjL73vrb9KwZv0Cq6b6hNUS2gxmQWzanRD0juLB4V5SL2BEE
2FY9IElHUcoDVpzaGJmfX7G0lpVNbjlFD3lu66Xvz4SjhtCVHr0X16RvO/Myfrv9XiXuiabJYNfk
uQtF09PaH3HxR4DOYu2dAevlvWB4oQHr98aYrYMmNDgiY0qRigwlOzouGC4X5woJ71DGQQDkGJUm
BKj+wmNfqSzzMm9kJEg9QvIfw5COy/Q3SmJlI8ij4GJViXprwTWu5XqAbVg27BTh4UzWIr5jAzn/
cNf9+qLzvCo+VYBGOqCeFNJQ7gKyekBVv0D+lUAGYneqEDYg2mEq5J9TBPscnw0Nrp79crZoYhOJ
9EhM113t4B/00On+PzRftoo4ezC/yKIuLLJ7ueov8xWfYTo7PvrnW6dNG12BI0mW1ZZ0dWM7eZ8C
xJxDSsrM5C8+YJy5bftL07v8vhcFq0+Jx9aVXcaJgMd9aS9cE6ooeoVjpuG/NK8YfV95Ua0uWExB
QPfgjTW9D1lCrgiD44BDMkbkBsk1i860SBhMt+/+aadfxYA9G6r+A+zNjpmnSWLskwP8uFvohzZ+
N7DeWpBoCC9Fu67Sbe8UhjLiCeDXuCEED53Qu6PdCj3yGlASO/9++S3yqb4DgCJjnnUN6k6LcvAA
xUAGo7/F3n9lwoVTSuz4n82v15Cl/9qWymRDcNNLmmWbDtQXVlTMenVA9GU7T7yTrA93F9C+8CjS
7h3NaSOQ4sM8uP5AAuswxPd032C9225ieXWHu93hmUtpLUez9enQPRVV5Bx264wSwumg13plbdT1
4l89YWZgyq5GM8+VSP4CLanCbAvmqrUuL52YBqtHjt5g/dnzGQmXRFPtUZfd9ijVmOqc3m6aH9EE
GBZU4vpD2IqM6kaNa+/UZJbouD2aunLYNo3Lom6abBJCjMZ0VVDL6B8DOIVMRmUKw0AWFIicXH42
TN01silsBgqIBzm3vZd6VnUP8eK5nDBZYd8xZdj+JNFxUmwlI7wcI/5Es5jpw+9FsnoTZMkKaq2Q
piv2F5tXplDxaTBR0hnRZ28wW8VhmeuA9jOyVKRsdOvvg0YdZVeRVeZlBMqHBUsWSVfQqAgdWCdZ
RZqef5q0Tw7PK59QU4BOXoUlIMlqCotMjZFZ26Tzu/bEWFUarEmRi4zymX4xNf6b/HojFtSMA7zn
+56ZFYYJd1yutn97P+QPS1BbDsqZa3f46QaWC7fIj8DcABRnwiWd/lxLpScJqUiYiAn5nhvLAqXf
oxJ10SUhvAg4HttygKy2ITRbje9KV8cJqVLVOxphCgmf03RQzOqseUMG6Dehpq+IkkNGTdnT3D3P
i7ASpZIuM27W9rcpnJ7PJqjA9XPszHes+la6Gvv2z9MMx3n52Ll+FksUH1ZD89Wi1wDsPxIA8izS
iS6Z1O7R9ncTsHkneWcyPJl2Hdv1xwf+k5HD+cusFzXTUNXaNyzrA+RAgg/gz86vFmtaNtw9gegx
et9WfhZdg66JBVX3KNDE861K6m4Yv0/fPIKR5pKYe2t/RXvt46Q8lHcaUhUdAwVfGC60+ro7Uizc
98lTPbWM89hWoArGC13WgISQND01a+ZvSqaHSTH/NMlDsE5kzCfkPaG5l8NoiQLbZEyO+geLJIfc
5mcW8v5OQmmub8B+ci6lt2OWdY90p53IccsHQmauOLj1+3+w9pKNLoJjuq5MgGwyfYHuiD8nOIe4
kGRQltDHTwkzVwSB1mV4KUgNfMh0Nqc8VNRGStAYWaJfc2RQCujmVO2LEPc7c4yQWzR/6Cm494w2
/T647y3jLFxR/ce0yepK5ZH3q77GzGoB4hyrC7dAQf3eChxzwJEuhHgfsOtXPlETCE+JVdYuWTur
go0iSRhsFwHmlWp3rFecFH7B6xbn9czXBljMmhgn+36+w85qeRNTUoBlrm+vLpkr29pg3IxcBZYX
W1fIJb4iKdWuBD5Fy3xZ/fWiorYKRoCMWaD3DeNjAi3FrOrKtAsMjA84i1sgsey347BPcbMIZQGW
+Mec4Wvfrwp6ZYPOutzyh7WK8kP82bgouU2nJcswg+5ra4gARZ7k1Q1HhlcxOcCZ1Ijay9lWxB85
WftD83MIi3cWH7esBW5a2VWuG2sv+EBUuxN1fMiNVcwBd7YxyN6RIkPH4hKfRpPcWZVXJtPDHdzy
BsBQFEpYzxETH2vHXb9M8cZ/6q4FJqGOkFxiR6sPeQGxLOq7LFkqCTa2I5ZPeHxIraoT59psXqMf
Ywg5UGT71Rxa71kPbp3OMR2DUR8UDEwpyxHSMTmKk/ccRLA1B8PIaOAFWeIYty8o2AI4/oheeK0O
Te3UqJo6EsEt9wQtzyeuHCuD/fm6rXsTlWcgyJhcji1lvXN7Uhpndwhj2xvr5DB2Q2hlUkoFMVX/
H3uloPqbzXGIGZyVylJXH59kVlWJdC2ApZp4f4r+TSkCY9YREif+F+u+8lXT9H4S1iaoXOyIREtk
DJiF1Nprh7r0gFSNhQL3ixXCAs5RYXpHnhNnXYsnuiH/g5qdNDijGisMArc/7G0OiZhAtoEn+fuk
On7yBKGfkf3M2gOuQy8dR/4ACqiNVAdfDutx7F/jS50WqPsRzwQifwiiq33injvK3+ZTmputKCJ/
gp/gp8I2NvFugar8wDOWgwH8Rzn9gBebMPvIyECscGDF6IzAtwKAygppE0XsizPHWdGJc2sCZAZt
FEtkLrZxe2FCFpVNjlDbKG3E76sMGPCY00NhEegEUwnNMBu99fiD+nRx//Ic4885cGBmS3/KVqAg
VWUkBAZ9PoaMfpMUQU8hKGyGTwZbZbDmTMhl9/4mjK5j16eOmLlut5Vpti1/+tWnPKShlMfriZWR
ZwIWcC5hv8L4A67BZsOiVyF8A9gw1zJhBLFlDYg2LmPS0yuvH3ec0jmsnK7hERhhIg8JUuEGrI+i
Bqwmq/QASZba8w4gocP5uphwz1oCGYDpLhRXz6Gnt3lw2Xo/9akBWXxdLRaStrl0LpC6MYceOKL6
jEZjlesPI0VkO+Q5DAzEONO79DZrIl73YVnYS6CGzuCO1qe5vR3vzDPqdXXBt2zAC/GqBs/GAgdD
nsB4RyeYWeelVkjJ2UZ/OteNN5TlYh+wNqoCKx1JYDGnmCI+gSrWtbEPeL4+3yIym/8FO1LLzM3b
qvh9iGPKLO+sviYylGBWJEboHdOXkLGHvPOOogDg+X2edVt9LAfmYCmh/yo7EiU9edj/aTeRNPtX
sge0gACALvgWwYqdtalSF3w9wvlkyAwB0wwQ8AZiijXGpx4aK5ACGO1PjqA/WPa9YFh6DMsaZwTT
8W2fxkExOb7d5jtkcu7VXl2qVDQI73mpNrBc5CjZzBtHGFDTrUnqOf9TTMrVJpOiCXdCyBA1BqnD
si65ajIzQgOZdrlhHJ7E+rAa4reOXfAAQUDAsNFCRYfDW0kSjfBKTcZL6Jf3LGyrHCj0IFsYxhnD
yNk5HCnI/oi15AZf9dMCXIu/lIQaUi9hxvV1EArCXsXfe5bVzJERRIQc/fv71S+YiRDz/M9bxFaU
DNugPOjsTs1S9BT3pYqSaVLYqk4kGDjsV2bAIl9ISplY9vbRN8nFsvUCtK5e2f9EycTTMDGIv/5e
LTzLHGDu8WKl5GfLgWQYN2BExSwnk9Z2f4xC4draM6mnyC/d5TJwIL+99nmQDgdhFHsrV0fs3NRF
zUVCkgRMj4UWu+/kSWxmLQOwcRrZQ/+b04RZZhszFJf7gJqrv8Ay6qIh0Ns8G3bm6pC/e3ZN+/Gw
3czMJ+u3mk86UIoTTeCqpwzaAc8pDhe4SWC4o14rp+WJfRYY6tXmCFMUcpWqxWGGiePFnNH2fr/j
71sF1f7/kyk0SkYWCxyaJO1b0WU+e1HBHB7RLN3ycnKeNn0+/5/YkKnHRbnNkDGf8m0W4XlN1hJ0
J2MZYk3OJAvv2u3MWhSPl+6Ig79hU8yOi4i+81cHRiHniwOzCMb2b/RtP+Sl/wWl6M1Psl7/b3fQ
WiCalf8MFARJJ11q2pMm2f5mZocbpAWksKhDeL7O0pljizUk7yj5Pe47ppsDTyj3yqc7kVo6hGgC
eQ9nX+w1JP1Dy2TJ/cy+zKSxKe9REYObLxyzZAfYYZkNvTqDfliOQYzEJgs9gxB3pgLYbeHFe6F3
tLq82Ybk0LkWP7aHJHAxpSZ2jLZ2O766+ocNTnfd+2cA5p6GOzXDihiAcjrzNYvtpwjgd0I+t9Gn
BXgKa9HjDdnA3vu5+tDNqyHjmtSB6ve7+WPD+geWAr1oqcsCbTwpwaJipZ9uZ5eJp+V3uZ/Fd8Yz
oYEJuvtHhkpFT96kdXEaEfoehXdGZmgQ+DXCu47CTXcpzouYElJ8zD4OGyee5EBbnTnqDJMuqYgL
Yg7y6jXNBl7YNc8L5qGd0QNBmdBi6GsL+Rr98Qt7h5DhFZk70hdNxUPihQ/+hEkSRp4C0rfopyXS
eEuRdEbg9upGkAqu5/mNeKSPVkdC2maVZBD4tGtQvotNu2w4TeD8qJiMPiYtzINmkBKFIwD/mDnJ
quVKoPMeULzFmpfV3E6YXdSB3arUFrYbGaO6j9F7ss1gxZhVGFHufSZeNU+mqpRpSWxnIB8gzz8u
2m0Rn39PWGJdJ9Jvvfx98djptPW2BBW25RoC4oZDDOBZSIJUMkqBRJI+1ZTLlyav/vPUv0srvDgm
37KcEubeyigrVDh+lrgGHVwI7krBrv+KHwsmSIq+WCjsUV82AO994MaRHrpT7WWchh0iJudX4C14
p0VJWPj/Btc3qrlyOWN7Ob16cq2Hhacz5mND35NuoULhcwqYlOEwAKUYzqVm8MoStRdinfiZm+B8
IYFRhbruPpLyJnTX+fu5Az1ZSqOQ51CW1OjsR8fCIN4G/Btv4zlqlA+vjGMwAQypKQ+TBxQPIUm9
abIxXXykvpGziSMTN34bA9a60ocvcFemWUINSk9cY/hRuWFFQG1NC/8CJBFk/hsKl8pQsj4hUYUC
e+L0HKsiy77oVPhdwDbqGewaKpPNsWC/1ekaN0dULoM08arr9tqQHljNlvBLbqNgp90PTRWKI3iH
SRJbiqwbajQPwMZ2xltjtkFbk3YX5trm9cW06bsZvf+NnrsQ99ra9L/mEFEsOUssHDR6G2LoNAmU
lsMIV9TyL4JLnmR4VMG97AYibEWlPpQTcYJwjHTM+WJ00h1AAG/YQ5rI6+9jIvnQ6jjrSbH+5B+j
mN/pYffHaIf0Hz/P56gcxccE6lr9CtUByQt6V9ebvOZuOzdug01tQ+76Vz+o9wNTEZw0tYSH4DUr
VsXtsLhDYDOlDDnaAG23uWXLnXF99r0sJqo3HYyUIeClD1vAJGB1uFOWO3rw8sGzZXMiPEQ5zv2B
XR+DDS5zXCHWYkqW2qpFQYBJuzJ1e09s1RTIAxyIy41+H9o3dDHHBPdPrJflS5Ddk/Ai7w1BmK13
7KaFZCrdjZo5q0rnZ5WujvjK2H3RVJIJLmQHpdUw0lb26oqXmUdXWYpvNJOoxaz1ee2c1ThKmWyx
hj0R7o4OluvkFVtLi+anRgOmXH+fbVu2/ktfLy/oDyRJZaGkLQcmoyE8XCuxM6btD+zNG6cagEhJ
RWDg0D9WkYgg46MLbhJa2gYl8ZS/kuZIGDQvCGZ12HGLVsUZBobSuxx69Neqhy0TVqjq1clqb9OF
6P+QZG6kRPYaYUOpf8nqge8BZA/FqLQNpNE8YbEDsFHS5vctcmAHQHkmt3/AkKg6DqVaecPaIw26
DUthhzgG8b8g021HOXzS4OawVFIUo8K8VyYxSpBPUVb2t0OlytrhPYBGf//bgnfvdYcCKTpQ6cLv
c8EFodK7zwMyDTBP+XJi2+k1JkbUd65yg7H+WAWdwTFCVUFtLXcpx01J9Qy2AfoK4E8p96Z7pAeL
kf+1rj4e67pYQqYXqv/Q6jnKnHFHr5qVfHAJcK7ziw6JgJ+A6F61F++FdvQuwcEgz5Y5NJy6GWp/
fkQwgeGy0snUs0HBglt162d0wmajM8nLFVCysMBKUcNvQowiWonPlk+Ugel670/wI49Y4KYApryK
gu7hzFqfATmDnBNsEohp/ilkFUpSbMUktZ5f+RzvV4b38txII6yLU74B6FgTuFh0vKTc2xS8ngIK
hQIxBerUfwFBQKDbCVSdP62o9OCZNJgrpfltuEaUxibq5loZBZSxuK2+kQSN8lb+eEjpX0PxeQRb
2uXV0wZ5XjIm1CzKll3lvNZj35lcOcmLo7sCG/YdY8WGXk8ar8UpkelPsUDQETzq7G0PPo2F1Hji
U+/N0+jzr5TRXxhb5HgjErK+CBlorWqfRNH/UoJzmU+ggchZ1JPQBbH5l3Wi8btqeKkD3xntMjxj
1sgVXqTmpCD2mpVmEyvIMwszOyuffxp7s2fb8FXB/og/d9njRTJ3CoDreyw+7UAiPUo3KqJn1ig+
1gdpnULHAkHietVRpWjFkCgFlSGh2M/0wtAcRPpbuhynOzouGYJCh5acJXTlFD3ljYUfwySKQwBq
l0h9QtuSi2FTvy10y9D3N8ZJxzpm1q3p2Agmp06JoL+U0DxxhdmiGxHLDThjruMEr7Tb4QVIEqOS
wWfnmlFu5t80jJU/wJK91j3wnLInqy0xRDBA9km5LykVcF6lyPlulh0Ose5tGET2Ed7wCxeHgPy8
sBaPZBnBaDsrk5D++nFftnY6zhD4j+duYBS13aCkkDa+67nNH9LYWVV0oX/tV+qXPhO7yoy9/tvG
Z9fkYkMkFUnq+jnBLVX6eHSnTSpVrjTgtgMVZIIriC5/SBXklcv3aHCXBD4qMFqXoEznBo+KWMUq
oUc7pDBD5p9+6/jWqfDRX8tXf/h7caSpBdKT4iIFgy0yEqJhamvVfzN0GqFMP2lJdhx0DQm3p6CW
RGN4N83aD0cMPob4j0/gCyKQFgeHEoy80tIzoWJvjQQsBeQEK7FPQO+Qrx4BTw7DZQNg0/44MRJl
eMgRmX0iPhVmHI4aelwcopfWodO89ssR2nSLBL60a+GzH1d/kapjedBs+k9dMI4ICJuxB1kESAi6
Nn6FWoLpRLJmOIM5qLNEVfrQpqzTajFCIWdvNWnTeIBFUJKZkgdh9famAQcl6RzcIktsdcqO+9HS
221RTwx8aRfanPa2Z+1+GEkPsjns1X7JEtAlZIlgT75Klc01p3PNXKvRSVGTYaK/Q/MRXaYQ4hZA
l33my6HK1ejfZXDQXIUd95MH1TVEH/y1704zwYB/E6xmbyWyf7Gcmu/SgwHvDQC0UF3t1DRt4HHs
2H/+LxYAfH2QXDKDPb3WwaeVPOFFZzeZ//ZaIn6TqPORdiJ8a7Kit6wkWNMf4qf2PWlUnAjecE0o
UpZUmuHUMXklAzIedUFf66Hy2mGkNU5yDwVgxBO6GBI5AJu9dqHPBKhSxn3Gekt2iaOACHDPnqeN
3TEgQINlPJWTwW4x34oMl3OKY9ByIikhOHpoxBNtXhS6Gj2EuOfdD04tcMFSaGhVC8p6rZUP2cJl
cEElg3PikgTxHOHDqaD57fXpaNH/fnzkclGAysrNE17U3YEhzjz6oRaRFLyAPeA4LNtr5wkRFXqz
KmJPs/HsyqoJ/NTXfGaXw9xPxpFpd0+V4KJriFUiUpbfalisOT/RB4S+pTsURaG5vnCWouk/SiHl
Fn8RpAmeQ1RgLvCTrIsUhDft5+948k9PYMztTm+zDHz9kZxdy88d+0weY5UB5LQkIsVgmxjQPIFs
QVPCGcBq2c7RVKPx0OSKMLuAJ7v/T9gWlCrOgttTclI/zUN0eTwCJaoOhiAS/tgccnH2K+4RS+Wb
8vSLcYqBgmwt7fuojCH6GxGTGSheyJkvtItPtzYbXlF7vzYkzB5toZfwYWMjkkeUTy9Ej6XY5Dm2
ABRIDXe+F6WPA5h1aTUfQ1INiJp1NsRsy+ByYYKL6vAQjE18rZBhGv+/BgS1SmugZub9oEgef/Qh
kD3VBZW0fJogI033OlD8+KZM0ouq9idKkveyVkQH2gxNor6GmRtrptREtefKyXi5jttHSWnIpDQ0
XpCKbunYQkBffRTAt56hs3FG9rbcZ5LNXSQKtUF35amVdWnkPl78FV1ntwbSFdGgwbhizlxxNBqz
zBHlpsaGvMLJkh/BEq7BWSHbU1rbkvwzdNF/G6C66lxkf+aBUxLb6Vk5Pu4tQ8WO8UrS8ay9pqoH
5TNLdQ7oJn9OIQ93HExqd9g1E5sWIO3iT2BRYiHFTtKRGw7WSYFOmU77YO4g+IW2g29cCMKXKhED
PdD1p/Pd/jGCQ1BDfZH+HjIVJ+SDPbbuuiaLp4e4R0Nz/nvrr3o7FQOJ458zV+Ubj2JFPJLoN4qZ
1fQiQKph3tq4T4qM0qNo7spboxkEj/iYuDsQLzfeO1qbsCVdoVPRmiVSjBNv5P1VZwcmXkh+AJgY
QQTz4GsT3fheFMcpRSs4Jls5f2h1YhnnNW+Va//pINGYGn67mla9eIRSBX1AmdPuOEncvrk6QAzh
vzcBrDZDCo3ONwgdnMHaUjN5eOoBFTwZonAJ5cdMN3fQpi5ys6rIW90xmSyDF9HXnUWvu4mpUaYQ
egUGg+UEMAC3od6/7uhVhi3fO/dLygl1ypHDMuc6I4lgM/IWzhoCOObl+y1qd+VLiMxWrR+pBX5+
XsKe/6KplJ7TpMqT4ipBaVPbsSSB1eAH1hLkHAIJqbi1RLJBRuNwY6YOPQjI9YPyRyT9pBK0s9yJ
ic46V1Iv1w/SFBhVasIDZFzu9dXHG3oIeQxttJNGc2z+GM1XS4a8opOlvbOqYj43QqQU1g2MGRY8
Jpx56m4nKeXl+5zlhdH24Ge9rZUu3kbOj8U8RzCniG8iGKOoXwrzHXtTaqkNsyff2hulCA22e5hr
QieJIE9u8FLZnZ5qTfT+Amxx6ssm/JP3EdjR3dje5b4WKUYFklRv8iUsWiMq95hM6rV6YXGSZnGd
7VMJXQvaqLTDNR4oBzrMcHuL/PKF5vlcOOCkYlLwxV4M9i2BjZgQVj6HIEv5peOP7cDkO/ThySTn
yyRcbxNagfiG6/zpVb1drSwJrwC1MiODrY2chTBrfoFZytoIStpN1Q8oHGafC3fYXzGzvNpNDuBf
83bCpfJQEaCu2Jije/hIHzypzLuLjRJGQcL0+OuHDP6oLibpWE5aFwr3pkzA1f8VE6rncWVJJMeg
t9vfCQqgiVvjvjUczSNSJSnBLOUJ35w+6I6eTiSV8kZ3fAfD84uTG8MvQN1zaAeZU5hjXD25+/Cg
Nb7cy+cj9mzFPFYAKhA4R/ZoY20AacjtLR+61ZWnnO0AXf8y9WNVx2Nfdkhyo+D0DOjqXhUYzZaa
ApTBHMgAP7rFSQ+HxpYmTZKMWhPF5UhgNBa7AcTZcuEk15H3VYs9NmrzJQ/yCcPYNJp0x57xeDhH
BaWEw7FKw/V75O0om7IqJEFVobXV4T3s1WpgnhZE684d0GyY1nMEWGRtbT0rR2+Y4y7f189JCN4I
uQ5MNZlFGC5QVYfMKhU6tEDM2NvzYiJ8za0cbRED2WIDxuU8nrmGXNwSHIQy23/g84NnPhHP9CQb
hOWCdG4/nHTgmlt6vdhOyF93txVUUH5E+1QkSvSDeKWLH2SJt0lw+e2x20FXxMzbSOPjizOVGCGh
KlnJDjNyol1RQkmw/MFPq5xFjeVTRxhk8DRGc1KxaeMPDIlgxKdog8Gq0rIGBzkB8U6zirQv6US4
V9xnpaXZ3amQiSJPXnK2OWwueJ8s+5StodmtjPNGeVhh0oCbsURlg3qus6vb7qdtP73ZGDTcG7oG
c5Tw0u6u29NVsY45KDVjpoJHlDJ9Gi1Fk+82joY6ZaP5HpjVyFDHfRD0fiPLePaZkhVjts88dlbW
lD7J8xJMZ1JbFByrDtu5jJ8gOEc+7Tr+2ruhqXi8NU8OtgDslQvXLV7UcLZWqgjQbzkTq2OpD+Su
iP+ArFgQFxyQNt37QFGYin1R9cN4ZvpQKBVbN/Vfc/6VRRDpHPwTNgUC641BFiTU8/gXjxEaKXir
Rw7frgGlzYyqHB34u7l6zc9CzFXXT2uC8PhHza0gDY9eY18vquyoXVeJUnBWAOIlsuweJlqRLqzJ
idpbK9CqJxLX/V0XhZybGJ6WbBOsGqIcvMEaOP0zuEBpxyvl5OAKmkZv3fyphu2oIuwhqatjYVbI
nAN9GyRg8yrua610W4oRYMmxaZImaoOjc7cUXFcTaU0MiiMP3U5YivxeR7gwWFPGB5vR5t5n1Xu6
/IxjrOvofPvULglJ9rJtVqPbMNRgyych1n68gnoFw9G7H4pl5rQlXxzd8xtTcEP3DG1rE+/6nBR+
C2HWx3nRNK5ERb+cIKNO/80kTAUzmcSLzIWLBMmVUBoRS31fEeStHG0o0sv9C/EBz5iZJmlh/eUM
SeHyXqDqaoQaq+HEjCvF5OJCXRFafU0WlbQYg5wC7BOuDZ0Las+IPqzLKnOsa+vKIk2mRQDF95xu
YKj9SfwH/WHyuBRAZBqMO1Kx5nzFPZ5MlTB1itafbXbA5ddKOb/nmtT2aXlMOoX5zWeozZolbRVs
r1yjgGp28NT9sQRZuNwzzAYenVMnrmdRKvk4uMln2fF/JaBxhpXKjBijAR52In/uf4ZLcXrXMdjP
KKeMcWwUZ1Whoq4h8BF616DEMhWm/KbQczij5OjxAhvij12KW1pCxqvx5QFN7YGxzAjJMhKtuLoi
QSfoIGy1ovHQe8pPs4ugYIgq6lN1D5ZwAk3fXkyyfIWOyE2djNs5KwgM/KNqG8kzYsGQtw43RtZ3
ccC0vmy6x2CDuLq5zM6xXjcbnsvkHNKuMm5hSym0f30gntm30/d9l75rlpawkN0b7/meSIzi0y3w
schxQKGVyVO5JLkh0xGTH/iyVM8i9iz+4d0cN5qVZkvx8q2TQZ6Lk/nf/YYCw07egzhqlc5zPOjz
TfOisx0t1g7i1MDKJ08n3qimQJgPbsIXhBESwpMEDSwrKnzjbzdLntvmluiOIWaIU+Mx/X8+ST4d
91zfSc2k4neYYRGtzEHQHalld9Y7/tuYBG4/2If8uFB2ZwX8Rovl1vay3BWUYJ+bZxQ6UhYWD2+C
WYVSp8bcffaoRzlxK6oCwSlFh0pQ5eodhsrsLlthxM/Hht6hgmuiiPwRKXetk8l274VSa6/aKBkZ
/n7SW4LInN037fS5p2pgrPG/s/qvjMQZ4H+zqp0qEgy3roXbiU7T7/vJkagKrFVaPsQcKpx9V3co
fOun+BHNKm922MBOG+GB9YJ2Y8XAk6HJFx1ewKf2NnK3doD+Uq64hm+Ml3BwlFSGpuOtXQV8q0H/
1qZTkIfFJC/wRHDNsapt+Ilpw3DGnLAzZV9LUQFFH/d94ZHKGLEOZ49KYXgJSPQS//ZSGczu6G8f
ByrrBD2NgdUyK6fLo5REZjz9JCRQv2HVTwivNm0VF6c8lCJ0gQiUqocsrCHKm+awOTZhQntBkHxV
hyyWEhyFX74YF8h1Cdt+gNZf4/7/DzZ4FGsrxIJcfzNeC7VVk5RzyIsLHVWcwmuW9AgMHgLqlzwh
AmQzcvPFMWO/PHErNGohJAojR6teSiFrr7GEnaFGonp4nxMQBjUqOFNppGII87iNL+1+ivwlgL8k
gm0KHtvx1yLOD5cv1+/6d0w31ZttZYksJccO5AscPw1xax1nocq79AxtKeNfzLNb6eRJ+jiP8Qet
KgVupzr2ExtS+GZz4WaK2lW5VQJ9srLxcz3ybvW+40XUXpfXQS8wrZDOuypuejxOtzYN7EqUVMWp
ot6P7jV2wgS0Xd5B2ugR5SsbE0Azg8pHyDF7Lyd+KCp2W1UUFqhKQyusNX8UrbWxatnb1YvOnnha
diODLmAiUKLwKaGVqHpx7XnYWPIK7Y0RLIvlybOsC8IcZLUorgInM36O6aIvNOrZwadi0iLO+47r
kYnXomvwXLh87KVHdoR0TVD5a4Bj9Z5wIAxSbop1Gq+y7J3pawHc4TocmAE2NXpNTngoqw0RQmca
vEiK81nvCZWCyEzg2WhsUCDi8NxX8cdcMlL4xyg4gbYviF4uCNGrAWZu9cNHsTkZwWfCrtIuuBC7
BRvImaM6XnRm447oBiJxJBcdQZDSv3Ib2+rf6gEamJd3POJNgBp3OOIZTdljLPvoct4AlcoP15UZ
Ge0MOCBUhTCtL2Uep4aT/LRZZ2DKhdbU/felOUgEawoin26JEyCIS72MoUqxv/dZ/vTu4NgmfuQC
Gstf4JTKFClF553DmX6wDNC3uxjo3nuOX5lSBhfIt5k4N+//LDE9xIjOJRGVYfiilPbUcwt+18FO
k3DHgnBdVvsmEPCn4fX8f+edV+DigwEscWmelSxN6dde65CXjVT4uVy0swKkU3YIZn8pjjhFLzRg
YRDvXARYs9g7ZE+WcpMCTr5h9Sj0FtIs3BUnz+is8fnYh8qF6h7oQLz2V/135L81ajaGdtu+xQoV
kykD3MerkSImbIkZaTzRL/PR507oO6ZZxrt/ka0ak/0X3PgQSrDWINxU4RBfWSQyXKXmHWFm5Kdi
g15yyOFsOajUU4jj1XJcZXNZ+BwfafVU40b6wgkMLndtb4ocupbhBdYgagWDJeNifHEC8FoAhaRK
NhsvspbZdGOArvDNmSZ+RMlSUad52+LRysXkR8uYwMZz8pj6EElUnc4HPV0b6mRb72fu0PBXETSw
E46lA163iOunmCA0q6kSF9SACLw3g+EKxroC2RgPG2HbkB3vgIF3g5GxD0u5WvHpV9StZZjsC+h8
i3anhtlbxaKPORHgfFFGl+ul3+f3wXey68JxT185s1/nJo87MXkILNbKtSYsBwLaq0Y1D7qQZVvh
HwhkuceYdVQVsf+rjKgoGz1aQk4nNCHAiYtAvMGcuio9IIpOrYj9rSLoQNKLt75UnVvduBR6R/o5
gZiQQy2JG7e67JZzcnoETl2Ed+DO/wFPI983H0nSgnVRxq2HirWKsaZVABQUuT8vrGUAqqavvOPd
6AvlunEDKhO0VedHxLXFa7yk5kpprN7KOr8LMUUnKKpVp0NG0x1CxKpEwoieCTgt9S0c7xbQQd9J
UkfE/QL18beZTXLrxtYZY8WZjLuGOHmZvLyUcOOjvtUtaIb4gZ6GgergmoSMSh1qPJDlX6B5g/sO
t/ADtu09ADrp60h28AzzykyokWRgb7+2wXSOzSxx6RXIGRn1Fx8/3a6Ijfz58hfUMDFCntu8cxZ5
S3IfTm40gWTBRibIgLs19tCJTutPemkbloDj7qoW1JFlhgKVJMccXIIJNWOPelWO9obW0W9ja23S
oJMp8lKqV6iMR/eYpx62cvQOhxFjjgFD27od4Xa/piFhFdFv0c8ik4klXuWAOYeSXPMWwpWgUiXC
UqRoLzmOCT48pZzt+BhxSGuNlI8Lxz5y/O7KhPf8D7H3VXPurMks4yVqdNrrZGomejwij7y4GhjF
3jE4Iy+ZYWY6w9GF515AvyRKrUkV1sQfz1YExUfyx5IKo5Szri5dIHxbg/yc7GV0yWBFq2Yu1ngD
Sj9Y1AoVgrsskGYH1qnhqD858oQQyxXWso5jCHdKK+57nQj/orAZusR86LNziaTai7IJAZAA+DvQ
vTlIUYSTA/MaPuWGN7soQljRj3Ytdb+8v4L26K3gT31xPquU+KHhPSkewZQSUUBCUuHLHNbG2p8h
bbzr/l7seDHEWwav9C8oYuFCNnELMkXBDz+XTDpWFW0KPm56jEe9/GxD8OVOMbo5V/xJSVgfkqUG
Iq3EFI3JDu+/rZ4uzvY3uY0qldyok6OguH1tskf41SnIV0iQRvE4vZp3ffpuBm0K+HJPCE6NiU3h
hV/99bd73WplfPxY6AquRWRIaDWQ+lgYRZdx85uIWhiQ0/MXeyxogxcNf4o5RKiOhgD++Qm65Sf/
XLj1hNeOGTXqLdOJ9Of1MggRDO+QVwU5EZ894VtyqBlv0/NWWtT6+ZCQJaHZmg6yi3crSlwkT7kq
R65z3cl1i08YMbHgNXTXatlypanh9G70y/CVKLyqhzu1klC+cyE1runlFxjoW0WYQmj34luotAD0
us83abXDCO8hZ7DY3qmYgHgwKz5T5GXbrQPBKLKVOosXWYs2dug+6qabFAuF3rdT0g96X9OP4YD5
9+Q585Gwn+WVU7xtnD00Yph6vRcJZTgCnzxL3WKWyGHwpnKFXfdtzFfk4HBzzBuaCMOMur14C3tN
GcyIIx6Kri0MNsHiuQOh7/S5PRhfa48Phm4iL5lBsQkTbqkNmSuYVbYL0lz2gdOUiIWmc41KzG+9
gpseMLbKgoFrTyhnxoRgx5fCX6u1HK+l94XrS6USm0eRNLsJMdcEHga5SxbRZppxwgprQBsIhp4w
+t1+z5SpBOt19zBIdmrASczyftCUkRtAZ/eEOpi3/AUGoYfytwQNgEWlHCafGrDg6mgqXNA7nks8
oiLiMlibjVKvkTluzOdJoqNy81Uld/hm2LF7F9j/yguKwXa9+uXr5ylQvoemOlvlPuwPNwBpXgxZ
S6gG5jWvdzWMfTe076OYg5PkcTtuZIIfceJrzlpPRHvWRAaL8911k5H041eU1ubJg2ZHLYRKs20X
ikKTpEuyZBi4jdcXMi5wefSScoyoff1dHybNNPT1Nrdg3KzpAYzayBx1Gy220gfWMSbh3ojNREhc
vRwykAJJEAeQq4aWqTZh50CTPWdEDg+dnJch1E4NXDOhxtqvCaR8w3YP8mzO8Z3Iio9jTHNZdW+v
h14QpUz+Dqw7iezwJUL7IqpJeiWScZYDudegdPD5qWTtWMNHIstF/2uW1SmeJMIS0OmdzS8DanCV
AsUmHak9gLGXifZIRD1v/e/iK3Fl86GXxHt2VWF9IzUEYVecUcATY6DxEgjqMB8FiF0cPAqUc0zZ
WtEeq55TmQCeS+LOnS0sXf/HoL1Sru4yaJqDvfXFWfv58+oHP8y31Hq0DUCfQ4hqYfcko2MOwjBW
wNe1mFwSIS6yar+vNpEpHjIRQVSSvsLzbWuOBPObZ3aYJ0OizKpGvyR2LG/lIW2e1TRc6C058G4c
sCmi9w1Va2Gmj690QYr6rOd156dl91rGCh1tqsI11Zghb55WqkTuzpuQFV6y/pzJUzSyiqblrYMt
1VjExiKrxOFEJc9mBJL5VRkN9eIqelTtcmhY+TQoJFpFAUqNHWi7nIel74/CzVm0ZllacxItbc7V
rhGB32z65MxCL23AicayL2/9jQ7ftnyZQLCfe0DYVMDjAS2BaD8ElesfTaeN2d60IwZXN4iRLBOt
z0zsamVsyG9jSkDQEgDvZOGg5Oke9oyRyWM7b3Rn5TbKmwiYNkPB9mrHBF88MolLAVbRfIOeFKqs
rZo5ePn7wKjBsG6Y85eaunu/XThj618+PPq9EErRGEfoRNvR+Vlbn+5GHAPYdPS1rJmYV+y2awd4
Vdbh+X22WHj9Y0n+yPvQYUWHjLtP0VZWgooIe7dPDsOZ/mkVYp122Dtx4kuaMAqy+Qgy218EjF8m
OZrhjn0NwCGb5VlNxItLfIVSgABI4T2BAhBnAN6JJFwX/6ZWy2s42ziNaJg2jg9+Apwuec8FKwj1
O5IIMk5C5d0cK0OPA71fBEWlFGSmCj1fbV+KavUdmCakUD6c/PDKzsf19m/Y2H5pnAgv0dxx+yEG
BU9/OjqT3zeKd4G6XI81YwtBvNw/egw487Ew2s03eFepB7HKJemCjNsxXEFmR/U5qrb27TiMlPwh
WSIJQHAdP9S6AZIpbKzoSzZg2qvSwxjU92DT1q8ZS6sDA1qxOvcYVjltQFpISWjdDcVSGD33BkZK
rB57HDQq2i4+wYMredq8+dWfsULE/fS39sDKsmd28vYEDVP1eKpSTkQcHW3kjW33V8GGQAXle/XM
LgdtdKHXO62EbR5+wusSkKPAzXp8hif0LfJmF/XyhGhuQRhGrRA4i26786NQX51/6r/AyosV0xBT
crTdJg77Mgwix5ZVSqdxI7i0Sqai0MLUkvv6iTSoarfc9DZJQytei9m0M5DO9BNyrqJOKgqLuXgx
qbSRj6sEDY9fw/Cry5pME9CIwDqHyqWHUeL+BSaRpSsO8yGIVpnZZNXQhSsElEbtZCqTxBSpgV0I
FxVDpGDiSIZefCVDusVYKOKT0I3DCX9YjNymRJKaGOftkHjGztOTLaIk/7N6KffY//5AGMiEcPkG
A6tZvXjBNNkomi3vXiqUVQEoGJqJ1qiYU4qe0ues8l1/H80U7/VHAdR6UbUIwmHwbdSAilQu+p7R
Mk4eIsv4wqI0GtDvcUfx9KsjTU1966nu4QkPdvVXYNKes1+hZ/L4tjPu9Bpj8IZrzn9p+heHv+m6
JVNkfsO7g7OPmANt1lR1xg1Mz9TKe0pf2ZVI/awvIjffC0v9h1PWnAQzs46R372TWOGAwfjReZrs
pWQv1MFJYOTs4cGdl4RENAGR0qU4NgIXTJJpj9yNKOsdvIt8LRonpMfR1RKIfvw9tXPtASpLdgyC
Ea7+CjVcEyAPik9nIzSQT2tiu6rTVu5ET5LnmS1l20TG7Rx2BJR9hFxKRLQtEZzfDHmCznt2qO1f
i3uzHSfi53DrFwI9tMo4bnR/44VEOghMwE8J7LomJUZMoYEelTJ0q/icXdowz1b4gZrHjPHZO7Dq
AKMGA3Dz000J5bgbz6qZRHsOgPEQI/eJEnYR7rlORkWK5ROdFEHM46FfFaubLtH2q/Hsu22IyQxn
KvP8UIFCkmp+jwJ2B5JThlY9o6pZIboBy2Y6OL9vE2GJX/hTjN2aaqX3gOoEIwh3sS/3JK5iuj3d
+6wqWmN2RoL80Z+fo4lxoSQuRr6NXjj4SGxdf5Ml43123h44nKIZYUbpg++EwGN4ZzK4b/voME5C
bA403HWBUcp6wNg/QRjBtkCS8UNh4QnsCYAi6xrTyqmiaeUbwVDFSjJRz7Nb70fch/KEIQO2YTrk
rqZ9hyiTX++MnlqAGJU0FXBmCMFQExy5PITnp7TDX3J2rDTyTcArf0WQFhKSMCWMWWtHggVIArKJ
T6DPlbPaYsC91kViyUCZsUMfZbhuB+6H03s+SLzbjh6E78o6jzqHSnFljeC3wBf8N55vagjVf6IT
0AfMwupOMr7d5o02+xxNFw2KdJG2v6j+CiwN90jKBq4Mi7Op00VYPGGgHV5HNFb6EY6zp2BEAoWX
pCICjLCnADSbQH5sGNxHQD32eIDP8pYM1cI+RvU/1reSIZGKR82OWlX1ohuRjJP4hFTB7HJt0NBV
rI31k0PGKbAmM4sHEC2tsbPOtu8jJ/GCnxNi7z21ZpcJYTRjkGuxL9Y2WgCnj2aky5ZAWgyzgsWd
9obLJxaO3QnTeFh2R0OU0fev7d2gIVuk6qLjOgxoD+BgfC43v0kCFR0i+UYlvCgsYD4ILOwRVS8k
K16LVyMFbw7FDcrSiK6vQVCIOQgtJZDVRo/rH/erQA1WbV3xVztUVb4GujJW8qK5tM+xTBY8OwOm
vbzNluC8j8Mi4oQ80qANsmVjU2htFRgLU5v2PkDgFf/naA4FPdhMssRsle67mCzRDeiwVYVVoS6V
DL8UgUMvDVQBcXCTPL7Sq9wGZw9Onl3ZZl+jZOu9D6IewpriDpKRCX5UF1TgJTxfJHYPyoqB5vSV
/8OJSZeVZMOoVjgXKT0R/rNKS6kjg0+VC+4qjMc/6p+6xJcDQ/lh35L9wspUAV12itepE8qcoJfW
z6KnTlXPwbhz9uITVVKHoQmfsjMOMhOU8HKgxZhKekL8ld+9CQdSQt3U8ORy4GOiv5oyKk67RHzS
DUaiU6psP+K3AG71l3QesBlkiFoorw6n91o6WzcfW9pb+SLkECOY4qB0vWZRXTvB6WfkA768K4ht
iNQkld2405Q4ak7s8moowVdl+jXc/1ykHjVFQwRLeQ7AygCb3rymlhSED3R99Y5SGGVRaeoG4N1n
ZSCgvUJTUSaQQSpiLS+B8qSgyQuOMbQGTcZe1bO6a0nP8IKjy+g20CdH1Vhu8VMKcGjcdiPxFu7Y
8lr+ju0rDN8Z8mbsyuPN+UHgsgIvInxVB96rATVZEeLtVNvLqV/EJ/4WwT1TvwyGwW3V5nP7+MLD
lMNx7gUxQ/0C5cmjC1G2wHBBEB6r0Pi2g8m9M8R220axZqvNmDcp9O9klzGY9kn9aZAc0sTNQDkX
Z2i1GepitFBxE6rSkHlfBnTGNhuz01wofZaHGiifr9OM3rf7jvUfqQsxnarDna0ILVy7KfcN9fBf
zklcxGBe/9NS5PxyHXuA8Pl8xp+A2T1ozng6sA+OKWs/9mt5VmTl5muPgN6jHdqIre/PioXAU172
pqWZBXE/16hRxVTXcgfy6FOXZhZmTR92tm07z3t3uTHRePvWcMkV8wETV4LgDeUhThfBKwZhW60Y
YH3d53PBR4EPHK5t2ky+AoNJwTxk+vOLeCVxoHdYhehLUSaPb17HKInwAUWHnuTH10Do52Br9Ugf
8AlULVwWsb8rAtvPSY6wZvn9ohDpiWSdZZwBOtji67BgJts7twWXOGYWqqcqgtfb+YcMW1V5/4S0
zEZ4U/FGKeckP957oXckACQg44EkFyTplEdsUBJfebQP+XgKFAu1WWiFG9xsIAtIV7BS0rIRLhUh
0HabA5eOJJbP/nE4SNe6+XkZkgpnqD5J5ZzWwKWyGfvofv01JoXW+IbrGm5tTO7TADVdc+wriwgL
YIgKQY8BTsr01grj0tQD8UiTKW2u6vBo/OQ/9Q3eobmS35cEi3nevIFjOgDOa040gmD4yWLk7E79
jL4egczutSvMpL57W/Mim9P2kEuF0h7/KApxnwuCQr8ZLAEgbmlJQUVLTSgmfNDFfW1QYf6znEvG
8BmIJPRsPoibsOx+45WAtpiA4+hfrhAUNC6GEs2iE7A8UOvhqDB9cheFk8QNperdJRoAsTHdy3az
aSoavGH125THLc4cV3hobQBJPEJWTUBnZd4ngn0yAhKIabbirLlSMbrVNe6WRiliJzpHlBdjVtVv
0/kP/BxgUymg6TniCDkdTzzWHnEFtCr0ne4IfNO9pNZjJNNZ28z0RAY2JqoyMyWl1ei4RPqHNw0s
GoYlVGHJ6ll5Y4442KeQIRy3mfM4zn2BHGdzZCM0cefe3CaWiASdxislszQ2+2KVjxyrTNHSDgif
mm3hDxg1Y4jMAaccO8mQlBAj7DNYYAqQtwkg8cvP5lrJyuTxYE7/PFWNN+7sAQmks156DfeMvHAF
TXYuV7AF3Y8pvUFMzIMbb1j+H57Ep34zPr78MzOyN3PuV1ZBOoLa+sa1YkNGFE4gl7DRY6J9K8lS
P1rfIWzenL9Uzhn9tt2KGPUdde9OdHBeWL1sLnDHNHpN0Dm+TFbF375i0s0fs1GSiT7ijRiqS6N9
e/i3MC8+g+ru+JJ7XEghCW0XHP3wgKGFLCacMv7PL1Zg59wUpUXAHZ+iAAHmwUUn0K/2Ll0YnPMH
NXiHHdH+/02stjLc0oPkGfA+UXFQWSUZgoci29xtxvtZHMerWy720Y5k+4S1+aedbJ09RsDOTP6F
Y/9xy5aOQkI4VSr6A4O6QxH6W2zx+bKMQ20NPtO8KP8DXaA7+MPCEQWbOj5VUng2spHTA5HnZCQ3
Ss9gdlBusWLUBTbS/pZn1KQJVPMenlNcSM55VNY5RI2R61k4pGGs4Zc49mTuURJYqvAyrse1uO5c
e8Jc4ab5NtnR3C5w4a57RW8R7gsvVTHbffW4Z6YU24YTWcddm+/MC9FlCfDiBA2Kq2b4hfITY0yw
AzRmdijNsbbvNUFpyDs7PFb+/Mjp4X7+NB+BWN6wTeJ+eIxU8U37NSMoPVXrIRANM5/9vwn7W7Xb
GzY2q8lnAMYO7vL+xZFoBcXmJi9hSvNVS+n101TMFeL99SvBQEA5Lp3jE/dW6fpaeLdwvzFoHuxp
RAofONaXGvuDcpv4RD2HzABP5Y1iqsGHVGwfScwDE/EVgUARVTFOJDPwg52ajJdEU9kMqS3Uy6Zb
2CDlwq6ylLciISkgKh4rCCfYiWuY+/RFbScwsm/sHG5qf1d/e+7cj6hsexq/Wgeb0nhpyX8aQl18
SZbNc/e35p8NriWjubVsEUDmWrlRZi6nMeNtjm88Hkm7CYW2VXUX2vR7Ki94C3QOcAfoAb8nBSXr
8gYjtxfZo6g9yqSCcWot1zc8cf0/DYo+PLT9qZeDR8UkvttrfNDIV/CNkjAlczivZKxmvkS9FGys
cou+mT6/qwnO4/NxAOEuh+8niPrfqBgEqumfhkmV/axGP2JMwsQwFKWq+RPu6rZsXpsSZ8sZMRC+
cpMg6Z2IQixdwD3ksDPAFwrTnSmnZtkeYc67uhx+4paXb1afRKll9rpZw+zQ3mdAWgoLqyqTo4cW
DqjZ8dfJGS8fiKebktQHMdmnP0S2+lO23vjdA9rgZHF6ND06IJaMgBMG3+oNhJn6hdosj+qYzCQp
qrJryUcwUG4OKEGtGM0SNjMcPr1jLC9y/OkMP2nAQiwtXmx9HWIZ0UAoSlki8ceNnRlvjRtEsta0
s7fYOoIQu4f0mQIMA+Htk8stFBxMidywm1WLRLw7wBzZ2ictHcH9j68UJCsMjx8OCeeUpgZmFlKj
85K1AFGsGfi6uwx6KB5PkqMShQLDTVFM+GNuTxah8LafrHWaa8GdjSnn/nMLde2YhrlAZpTjcVc2
vVq0Re0VmEyqLZBW2mt8tsxt9lkP5LQs3LK4h9xqWUd2tKyBv2DHj5ZB9VEVq16HmcQBVmqVTegX
686+5Bj3eJGY89CnBuou0g5DPDSdPjGZjb095xCZQrLR9ggTwlzq9tZgAl9iU5T9hjquxbfXlDEa
/ztS8DNBBSSw3GylSNlCHgis5NjLS2CFlY4hweShO/l9iwTYPSbj2WG++Nv4pNghpy9PeSRWUJ+A
5GkDAX0U3m95mXoSqWlJsccwuhjXaRIVx3RL+2pxh+cpTjF3xDwdmmG7+Q4ULumGbBlCdlj/1QBE
pebR+6XCY8fI/dTu0g7/4mE0m1RxPugrjYaEEM4Uy1Qkf56vmoQXj7D68X/aqEL7uIUxSKhACxIY
rLJ+nobUh6xPoZN99/TAeFgNMzJSNT9MsTdDvQpwN7Gug5FkXHGhBp8Pwxmx/Nps6np607uxKJNU
eGSH3SPK9AlMSUQ9lMGD+oh0EGrjmgcp/nDRWVvg54KDTTMQ4bLyT74N3j5JsTV4o8K6rWQY0Fgv
iK0VJYwMWccwMAJal1CGnjhEvq4NHpxhfOnH+/cgIj8K9MEQmcd3vb4zn8hdrDBqyVZ3XSc9K/5D
a3mhZDNDyEXemx4fSxznWxrdEoAILN/sGr/Wzfll7EDKmBpP3qDeyIhj9Y2N/jph2Df5kSLwz8Mr
fhxDP5jQ74d8L+CuU23qyjXbzZ62h1YreWJhkE1a2R37IjqtO6xoJbbpeCQiRu/cwlh9nnw3eOf9
oyGxbIgvPlxy5mpgr2JU3bgOv8VfG+apEWrK3mpFybVU6vQmjwBWebhpWtCn7waacJqodQ1Q1rFE
PW6bYc9BwKwo9HT35nwHI09Rm+88lqjsEL/fwXyo0m1YFf0aobu85C9pu6tkSpTkOGNjVma63QJ+
JQ5BfQ8fn+Qn6fmTNeu9jUMvLzmaxRv+q1eL2W3qpxGxw36zrcKE0i/s8QvTEBmjEjtOrU7fwofM
m0V2hPT6yX+EdGc/x0duQzMiiFv3K5apIGVTKqaUY4+XQD9r0O6laLmS8mUjho4rEHwVTo9JcRqu
s1H54FrdwonQ1RHNIjuxAPQTKUtlHTL7P0qHYP8q43ibAyPuhqIMHHzf7qMFDNnSjwGNQNQZvvRk
R9P0UuH0OSYbEJ94sVSEQ3f+P2lXW4d3hNxutWjjmXfzWQZJIZbQ9iw0FwFvjrQpkfybgbXu7wvT
GGTyx+hvau17aNOhGwyBIuce0R+l3XUKydZvI//NLQsBnrnEPEwphcXvrilykxn11r4v4mUt5YzB
y/hMtcAO5WDzHea6rKxWDO1HXgNJCAu90Vvw6oEAxcEWKmICS93ftth5ItffqKTmcD5HTEHHLz8y
GIVtC5Bl7P5lDnACuYctakHkmV3A+kS399/VENNZpngzhdzF37FyLMsqoT8YMBuOdfvGMQojt0dK
ITROWIAARF53ksG5xg8s+e+bpQx/JMoW2pGdP78KTDCMyBuNtdw/uth6qUbBTTmRJpLGgnhwDXGj
sSSizLhTIoQiigbA33eotBl0GSYMR6Xr9PqNjqHKOunKKkta2ZlVV4HqWBO9I7Va8jARRC4VKTR7
sIvmcE8nVFQ8Ej9YZQeOUba/9snD54XtemFIqmanmns/e6yx30T6qSabWN9IPVmZkqf5lU6fubvv
7U2lp4w2X5rPwmQZ+l5ziCWh/IJIZAWtfVXfkPQEv67r7wubm1udu1YpbTKZeVP5N2d/3iJSxdkb
U8vkl8NXI2k0kkAVaCTIViijhbaZn+i0A50M7OdaL+nMUcsXu05Oger0yjRNa265usdEsUqFdqaL
KOO94wQ7V8RDEJJDTY7GLDIY63BQl8Bg7kHYg4lTzEWXk8zDRbe+NTgFhPoF5uRn3eiRmQmTO4S7
rk1x1PXeNrK8z3MvibhLFKMaR1/1gHc+WUnJAV2JFGslHTlFtoJ9x97BQS410DCcns2LwdGEiflJ
BpXoiYydXJuHL0w3HvAx/Vql1yKa3u2R6fS1Slo4HJxzEYn/zlev/RCEeTMo6GbfPKKEMH2NziK5
hKzneoUU3lfqwDwVSCrQvDFr047JiW1Uxk7IJ/SvQyuEAJlAksb156/CLmvADVyyU1CZWgY5EZAs
Q1d5wG13xP25LEW3TeTZkj+K0LX7atKqj5QzDeCBoq3od31P6D2Ja48dC6/niDbOkIlH5rxHWxKm
xSZPKCnY/d/jeA41eS26Ko0BnTyISVOLFxhVeQ9LFDt08glL2tZkq+OP8/74U8Ndp/SyOwp+HbDM
TVixtSlPnUaJw7fF5EGGFt6F+OadU/DOxCg22rTeZgaD8uo83MuH0Lc+/yI0vTaLGxA6gPzr1mTZ
dqMyiF/uO9blu4jq2TLgWkhVRZ/mXM/XOAxr867l52t8owOhWqNh6wgAHek52LhJzX7+E9InsnQd
3K6sU/E9EHFhVohFLtNvRDKiIZAkxIOWwauXLdjQY1DpL2sAs0En9fpcU/jLNoMJHC2K9AvqE4v0
mLEzPmN5HDhI0gsLZ4OFqR2kMljX4CEFen7tsm5lrZF3BTZJJaffijtLys6KavwBdAXbNcXPht4D
9QonSHfGOl/5MqdQ580cvq3b2NPlk3trehMAGiDw+J7RWHzmfj3aEKnhj39JXBpxntjmRD0Lx0B5
9Mk0p96RKgRoKG/QhqzaCGTimqAJNpVmoCUJNKih8t+jHiX34WJUhFPADgqDiRxvfnTdnbdnHvW2
V7kXcD/iFQo5PPKCPiULt4ndJUM6jXihMsdxUgmo/z1/9fjxdjF4kMdy37XEbUDkPG4aI/HaoKQr
VXRXiqjKURcsHQntSHfP8cM96fvP3aJIgZbc4OAfPpykVpi3xtt6uVfj2v+4ZI6kLYGG6sS4F8DQ
HxSjB9yzv9adam9SYUMCaYymcXvLpbR7khp3Cm1Rl14gdBoFJZJunG5PNyD37kEiTXAslNajw3bC
6bJroLvbwdEJQS+BlUN+/lLEIPBbWNKl6JoLfwncQp4F0Z9EQa9fgjDT5tLwEymG4W7u0ebCYjmL
dyPM1nnIm9eSOmctFMf2eha7s61KpwDvsu9zQR4vROTqtuze/qRylel3C8EDmhLVn0UFvNthLxaj
SfmhJ3jl3S6dPvF4/KiStn367W8EGJao0I/FntU0NDxKlgVKTCk5U0x8J5Z/SieQVzJGe/UY9gri
xaSXD0w5drMe4c1GkYkug+SWHI3GD4fKs0MTLb7mtLdGB+sPlzAZbJ6bR/VNbD8XOec4kaTOcYQq
w2EzRBqJZ9OlU4dvEeOTFM3c0xePIngnYXNDBgHDi/m/EXqFSn8b/lKa/4Fg/MkINtUd2nCtc7km
svBh8q1QUWrfed8mClPPbQFilYsitGNX/TkUUZxz3uEqF3TKn64DEKGzYqL6oU743D0RO7T1pj/f
hMKl+v45fUa8A6WmoPKs6j8ou5sxnj5n86Cu3tInnkr6WDXIuORgTAI+cCfEfHuuW+JQ+zzIvyTL
qXWVhs73MzeToxNefACDMtWd72JinEsvtIsrlcf6mEZ/k/GMJQvcGudtk3Y82wbjv2tB4mGeMf0N
WJ4fOaVWiLEMqt9WMGXzgtUBJDIoAC1IBeFzUNXlVHXgsHPWUIY2IHwImErxIn5PBlbmGE5YLn2Q
jSoSeXovJ7cTik7OGmjsDmZ/mEi6R5lNxhXa/xjRIa70QWHvhRjvjy91XGtz2cWcamNHWtJUwqqt
9KLQLks7Vuotc9XU46ts+1smgM9D9RippoOZau92g1UX2iMaIPIyrUI5tCpeRgvT9v/NqiXfwy5P
obrxnvePhDKJPZxPDDeqqCV9SUi0wXSwFrJIShbZTB2Pa5zzrMtNerj6x7zCBL6GIxNsWErQ598u
R3gsSjXePU9r+xBDhju+J+JgSwWtqZ9uzlWY5h4zK1qzf+IKGlAlITSoYBc+p5ZCkhamq7h/Ac8/
vwDk2kBmaZCCl/wVy+FJTkRIj6GacqijWbPPad3tob9RHveO9t+CX2au7GXaHry228hcs5HmBLIL
1Jeo1poprveVTk1nDrjvv8gfpjoV86KCXt0aEqxSGsx5iBwB7eokx6Go44Dxg7a0+paQQ8uybb6C
tCyiMgFM+iZxp6tB8WzMp+A/YEU2wK+yjOLuOjF1K9dwgl8xZeF40nPzJKRBEshh6XYOUQjUdnY3
dHrvWsf98Yi2/tESJgDzqzNUQEBFkOZUxiSgcvjxLRXLPtlLruLzOZwWkqbOwkRMFfKBxbY/0bJd
AVPf+RtVnNRCl2uNnomWdKA7Smhz7u13sMJjNUbxTJkIvqHsZeii1/bNIZuGEZX7qDUEdUyjDVbM
w3rSDXHiI0YdkRdmBC3I1nkIlYqpA8aLKDKFRAv9XsS78WU0CQIGEw3dzML+MVvtjJvjuxRZjFTA
GPtu2uam+4akVxebDhhDY2raYvjwWmZ3hThrfAnSTP4Zfhf85EM1BXetR3o40qA4Pf2Gyg76Jaz6
22+a5pNrb9a33tJDbgrqbe2XFq8mGVgsTKiQKD3Y+waV8My4Ok6HAqBtjHMyE5BtUAfN2pLEdtov
TNvkj01kFwlm6cj14fFNAmlbHhcpJ7X2TFOAGkVHXyt7Yw2tZHqQfOXn0yIQmKE5TdgEECGVSeOF
/6YND3lxkmLOQcHtqA0qMiFWOAkWngaLezxEp9Gdj9BkE0Mr8GiDtkqkcsB6E0u+yO3TT7TYT3+a
fEGHW/Ftak7fLHD8feLxNBudJgPm3zI63HdalgFatmIDEpDO5G85eYoBoay7hF3MY/UnDzZoz0j1
NeSx7PKRjHXtSoJ/Mpi6JjbnaPQ5LWkCL8N1p+CxYM17kczALi/lOiGoy2PkGn5ovLZNEUpY1qhA
bSBEuDUFtcfrhoBBOBUO3zIwWWVVC0zdpMerHhNjvWmGjapj9CBK8HNBkbAN/zG+lPgw0NGEb93i
gITVfOerJe4VauraIjhFQOP77yfoyse4aRmj76etrnbGo1C8+tuZOwo6NYPwNbcMQn0+OuGggmw5
AZN7xtfhPjp1A8V6+9wPRNZx6xhxEZHBK38Z5qEjyOoyEHfW3xnnVwSbl1pcIYS2spt7XPsD5HHO
LSIZpccA0yl6lwiZJBcpkZWuj971oz4PnDbzS+advqEepJeIfM5QNRFWNv5Lf8XZhCMCpqBjtrZL
uq7vNpdGSmPZexJeUwHgKlsH31c0tJgwwXHgzqa+qH3kTDrlqVD2V/sfp0Yep0lIHqm0s9khv9pR
IIHwDWAH5W+i+rmVoKbLLQCyQwjBzVDfwORwpw+I3qG2wZB6Z+poPLgz0Ul1kbgTkjiuwt/z2lrD
tk19BRXI8INJxTcM/mwxQmI8JIS4nhqb4E+xHxcCoRlUB2LiBYaJEHpI2PVdhyWzBs4CvdFSy02/
KebjNio5doG4JP7nQnOHv1zylCkbE8Q/GIPKgdeIlfT9ywwoC9WSQD6G9iKIPCupn4YQ+ys0N7lw
KupyuEn/Aebnd6iXuMQ+aD2iGMdhMCEWOukMXJZkUEdAIYkeZszhGtgBYnQ88U0P4Z/BZ2ybHqX1
1kFXpN92D4Qlv7qG9GM301fEDk4M44uOMBUMXCAV6nl6JISc4tiZvW7fPLEnkrSR6Pntv8ZMHIrW
Lbza0LsAv6DkHXiTDtMYLh/xC66sCW5ZyIx5kaHfwgi59znEFCEmtALCH669wOEnVJ4ylZae72AR
WWjKB1gSYaBlRu8mz+9IayBCyZdabTuBVYT4kPJuxlhG6Mmr0FInB3lSnCWMAuRjdwNqwYq95+0l
nayyD9UCkBcN8TjFRUUeLDzHuLPXRe0enFOYGeWyzFk3ARbK73ahE1Oytc+mtx2d3EEZNQBwR1tG
pzE+TOtlZJ0iSz10kNWaCJszAFYjLtJkU7fEy9euPmsvS4YBd/sotdlbwtlGJUAvxU29kfccOHFA
YUBAPSlvARd8oVum/xUtSVadD8ExmSswHYkXxhPclCWTRg/ieOiJCtc1/jAPo4ZqR4PO9/a0SmUC
+ynjDuuDqKJpeq6rqYR4wZWilnjo6hMq8xnaCpzmHR/ttfpga6WiDCJF5YVF4rl8kmGWEBBRDObp
koS/nxJskAYEDKWN0A++jgxTzV2dZ5qwe70WuGnS8sTr7RV9D623hvBPA2ZUHgk8xwFx7UEpcksC
0Nvwb3Bct0Houao/HN7OnLFeUbKAMHgoY9wIpAEvOewDO6WVhMrUwCymDyTqVLVP9/EYCswjA+we
1dr8wBu3Co173BAHjpgxaeK1LY7W7QZtuJhVqx2EL+KypVoUWLqNf3YIGeOEie+qK7MHKc9UOcKm
meo3vmsXV5GlSL07evjMqKqn15NbrduydjxkD3Y8j7kRCFWr9zm3F1aaNS/PNEdk8TK0BWIaapWE
aZARI9psQW85Fk++HdvYpO1BLfe4Ijehyintu/o/CsNG3gzXJ3Pr/Gm7ZeKGSj0AaKWR1gDpvR1o
n5yGYdb84M12H8BeDnsudrwaj4tEIwpOpa5uLDVbmLL5d+s4sQCHiw2sAFQi+c5T9tSsHaGGdLg0
SnWeGG+e4AJPf9RB7UPvu5Dy/W/SBfK7BEJekzFnqtY+0xnnH3NgbMJwTH7zF+84eOt6VAwFhPxy
gNpUt2Oc/Oydv4bQw7eXV99fy/yVolCnrBpNh62XIqOQpT9U/0/tx6NHLyQJcbyjZHM3ztBQOcLM
UhjZMk4gOQ42zI3ItyCRLHGh6G+8dGocI1AsoJAeKZymEajYE9FuFJJgtX+siD6svN5UAjut4Vdt
LQMfdv5gYtevoRk5qubyfyKYgqL4EeJE7iL7KVYKak7sLik1z0futPC9gtyZE0IFryLBs6QJLekg
xzLUsOTTnWyR7zV0khIn1OzQUbSYMDjejYoBR8BSw0w0Gbaf6kYa1WEz4a7F1tN9ZuY2mR0YlmMz
8K33t7wvWEG4HUh0qUoDYitmARIwd7UH0fi/pTY2jKOGnYpKlf2ErRuKv7lh0aJpacIbVsucydGV
0N1Hh/YMLciQHhpmb2mJux5dXSH2IcgAMv1jrWy7vR5qq7BhZd+9Ylr+MA7/A1lTWvNpWu/AD/aC
Qv97H3LkSmNupBIDZ7yYasN19BdGeXwhSgu5KdQiC+bbMSHLhL/ASKlDxVbxvlzET+SttedQN47K
nV0unfA/bWkVw8NfEGl1r1Ozjd598d6Ke64VzrYZJWKlxN3E9w8frwnotMEldDjIIOK0uwqEcf2S
ng+9HRfOim25alHKtoTzYhdXAqIgcTxN8xj8Ph38/ewzVrkMcJQgawrZxNFgIuLgahVohnsfOfJp
bPrUvGAuJMab/B94aJff5TzVk28qBDUKbKSpcXvoEVamXv+HFY18QA2W2ufFlBxmT2NCy0IODkxr
5FFRX+up/2Ov7yruJ1rYo3kwTJJQ/8LiQPhfP5H8PcJWC0tEB7OjhuICMAVzKShPuJ5+oZgevM/E
+EekQgfqyW1VJlM5fHIoX8c1zLnKHG8wQLrsBBDfvm2qMnon5ty+E4GoNdDbZGS5C5rBQcpzv5GH
BbPrvD53i1HkEXDLVg1bXaT7VW2DJtOsVjNQ4RBxy1WxZ+XB00n9zxHowWL7PqA3GGoV6x+0/0e3
6qsXFJVwkXPEbNbJTs8pO7OuBkcsWUHvX9FE/45VkopmW07M3yC8WA+gqc+om/DLuIs6abqO3yVO
TVaHEUK8butUclVIu8CFYST9sgjtxqTM5Yy0//xEOV8Z/B4GcOSXa4DUY4N0ntc/ZjCvh6/x3Olb
oFqagZfeh9pcUFmzKovS8BAWPdUtg6SJX5rsCdnczvJ/ZaWLvMRCS1RCO5o8oXnLmspmFNFoep6Q
3yC6DwfcbvX57w1a7QIBnpbA7w8XPI2hawZ9vUtJ3u6q1pRkjzN8MhmUJw/N6+x4Ck7TnNrtr9Ex
rO3dmWvP6+ZO3kgdTi0z8R3Dxaog2Cu0cFteDSGb4pop6Hq6L25I24WdCI+wLI6g5zqpZZ91NUKM
r4CBm6obok0u0jqyQju+VHNhG8ZJidN0EdHcP+jdOohYJJ/oeY9I6cpC7UGg2u9Ac2fVKqScoV5U
1nuAbkPno92QJwqNhKPPnNUJXe550RMlBdpzId+TB62DweSmKy1HV6MP3Ph5yvhSHn46i+72vA+t
/HeBzhII63ca5Xtf1NZoynKMB2GjBNcNUAiDdKQVw1fIwPG61wEFySU+LBN7TvuFVnkEHfFPRmpo
D71xfEhaoRYCDBMy6JpT4Z2OvoY1EJkth4IEKdX1fhbMdGGIO/tuoxVHZShQks/31KwrJpOxQwu1
Z/GLYRawFf5urfMHgHt6lD9LD1TFTJvobEtVTrklNouSJgc3Jrn8H3xmVW8a0ffjbpEHiSq8T6ua
tfNhS91Je6HaE+9iG/uZNHMb4klH0xYUfFCgd0d11LlcnE8BbcahM0DwCW4hkPEjzPG0WX6lW3g0
AKC436g+d7J+Tn7U/wkoQ0FMVLKwNZdeC3MAsvIVNJCIH9TDNMnvPFHVCKBNfdrDomssfpEyNiZT
/9qEmOYGvWV9kG9qOmL64a8ZV5Oy+92Gs8AwvxfQowInVbylP4pHbdia1Fn8Kvrnh8/7Wdj8PtQh
4UtMlRlXdXHeGZgdrYVic+QFavIaUQHGf/oa/Nk8X4r+iqJglysNK5I4aeJP2hOSry9byGp8hbzy
p8L0/2xRWJWIcRq8dwzXZ6KEWorNcjsGM1p4+lhNRogBdewOrmqkXYEGlBr+jd9Y2c4vlYPcAuB/
Vuw8zJC4ZyOIpOP48TksuI8jEDQZqOM6Qwe+wBTwoZcZGvKhGAFY90Sd/UDOJ5VT8D2yJZSWeWyL
vmy1tH6xcVCQ5Qp/sByxeTC+Y1493Q9xu6A6NxfxuJ8c+F+jBEQJTEIjKxOR0e1zNjczXJ74/LMX
trfzUQ0tLxRc3ep5qYnpNBZoXiS05ahpilcMQAgUD6Eo/BZ6oNgaBHu1i3BypnBX5a9qLZUqSjVt
yCq2hSQFENFEISLezSO/pHk+k+vZcz+0REmq9NxjeHO/1DmBlqN6ZpZ98LdNOqeql96eEsgra2+t
9yrMUTkeVElcbakkDVVD+OHY4DmTSx+/8FnvE4a8NW0UNu6wddjCo1IegrAzb1QrvlDXk/gGiPdY
y5YPr9KbLtRdBg3v6sZk6/ytSmgnAlrcxjhqP4cWAsEBoU6VCvMzrycfTzB6aWRz+OGBcVThQn53
eBvMt6xgsohcCZLrvMksA68UsHadAtNIHq64j6POJnRAh6+88tVDLXVreYYbGA15dYv4zG2TUuea
Pg0uhIvt5bxNLiznxnClGoOp05NJ/I1ngrGJfrpcH1ORcD8c4WK8FUD7iSx+sP4FYhLLNrx2fQqP
++ULPADe/PhcVzXqt0lBYL1P5RWnmr8Dq2U1+6JUzDMVk0ES9bIt2VPl5tJvOKh6Dnnjhuv984b+
DCN0PatY/6crf+UeTOb6EfHc3drP/YwH52Krp/guoLLwVJEUniZLMtx4VHf/No6HSbVDUo//rqbg
ytV5j+4b9qBEfF2KtA25uZHhPBwih+M8/1Fkh6Ozkk3T5WsjX2I4B6dhaXVHV40LW9nJrJlMAqpn
c8EDd/J8dJDC2r+RQ62HFSERAbWx0Rj7mE3vVeHbEO0iysyGVSCXh8/XV+ZJ3Zvw6PPqRUwuIMaw
P7qBiz+b3tAbN12+SI4FOMl+9phBJJTBT6DSprU6zPnS4CxOurCsWA762sP4+flvGLWbckyIFR67
7ejElG8Ovj7LdJ8fcFBRdu2knCc2PJQE5LVmYL7clUrcS+Vb3Zys0QK7pKVuKCDSycZtuqH3wGTP
JulaAVD/LLo0LBdgGQwzlimYMb2c8A9VZae5byBPu+Y6rwF3z2EeJqMSCKfmgad0Yj3+5zCMS8PT
F7g/GLsBR3Ss95vj54tRXJDxe1J+gTOfgsV5YLhjvBFNM9k1fjXu2CO3P3Fd7anPiaRj7I05pstB
gStnITYh6BKO13Z384uJBLIgc+7lKMA9hPLN5IjLz3S4c7ljVTu/PmKzfJ082JwhgdZ1qsDYaPE4
1YGITk8cHR5lqLZa5ICONPhjbi+0ZQV/R0rmeLJME3NT+DyinbPvnfGURB6FOs2lZ3AFXfHhgnnq
AVxF/HnUe/4c4p5/ZOa0LzHD2aRVr7CS6ksEnTCqRHeubHEOYyZ70h4PeQNmwQEiHuT3lton2lDw
j3odYvHZp4LqCdd5drHcWocfzLY9T1jYGYx8GqRAx5ewrH5ppubjea6hDWNEryGNXK6TIMqD71uT
2F/epkYixA4t30dZbBJ36/KVItqV4JMkzcxpDJMcPqmZEIPx/nJCnbAscWUE1fgk2UQZHAa3iiWG
3V6w9gQQUCOq4+H9L6FlSYNYnuOMrnMs1DXR1l435K266Wx43ZPTTs2gWiS9jD2uV2swXlXv94/c
r8Gc6J3kJEsAf0RNrT6298TGVa0v7CwSWFVlFLeNNEQNDKkwSAH5oINLEQZFMDWdD4rjx5vHe7cn
RoxNGs3rw6ruw+UgbhsVY+mn5qw/0t8U2hVgQq7LU3nS4pIeQAK51dgU0mRloh8Ekb0ouvAqO91A
SAjavYTkzL8D8Dh7GPa4VTWJBtTAf6LOoUjKM6m91XhCNGXr3i251NH7tFUKzYWcxOepg2asLRcS
emvLIft8agMXrFlIDNd794/lpyC4KYrx3lq3svx7pukyC0zkeNd+cNYEmbW8hr/RQ+pUF9u4t8Og
gaQ5F9ia30rWWHJ4I5FilXt+7JhXPxviKj0ifEOsgMnm30ihK++Lp7W+QGNAVQPy+90FISDVh1WV
SigqHzHcbXXbqPG0msamEb6GfvJF3xwepR8qD49rzPo25NxL5qr18yS7379NU66yFSJ9Mc5Rbve8
6gfrTia235dPv1YE5onaLNC8a0SCJSRUZ3/WyYRU+fpdbsX01qKdboLN3JJugx1FbvEhUJXkc95z
hTG/kSKbyTtuUjohk7li8l2lJqEiwJOuSiT5XWWb43h2CCyk6oxDTjiu+hRPg7I7ElRRTFnxgQ/e
Qumwls4ZJsPMlL1bUQK56A8Dd8bMLlXk6UmFwo0kd36nYLhXOgnvkiH5cDEgtbBzdWNXrTd7YFIO
fK1GwPtpyS/8S+Noh7nW+ZpXRL06rthoAhz0+uk5SBPMaT/2hGOiv3c+ploRXznoMaIp+eRidXNk
NnOAEGDyU72ZoSqEJaOpA3hMLmopcvVfHJ+AOtosDNvI0XQ+jbb4qoU4h/zBlia7BQ5UejHX4/RA
I2mgi/y35rJm87Z9ts66TPLkUy6T9SS7FIrUzHBqUE3PDvlX8akPdQSAPZ+/AmgvRVeYvag+Sk37
tl8pThAYqMjRGacEta//r4nZ1qdKe82/fsAw22eKzMvLSxcvc6kqMnQR4XkjZ6zdnngOd+SuCja/
n4SMvt842RLF3Smk4cJgC425Z/2G7+kXn4IUrQbKP4yhPbehNCI0J5gvivrHT9jlKpJGcQRWEQtY
7Ox+x585YkKuXELKGkxxWGRgkhdo3BMSvNJuL253aDbHTG+9/F5VWhUWeGygn3ua0TTlSBf+/5P5
EbWodfHxeXqQZHxKIDcSKZZio/Bk/naBRNmbrK4thoH6Nh3qDBo6fvZ6WBKw7OZpmkFPR3QrRBOI
sI9o4kCwld7Hs1zsxsKLPhRJm500IAHN08QzBda9SDBBjIoKS5ZMWRSBbTxfM9y6Cdo4DQjP1SLE
VbMHmgbIh6FRjHvwxp0eHxGs11cJkktMi6VDmFdoKfYiB11iKkpP81OazUwIX5vrO9Sj/ARIlJTC
spm4US6QZzG2aMn5w9mt+rUVvQ9XSnlN3EGono7XRHO+owZmuF1UcQp/ozYys1iDjoV5alJASkVL
lTAbIPRg9lEj9XsOiJ1GECxoAXOAu03C7dRywcg2Qi55hAFXnd3pVzVq3kuPIfuUfXQOmExJM0fz
RIyKLmTGvluY7qazV2igIudOJWVzTKT4sCBKhfXqbzaFxAKDQyGcLr1+Jl4BinsYtFqqX3K1tI4D
Wd7JO+0QyWBgbkal+Zskp/42cMZJ1pbX97kQ1ixzqh9skYq1s4NEed0JenvuSSUs7AMftXofxlV1
Wx8c8k+Ttmnve+g3qbN+r3wzFaB1BE3IR7QrfLi/bnfQPrjfCF2OjEZB/RV4BQPp5z2/iiYaVXMB
ff3UjmE83HE1smOVLpoh+woeob/FbtOC3TkAQWRn6HyDvWUXgtu6trkU7iST1wIHTFTbbj0devS4
CoDl44qT8R2bYGrw7A8PEjfLr1oTcIBZBxPCnSNRbpQN7S3dG1HPV6W6GH8HQpqTTlE+rcEeG0Os
XbvWQRvmhr0ZvBWYInxzjv4FRZ9aI2NulrNfivgN59BEECe5I+Be6rhMUwlIfGf1tl/6jLAQBDSx
c1LTsMC9O1O8IsYvNpvW0jlRnx+GBIn0lcL523Y87FrmOD1zHWoWZodHyRl92SGYjXqltfGAEzrn
xIXz9xci3g6/Qlg2ySgyQ/ZnoQuZ+yR7ySj/Rgk5EHdGr5pxsCj10ntxUNuVy/6EslT7Hhl2nCqK
4vMGfpLZKvUO5l6+VGKkoUxfQGeEwLDlXEebqOcCefNNfIQo2m3RirtpAEKE/RbkOQ1gAd7nXOkj
24vHaWS88RuIF8KnA5FkxUXQyFbXb0EMeiJui5AxewmhsTmYkej32Uq4FieD/tOd8MVmHX/z3TqV
3CdHenOeQwVvuiWbx4FVA6LGb1ZD+JQrgE087CTWpD2k3BLgfdOFzfpF1u6m5GVvU41pLzVs9MLb
3UBkV6+47pys6j2DkebE5cZ/Jof0eTU6fbnJcAd0zyv7aKyXzq9xYDebpadR1Rj1RxoX9KCQe4fB
Hs+AdTahncwdcpa/g4+XQSfkoPrBF5BWvV0kE6a2oGzanOCuoqzxZhztX4H9iMVIvnDHqllrsy3b
4ykH4y4caW25i2ePs1NfqePuo4wSIzW3uYgqTsR+bWCLiSnCCbxDpgZkINFHJ42Da2yh0HNRmCnU
zF7fRi0XyOQ3Z/iL/KRuKyy8OPDLteGP4E93YmltXzPw1sN8+vY2Uw9RdHIjPfnOD6VvAwMN6adK
ob6T3W+i6VzVEdhyBGo6QS8wllej3w63uS1l3bcRPcdWuoHqFA/A2f/KinD7yr6Vn8aq/084UV63
nVyCh9ivIaZ3euWzm3U0jheWAvJKeQm74J0EP9y9oTQg0zJapdPL+cyjTf7EIAv33y6eAX2feUkA
XNmPORM7wdmMij+0SNFFmwQemCYB1Ypy8le0J9BfdEcEWWl85JPCiwz92spF4/RkjrBtW5ALaHld
kMbUiDQvUtjNR3fICjc1R2xuuiMAXdbA4DgVvBJg78LEtXLQlX8ky+UMxbItxrF8pcGk0vnaZz7F
/zHv272X4pLj2hzmZg2rEa4h+CaI0CqRoLS4t5s4m+NlM6VSXf1PUlzRT/lg8oEW9JQfDbVKkk7I
2iMU7yU5YQPYk4nw9zNSeO1vImcIN4EoLKzLBiM1HUVTkinTqHujmNoHjU2UGEyqDU+JNNXDxir+
KiQz3C5Mouym7rWpe+QdueOzWB0ngEj2sxgUt3spJbo9x7l9mIEz8rCyDelzwqc5LkUtfTW7Th53
LRdsZh+0oNgyUYyO95KdtTp7utIolhkvIxo7lFNCHCX75BYErGQhRxJbzW/kGnN0ZaG1swH6G1OC
sUn/bEd4APcv7vI6DOtvUmRQ+/1rFOMU4Fo9cwnA4QHsg8Eaaxn2fwK9Gd3Y6bXKzGaU6gOU/VXM
Gty0NcDEo2vuwgsVT/SBmQt+Z9dyaWLpKaXvyg4EfOZy9gix5Ow7WDCzusGCh41VXkLMRpxAQgI2
edX5qL6c7ztVdvjN6mI7AvdKQFWqfU6oAuNdymX/RCu1Sv/MLaMKijiow2lbbSMHj3KBYRjLbwBQ
DcpCOE1p9Z23I8M2lJsnbR3+21Zv6aPs6nYU4++LMGt2ZqabIAo+A3cE8JnaOUuMK2X8rMkRU5bD
i3D9Hj3d33kYLfJAXHAfSwl7t7zYWQLBNhJJwI58JS/aaUOYnx9g+0pGcYq8rMsK6ADI8HDafgvQ
BEpYC5s3v4o3y0R5UO6TWWis/7TMR4ABP/rjk+cMW0xrF6yxHvKDHa7GIr7GgswXonnw4DVg5HRt
t6gi8NquBlt9k13i2131i4L7T36xZhV7TPcmfCIUEkv/6LLD4rzdRemK0jmBYptsVQJONqviH2Mw
6fl0a7ADy5xIWc+/G2JpINm7md4U9aeAXRLnVish9/xxdqV1+RNdRIag8g8G0QKTh/kBVq5IgiMa
9UhiAljZEym2meclCbTDsccYI6g5dC8eVOv915T4HQocj6lODzFdhbg/7jkOWgeAaLJxgcxB9HDS
prhi2Ev8ywPQITrZG3Ur/zUs6tIUpisddFmWtugWM0j9CLj5scJ3jfPQF+ok4CmvVVgcqPAm4G4g
a2r18E/vtvYbUlBmsZ4/LXL/IOwrFJjzpXcykhpAu8Scmi/bSmU8+ZALtxurWiyv+MqqgDfZFun+
Yi8HILg3ydlp/dWyuGFZGBe0Jn+8tqYd/9rFjW4mQW2JTjHjT7gYr9Q6QOlEKQPtkesZRcaaajTw
nPI1xlvqIQK4XWCZs+4XGuiMzoSnD6ABMmBAgP2Oiykgo9OonhrcGg+wTm+LctcyIKIJ6o17ikL1
Ylt/fw/hjTw10CfACw2mFeCKxpgltAwp8zrR0YH7J+TPBy3aitVrlrv+dXOkc8S7EXgl0oXJ5DxD
8KJuVoh+h+P1ri9tgbL0ETk/5d0tM8+zLNBqIit3z8/ja0fkaAKW9dzj8vOKVuJey9do1hnqhp+3
Ao4UvYmeCwVqPheFc/zgdaj9DMCJ9is29cJY0QR6F7rXc4INRB+jUHaws5waZwxzBrQ7kLmxtKQy
G3S0s4TY9Y+3m2EpFtS2IgNKJ47/DqnfcVmc5mihe5oTVwZ11u3R7R+iGxib0rhkERDPimsOi31S
DXrlsawfxjKYQcV1UiecONR0Pjn79ftR7fFm5dvBLg21m3DTGBVuk+2lKHDT0KM6puWwo9UaAqr/
99+2xTZ5dzG1FCHDSo1OsV3eMY4hgWC44rxFhMPl3WXxxaUn0jTzF87krrZ9Zf++23LRnQHa3VME
kAuYaXiLsKIsMjViYE4tqHV/A7EHexUxxSSmbpYUGzbMRUi/b9ZT/pJYC0KEUk0Yh6F95X9KgTad
9Azn10sGkdX0pweueHghw50U7/Mp8GLcfvFvUXthsjuCneB/PLEy+gpkpdtu1Pjek5FzspnkknKg
HCOkX9x2BY2XJZ4cF4RhToR+22LN+eeNZSAcvZ25kphKtsiQUND9qTVp7taKzb5m54W4hSJO6yDl
S6z7r91eFHE4Mg5FE6Og/h6MywpCVCRdPZNcRKGSVV+I1m3RqJuypXaJsgMJAr45KsZU2PzDDgTF
lTACI4hXMrQhc+0UUJhbbHW8LnFf5sxNsGU+2MQ+2FrE8XYkLAYSavFc/pECPjKIASNgsfnZzbdH
YcdSoDUe1TTPAB+efZ0kDXGQEu28czr30v5/f86TiqFY/IK0gsU89iUKKIyzFN0UpEcJQ2eK5654
3LZnSrIx9yjAfrshW6ZfqWKqCmik7+LH9IDVrdmT011BPSQXUVhnqCfbxatcOUihksCccLxSf6kQ
/QXk3k4IlxT/OGt/dMQa6tvoQhkDihGGMf66gUuFP5Rz7ibnLvV2jjXEdZuCnZP0nNJY3NxSRsuI
LtW6Awxx7/sJeWoXzKNou6upkGbGsoKnxhc7ShgO5eFkPYIxDzmiiRQCxrf1/jhXazcaVxJi6YVk
DtcrzcFgg2tMtR7t1pLB4qlqioUOBJ550xNVhTOr3s9DGLAli08A8xbHyhj0g8ZgVYnekJFUveZy
EPs2nNpv9g0Qp3891fhY0h412UixZVVjMOXViDL+vgfYrimcBeWjKsnDJSbH0Q4qcJl/TLFsu/zE
oXoZ+1n3qaw3HwWibOLPgmmnmWzXuSzdr+y/9nOpSGYeoOLf+LpKr252M3UnKWojNk5AQVdqWrvB
lVhBUG4fYodyPlVd3WBZkAZQVhZoW4STn33wYFCQb0KqAzELb5bQJWUi253I4w2mIkKLauQLcd0v
PdO89udD/eb8scvW0A3qtAzUAlMPyTOPW69p1nDycENMq24sjXn5KkiowqYR77XifDpeyOpOg29F
BrvS1rt46/kAQvsT6w1Ibc/pOz0smbSJPe/TBVq1sAxEutnU3o2oiUqWWSidvsC1kJGrAj636ymG
XeBBDVcNJIxQtstk9orbd93m3wpuxdXoIkPUxd6MfZRWxQ6W6Z5V7x/uyTc4pz+DwmsgCltrOaAT
sMvdoRsU7FRFF5ALCVv2imRhlK4v3cERAMkO4L0yGH6ub3739cJR3UI1/pycqhR5NH37g42WQ8kk
x4CefE/jOYdRdg3fwqB9p/Gc0HcHwzXvCZMjxLlUQ7ll5nN6vdh1M7bO+PyVchx0n97TAzLo/TS3
hjLcrNwRhrzKnrDgzkqtyrmi6PwVR3fm3eU2+tSfS3mBFoYpHQOnc2z3Kyn6X34YXfi3Y9XBi7X8
C6CMIRD4dvwHyoYu4nVcrVqBrc//dPAGc5AghFGo4u48YCagVYTl0wXBVoEh2urwpjuLVeJR+bUZ
zK607onuuzyuGyqB8Y4srnclaeuVuWOfQ+KnfIRzkMM//SoeDxWM/Q4CDTwek3qXIxDZvd6ULlF8
s5fiF8Pe07Uv/76WA16zZ5psZh43WI8f+ZeZfGITuCv89TPSZfLMXeZNRM3CYi6qBApQL+GlGHFl
31ZrcurBMhUSG38x4MO8dFRWl28WNX4C/q/ewaIhgtiuVaprh5dB0RHCr6gnqR4mbqkprGcl8dUA
0dxEz5VOqM/vGfla6OYzx6GbJ9LMGkp/Y29PRVpxu6mquQ2nnO9e08VoU/oB30uvn44YSQhq3uKx
AAaHSgrvTtusn1h41VuSzBOFI5iMLyI4kddHkUzJNQwpjhq1nVRu7pGsdlugJ2rDtw88CyyUFmBD
Aa4L+Iq9NJPVyWIM7bkhir103cB7KGw35oSFS+UwFuoXLbQ8qYCx5mFZCF5H0WE88e9Dijs5PWLm
jjeF1D3D/3Z3s81V6PCGi2XIa3m0kVKkGr2k3ciGAMMcOtU6wqCaI1C5fdXOFHGSdhC2AdYug1xB
xFIeBmWRlsCGXfzI+8NuwppHkE5hYbVN56eusuyuY/mYX+eu8wcBmY/9bWGQCrjdqO6X3rSR/iPE
p30icPNMRZ9Jy0ZWkmi96ceuloma2CM2uvyYsiNnLCmgjnJx6Pnvebm8DpTFZ+Tsnn8S7fE3WmBd
W0mPNvI/VVJ0EU0sVfinKyjut0S3zg/EqkKz5sXeVfQ25nJzUxAgFdgx3RVhdUPrLyCSOa3zjE8R
YM52v+IS1I0HB/WuMx1BFyCbtrr58MsqtILQ7cIwuVV3TU1WwHz59yPsdWtauNY0k2KbS1ceg/T0
5leAnMFaePec1BSVQ6rYfFgDTP3euDkNEMA3vciTwpe+9bbviyhbvDRkDJ8TX/LPSXNKQ7EyCjes
0V+GeqCKGW2t363BzcPXE3tCFIq5HLxB/fMvUkSGDRUP1389QtZFk3cHt1v/3aLYbGOFAm5jeIWX
6e+Z58MEdTUc6oAIFtU0vkFbZzRBgeizpJMsG+VXvHjiRAhgsKsdTWw+aKGOoYeh+TyXQLt7n50S
g/rTcSs0+1I2ntr2KiX4mD5mJ5xDh9KeENBSxorAZgfTx69fKA1qmwIj9HBhWVG6URAVlxOKwmgj
VsMsLBkXSdEkwVKcFlA8E3PU/Kz5fSEVZSUhyGof1cqXWZlc9n88jHfggTGYIxtk5s3kmN/xncQt
AjaQXVZZ76kZhjw/VNRDMWHZSHk1LDuvQ27PukRx60iP9AIfJfq7+whuqAiFovFUKin1w6pBKD1z
AXUsYHXhqlGkgj98GAvKS4B7IkY5ILn7PAgKCR1ZSKnW2r1oZ9cmvRCn5aA7hj0s4flRosrVH0JM
QqVdA5Pnf7nfBLtjUo5V0tfKczKhVU7tR6jx/OTuH62p/wx9gWQrXn7Y27Sw/LZ0LZJjUmVx0GqQ
7ZHD+3No2de+Uen8WZDeY9keap+N7275po6WIYuc1mYIZ13qK8zhc3oEwvxi07RA5LG0oZiKKNYZ
rpY2PfZ6vn/pUWjXcW3k0qaH/j8K9mvlXyvX2LFjQCslCvvLzL7VBZxSe2G20KpRz7j2KYqw5I99
g3jPBN3jlNBaWuh/HeDeYPcxPEh9/LY9EgCBA1HMItzWcFPbc2uyokbcNeuRkFx7Av4CC4abjdhQ
riRfmsOf6aWdDHAg40X6kwBqHozRmpQPpkEsqyYLCRCNb68jX+Ueyj1TJP8ikjlyHKs+ABcHbgCj
aqdRa9f5fnGO7Mm99bZaheKYrupZQ9oM6I8VoELX1PcNmXuWCWDrZK0J4YFu6ZF2GdBcdqU894Gs
NjH/rQcI3BUo/2FxyrEs28p51aEOZ+YWiAzHOPSjySdLJqYC7U38J8bmlpJF1wjeto48BLqqbQjU
uVxFzWpDKxEz5btq5wAXHWBQVVIdpO378VKrERDtEN3ZoyYM0gBR+ZOvwnv/O2InnHg04Njm94bL
Ffj7V2ULzikC1V/TmTZoiGQVo8eZWp+juGoxjYrtgjIs+X4EVXB6ogdpiVaMpSWv4+vz42FYdAxk
BOiOk+7gyfaK2vLIn0xuuH2dfkGTj/mQGr3vTJPcXEfVeZOTaud8F/YyZbzbpuTQPFN1UATGDN6y
7+64r76ajK9V/Rkq/3E20JDeosuNIz+yc5s+Ygi6yko9n3q10SjSlmvrjqiXfV1GMPoSpAFE/ep7
BvYTugPr64rlu5OYH1Ah5uiJ/TDmhgGD9ODvQXTw1OwzM8+5QgB+qAN95y8cJzvxqv/hCmMzwM9p
uKRTcKmAl1UJK6/SV/5brbtRUZRLW+n6aPb8Waoo+aYWJgVVQHwVhszsCAS5H9qp9udCZ7CiLrQR
v8WppEn3sEplsGDL90U46d19/yYTdCOXFoee+OgPhJeWT6CP4ZaCKryqMFIoXq7h/8VnzTyfbW9t
yLaTrxVRpxk4XwgM+lQfKq2IfYY9kbPyWxnev7afZ81P+eLY3G2tJHjhdSd0jcZ1j1taRQv7CRUN
ZObKKZkqSvaQ+ButPCooairhkZ3rGAd7tWXgBeqPeLsCbg3P06VOI6+5wsd7KKUais0doXyeEBVu
b6CHheCLZ+frj6wF2uID19F31nL7RtALwH5hfFDzC+nntGz43cjFgnqr6PiHnlki3IEYqfMGpqrd
XR80wdj7Pb/vdaA62nFI4+bBOIivr19tSs3W5AX5TWf6tGOf5FzkERauZDe7fQzz8SM0k7erPeIv
euVVBZWRucqJA0MAHSMzdzRoljZXXCEmUTlCH2xVRTrO4wpEXmJ98hwHNX2a33JYc4IsbLCrfn6g
pBRxJekpcfeGTC76+EcIms+z0uugxK5GvATFxALRn8AAnNoKqC7ImOrW1Ljp0CtswxzPVue/ydgM
phbP2Ck076DAp3Ku5L9N3QnQnJzDHtMyNpZ/KbOZ1zBfGdaQTcLzyG5LJImN69duN+hHO/kLauRp
YzpKQVsjvmGJ7owx4HixtDIcD49npwbmfQ9fnbJ0OF7OE6J1u2CqquilyD7qs0mPNNdJqKiIAaBy
1mCU0HMW3YnkN/aBfJ/9MpQsb7PfTlRZbMyDWH6+vU7YTgu5PG3JGfVc9zHYidZHwsmU8kYsS3cB
5fW/XFy7S4LcRvCiutCSbi17cFHJ+HCwqWWcpOteqcV4JMsCONt6L/EBepY5fKhwgYQIjndjbwP9
qBNLjvKEpcIsM0lzFbWwS+biUqaJUu+rbj7I/gO6Vvz3WwJZhmWgmWDeD5pWYbU0wATgoQaLUPdn
vQ02bOieXky4LHqW4LxVBNSlAb4wZ1PQNa+aYL4YXVP23vb8cStK/d6N/tUuzqOT7IF6O2n38bBd
zhKwzRLzp0QOi7g0R4o+E5abAfYJWUUVUOgV+HoPfL5tUHn3cNIhbdJKTw83mE+WCca8djr9enXy
c6LnMZp2+S26ig0itnrBSaimLPl4eeWAfk/oI4926+5j4h/dSXc4xjLRgmheK2AAgKtteQmnuiAf
/cPud75NyllUmRskUBuzsWHcnI45Ly8KoA/7ByeI/6jfJkhNoqrfOAjX6XRBYk9HkQtvt3sVTko4
GaBDKEUHkpLsHXLDZMPtjJ1Gi8TA886KtZyfBs4/q9PjiXMkWTSHGCS69GWC5a+vgt+jEsiv2qJt
AE6SfaWmDEIUSB0z9u0kyWUhoN3rHeRRDDUNrAHSnjWC/lt83dyw4J3TNf6lky3zTxK+QHY8orOh
RNUWbNeQZdvGfqqMibmh4KLjrtYV/as89N+mb20kmIj1ypR6Mq5ouLSShURq0w6bFTrnP0xAY6D3
6CiDgMwLNXbxwnb2ixtrlpk98avi12Ya1HheFB8PLkl+SgQIFemIWqyY3mx61xFDCLsclCJdXtOL
A1atCKyvM+4gqxMPoVajIqj24X6P3iO8Of0C9lo92V2tQPoa/w8g/Qb8DASS+qXnQMjd41G73IY8
gJHLM3kbc5uiJ86uiO05P9cMuBqXQ15CsvCBgS4+t5iUAVI01RNn3s9Qr08drQA4A9585XvhpDvj
OwditIJfbaR9mzU1L6xn0zTyjWwl0ykFKxlKhFtyGygoDYEb1FTPQ3O705UvME26ektbBzrlztUP
zTRjhkqFUTzpsX1Lo+ft/mCPaRjTXSU1/djy0fkYl8y1BDnm2gTG4Ms4HEjbmUMd3XoLYBJeI3qz
/r6SSM/NW/ksiaOGZX0z+fqkhLP98vrtJIJKbBIWVn9qC3GW+TXVGuj+yHr7FLH73ihHL4jZaZAx
8zxhEtsnTRGCHsVwV7U9MLJMQdQkNq18Ian5PV7jeXKuyWlow3t16bBVPUzSaHe3BhexsfAZLMYg
lIopPfxWEKtKPxG0uOYs7FnRkBayRw96Pjhy8YbpSE3xUPOz8R33h/kVZOnlbNqlx1D/CAggplWR
WOeLRKxr8iUtPJT6DMF6hFFwylTce4rYQ+BIQlKp9cXBCX9vPkDOjEsEo4y7682i5S1+s5mrVA40
C2uFyYuIPfxECNoFHBW/CVFlCSCYhQ/kOUcNYb9WnjqtTkoZvPRV9Kq0EQWdS/kYHJGYZ60BEdct
gKmoll6cXYgaLfXukIFTRkmqSG9Qr5HYvFwOEkMcg9ZutVjskoiApZz69eCZHECgq21umuxUO7pZ
B9BKZvISiFfJgrZlHNGO8zjkdpwn+fJZyLwysEG4VAMBPQ3sYjo2BSH9ssJWo1klAemiT0givZGN
ptye5oWkQ6kYxvCCfLyE1OTUr9jQDVr5QJ7Ms3b1ESOvMAIi5iv9vpr7OIdgoZCbx1HFKX250I4o
pgejs2yeMdE1I9nntHkodgCWFU3vLqm/B+EKk9xtjBq/A4OMuIx+WuS0x0Rqriw2gtrgzX2sASft
4UBL+/yazR+9JfXguWYDVkc5Ov+C3LBON/92Z62z4HByCegsy5f172HPLk45oz/2MhgfIfbKjE2P
+Mi313jppXGMKChWBxtwICOz06rrj6+scZ3GsEuPMlo9E82wftr0IMl0uymBFP+IzTnp8oLHNHFH
iFLH1vlW1WLxdgdRsEgLiXpB0bC9/TM9EldrSHnXLbe1brMsYmnA9IP56uMl3deLHqjoBIwSr49t
b6jKXmFX+SVKgstbKU0J0H5WmyzEChV8+jIn/8wVh0bA2ADp/ZxUapcxkY+5jCyajldIMMUdQ73V
o+aB8fVJ2hcOZ22K3oldW9MeKFm6SKSKVqqUqLVFTvWkFVqt5/WnX7YgB3UXm2jUBz0D9ZtWIK/U
zWitd4sstMG20lB3Assm8P2WL/dBCS61QzZast8SJWtVayYRMusCzJJYD98gZhQhD6En6D0g4UYE
3tUc9cShbWSrbJd5hT6T2GUVJhTyTNYKYcmDvSRNX3wIi9njf4TLkYeblfSFtkmmUN8u5TNWzacv
nzgA+1IdQMRePCXWl4q7ppM4ijSVWWCXyZ90EXuaqiNB1MhjnRX2ugIUTEsFk4gZTeebwf2XLz01
nHz5qQeX76F7NIsvD2mJ/c81jqShlUF1g/9tuFpV95QoPQMtUkRoMrxljBLM57aNIl3GSdFfmKPX
pvCUmvKb29VNChkZZDvZwP2FzIT6G5fmBZjJyOipu/RLWpFtTJMVDdX/J69p/l/RXPTIGceBjAOu
mkCnhGCe/Lqk3pQrzrJ+e7+cSvKi6n23XikDm15l/h8qGXTZMahm5GIEtU15AAJXrugX720LNr7k
HX8aGuAQuSLzsz2AEH04S2sAuh1Z1sbL8v3NIC0mumZh0sAm3sxaX3kq81iB5YWtO+AG8hFQBFtg
bcFBKbCP1xXh9L+eSeYOAJu4A9cBiDhhRu3HCJlez66zqH1uPrPtRAprS3SBh9Wi9wKiDq/W8bYT
uWrD3Q7vKAHK+pkfNB2FmkABOyscUSI+0Xh06MUKCk0Px4fE3SpoHivAubuwCGmtUSXFXypB3rEJ
ksqe5xB0PV9Kj1fNtod3+6TKrD5QE7cW34IheqAMiDIfDPC68Bq99DtLNQeB/u2t3m/6h8RNAS5n
5LQTbwKnR/XV0VCa1+Hc7BIrp6s9gxrEjmR5/G1mxgX981jzXOlYs5ot0c5l6FjDXR2Q/zkSjeB6
NI1FeA+JosbfrLhyeutgg0SBG6d9Ke7urcvexLvti7l0me8s3f/5PSyTjBMRva7ZaipjH0ZTxoAS
IngnbQLPMNakT8CqqQiIGBi7bBlD/sBrPcLY9C6p3QX3/hlAxSr6WvwsX0pw0wqj+7RgFpNc9xKL
9FvED6jN7OBt+wEOYEaaXvu6ZwVIUSZhDEs8P8bjp+oAfPwZXG0mgkA2/8Y+YFbx1bcKmqcHy3NK
aM9b/MY16CKUMX1M+dG3whlFwTWDhXqWC6tRMN0LK1RkbkzYQYU4a6kG9Gh1SM5xqQVgjfk4tV8u
NQnrdfigWsy+fGK76505EoGJcsMd/azkuRIbvy6tuhKVwtgEeQG7EdAqFKecnBlZzd99aZwzCMvh
fcpFpG0GOqdi1j+ThtC+z/gJeOBp4BAPD+iXC/X+Pe2YlI0CsDb36+QxcQGrYYvN/MeeWeTBX2sw
TFG5MxUYfEiVzjO1s+vRXwsIBDmaAecmolVlhbjqCFZ1BEpJmAKBtpZFmS1Yw7/VR/IfPhwvcGEf
WXS/ZWA/o/ZFYlInMz0w4jQcKOKMo9fM00/2kvKugfSx10EpSGY4NevuPcC86p4r4mTXu0XnT2Hp
sPSjydoAF2SXmPFtPjTIRnYR+ZlosFmuVwg6jiFGF3f/tgbtw4RZAZtYUoeoSnBbUGXAczIZewDA
cXtNv7JkmZRqVbgqyNYMQFyGuC3Cnl4gChfNvBr6NDMSSC8OLwIWHbNCaFlGL1w54M4iykvyHUx7
sHi5mEBFVlRKCHLC5GQc8Ux1nuobtnCSBIIAmj3JARkwW4oDiGcOWgy9Tf4O5Eias+3vqw0Ye97D
pY5QVd92yLz4Yz1/uXug09T4Mw6HtzWhWIrMOlCmWjl3E/FWP5XbBQ2NTPS5ma4w6sa7lCrnRCQu
YIoA8IjDlGPJCdVAp+X3GmLSqeqVykJdqQbXrF4sWRi1VF+LVm9prPNNX975C6Z7ITrCV8oS9O9C
duZCBCmA4NkQTa8Ua80WDsVniD5/xfzpU8s+gHO1xhVnKjYsford61gnXyjTYSAh/+F2xOL8woFe
pPhBzRB+6hvBzS1YyBfNLl4L3TfXtUy1Bkwwf1H91zJ8dyR7SJMeo86S255oSUmZspAKnN2N85T6
B6IW5Tniu99qnG/ntedgXoabS2yCOOO3zlUfsiTUUcrj8b7im3xN5uVzcQrhZ9Z2r1B995GQdSmW
3zt4EYTV4tBIzskEVba6MsmyERBvQPTkfrC/8GJlUlMDL7TPjLojAVzo7Qo2bXko1IW4wXhXtV2p
ImnipOUYcvd9NBfQSNPhAtMq9oxMKfiFpo3YGMrX9x1xAsGyaDo6idHwFaH0ZtnY9xG4dfUm8pWx
Yn9oCGYSBk6GPmYTt3OfnBcy2G+XqaohotSu0ZKZy/rQdAEX1wgZC8S/06YC5mGK96fP8CtaD6rP
FaAnyYZyrXGAHg8hLIf9/mK7GcFSak1R3a/BdNKP5wqF+yNOzvdkAOza+szFyi+61Slxr6i6Pvh9
1+e9lNN1umBiuV9nTVA+NkPt14v3YWjc+2ob7mPuDSJisrfLyj8nncMQ0+hW8W6nH30KHXMYY9gA
CVX1NdwE4IMK8qBbXXGu29AUIM++dTMutdAdvR31ZLvk1NRfrZkOH3+T7Y87B2PDDPbduLv2fLi5
FZOFp+ofRei99Vv4FWpCLaTRMRso4WToiRjEbGUO9VakZqkAa0SKqGBwTIGzFrBy0eHxOybpRt1G
8J04WOO6jEzj1LYDlgtWW05K7389aBgeSIXGKN8qdzeel73CeS1+dZrBe6J23qkY7Wh20Vk4ExtY
QYHjljkYheO+dSh+VIZ5MGIi7D0PZjKDIlzgbxvpMjIdlPN6lXOJ0CkSzbQk6pi0gJH/NEBvrOFR
eN9y8ZU5nIzblilge4E76XXycTNRCVMzQta862U9w0UYbAk6h2g4A03p25Mkjl6Wt7jG5DlMUyUE
oepaB76PZx7onVDkLr4WOL5LHmEigrFBW4E8nFUlPnd0r/SkxQWUvm61XSXtbgfEVb6VvEmA1dYX
83NlnvwrRUvgi5ocKtLbbVs9eBRZBxIHpbT/M7NhEFfFmxM7TPCv8a7ngrkTRJi4STfAgTQnksvT
5Bj8zFKi9KmZUODTJJwqSYIGYsOZ7r4/n2+dYnuBRnXoUqeb1ZKyqaMn6Pq8m9b2LF/vKb6We2rJ
uESglIRGH1g1RTY2yW0kQSu9cSM6Xz6WQtftJH62XNaqPgw7j78E+ESn1L+qmL4U2kVZfkHYt8cn
PP3oqd6ACVeCB4Cnt6aVE1HcMIEVIuylEBybaw0txUMrt4GwdJGdmDeEDK5gGQEf0WsTq887hVRz
TrL9X/LqU21+7h+KsWXgztRRpP6CySf4Lfx6T3/9QZTAkux9o8HbYgqykIYijSMsAOLfr2PAcifs
VvuEibXXsR2JOFDcgV+zfsqRQIQ0xd/72FA53Qqfabpvzcu2AbH2M3AsTaB7/FjUqnywXu67kOWw
EB0t4RbY1guQg4e7rV4ocTJR4GsIUBEfQdIZ/42xNe5CZ7Yd6T8k8TFhBcuQJRlGuw+DpETd/YOU
yfzTXfYJeasEertaU5kQEVmo3YXJ7dH/qWFkC0xHG7tqKXRQMUbCjx+fxv93Oktsogp9PhiejzQc
4DHaoTVLY+Bd92g/or1ZpHxi2GQDfY6BY/MQGUf5fD/A8LMLiebUORm63pDl5oRoh15TkK3lvMyD
4WE32woQ12mlqYkXZGZhdY+RVy0abB90lPnzbrtK/2rkDYgrEjSeBShuWqW0LDw3ZS4P5SJ21RRQ
PoodQmtau0hEq1ulkDCwkeiXfTwYXEWhfDlEwJ+XszFOP4gZ8ZbA8G2FtuYbwYihKoFKXJdY2Odv
/6MkNJ8T77rOUQZH0I4spNOO72h7wWh9O4FhtHZx/cbqsnOCaSFYIEClLOkDB2zneNpAN9kYggcV
x48zqcYxv+scz6v9Q6h0f/cHisyF+9LT6seViiuREa9OYRQhIyWRXY71NiXacQVpNgH8cNyjXzSC
TmoJngG051QWMi9u5eYaLolJ/qH3JIjnUdUgh3+ra5LW/HaRdEnib6pWxsRO2J7KYcOpyi8JlJvz
TFMi/J3jXBcOkBVi3nUXo3taEVeAJXdWdFVwmwqodZYPkYo9WuRkPZiYYVeNVNkssjMM/6aY3+HW
yc6XKieiWZWSEWxJu5Rw6PTi8gtp3jWPHoLSHZd14okIdNeKTJZNznvyAN6Un5eqdPLx0FYjYhLU
9nqOO1D5uakFnLbDvv/qDxlF4qDQPHdDOAwQgCF+jCaJgeAja3y/hIxYhnYklGSjVpiypEpNtAen
ysloEkPI5U+pN9+rP/MGdWyc5RACxxZT3FUwq0PMV9hNhMBKFacRSZtE5Vyl3UkoBPHbdRL0UUwj
HOBIbyhE0ZnbDasg51zi0F8NbQA85NOffOo49WFNV0yjTcdWQsD7T0neEHugWsS/ggZaYqMMNynb
dNMvUcsCtHti4uHaK/vN1A2v9z6844iVxr/2TQ7+FqcXw6HAjtABBhLdvZTrqFG1Ype8PvTzg32F
DjfojZwokZoATVVVVjPf6AP0SPDh/0y0XXrp66w5koJf/Vbh8S9APSxN/8XCknpnCfs8rJ1b06kE
k1llnCezZmKlWgk4Zal4Mwtrrne9zMYs7kJRN38HLlCwmfsBCl6ggcdpBIWIWv71z7wGltKv2CNB
8rGp8Ef4YnP2DOV7XWpUibzYETbzyStUrFFNI77bMeg59clAS0Bfoosi3CZHu8Iy7uUAz/2wflPq
e7ESp3lgt6Z/cWIWSJ/8GSCYJdgM9MSJ0oETNanuIT4ob44Scdv1bsSVH3D9E9khn/EO5yxYbau9
cR1zuUcazT/NVD2h27fn4Nj3FKlY5m0WMEuLvsNAY9SD3zBjBtccw+2upPIy2oH4j8aKu2rwhPSY
C/lYAvbOASi7Q9jxuQyBY7lqhWkMt48ExQZGY6JVK5VE5lYa/Qg8aGOzKiovbZnu2b2N2lGPz3ku
IjEyNnMouGFNF+xrd7JPeuP+GhHvZ3Z184WVjOujgfo0mgK/uHK7BW5b7XalUA7m0PQiS4oUfIal
awmWmyEVajQYBAtMcniWWN6aWnyOoR/7n0N+B7uH0OC6M7Y3fmofxAU44LUCsYkZjTjcakBKhHQA
1W5uzkkfgYc8zIq3ioPa5Y71hkofN4tGy0BZZHPprJwzRGwDCbP5DCOKYJjX0IVRrgz8f8Vsq5XE
MQt07c2/fvuYg9os3+ExPj/oSBXhJH+GdZH2ifV7ahyZ54E8am0seDf8BceenpBHofawpVk/1osH
pkKjsTvX6Fqom7ke/gvd2nR4uwpWAVE99mylf6sxg314HRH8377s9ga8JBA1OvpBmTEvmWtkemk/
f63o58FPEH/nTmxrrQ+yYtDfypRMUtZf2jE805D2mEb+JSWI1d3HFvQB00Od79VZuol3IUoWZGvC
LsHax2bL3jJsnzo+8IXP3uQ2462SxB6iBLg0cdcGeC3C2seRU39PILKxLRRMBOHfp22odip+YusU
y8Et6P9ho58u/ueIx3XxqBCXz8FqX4IYmretKNnAkrUBgf84adOkqtprgpDWb2nSzu8HdY03k/5c
qdg+mHyoIkCJQEMeSAx9AGQpNqxgWBZxV2e2/gTBmkYJTaFQ3dz8h4prBQNa5aAyKZHtTtKOCVbH
by1uUAXLD6AQLr+UFT7bk9TiLMdJ9ZCRXUJNxAapxwm4OVaeBsIcbz5OszXkerXglt03fimgTbFk
q1JejQGFKeZIGC1gXZkLhsjbhXs0sqy1xrv5m/emrMujNygnnhKdJzr/qo1qXhZQPjOC4xZqctpH
vgp6WB58qNAUI+SVBoU5mOl0dgMsU32hiXHgUfbI2BjPvK+WlXjWpgzgeKnpkdTjZtl1YbFOeHmS
LzM7Sjp9oAQgFjpQsCoFYuqsGmY1OA5lTMvmd0+kZxA89mOeXdSu5ILqhY+ghCQzbqITgWGv8ZBJ
wqcx1HsqpHy95/y5XO1NBM2WWX4JxJcQVLcoo/bIw2tTwu79mgO6am6mJlWN9As/6/8cNZi1gPwb
9FPNjhO8ezhCG8foLOoTdPJd3XZzXf5dac4TcMjqDO3QldiFcY9VljBDTvMHEmd9+8P3uJudju3B
zgFdjxPR1WY9TZTMYcS3X/5zNLiLz7uMcopUnwf/4/QeLjlMlAAoIXBNN9yY2ROYDOcd3oZvn5u9
s4Tt8e7vL01R9JmXSFwdqZmC7tutS55NYxQkY+xTpUVSAxIo2d8ddJaSp6GHG+kbsJEto/Re3H5m
ShaQiGYIyHOyvWUB83pqnYwsxhOwd4jW6C+ayLPC+ylfUsTEpzBnanJX/e5AtpJ1x9OEnaEk0Lb6
tBuS+tLut5vGQRdSGFM1F9lQ5Vbc1RdHQ6EcKTicd6NfdhfylDmPFoVmyfTNAGZDhxlYOU791mg4
83qsO8PSPdulR+opvB5rnNR6qv07kDGb30+efTYWLpthe6TovmIjroYsJoNyCWPepE4K+heiaHnt
A1hOQ263PnFDAw5ELW1h8lk+MBDWZ3xXvTP9FJZ3VkiSFNthtYy/g3uzfu5NY4qjZ+idSx2FuGFu
Skde1kNxj8tD8o/yMp2eZDVxs2rwU0/kYNMlwzlLPsa4EzRT7zTH399YNZnGtoIk1rdQuAxddXG8
J4y+kt+sXHIbc5LReJPG0LDXp5OhiwY4twIYDUyB8Oxbqoh2wOuHVsTe+X2JEzdJHc6ZvE/Wwwoh
BMD2j003AB8zwyVYeiS8Pv8hH2vE2EuThTj/HqCjjGGNyIr5JPB4sVLg0oMX5ImqZZVJw0Tqp5PH
Z16Si6W5q/Q47nu+5467m2Ac1t3xqdUo3hvRw6krKo3tVLOsj+Oo/yzZPbvwwnyntWGvHQ/Ei/Ow
MG6z3giRvEhrxtPG+74Bco3wDE40U044yU1PR1nyS3Nh7yq4ZD2MXPaV/lFjANhnefLR3S6D0szN
cG842Bvob4TsQHxFQZQ7AS/UQHrfMK7SvSVMM/F1cp3eqVpERORnb5I1ZT8oo8H3VylKSgoysuox
xW7pG4PRbnxvFrKzgUjmMsFHT/R0pXEw5iY0ScPATWK5aHRlum8KWJfyCy90cI5GtwJLBHFcmNJS
uQxkq00KTxnNyPV5DjxBR7gEjPay0hVjjZijvJd3/yYL8PBVOPrgE5btKIduqIWv4GMzwiLGoB2V
+sJH2gKGx5DBVIxXiyozAQytJjzw+dX/dZvQYl9SerKKNA3UQEQ8Dh0zIn8FGdMXSc8Evjp/+Jb+
f6QQMKgGLFVuqb9K0H+nWBJoVfH5un3MsU4JEEeDvZ25yw+wXq2IvBpb6L8LOB43eAxMLzYDzqAF
v361DZmAv94iDCdHJ0AKWZHfQAMI2ZTQ4PzpYowF9XD2bE6IQ28gdanjtp/cSBKF1hAp0KJjXll9
9IRyPf03QNei5mljeNT9dv9p4+XajYqbpMyf+9Gg/tb65C0oe2+Ik98BRmNNiGlvZ4Zc2aRaG6wH
8o9dXvDnpIrqpe3q+c4/t/SsJG6fiSrA94mIjVTn8YpjJsi7SEa7mMFjXWNWgzcBAWhxW1FW0GPn
RnwgQmk/DaB+gqFZEev7biu2dnN8QOxQSPfGA5uEQjumiA7RvuUyGP4TVmCzzvnGmnfB3jUXARXb
fsnwOChQ31m5OVfP9dJkBm6sGYKXfX+j3MRhGkWYSQSUi972PukW/FR6WQsMK+60xJls2zQ+1Gtp
q+AaIxP2fOFKFk/FZLCozuJ4N2K1KPXaVT4EqBrlVKylbEUmZGi7c2wY0gVAX/XF+3kmlvI3TvZw
ePUENwyVyQM18ytNX9cCc14qb8XOb7Bwzx9cUwdqOcvoJBaH040YZftTi3Xq61PUzoW9pxiEzUsf
UAUhdcDO0sHxmaOPIJ14g7mWkXjdnMlmMaYCbOFuYzr0RUKf5bkCOUvYiXAiOf7ybOOWA/aZLrji
D4gZY/Q4CcEYyxUimVezgRLNGoO2jZOWGujL9WrxnFsDyEwAlZUc58wi5WfIEmbBx7ytHMZOjeLV
L3+ALOZMGcERb1O1aFWhQszyW/NEHQXRTC21BILbFzKYdFXhBcRtqfDoOvijbOpwxeVBZ0rVkPA5
GZujhBj4g0iKKizCLXLI8HiUPT1GZxbqQRCYggEFcdgIxdOY/ifNZ2wL5RGmAfbB7p9YGr3ArOW9
qxI+8iAgt5taufkkfzAqg5TXL5jNqvD03sIK4rPCrPCRfINXjQsBZL4tbLHcQbLYR0S4g+SdZ5wb
/7Y6lcSEarvoUEWLf4DNa20e1jpWqePH+Kky748kHMOSCqBfgkV/+iYXcOGYrh11cVflhE9H1IAE
S1Lqi51HRmpZQBESBrf0IONOcSS35uZAcxtHNoa1erEOkQ/qqhGyJYwc3atDx+wyD8o/LPSNpyas
72LCHDs+7Fe3EvRUMueCLg43Yfq8WyCMhqzorjEJMFyYvWBvAJw8ONnV11RbdRQWbf/AZA97sPxf
qKKNz5rtJqwOyAP0S75nk4BS4VIqAuC0uBSkdC3aA9U2JkCJjmq1/4V04eXN2DTR9UIKO6/MDyg1
Lj+rfv4SAK2sheGJi1KTiptpTybL7oWJqFWoCPIh4zFN5N3q+moa2Nw/o/YhxGw9PS9hAlaKEbjJ
GGC+/eNzfiIlIwzGYEkoTeQIt7KOoAdVkQfds+sUk2MYJKZvP8XK9cfMLCOJtpn8438eLOTCvw5s
RmhESoH1OVz0PO3wIoCEvA6WuxzJUGBkscmiL9tG06DbN3Z2ORuYS0fbiQ5ZEzFhidSXyDNRoj+m
PI8+LKurrG0oGMnNa0j7rdi1fPGYgoRLZ08w1C/w/1Qk48pRHDnArAAN5xvemv0oACH8GWCWBnMr
5b/Qz/ZL7oTdPWMC3i3/MwhHWB79PVeyKAMLd6Hy63Vz5t3txozBGjgnF3ictPp7itLlXdDcV0Is
j8hlUYm2TOeJrB0UQhVErFzgdLgwCFbW6V/yYxxtbonv2/DRZyfiQvbQvM4gKIvfSmNVxgPuPuGe
eyAIr5bw/FuCXpwLQwyPp28q4Jkv3BsXs1iK4BfpDcI8tD04mD5myjIC3adKn6dy7aE0mqEoM28+
SXWGH7qovKQddMAZrB31U+AbCcNtANXFhTNVdnPg8sNxawHialQVh2m45FDsdgRYXFjNAyb4GFdz
Bpop4xYTWyGLItZBRDHIq4OCTDVTuP4fBNFrhujjRM1nmdyUqJg1s0fgrlA7tG7qsIwCsCiLd/YN
UB527kggbsf1eIC1iTey6YVOx2KY/uTzIWvslkzQ8Pqzxdyfu8FWKFli488HF+Q4wKP+oMgT/bfs
FM7svMmZ+iALNR0Q4PQAXU1jKYweiGrA6hjq8HiIslNaMcfygv0OXvSkSVQ7jM1Rn9HklIMb3jd0
7x8enLrQHSApAxoTC6rdE80TpWxkufipXcM5YMm/QrVRIYnrmEvUb2tge394hs0vWopNOF3cxp2h
siUG3/uL9PjnoUhcUj005EbIs+hBAuiNwBG5BUmOsD8psBTNEFypLs5DouXFmu7aRFaoTRpaZa2+
OridiVb6bgDY0btjA1CNP43k0N6IMcQqW1SvLdwRGYZcV6vgmsKYm61OD8+weN6tBUqi7v3hRew5
1jpVREEtw0B4sNCTFQq/8d3k0DxrjvZvgzY2NhPBMMlqI4Ir6wHvuwu+H40L2bSGG9PhN/ot3fF5
tkA0/AS+RmseIAExvrTe/KFxOlmRsotVoxfYOZn1FJ305XBedGrxhix9TBNcj53e0GsuwcJu5Qyu
9REzaC95OXkdFznaJHikQHRjFcHFj74DVFP1jEnG+Uk1s22TZMWRyywErAYbLS/ebB4vEG4UkMaH
yG/wALNcMfa7q61Vct3GSFtDXHfi7vdE5amE350KT01/CDqHNePTNTVW2C+X6w5/kdL6/TR7mD3I
jhKhlv8FF+5IK74p9Y1bi5yrpPrU8qX5YGPj3J+XuLrG+a0fqJ47XaMAjiNqFNz0o8M+6RNragZ+
PT7X8I0pRE8W8029qY1NJ+fEhf0ou8DUh/J/9y8TNMVH2VXvlk/HT77vFmcEq0K1B5ita4st6Ej0
83wluMWX3j+OWUxIWIHi2YTBVEAZWtvB+VF5+SBTFuXSQH8A3QlTdw0Z+GnWTLWYFvBMzWT7UkMd
RUmxE+7Of/AEwOPDc4VwYXwmFCrAuX6wZi9lgm2ZaYNyXiQKlB1IYJAAldRgmKyx67rY9y8sYUnz
WIbYcS0GhcrHeAOwFYWDyb2G07GEZt64jgiaefB7Qy7UbDArtmi4m0pO7ij+XaEW8jPcuBxWTDt7
usv2qLper6jY1bquTCOGQTjQxsarwxu7PoSHvLc0JlyrI126OPgk1EiJtaPkuzACduiF5OyEhehu
7RyxAwmg/yBAJEDuzpvXV+5pfp4TC2TxqndhMV0IDxp77pAm3V9LdUzD8E3F3Z10YXN9nC4sXRUB
c8dmZqoJHJavxJjPkgI6TiGbmPqgCe0w9sejJGMnc1xkmX9Wb61k4weEEYIfrQPVte7Qfjh8w/qm
9oVDR3qQtZy9Lf+OJoUwZH1cLUaO8R3GPVAUKH7yBZFQRgtO06PZZ6cLETfkBSWlOGNOD8Y23uNG
kEnbv0D5SdJGigtWExjd8yn0ft0TktWp4dE+smcs1R4ErfYJYcRLt4ykrNfWgx/W/1Sshk3vc1kE
M9vIDtr1uFfX6KzoF0uepEsJpa0Ipnixj7TB1DX0yfsy4wjmBK6ApNBSAojJpUKSioD+H7k2bMdD
nGvb0kICCQIuKpVKM4DxgudoDmrAK1PHMh3gB0zUrpjvQZOMuveN4Uuku80zrpsOYyDFD1nnfTER
cUKLBRdDxPuuuYwwW7QdP3BTezUHEwiC/xg8i2AlROqeGI8J6L77dznllPqe92ViNSuiaG8HrHp5
wXAXBkJ8UMSkzIZ32cZdJP7fXPR0DL1mnlh+nPKeDOQM37N9w1VkJilnwAYdlnvtxFwWNy6bKx+0
bJgIht5vOl1phKzaUyK0JsG9UaGRwRluPuWgqF50wkSrf3S/sCLRnSo2ognVODtM0U1DPrAD9piZ
XNAmV4cnEfiIFDZNBAQRQQO/UqhcMHYRHakqzHS5Er/wsgwLD5JjosyzGQRzPEjEeVVGqTyi3/RG
c0KbrfiExWDN3pLHPuuz+e/fVHWIW8PoJpYvepje3QE35p2PyCEEz4BKy161V0ztVPx5hRsX3zoQ
0ReJd8ZUsavWRv9mmt4Xv/ONIuLrDG4DKsiEv0UahrS+sg3SBNEE/OI7bXEhnxwNHc0XNuAPqLrg
rpXgd9QbOpth06ibI+sJ6VVdKbR99GdOWrEJwKC8nfKEaiXt8/aoQJqWevsZGpi4LjKVsyIz+6mp
touhFSQSPSkq7Ilmhvhhd8IaWAdHKLK8gi9bsHF11kI+Y9AlVZoAfHMk9xm4ka5Yt1/2ys3eAnPq
muUJHamMyJSx9nR4Hlgd747J6Z3ILs2ugn7AtfeuBCXJ4fxDhcwxmNgZW6195Es4kr4qYw6zzR5S
PcOe5MDL5mhIB1ObkskI2c8l7CCdfKI1A0dIflcZnLwYM3FsP/hoE6EBB2X5iRUTKxwuXHM0otb9
PwSr0CR4oS9BOXRHTiLMf1g832JDwpZXVLIeMY0hh8wc4eC2qZZhdvaqEJXJdvQtyBrxy0+q1xPa
Mrw4t7OIJvIfulNMzpQ1SOrLm/4YgUtG/vzJymS4pK3rXXYai9J54tYCuNalVmaNz8DewxYYBywj
+QYg8xVUmFAW/LKxaGgNMzRr5b4VChQkOjZXEUvMs7O58yJtf6EdbG3N698cQTXoE4tnD9mzQ8au
UpgpgSnuMO2l4KVRw1fWdWXehER9+hn0lx2qq0js2yM6KMOgtu6pNErdKMCXMfXrbCn0fptNTd2L
pyw06GTNar456HetyAfh/Xi6ajsZKixw4KEaJSPzDBQRuFXEIpGPjY+41NC12/DuazfX7DVi+AS1
rfixSeVB3qPpa7CoaRexO5Jwhoj/smnLB2SQaNiIEEjZDQKj6HoOTtnUDCyCBhqxH+JhsbkOcT2w
j0e1XvPVV6ugwWTl+tkv6xYRh7+6OPILT940F7jW1mIKK3+YZniLr6beFksC+A6RTUA/54bDwxDF
1LCAQL07ZxuAFOnhx4zhbeLJEPLoG7xyoiweqLVp20CSVRWaALXMuUt43q5ocxEX7Yu5QhvzjcTM
zAaLhZvE3afGENJeZysGZXWwMAveDyvndYLkf59AD7TNgcvfqQcehag6dCx+6r2beoP1b4c+7GUB
z4OUlPV/6QkeXTdTJv1QfXof79XpB7lnwigAuAtxs9c1wRqUMqbYdQSkZykT2/5uyet4qGHtu+M1
LMl2teEwwQ8boPLrMmNDDgp8rur3rGnTtRn+F8gDbvNzR4rE/nMxsxeR1IIQfZlCkHwD2Lzmti4x
36+i0QMUqOVaSGFCR5CDF+r0hZqFWXBAKyKirC9vFSBpE6S8wjdGar83QDsn6pazdcqRnlxtaMIV
fcknmkCEf3qAeCfpXn4eJg9PK4U+Li6aKRINGCmfAZ5Y5HmfduysonYQXkvxSlQJGFb+n3N/VCUz
rowqybFFzxE5djsEU4yQg9ewz7oTdNaSgMqrMerADMFhATYm7irHddfHpceoSdXXmYViG4IsWy5E
0VAOTvDkDMBcNWX0N2Dnyf34WWzTixKPArPR44AKKKMDlkWxRUmvzDCYNWnYTgVSqgMwJVViwkbQ
qPaI4xQt4/BPI5UlJ0gTRTSqf6L0jsHOCNwNnn0Y5PtrVR1EZ5Dhc59CsIKGlNTBLAmH43C9f2ND
zeSAmfLcBE1ROu72NOdg37whdYpo+Y9Or0+5g9653QolfAGPJfjDij7xc8+GFrViL79tiwLKGJts
qC+MOECBgK7MAmA/MV0Ap2LBzUum1wokZQPiln7/YMBD5FtjLB2m3ppJQE56J7mqpmzlYm4+AbVC
d0Kz4VkQSGsJcRSqBZx59dhgdOd21d3J3uZy4D0LiIZ9vmF/zc9t75xF84j0WzAdJszMe9p/iEMO
fq3Lcji6Hns3JkDDQEOdbpw6rFgSL3d1jujszLsCfpZCJuSgI+8F75Q56hS8CXKJmj7AK8/zQg6C
Ijw3PUW9PQ/9WY+bEBTXzyRuqgJrukHEokagZpzn2SFGe+oeruA38uS1F+x3orHAYESaaeF2YA1C
kIfrNNHcQ97cqte59WZiUAVwGyu06xqW0g3b8iOhEPDZxQWYp1CQMdLnFyaVFqTKZE5WxQtogK/6
J29pc9Rr9m65PYmR/5eBB+yTiQ9v2BIglLxxZNoNrQ85M7iCG3kJAw8LIhowbd77XqRo+IkJQ1Sp
4IB4vFpwHL4bWBjlcrd21RgCnFq/dL/Id0iVFf8i9O3g31exPGITK1pG2fDBHvj6wSpgbhklZ5Fl
rkhV3rXGFkhFD2O7FO+OeGMyXWTDw+iLfYmJep7nqeOWQrMv/t+jcFYmEJVQWgyS5KXyTqIZ6yEF
+95ZWPJk4bAWkpRxsFhqFU34ag74G0NAycozJGfz/GTJ6l9SYL/0RKE+axKbFH2g8rzbWuP8NMIA
0N4/pfNEehchOImi6DlW85qtN6y2my2S/oJf26pgtWckXCo+1Rawb3RoDkvoMCnPjFjhByRcsjpD
YxX8LlikL7kZ3sAxdr/DpwTDVOoPtPV0EXtNFFlWp0TN8txl2SElpvJvh4IhKXEK9c+fpBlov5vL
VwNFdCI8giJAPmVjaMnHr93uR5OzhSQOBQ0oaatFyKvdgAoVsapLOeKqvXlw2auje90X7qA+gseK
NnjP7TOCNPv7BV7MfbdZ45FLRAgc580G+z6xzTNR2JRS5BrqcSml1wufF6h6Zox4m/TWR7Y3R6bv
DfO4jJdCsbgYcRI3ETq0rEyPoyhgPDny7rIN87Cu0+DoKJEofpaL1AYHzFke8u4iDvDrGBY02++G
le8e4IOnO2ZgJ3UEuYZ8rcJsuLSMSR69/J/Mus1Os189fomJ5jvxMcizWOyl26NaqQy0xtfJ3JBw
54CBDPQ89HmEVtm/PU6QUUsbg6NN2cZ7/DMb4APqCn8W/IXqAJX0u8ab7Bsv+hAa1KS3ILjym6lb
rMX25QyT8f8fBJ1YhYZvmSRXNmXGQJCUZHkwGUATsZX7XvRD9DZluR+JnYIRcJJiwviq40WunQqR
e5LZYrWEpmfXY8LSRvlBGZIILNcMLq1yz6Pm9GASvnzX49JCQNmYlwXRDqpzQshFwEA+jO9MArxm
+x3mRYeIKxUYPqGRF5AuYTyXm6TdqoCA5voFJTv577Mveid1SbMlvLIziTi9/YkqVcOl+UrtWJU1
KZRAY3MeIVfdFmRxNP5DqCkVSuiwvj0/Drn9CcGC2RU6dJLO/qNxTIKaEamsdiC9zT3US65BrMMv
F1HVGz0Zx1tHwBDeNJ//1rP4JCmqxoV6OHpt1pv/EjBtTlH5KvYC42zPGBAXKdv7ZIcURy4+ZuHW
WT9MSYyEVlXgUV+KbJFRWLxvJKXtUqbOoAJG4n9vmcupj4uNoDJ6R9O4aO32BPFQoonuL13E+T1x
wBZ/HpF8tW8hS8TcQ1ZimLlMFhMEY0j75nZ1BVQXaEZhM/yNRuxBDKwRMi0vv/yy2JX1L1IOD5er
LjtN1DjjmvuFQym0zfJOpU8eLOSXchOGP0JdpR2HHIYJzwVHcwW+boK4qgPZMJl+jZgrkq0Mkbts
sZAFvMO4XaudywoYe0BME+e/FK0f2smGif7Q5I/wuhHQ0urbTUqe7zbb5SYK3EMK9t3tzPzZkj1f
DkGCWZYXYjuZPXby3ESEPilpccX6fTU3TBr+tbNvXBc9Q2i+QwXTWoO1541hPJLbcLOniAydDXfm
keRinAVX1THcwNv+Nfbi1FUe9ajav6KW4ClcsWSNjj4nEZNfnqX9/jTH7aeuLo5fF3xMZjWf76E6
TAsqGZSmp89Q72uo6P0aTd13WAaxcUdqEc9AEvSsgXiZEwxYTLK5hEdVR/WvzbZkaMj6xy2z/zW2
PeJpTjYvQDhobYGI0rStEQ5z34gCVvmmaSvxsqSwxeDLxRw190Esvlta4a/WBId+AxhUF6TTMo1u
UvlMQit8DyX0CyXTympyax08sG5yRYL1j59aXYBlJouwU9cPL3hHwujqRzRPJoMC6kwcLnjxh/wU
nRcX04vNejgr8zCnOVx58yjAGjLO4XY0FtXAMqJQ5486Yosd03YBtXK2IMQIGxjQHdYHOvI0Vlpy
n4vyVPwEZ6+KbzJgndMee/mmQ5XFVNzoj829v4DAAPo+ONji5edULis3PnSgsWP2jMd0g6oMOfrQ
f0TaDjahBsqRyA6M5X/1wLlQTjCq3rowE5UZz+gw4IDBYaGJB8ynTGLUZEgd+2En6Rf4HKeP+UKt
RFSYXsL6Yz4YLA5eC8sOIZS1E2dg7BRQmbv6fhgqc9fNUaUfrJKteaA8aqYrA9DAP0fwAqCRrrLH
yUFKYPOjJXxWr7UPyW+FZ9P640KfD4+rTQ/UvM2wBNwoPqFQ7+xacnOhOXOa8F4CoslB4VzxxX2g
8EKsTBa+9cYl7RIbfHVKLihJ/aTgAsf0g9dla+p0Z880Xsgr4AxpkhkI2B41lVIWwQdZ1unJonas
a/BA94x9SSDFh0NS9H9zL+uzt5CKlFiTtv4qIjRp787tDUWMBd/wX7Lwy02zjK0X/itxBaCNLdh6
Y8SpR7o4EMfVmyqnJhACaMuo7A2Pf8ryxXHZ7mLW0OfAdrcaUUFc150RRmTaV/rw4ewtxUMq9sII
Ji7ttLcQnjKiMTTsr2mPBUXIoqXcj03CMsLhbEcc8n1hOL0bVwdzMzRQZv3jCWeBn50QxE84kCJS
irrNLp2Zh8JcE3Q6Mg0llHtYCFh24RbPmFFIp+Qns6Y8+mIXisYv3kcZG229dGaZYTHiB3hlNCMM
cDrvKI6cUzh/LBMq/q6NeFDubHHbg/aevtsPOCJh9L3R/ZfF2NWjW/xlH/A4SnUwjzb5Z7uZstZw
zqrgbFr60L51Oytd32FGUZj6x/4+gMIL9fDeWmEjLkqvI7xK7PidB5mLf/+qIbISP7V7HnVKgXi2
kYIab4dePVtECyhKyzsbZZF0Y3cUZKllvQJVfzAZ6M/SiBWg+CGgHR+Ivv52jbooWk7qpYJaV9zB
wWxTJPZbGK3jjKw4RtepXtrqX0tbxD9uYC7C/snBpeh19aBAukdDoy0P65JZsxdVqE53PyvulcQz
LQn247UHjcXZh9JaqbjHcVM8EL9/diu+Wpn9jofY60cIX2LbWBmL4oAkA37zKBXNr1QIvgfPaUSo
kuI0RgiLh887gNV8ztXHoLnTSG5QcANYZhEChpRatTlVIQPUhWSTWIjOlo5cZenpl3zSqTJyZ3Xq
OcoJ/t93jCB7Zxe98arcnCWcDMjOS2X+GNLSdWdCB3KpsEIh22BIMo/BmjfNq/LrFxBXXD4jSBRP
vTKyLgfC0J9tYwbEpytroERMR17eZyH7SMvkb8hmL70PdfMkYXXhgRUKACxG7BjLRB4aetYLy1TD
rW1DTYMcPO/ps+Oam7Dr7AXZdDPSjk8FcZ+sX6NWCmyOdxv9gmfvSQ+OFsa0ndu521RaxE7xqEz9
nx2eByCWDy6/neESx0KOENL4r1KuSMbni79KqMz/LJqMP+9lqDCAmZalBkvL9lcT8FU5WbYX4u7M
txmQ9FNOgGlp+ykwqrWvdTLxgUxZkC25pRzVfgfIQZbHyP7olOGGBXblB22UcRsYd4pBw/CIU77M
fUWec64v740/1mYPldKZ3DF43IY30PYey8lpGDeXaO8e2XOzR1EAjxjw/xVpzGWWbVoQyE/H4Myr
T8KTmRExAQkId1Oznl/WOSD/97LtWKLH2/eC1aF6FdR88JgjfFTkAu0x5cDZm1855UOhYw3Q0D2F
wdxwtb7fO8kQaHwAfJq9hSc/ZZE8oCJH7ZorF98xpHDdZYhJTVc2KpRoKY4xMWtA88xfEazey1Vv
Xfd3HAFAxXzt6jPV4Feo3WE+LSDb3cbMLB1P0YcLL3gCaDx54yTVmFR8AZigAQqxpf6U45CSGPxl
9UgaxFiH2Vu7ibdlRkU0qR2q7PZiVtRH7jnfN9n1nqviMfK2dk73o1sXdaNdSBDqNrMVv/20nhIh
99+8T3eExMdhQjEOoWN0xMaNFRm/EKl4syfQE1XfcynuLVdMdrMqMrTJa6QuPLAMCJuoD2EDW3pR
/85ZrI3LhKOCJHVB3vPd1YK8mtSsGkwz/lKdMMzTghVv4OWqoLEo06Yr8mRg0gTTT0S1Hl/AbDbr
B58iXJ2hUP/HQ98x+h8p6ix6uMUfSxaBKdwvebVY8fTQMfZQLqyvFlUmLIxGSF5XxEeWSv5Ae5t1
enc2xprvFvsuVC1AVixUvgDiGVQnaFoZBp/M6STeiy3bSjh2u3Dn7b4XTekuPbHLo65bq9oOc78m
8XFsH5DOrOEeEX34R2UicvCdKx6wM+vXPds+2KuLN6csT3i+ci4s7Q9ZJn55ZMbs9Et4KHA8cfkC
TfMySnWiqcpLLQjfA6TKihdWYP77IegucxmwMFEDJwrfEIQCtZn+tl4MBVFQwfKGRYA6k29rpUBF
jGsCzEZJtRMXgN+vUeRQs0ijBzLMM1Zli/1hhYV6xWUgi+3fQGNsd7uSHJy5EbI8Rowv0oWGMiIZ
d1hVOspTVkQcgJaD49hlDE+URuc17P882jk39R1sPnQFwqqTkbLL4JJdwART1XxHpqdGWpd+bZH2
dZLzWv2tqg+rHpY9lal+Eu08j73IQK6yiHlaKQgMGziMRDgkIFtrYL1fLZhDmAuR1lTvZY26SjNQ
j56ZIc8PwZqeifFLU8x04LcWKBUITPaf0DjZ0qCpQBpav/PH58CoUebSKYTDWouhi0Bp7kpT5Vnn
IVhFiFpjGd8udtRPeOZuU/+axB5JTpub6M568NUeDF30X1VHuUe/omG2mj9vRNuOJAYx7e7htL/+
R58U5m0w1slVgCVWtScz+YjbdYVjPhJS7vdiGldkCjWVcTPP12UBFdTYmv8HhWZzegjn/+jBFXeN
+kiifAZ2SN76/hK9XPR73KTwlvP5knfXyApOBsZlvKeETIHM6kAh50VCrAJ65yqVWdjY9MQwHidc
J0YWwDiBk3Qda0JZLLljj79dkG3fZQlT2aqEIAEJ1NGKpl5iJLjAjZOeZab06kmASiLM4CS8wO4W
5ubHJyezx7DHPmZppbOuUjAvE7T+hPcPrHRNpEicqUrWRgkDFlXnjNsDkXNvFkaxkV8jRstHqhgg
/EdJvq69hiK1wpD8DYhcxmg4DrQdFgpuNSrChnYakgioCM5cbaY6Y1GZV6NMqRg3DajgncXgY8BM
bmQ+zCiHsmqe/BbHUMI0l9ajE5sVK9JKg7RtKnG5omo1aRrpml3IrEWUJaArCX4Ewf7i8J9Tgqkt
ZGqVoq6K2IIsmpDfq4h8cUoZjmiZWc2RaboVwmaw1WeJGIxEKMZu5nRaQ+lq2UQ5i1UBgdJQs+wC
fLqv8ucEXCcZzn1diWgu5LAK3V1AJUe+MDSRWeiBScSzgtOg3HeoQldCgIz28cdZktB/xJdXSp+f
nDanq6DTJ6DZ5f8fT2pC37mfiUycWbYNniweW9l86gmav5V0YFfkKrz/QbYiCtw9dBn6rW31OrWg
bpAe2+VQrQXbkYEbgyBLP73q8jiVEL2/bqC70hmQgoMdU2Tz3eftK4/GGmo8sd6jdh/cKnWDKl4p
zhKd6PW7O2c5Xty0h7B/s2ry7z/tseSJgMvzXt7ibHAMFJJl3hHWEtUETJpVBv4ClvAW3/bDnj82
S3f1Ew8tT28Yfu77LY0TaPJbmI6qLV50O9RAij7CIWCIMifWpfOFxQkvWYHJXfSE+iOGJyOKOhj3
QWs64WGRkaoDFiHZe70rUvzP4YDM/RfkJWazfrd+8kgtYwKYeDZjzZ8WwRQ4pwo2Gavfj8l4YT3f
/x4gBykFhivU3BxJkBIiwEX6wG8MtODhq+cI+J7yaG0Oq+zGqbd1MzylhGWxz3YBL188G2S7rJ89
l/FzAxnOFgW34Zr4FLqgnfcnfQyKea3CJlhQkdiRTAusjaW8X9QRcdXaPcpUqaMPPQ6G371ximPR
Q4+YA3fjeoKMp2D3iZnGnI487Cj1ES7ZRjy2urJ7gz3g+lD58/CepyzFTKAbtwA/eZQVgcVFRerp
0Nr8gMgLstte4GyclP4Uo6yWl8WYC6LSwWkdPobGvFVwD3sPnvcT3+wrT7PPaEsK7ZbxS0nbt1ra
5cy5NMHRb4dTUP6S4tm6i/0snqqc4oBYP+qzSRjwCzEulKovAWuKAGRl1E6PZjk3vQtDlRmpsbE8
W6GQQYDSi2ATvculUs98XZ57rlN9Uy3SSfGbg7CDnQtbBc2NW2EA869PHf1KrApxfso445f1dpDZ
5AjcovXosHCfXLI4uHzJFi0XGbc2/AOJDHMMzVnV5KtRJFjnzXQY1s7rrVBm2f0BX625CXUSol+G
Rgj0d7kUNlwTIMTC37steaTH7MG50DjBWsEeWe+b63ULVfftSuM+hAlfPv88GKg1AvzE4SyySSRA
sNZjnS/UpxV3g5WOmBLv9ky8ADXPAFpQ9g2JGdfyEH36Jwwuh4iSuTjbySQ0rTcdbw+phL4x/0sd
oiuuOM2276o0xd1DmhaalngR1KYh9wZZKJ2fWhS1cyxcx8hCJKHkyNUh86sgPt7K8u2dJUBcszK5
2ONgwT6l64g/HcWhykPH1TwNa6PE1c7TEq6mZlnTIFd4dpF5vfTQ8EwDuQN6UwxkLKR127IgmZYZ
HDkIYBANdj3IdUFnl3+9g6VPyYUgKxFmj406cjcOHwMp7dyx9VVNuTOmgJXtiN5FWgLo3ONbpUMU
yjstFjP3Qb/I467q4giSDjD3xQklRGSrJ6m0h5nV/GXL+ou4lGCovF3NZd7oNNG0aMgRh6SsB+Sl
oHVLhQThc/adxPeznOhWhgTMyFOADx2pwAGytuXoQB3qElqakuEOKQOddQ6ChstNHQyVEoKA3U28
vVeuQJO02HyaCpdE+FPWKLjA+jzdHf1qpNdBV4FBKTVXvRf/Rwmz4Fh/mr1klpcXCepoUt3GZY6g
rpq1BICm0VYOxHcUWgHVJtxgKm6bjF7+1/RxHlgzbjXDRWel1e9YL9gkgDnj6jDjEImtQp1VL3O0
OvqYjMTYD6OZQKSDOZb1cCrBnclBCC8tP7MvYnS19UX/3Xm+in+gmrms0ES+G1N0kAvNyGLKARGT
iSkJS/pr97LTzd8jU+8efuiwHWJnJ+LxZm5mI0sp4EMQcIhVp4ayiNV7/4kTfPTSBpaNhlBrRrqQ
7HgKTy4geUNw6QCKnvFQ/thjMLulSs94BEcpdlBMEhiqWXq/WMme6Umv8ZdwNGmVx6oyVhv1ckyk
s1O6Jxde1QlhzAM0Bz3dujuhTaELAHcpxlOVoNUI6rziRUrg/oBhZQwflq6FKG2nAG8H5bKLlLwb
YDnCek9Y2/JRJE0cPw34b3SyRYaFvzfCb3GGrvMRM2u+SUWtozTCMPyaLJU0BwWoHjZd9jx2GymZ
97qY4ZF0eg428W5EsPpqcvfpOTfQEwxSeZXQ5HIgP63PcTALaZvfwA7LE73HMs7yWUa3TkrnEwoQ
UVQSg0yODT8QRHdn3/34jJo/g8pPkETPhzpXHWZoBlEerOuHOnFXCe+TXJOwERdwAVR2S2BjADq/
ISzoBDolt5oCLavFsJJFpdQX8nGGmaoZiTm3sKtvqGTDfjDNO9lyDOmqdkHTrs2s0LVV87ucvtZo
YmbiH36gn3tD+Zwzulrt7eDArL4QOuSq2Fvs6uChKy7ZWyrFXFztQ54oJRhX+zSs0pKXVAql83hu
VUYb658i0oLFMUgJ+6MK43R6WE7RtMYA/so02n8w66WSqX6NDPwmN6eR5S/6YZ/6S2u5Efae/wHE
VaJOCyga6cslRbfMd44QAChGaIyvcrRHetwwSaO1MzGU1dnlY0VrNGyDpgVqipjjAoUBkR63uHyk
Xm+f89c5x/tfxuiMcsOxQbyufgo1Ou6nV7llNhkRAesD4m2ysSpXNow7MysJ626ON8IuYDGIdu5s
1okFPaNNNSikIBKSih++l5+UZxm98KY2n6UCKxLHwABen2u3kRkJ6gk45TpanKCgfXtUhQn7WhD9
UkD4rXChg8kxUiSHP1zxK11ptdl3VFozim+fuB06liDvH5vCf4rwSZEt+MwyzWNl5Q28ilrK6uvi
wPM0jVombQtd5ZX6G/1mR6RMYOZIqbpN1Byx640w4bQ6pxG9CSC+ZxCjcZZcLaHqJHT74tYanysT
r7i9hk0Y0OEKQgUVlIY3c31d7fzabF0jVl9Ktwpauto1IWUiTI3vvpkiS4hf2It98NUGx7htgCHB
6djgR7I9CUYCT5aIkMVOImCHVp5fCM6Lc7X/Khl4VSrXKXzVcFoD/G5F9bwQCdC8TVR+CjfvZ3kR
CACGmXgwAM0d44wTxsecd8MSZPHYDFSLScdPTQ/QC7MqltdHyb3WySTHDvTFenJvaGRBvBKvVi0I
+sBAUw12p9E8eZAuYAB5jAmymjAN6xWRJ7ian9igPkA+mGyOF9x9tKPeI9AUmYDndcxEgFp9n1WF
HRR2eJs33WMpEFgVcJoGkh1K8RyoOMskd+0yyTX2cHvfHCl1IrPpO3ZLmUXNy6MlSAF3Sq5A814O
acFKWaj7a4dYMJp5QQNtcpdRDGXcPuoctxxom7ggM+HSCU0Lb0UbFfWpH5tLH0AOclRvPJA/kI8i
H1y+SIQKZ+GCxVCILqSzKF7UMGzJqZ8USLJyIa3mrq5F79AsEy4HCIpX/ZLrrpms51p019/7KSld
CuRErBDSkSOb8MCjZ7cm/4HR6X8WH+qlcW65KMHwLqQm5xvvquAISwA1oAfi4lqdWJ0R+UGrAOgc
h4TFLmn50gV3KarByz/CiNRuVD7lAa/jBXvtmO38Z2GVgxxgw0rwU1qVfuWhpwAAv+rStl0ipk7I
V3P0zhpAv36bTEIneB38w8HHGatRLYLCFGzLejyEeCpNIn6DpeejQO+2cgwUqf5zd/YNm6qLRlQ3
XuCAV9vvbL7zUizmwzTIz1u+ohMSF9EbmDYEXVpw/wrSZrBuUtRAEZCtoSOFobSSZ+3T6qN/+JC0
2KYVvdeP8nXHgc1SdCtNJg4D4HAbFxfpOwETcSJGt18qh0bx+beehLd6IEKCr3E9Krzbnpi2uo0s
uSg3YlKc6kGY6EOfzc8rM04AWjLqLzypptMmGw0ZUIbE0fZvY3V7y1C+71WMEh4PMxTHz5SCKjKR
FOuimmq6/eW7z1Yy10EzmrtLI0Wr8mKks8z0vXIEyRN/PFvKUEjILFYLYmLvfejb1CcU9frg71Wm
OaXgJ9P/9YN0eGtoyJ5OGUM5FpeiV4rbQSi4figJdaGo17eCnGlZBK/WM531lTGCQbPqQb9I7xDp
ua7pzIRC2dL5K23txJ0IEWzJ3Kpxb5cul6E3u1DwgXKecNpvJcO4wxwVNXwWQrexUBrYz6cw5qHa
WLOC2HR3/Tk8yF/8cNjHNhrh//4YlDnsRZnJ5uIQMWP6JQ5myUUfcKOffUBwHljIWugoTd3MGA1M
gVtXaagyuCGKM++NGEK/CO1E9/RTVeR3EI+qAO28sh2ZCaPsiwK8Wl1V/hCpxd2MDOnvwR9aI5pa
JjPzPWOA3y0jvpskWC6KaMVPq/E7RPfmImWzqSwujtxl/lu+CRkrCqanNszkvhFkRMTSIedahj8l
eeCixyxb1c1pffq2hvfZ0OMAV7UwvwRe99khhPttbElAL0d1lh7DIC2BGcmfKjDpJhErxsVRRtAw
+9hrYBloq+IoDR65ykz6/8sfpIzY25g2bUsZ5LmvjgiADQ7W4R4nKRpziQKUQxRtele47nijTcHc
euigXxpG+QFeghBHEaGh6qL4CSra+WCREZnaX7biIllgoNggbChPwc/pK1Y9qOpjKnmmPvZIXyRf
YnR8aKCmQCAFVHQ5liZaXWisodpdaICMqY+Vd5nJHGdo8icImd0teVtvK5w40yeiCz0rb8ixK+BB
qvOEDYhuxDbdN+HCcCOmqeRevU6PXQm8OtjnpxSr6eYpdZ+3noXTTFBNVl5zATCBNzG3SaWr/KAM
2WExlneCFSPjJ2d3ChMSTPm6RR2dA394D90EelcyQU4Sp9Qk8L/OrgD0sq1G1bPSwtoQCKnRzREo
xgsocb7V0B0Eq6zdvhkG740Fb1hZNCXgioIRh7cuFQPzhTn/K40V/HDuHhe9G9gCdqggo7xPA5Aa
iUsKbJ3KrNbiq7LQGVbFOWSrppOADvep2MRFMzfyaroHiVwS6jT0TQiP/tOYWLOamDDLU4nFAOgh
2sK3qJglTkVkBfDJ2fRMcNq5bQu4HTv48dGIqhAcUrHZbMA2D04PetkM7t4b4wPcooP65Hs9r94G
pI5aI36TrAXuHU4o/b6ob6EtY9yg3Db506xZ0PSfh5/So+P1xXhHcfO89kkH/ctSmx3aAhX0z8At
VX779kGdo4I4i4itV+PX5sYKvFzlT+bpipEKhOqKSTFgNVI4mHdNDFSGt1QEhzgQzk5QlTZRqOgG
HP7eyuDK4WZso4JKIaHitbAOzSl2NOrNyHJ0XZGDilTDdUVlm3jAiAGRHdnna+95E02jmRWoAX5N
kfbWOhvbfxz6MhNxf2/rYhyoIa2L/QIHFaXJpI6/SrnULAwqwqIXyHEv+B7QV9uaPN0EDIF75tiJ
oCio/tLAS1UTuJpL09qAmYAH8vq7IPL7rDBGOQzeFBidSjgKXsllIU4I3AUIUnSeNWXaV7xqSj5T
BGwXBS0gKt1lLnBIu87t0LRsZmc4bbonzR5XXeBiV13HwP8WQw80BKKwqh4cscK9/x+NliRIxMFq
O3rXhtc1IbVuF80MaUBKw4Fqo1CPp2Ydms9vdMyLTqhr7l0iu/Y+xnfB+pqQsOPYZ1gIGNG4WJOv
dogMY7RKeTS1cxjbcGvjg90acIHtwY2+zho7ym6hfOZBsbVTPwR9h97yC2bEpkfCUaw8rsRoh50Y
/npzkoF/Xau2mx4L45wZ+M3rvO24klRnrn/PDYiZZbdZ9n/RF/EQM1F8R+T9X2ec7+NyFdve7DUT
R06LGBZj26Dl2GTOQFh2yG5U2FvQe9FPuC+N0sqIUAA9Bv+lAaZc8B8RuWGvID2FmdW01pUKJEQE
6aVk5g4PJuZHejbXJtv2CcTGh58iGP0oqwE2ZOsBLjzDuPQ/IBnOHiSlk4d2ojCApMTUua7KdwEv
lyID6mbF85FyAFaWFMbDjkSeCoZmvlXu4zRbvww05aN/r9slf/AlhCPjfjG0dC8WZOzeEwoFlfyU
ZAETcChd+/lZ3zRDg5dfNRwAj4GrcjUgcz8gf6PumGEs81iLY4tZcDh3i7HWDQ3Cd3VQjm0m6PWt
U7tPjOcus7Tc+sXB2EGI55nFEtww+PlzVDfiETnsIxvttgC4oGiextHJg+EJexLAOELUaXD9xe14
U4xqSMiluLy4qHL7+/6wk3pNbBYhNZy9G0tzRk0giyXp/FDwD5Zj/zg1HJKJF41sf+h74qAODqZp
0MeOC2EUaAMPFL66zW2bbHh1ZWhUw86tUx0gP6bDsWMSF9TCplAO+BRs+sqX7fRI10eMNzsuOeYD
3jnf6bJuE/HZXqYFa+8vII3XBOVzUJzcJC/iTazFRQKgFmMVKm45AzAm0MLVG6OKL6JiuZw5JZam
F20hnvaP/CB4xD85CFQZjVoe3d0thO23S73E2z6DhkOwB0m+xoHgwK1ozZOdXF92s/O/QDYaPHA3
Bw1gP+0hDb4QXi6sml3UE8AjUNKG1PosRax/aYK/V2QoPgseGuebZi481uXj9exCd6fsPfk1JWWk
hKWck883UmpP/up+ln345QAibKJmait/xd4wB23x12oHKvQkq6C4N4eHxz33huthEg6n+wToeQAm
MH/hOiZQXACD/PlQLBh+Qy8CcNqO9ixBh9keieTAzr9ReAmIDch8QzaK/rxFKN7XUG3QdTT+rmu6
Dgd/lA/ZnSKWMcwjN7APEXo2722PM7+L1PBgxE+twf8yU+WmAj06XxZcIxVsIw2j0R1oPEqlo1Im
rIl2Zyn5NTpUbNq11cyBP4jI8EaELg9tf5ub9FrL/N7JSkKXS/UxiEPQRuS7n6FkBZoPQZT+C5da
RgJMd1qL526ka5hk7pgDQJW8mMUuwjRR3IP4WyI856GKoRh/c8DYY5n7locSneHnPAUlCdOqKOA5
CGA+o5NNSCOK75glHNx2r1IewhoxyrNZqe+QCykKL3H642MuIUhHPmYS+FXEKfIBnHU/QEEAdmBr
HUTruYxTUMXawvyL/jjTBOqNuHiLebB7BOIZ+ARMoDqpbe7/FkZkUhrEx+GRBRDs0txiiLGgwVfJ
5tSQ5H0026mRtXs18VA8UQZ2PBSLEYfeSdjSvRc1r0TbcgKtSSDo7AM/nMN/E6cBpjbOkTmX4Z5F
4qY6qIzeJrK6oSWAMqfprKRLd0OmS+XE3LSjCUxmHkVX3sTVxGg0ke4oUJzjZNN5KIQ0uR9N3Ohi
wfwh6IAd2mvbkE6DqLys3Lm0KEL3GDp0TqAXSSw/bg+4pr+PmdK/pfElAPWsD0roGGbysdBwi69Q
g4I7K9i+OzSIyZynxBmzQsOdR6hMdFD+lILfZS2fOIqo2bqiJQGmj6VkxETVOvSWRmyM33fKdlyv
Bg9tzFOeU0gIOLOb1G+Lnooln1giwRc7JllXkVldKMLxdB7r9QJ68Gfd0WXhJbCvP8SPh1KvlVp2
Ni4qNRJG6okRCJI/iYuGAIM9OC3AaCDOXb51TFpwiPD5Ut86E7wfgnbC83DumcG66LEtZrHFZ2Br
JPNAHxc/QlvVbSIvPSNowuLw3hZnAlmuLlVGBWJW1taaCW4IRpLBj+oET8MhFIjr+2L83feaDQGH
f/2B15Fif2Dvy3TEo9bXkaHBavkmxV6XHWuxu8lWu5IQYK+VXIDdFlzvcUwZSH/Pl6Wd4w8KEyHW
qKOPDphiOKVEipMDv/dvbqhNCp0KKFVST4hLXh4yB8vDb7VfYdkrAo2jm/ho50HT05/qpGm/h51X
+d/Z9hngC86qMBMbPkb/F2ABf5Ps0fuP7cfiJMirusAigJ91VR47g3ljh9E+Qlsn40AVIYKYFcSR
irO+J2FoTy6saDKPFg+T0c8PziMwxqxktFSqulJ00W1gHHUX54RqEwZaYr+VZzN63yQnv6sCVU5L
4oP0+QWlESRYO/z7WA4XBjQkqkS92brt1FeApnYNBcqf+dN1KPDiWJQPVaYwsprzHi/GsU2Ne/4t
36vpM6y6/cfXLAWS3ekgc1kbhirGSL613F0caBE9FcpdzTswQUEwp/kXiWOZQwkPZZu9S3N+bb7H
YSPDhHOlk4/1Aq5SnCqsC9YscFRYlzRBM5XQKaALteukza59Rr1TGxECeRplVbdGScSGrBPZQWVD
LYo5fGZ6d77My8LtDwVJcaLPtMadcU6wZiZaRyGvdETQELEdNvZ8u4ndWwn490DplS9ThpvnYSPo
Eyt3iywqoqq7km13zxvsvSij4QrnTqBqrB37QiEb5SMEpsDNsR/1UrxNH3NB6uATvecrgAViI2ZN
AjbYFy/t3UGkxz664uDftLWGTqXw+oSa9Jv4FrcSVbuFqePyJNz32Ue5ZwmteBP1irRK3udZwz6Q
EEuMcWog+R6LB/w6ZRHnUiMTImpvIx/hGrbM8P4N3cgjyLMBvlvbYj48j33p1J5xx/B959eCKoGP
GsTjp1++7YlYUMjV0S+mEFciWHGh9Rspfs7Qgpsd9rXqcdvoSCKMWjzsKqp8VxbBPT0FikHn0SQu
jcAWkP0fl41GHwngk7HMh9G/O0CxNIClgUgw4SymlM7PbM6fVU0h5DtVCqX/NWW2/41PhOlaGfcN
qQqtR0W72qkFvukwIcZ35vKpdlQDePLd7cE1pRhDtQIXtn+j7iglYIWRr0j1008XZdBoKewjkrxH
caAR/+NRl+O/YjgfmH1PjJiRFqSy5nhH3zhhH77Hwr5g4rslKDIrg1plZXbItmojRpoR6FqZhZY+
KvjP6C3QMY3MAIEgR9fVPEf+BAjVVeFWEVfuVoUnscFntLvwlGutR+dcpHsuExn1eAWQDaJw/C6C
20aluzV0GQyb4/HxUHTLGYn/AA1IKpobCfhoS8q98P7TAw7x+uznUGv+3xfqbw97iCF+Xz9MNyoi
n8pCZjKNzLvtTOhIQLgqQz5PPjH8kZqn+9O9ikE2beQHyHfwki0jEL1NkD/LuLZlhBSph6t0GXVf
Jl/HdNVWTn2dT6zDSFiBOBoNyqTBDJL8yi0xKdbWRwl41zB3VTi4yNVknjvFZNHSN8oPZnasTY3X
PVjt5NNuQY0y40/+22lz7uCAHqFBMmzL1hObl60e3iT0AMIi0e0Syo0vTwV3x4Pr1orCfGvRZqlt
4r9AsBJaezPiGrjiNDB/AZU7YpcgymB1hO1cuFONOvP9s+WOEtkjDUIg8IENxON2kGqkMdZFsMkP
3x+/xuxDkWQzO7f6w49eJiuq2/1Ured89jAwja6gWsMwxE7aaycf6G4hVVV8FBf+iuyWeCgvWi3C
mhoetsb2lqovYjdworBR2If5MI8lJQuxjT2u+hubydKw56P/tdJ7GAzDerGe6MQySz/VgzJpVb5s
qxNIYGjBjKAXYA73zt7x1fQrMurDocAVUHhTrGYv+sjLMQupKcFAqgPAcYUc8e2KHgwZ1fOWXqcm
teCpITSghHCPP44A5H9/aC/WuhE47NwfS/fJndWr7mPxpcftg1dwrCnKlK9zDCMvn9/KSxHjx+3/
BgZjXo+siuGaS19L0S1o+sC70HZKBlw9o+zzu1OoThYmfSISiPF/IFmlP6NU4EEWLpmOqhtHT4B5
QgDBP/1fTnRaCNhd6Lp8A2Tuds27qcFn3f9ctDhOln3NBLH1niQvHCAl9e2KyBWMO6ALTZTg6BCn
rTejDGtwf92NrdaXXINnIc1ecDwqPboRhMRx9vEuR8iYqn87TRvKA2ijAYy707M8iEzhsVbVFamS
R2Ru5MbGsIWOlDgC6vjfwO+ExYTLWqAy+G5VEZlUHKND+/iRSuciCLimOzUz02r7n9up2vM5/2bg
YF9FAIdaNxG0LOs6SpmhhPwCiwRSWsNY30QNOa8LMkMe+V4Yx00l5K5TDP+WLYQdUC79kE/5KHHV
hO5VVkHBaK8R7XgLPAmuSy2jYYEGSqP4d9TpHDvIzB7IKCN1uknH+KGHfF1//j3BBT3Qm2nGKpok
mqDCpwhTflpKDkMTXuahphqiMdrEaJkrSkMm3Sag72+ql5r8ez5evtxAjmaheqYkme3gyTicLNPu
NXTAUabFFxPgb14+jD5VUaQcOX0O8hrgP1Aw5fdLG+eSY/GSomtfyWsh+SqI6yhU4di24E4/E9ct
AZb4eSqe9xo62JwD8doZcdNRnpgObYAwUjmPak4zVOPQ5Y5SbTF8BxBEAKayDHijurBcABOaqS6B
17W0u35WPtrvNwcPo1WXejim289QO0CPQ9sxoJbo+TM4BIAKNSQxY8HAJhAZEuj59hHA53ZurSVM
zGtpIm1WeD45MySRyFxqt74+H76Fol1FDkmRkjUQ2vUoF0V9G/ke128GnfQvyRMAgVvBDxYpm3KY
GZvq4NBGqD3TrLZKp5sHdBfFBAVoNSM9u/8xuAi8FR5UivZwYzBDfLKSyCnD9I6E01EPicQZ/qj/
BEYvzwMCSanb5pNmacLjvPVG7m1MjUonDOZHaEPUUAz/B+X2HGvcKKp6rb9aLAPRDyNB+m2YTRbd
YG5158ELNCiE1v0M7+IqVYWZvVmKe1zLzQQ0nZBQWh3PmvwaSWir57Aawvw0O3IDuYo9Qdnyu+2b
/V/X2a06jdXCg1WNce0lzo78gBM7sgrr2UxvNoob8LfefdFWaEMvHnWOgAn2PukgOI09ldZdJyfm
CWKl+Pm855aL9ZDlRyJCwRZWkffBrpxvfPQ9Xqt91obgf7NlHuN9dNiWESOQ8HvFMcrOZPNCAvS2
FtyE6rxazY5VDs56718kNL1kiMMWcGA5Tha6XWOBBfzAL+zuKCFdTE6gW+WV28ipZXd9ochW4bVM
IQoAae0cv4ZouOf0MZrHg/0Q8jDD6vBl7fhZzqAq2QGlYe7av9Cn2I5/17XJZIIXE7OeRTlURcwM
oOvsDmlvF2BH75nPqz1u6SG5JjNx6WWIB94FOqdXIpYUau0E7ZQiOsIcUg9nsiIhfod64xEIVICl
OLcxdCLosBT2jXpf95WGDuR9VqLemqrk/6w9oOJ7JjlXkkkL0s2g+UzBXIpR4/dVsTXqzV9GskpM
eDis6YsAnU73elUhiTClo9Js/lm0N2FOtA5HMANeZrWpvAt5j1ILjEW3sYPulRKKDaKntbeONbZr
LE96eZrJIZMbtH/I67fyMh4rXNMVi7CAPbd6XS1dbpK6JGaYijAMXsGoZ6qZDk1tS2x0gwqNw5Jj
qN82SCpWNUAd12hWNLsmuuCLYiqQvZnHC1XmZ5149zGrWgK7QaCWgUdp9TUEQg/Cqtno3v+LTnBc
1J3SJSxxWZtykg6n78RTNnoK1Ta/aCHs7jx7u7FPq3W6aiT/MrpSy59Ayr2UmMBxEW0834HJo/7n
YZx0xCLp36/MRhpAMGQU+KWg89CCFjYYEiGCUyWyVHVS05JI4j5zGs5AfqKnT+UH3yQ9QY99/bjj
WlB5pCG6MenMfxUEGVDxpYsgX70GphvJRMgue4tupp+/yOvPBAbLoLOLjZ9s6eJApHKlsdpyPyuE
rtUlu2tICSYxkWDFDr6IovRi8/jve6nQy5UKxLoUdtA5f60aN6SMqbAGeurUMA6SRvrE097sl/E1
ASGnp3slA3EY4asMyg6dj+plcZ6RVYpRf5GBLL3AHh9+VPjqUYV1Qx+1UBLnKwkXyT+eXrSDxXcw
NZmsEDFf6nu6BsVqpq553CL3hc2PPYJXqMyvXhTrkIqJJK4TExMnzJ7nGsDAcabxO9LGb7UWBeLM
Wt1AnqX5DplBh0zGVRnxDllFCC5M1qChulJ+f2Scmx6t6rlYgIIK5DhB1m23biXuasEDxcJiDU+t
zVoiTkiW/I6Dr9ntIIvC1isUEXGMNVcptmFyhIJ+ZFIOdYPqlQiATMvmU2aQOJiNAmsDAeoHMQ4+
5ox+v0S8WTvW/RzbjWd+tYqEZsxE7caM7fYABuvwjNBHkz+Xn9FYaBEQ+BUVasLNB/hR/tBR7+PZ
yhD97nyQGEBy3CKziHn/4YB/NGKo3TEGBUsAOgGkJxLS1aZksvLEThWJkVHmmG5UH1sBCNWJrJqG
TJR+Q8gTdGD5bSWLqaehlQ74xa5IQCCiJ447TtQWMl7CCpMkUiNczzk8CToBmYD6XPaYVfiNbAAy
0SoM8vBBzq4XGZws+nMd6H0cRWpJK7X4asPoUoSJqYSDcMTcTXH+6MwcbHkv3Pt9uc8SyDB/rCDV
Ra0HX+BhLpn416Lu857sMjs0twlIdIJeqiHs3ItvoTQgz8VVs1e7wIQo+mupwVdkblzjKlun/vb2
n9Fdm6JYuRhH5Vuy7PXO/jucDZ8eCtH8o0D+3cT5UvkES3G2ipcfJnr9h9/q1iwKOcgRxy2z2Vch
SO8rrEYigvK2FrwoeePfrSgekyUS1U1nM4oTetGY60bpFJdH6/J2+rmAJfzD/5uF8iNeChJpasB1
5V2xdmEjzZodl2sfgz9wJhOvwLXW7kX9LA9XFmPCngLNnkxOuPNFxjrXLFgtT+waZHZKvoVo2ho2
gaavSqyzuIyUfpLg/r7FJnCeup4+SKFRr/TCAmqw0ieofI7/nLKKFFGMK7aqpCGe57iQ7NDz6kU+
yxh5dIBmLvNUBhvzIl/R+4bISBiCJdjDuhLjp42AC/rk3ehE9+Kr7lN7SVQLuRtgnC9Z7dtzQV6E
bx9EyeJsCLsBBelxEG1E6iZArMSlkH9skmVSoKZAL54ap1LngaWuTEQI4WD/h3aXdtvXdN7yqkm/
IuHe+LsIlVjAbwZwlxsOnWAQn0C+83XR//qMQT2a0Bmk766c2KqNKVSdaVZfrTXz/iVH9gUJC8As
TcgHhpwyKbehtgwBcG1tZSRpyZHQOVXEgtpSANVoDOz0c37Bu0TsKO8mCz1pfZ5MrhQFK5NyCfUi
caUu26tHWuN8mxlli6DLl2DEZUWZGGJOIjQvd7CV0OKEY9U5HkPwUcgJWoTTiNHVnKgprtKd++Ub
SGX2F2CSaRlTnbeFOuRBJ6B/RFfRnj3HLTyl03b0O43Jc+x5aF6S/C1YXk3vTjGaKRZvg1R+AWAj
P4pzOtMApjRxciAZDbg0oOAEOj3DmQt7/Zy62JPlBitXahl9lHhQ3SF/pWvV6imjcLddw2oq5HME
s1UD/4C0g9EiNXy0gDxW5xnzlUITkIVkeaQONj/n8ENCW3RZejR2F9d4enJe7G5KPiqCMpljOH4B
4MbPpk77J3p3l8bjyk5csd24HNTsEvIiSoXQx5djAM5s7AIUqykAOb3PtpsKZ6qDJaHqr47CGE5E
DaMtDkt6bFIzZ8/opKHIs6az80lrfitGHJrcxDmWbvAQVBrOCRU27pRLAQIwH6QpeACN/rxqUxVb
LQcdwRi6SN/YAEoNXtx5ipWWbHcAhL8RHwHffoX1LI+hw5wy9DOgqpGcK96y/HO1aby/ym4mZDEy
KXhw3KMZiJRmmYdGOYgBq9U1g440GdZTKHcquUWV2nIpOcnXcqITio/ihiQo2UoKBXY0iVp4L5eR
zDzNkCSY+M+olLXeGy36jsvzUpRmAjOSbdSzGbcIJLGNKy91tc5dZk9IIFTHD7DcsWrvlQBMQE/j
EVcrvxZb1+JWAfR5Y1RX5Emr1pNxT6XVz0PqZoYKIdzJM5JH2uWrgOISMVwRbwKANLsXDXVM4qtz
qXFYxYTi3jtoFXNK7rp0JtErzlLAsW6G1xZeg0U+G1zOcTNTncNWmTxCTC6/mXs8ASol7IeiWAAu
ySxkp8N6RjMMmVqTvUGHvtRjd6iOlGc+rviV9vFF9waMOVIqfHRBzVcRaI9n04FGMsFZuMDuMOA1
GaeehS8zfOBGW2vJt2Q6gOiPYsWWLTwsDlXZBOAOyIDll0xDP1eQ0z/lTfxHcxpfTY0sYcZLdIx2
NbfL8/KPqqmP5Ctsjx6/nB2hI9QT8EmmKM60MUJlDfd7x9lI7v+BZSwM6OXUBh7YI+9Vel4qnsiT
+ctrTInTUH15ptY5XsjJehQEcNHEydu/3XtRS1klNiS09/n0Xi6R8/8qUJdo1nUMzExwtcTkcXJQ
mkk4lxO2udZd1LUa3yNhKDPXaPNhTcl6mMvFdWPvxY6sE3ic+y9afRvfhkuxGabG5SNRxREj40+u
fIGmdaE3pf9c/CdCIPm+SvsLZyFAVJ4ra9o6odRKkqqakqP3ZHF/JOG9Qkr9Z68OIO4T/ya8Ft0e
7hImDOnLOyqcYXIpETonr0YNf/1eCHuGUoSZoTw5tb5oc+dOvwCKSzAMw+Kmr8bmEVXeOsOayc2E
S+ylZFa4lS1jMtTKNzMNsmtFwhvmbOuUufP5LjTPP7DbQhUMKmMXDuic+uCckYefnTrZgCsapNqD
kGINmi649JGlUKuj6DLhqsF4E60ZdAQ6MxEkwK8VMv3R5fU3bat8HL9l2jxK0szHRoIoGGNxYvFa
RUU/OiLucrVLmWIbfaxPMoKR3PQZ2668Dvx93KDcECJzMoejZ+6nkiYHHnpUnueNA2IznB4IsHda
W0mgLGxKYIgXv4mvefK7fUDikizZJRmiTUBPToEAjkeMQs73xEBsj5Lk4doxyb5qmgaPQdATJWZO
oP0YFVIpOtWWoPaVdPRmZcYwod/M1DrTtgdLddqbtB/SkmWV1ZQvomc3ofzwuEjQks2NDhZQV0Qe
n6KPIqjy2unVqtGmLt/9KKbxCU5E9EIvjhGvFS3pBmVW5gZHOz+HK+SwCepdvhfjbTe/RsLPapch
O/g1eu3k/Jl2wLousl/AkTp1gISZ/P0KPSijItczI2rIAYVQTOrvhGwYErUspiLka3Gs9XD6GEUp
K4qxDHzwhqVvsL4bFNqJWNmice5EpRxHA3Imf2pdGH1c/cthDKe7SE93C1zgORXmPvm8iXY9YpPi
barRUNL0pDzfbt9W4o3V9jFt1HhpYMX8OXBzz4gJX8k+Vl+HOysLttviLMzrtfebJbMoVLocQCm5
31LLbPYCZ68YNBdDNQC9k9iGUq/mGxlwKeFrMrnWKs89sEPygQIvMmrBH3S7sGGewHLTXM+wh4CR
vWgODMlGnGlnYysgEPidjqEFmbG1yWjuSott9dKkYf4wpzSrMzfcq/xtP7nwMweiX4VLEwTmDSps
2OJ+ICq1AYu/VxGXo9GD1qeE2ICNFfWJY9fkPS4Rv4BZMyGIGKmDVnwhXVcdcGhqaJ22qcMAVoTm
FMryKakRvI59UmYqr+UUPRnS3wpF4fcDhmxzMvCfPam+ramehaCoWkhfWNBH/xMPiKuBZjd1U3BZ
sFhr7wOFK0FVeuTV/Qv+pEg0a3FhlysqI3b0cB1tCVNTEL0s+I4XYSxpJ2Xtk6RV9SgnWuC73IC1
dMxmSxaSEOUaYI8nt9YNM9xiZGRXJn2TaG+7ipKBr8rUmngv1p6QNzJxoEhVcdHIZ+Ix8aRMlCd2
Zonc2KaVmIhK46Zxfl+SjlmN/AsS8fA7+fI0AWyfiFrPILscZI7WugTO4DZ/ODI1IEdRZpFlUsHa
WTNdM+m39jjIlvPSxnph0deFkuAH7+k8sJiTY/gVqqG5K+qtmXLkV2dWYYUNHr0tTZaeOKtGUy23
OxuXwCGC4NhRm6dbSv+LbMpEcvu5BUipJGkXvt+ivtkdseOE3qsAe+ZDx4kx3wxo2rQAmXIbdr2F
PoH4xePh7O9tN1GLnE8kwNzYZnA+CZGaz/wilrT4FdJO5N27sAbw7hBBbYe50bYWTHZGowKnX7ss
jka/3sHaLH82a7bhYwmiYimez195aLzqukJI1GphWA7dW3a8ubqM/gxOzkYWntjRCyhPmnsU+r8B
ml+akqxJY66SVgc0lzhWVKTkKJ1+cqM6Q2h7FEB5/46BVk4S6udmUfkgr/1dylv7DzNZ/U/0eBTi
I5PijG9bYE7iR7nR/5wJtSisHY1uqwzjGh7d2mxBLTi6Dai0Srb8aiEM1l8NxCZ2U0gJzbg+eY+6
bix0ygdSwDd+f49lyX0hqqT/L+rbL0FT8hJD84QGydijvjeBeoeoKX+esf8PY40RPNGwjEwZMWND
ljyQ/xiRqm4+RqacEmbYWcBRsvrFdxaUvTcB4KFyp74OdCq/DPtWTECJU9ukUzd11PcoiOJ1fzV8
I0owYAkGr+oJHJSRhtxca1f0SJW9H/i6u1H2xrmd18CXpdb4ex2zckjm0+hXW+Pgo8vO/PqF0Tpz
AdWnf16SwYPmUbO0Tm2ndpIyAyni58X9TRHB4gPrEGX+pbdLaPcUsou74WS4sSkNqlpts62xrEdv
WlpcpMzHDeNVZ5gmh0d2ovNqeMjl97YcGzCF5G54r+LRtQMuJa6e6jQEJDvAtCAcQo7MvkllsaUj
OlGBrMyBZqHQZfmktvIsTBocZD37JsDELo1R2LhVb+lC/7ZvUuVsOWwfyterKXxQm8L7lsOYutMS
eJ7KZlA2fpyyPW7iJ1WTP/U4lP/4TikPWvITi1Pw92N3NYVmjFTr3SBwdKfD80jGY3HzjqIN1weL
p/C5FtGVz+upAo0Kr8ZQ7/78qy6F67hh18NqydO+UZ/GU9JdLH4tw2F0hKaRKRZRyS1gpNVuPe3K
dA35pKShmzon7biTbRhnAJiseHZ8scbH2FXApnQS24spAoW653JG8Id1SPzv37Gtg80QYNttl16/
PhOCPP09ieV9oXPEVOoyzCfeZ9pPSaKJjYasmRpYFRDoQoJyaNpmahgBTcWUW6Vg6Tdph+hIK/Po
FOMmsieuGDHHjI3YsBK+6mM8NSVs0NfQvdxPgSQfuQE7CMyamdCjvT0zcqfVdmxnyaG8TMXW6ISj
iT29CG6qrPT6iz7G2BYlukA/yER+0c78oze6IXzxD6vm4jQ4CteD26oNVlXINqYm/En3PfIwzEQO
dT3qN1g/j1OiTRNehDdHTxdXJgCmaGtFPIMb6GIkqF/opuM9UMWOlQpJ1rH/5dBaMB/7XqHy4GgO
26gGsoNr9bIz19ZTQqgwNr9EZKog4pWu+PuXDJ1AHqP7bTK7aQuAk2842XTzTH9dk1EvHGnbNvC/
QOMpPK5dYJIhnsD1DJLLERJJAnyv6PJJoJAf8ogiPjrGtNy8jjfeAJcKPsCfrwYDbphUdBbgDgCK
jWABGArUGCqAWiLk/jpK6GWWUThUIUdHsTaWvz4+HBGWsK1fK96HnZiWmxqrmjI38GVtw2kApfSx
s/mC2WpXFafYtPDQTnxo4v0nqGS91Uu6qDkDAC/N172A1yVHqCzYZtMkBQfF/ZAi0p9BLgDhglw3
5u5qZ/R6fUYZKB87ERA5I68wv0x8p/gGL/4vQR3AAl6ANwXxaFD6+JYhTZ4+Ixw4iYcEZzL4/sJ4
491ZznaUSw1oiHVXhQGHcvXZXn+dlWEOyDVaf5dQ/XKUpNIV4MDsBVPQTrr86+1ivPRZGa+3Tkwg
+MdR66a72GRdPZ/vmsGH3VIUK/31LH6snYbcclH21vskZuXXPCTffQr95AlnJasfA098kITOpKhb
qbl9IcqTSo21k/pyouQlHjuiB604mOrrlyGva01WPBGpAvtyNxtmmzAeCIcLhQiRirV6zyOfK2yr
FMfNTD9DDWoPn1MOOMtlgvI7+nkbFwxPG/jea+DWHRInQ0BGSgIQaKtyIIl/yMcmFrupUcZ7elvs
pxyNi95x67ZIDJe5UdCG/2qdoKqyDl9DnP7iz9PQmd0CRiIfjaowlBlii0Iphm54ZADQq2dcdj0M
bMhNiAwBEp9cgTbX6pBz8RO7GGEPQwBwvS5xcEjNwLXYD5eGFlSStbRV+01806p0ityaoCpbJoqL
E8pwqECgsGlGRY32cVulgfMqd8RmCzqPwbwn3BDhEygG3F9aBAFJnHgOxcrlNai+A3uRUzbMKaDj
yiiFeh167eoLDZHR6sXo5FfgsGqTovO5nny+KOyXO1L1Bb1CYSC0hZ+RPIV0X2+/sA2/eYCF6Tau
DAr2ChDHy8FvMLJgM+zDpIXWRTtcWEZWcvRFwn1v0s0nUbPG9HDgmy3KR4aKIwDOwTHFRk6hau7T
a4ZEv6tNIes6SB1Nh+cYzd5ockVlXkrejW7/TsEvuiEEbxw3VH4eGJ0I2lemD2DAEs35AqJ/4aSD
CVEOqj2v40F+JTaVEJDT/7Z9RHstDvqEliLpsmXV7FZ2qs+1y1YA14o6JTX93jugGfXyIme3Fi5j
oiYSC9LWqtJrBHQpO7mCVhoAr3cgIA6RFkWFSDBpiuuW92TpOWByKEGe+M/t4OAJN33dBekAQmIP
y3G5Ail24/6WdKXYiz4vRrgpmDZOG8WgK2lwIS8WOgnThusoMqNGap+vIPsQ4A1XSaqYKQ6DWzo1
hJmshX3V1+JeEVBIKubHkmqnEO5RcAghvtU2VM9jeEGt6JJYTdaH1vUKYj7PN8BpIeCQMGSs+hxd
5gVVOP2y23kKb159dCd7NtsQbGXpX3wTXiVguUQ5GoNf697cxuE5LFHzhE6yGf4cMi0mlz5PV5/B
mOysZF0z8T5uOMhbtO5mgscOIazetEirOIERq2t9Wf0xUift+aCw+c27hnnoH3Y66w/O2NUgUKDO
+HoUY1LLWgkUd6p7tYN847gJrpVGIX1ofiMy2fUvGtz+xLJDpiFAmieGYrl6O497EWO+EpjUMwAQ
u2QtcXVHTfjzn4YjHvrcUzhUZPPGKD1LzuSxo3uGbSAhemPgjMi7ZdJCigqExJlG1YvGYD84jT3g
WZ2J9d+5+8dHIqgTepJlpahQjGmMdCoL2uw5hntrBok2PNBZKQ6GsZNKlYOMqmAa6OKMdyXebjz2
TOJGlJevnqcs8bzml6DywggZrStvDn/dXNreGEfAmP/11rpSpEkug92Ae6uetlP45hi70V4+sA3y
RGAyBAWBNUBVJJxfByDBtevU5bzdNdPC6eHAGmHiEO6qNONpEFFJeOudGF3eXnQ+DRvC3KngSpNI
1gKmY42/kX5MNAUJTDpMbmCSFi8cpk/kdC4bb5Jc3BJfswDRqzz/WV0Azm+zRb3BU4hAPA14cs38
jd3ZyXhs4jDlxyH2680sfIXednWebGH7lHGEV+6GOXJSDO5WO2T7vrGrZc+NaT7flbaDORg75+Pa
ZLHnkH+n8wQN8TTUs3YUsEQf7/xUOU5tIXhia2RqgI2Cst1n6UoUlti2G3X9Yz9kpcrtXRGJCv0n
OI02s5M8bUlci1Ku6o28LzZ+LxpcSvdr+MAdR1i5R8szNqaBktoLR+eAzGBFMQ782G0B9CBGSAJG
aswsuPEmZ9ZtDk8phYcIHYQFOPmI7oostNsk2NvTipwMZ53cvrK9CIFyTYZgKHUFOCkPppdOOq0H
luavmHzAAy5zxk0BEw6MyxfvOPWDdYD9OWfqMOXu+XvAWN7nEWaTY6iNafxlkhKIMma+qucbz5l/
M9vabZmi4W8Q32WBAJvLb8Jf+5+z8aGG4v3hjxnnuV42k5Bdf7QAY0UyUueqIsoat00CFxRyNI2g
pfVGtSnc3y12bEd8bLruLaWYe4DI5dC6Rydhv84EICf8fCVHAhyYecX5ZLott4SSusmerqiaPLCu
JfaclFNsLYOCSf9OxXed3RfYbMPULdtbO+vxzzNm2Hc+A6y4HbSRGj47WqorCoX/DvU/HVKTFHhK
IcE31xgcmFdySS24nGy4d2ls3tpRnMQqaxC4KhLj0P/Z/Aote16xjuJYQCNZl+2parmjFDyFOKIu
ol6RlWIAOZ5cJSK6BHfx3fvwWA7yz2z41uP9yei3Caf164ktco5LfALif0+DAD+eB5WrGhlu+yx9
tToDoeXvLn1pxuVUofFoOw2DOqD8OlgPh3Vc2xeNxn9rnR19duD2LUqwe61HcABvZc/WB9jg+xKI
5LqQ4yHxfKN6i23jMfrCfWJSNMmPoXl6dDfg799T1oItg2HfZDTPx69CKXVKlMzga6AcVkLZeoBu
+d2lx+A3HCNejgRiaPiQzpRm6YI7bC4mr7jddqWoMEJD7sjajzaOlNxuR2MoyQkg6pIpkUYsfVAY
p7PneD8Kr/ZCRNYNEFYoin2LqaMLlmPxIHxZzsuSxfzPYHK+RWGs4nvs79s4p6UcLkA+kAEme0QR
eTaakPElEkUS9tXVm1DabaiBuSmrD1MsQSh+DxFEyFtIHJ+YRwaGXVqRMT5kkm8MnYFlUS8K1pSm
LL1No8MADyOA+O3PK9lIQ87w9seHYBAmsEr4OLjfixIzZtUYa550WzUlw4aafhn1jwBf/iUNfkSD
whM6iex6DvIhFSp7vo9Wf5KajLHCV/b3o98KKeK4dT9C9h7v/9wR2gWXOQ6I7UIE21cMUUVnFCGl
cSqAHCcDLQv/BDz1ZD1lanDfYu6BzZPlvBZA7Hv9hQ87/t/mC3g6LeeyIXTnmBiEI8CD9mdS4zla
cf5h3McBtu44aWXVcWMfYioGK0GskzE57pm61bDhRpyBU98EGmMY/htMnEzwPq+yct1L6KvY+PAv
2eMg7hniNpNr0jrAszF+P481gfRlL+v+DgzNf35NHShTTfPTb+jIHQuSDZrN6rQWdut/KyNBkjSm
nIFJ+nNke5EeiypXNb3ILbvlJ5E8AwznCdjpSOdEy7lbitjoCBKLUELGv0OhJscTHuSvfv/ei0L3
1lHzFMAZiFoY3LckufjW9KrDgcQd9MPfQX0Wy36rEP5uNC59pCFuV+cIEWYi3l3zDU2uy3OsiHT7
10yixfxrEzFqckIa2nPbUfRXlcd1BkloqazgHBrIktjVZ9O1EJ0UHU7jZ3gi4h68XX4wq7eliiLC
pVpGysvEhyViF1z9kgz50ni0zWVQ8eB93JLvyDOHxIfWGNJ5xw8OyeXkEiPiBgzX2TUGFrnj9okm
rMUFNoFW/DMwd3IPa2SHZEJgSkZ32mZ6FH4zKwkyO28aoFeJoSQSN/8CFcVr1bLcv+QBnVD1kEQG
AnpIilRhIIWqUM8/WVaVYec+VLDV9bXkuNqP9be3PYi59bMJUO45L2p+OGYA1BJDTtHeQgpN2bwZ
J3r0Sj2emx1dYJYkamlH2q9kj/x/msz8YGK82+vfVa1bN57jSJyljETwFtkp9aG5/wO/uyKAksNv
GYLzToge0m6AAbqFVI9ovKLd803hxxa8LCJey7Jy/24MFZM+zBtRgu1jD7NueGni7eyzNcGRR/Qx
qzcIQJmb2ufAtZANzdBlI8D6XozpeQjNJ5KYQSAgo1pxLaqAPpOegApn62RbNAPiLZlp756yO10R
GRhsHteJdIvtooOmhoDYUVk3fblHCLjqik3WogLTWplezBtNdjNV0KmcRi6Rg5Q/JVjsR2XSSAcL
gOWEQLxzu+a24UdZkw3rbqEhOXWdgH9GtmRDf1zxCtw0IYwM6mqo7xmmSDKTpebC0xUu8LfFpAo4
1bsAcKoiSJvpJx/ZBFSpOauGu4Uj0r7g6eflWHjzPhK0EjivbRERWc/6sKMpJEGrvcYsHSiv5GeB
dHJG1s4aWWZ0CCQmWB/qhUM4bbyaj0XPCyNBMMiqJLeMaah3LfgjxrHvpMJsNrEjKmZVowL6lqtr
6Wt0UiNYLm3QuOIW7nFe7q6JZ2BGxEGvj1XItOeIw5iomacNhAtGfLf8B2iGIDHXe5vB257GPKuL
O2GmLOZmsjTzkuTosfUmdQORM3hmsLOqPtGofROoMpn24yl+BFnYnLVDA3K0HezuWbfxLDev1hH+
UkNKBiIXRp7UTWSkj2K9kd5hlQbJAc2IPjKp1G/3efItIIWCMhosjRgjZqQGyR6bC0dGTL0wwhUB
J8R9Y0UeJl0zyUPEVta6lPX+UZbA9bTnlKiMVDvUXWnf6++CmYcGenMETkkGdhj+DwNgUNt9KzuC
EZDzwXinb5N39pFmwPfl+FsIJqFFpm2DD+tjqHPB4v/jFfVu+0UkctPCh40h+QIJXaET7l76sSIC
h0w0DscQFkDvtB+c9htWUJ2p19fY8D21k7XMbwh3QISgMdMRpLu08CSqcgrQ1JZ7MnnRl9+oDB5P
uZdUzvyzOrFXZX1uzps8g2p3QYQy5+xUw5VUvr0zPB1oaJEyeROYCDoYjdARyDNjFGHIcjayodWr
LTMF+jkKavlpR1AKxEAnI0ECorqgRk9+01IWJNkTHU8V2rYVA9eKp9XFyhR0ECM841kQBXJf9o5v
DZ9DrU7fowpIditlLUGTTokkAqkxhgTpZwIOXEG472uHwceQdHzaHQS1jTbk682s6qRNSPHLMYQd
uDHejWPr6ciLN9vVezS+FltpQHd8EmqctG8NQUkHxPEnWD8M6gboWpPhAH+DFl5l87RK+XxvyAwb
Xp27jCIwhl9qwUjjMOqv6JMP9XCpoFa8eQFSX7nwrmPFsBogPdHVLKi8gztv7vRQ37zynB1Z96ts
SamOj8fUp9UC0ZlCf4zq/yPiubbDEFYsLYC/jV5x8uwX7XoKJY6W0/9bYnggV08MhrPzlDzmK4Bu
ATlMcaQdgAxVGkgttrzuzoYPSVW8mRsS0tV6sgxjF5+NGuqse8VuNDTUe7mAQxcB4HJ2izJFjY+q
NRPMvCihrUXt3wZ3riJLT/F5yTqbazUlTR7Q6aY0jWP/UPecX2hkpyDoTlKTR1W2/1obMPzeZpY3
9LVu0kbnOCiLjyfBA/89gz+tDfTw9Or/FPCeXS9aC4m8Bij2C8oxda819ZOdqz9Gy02Ix24o+vHW
O864B2/nL84gTIMasOe/4X1mKxKZDp4Hq72+233JLWkuzLscRMWBh51aBDW0rbT2gaYJUg58t6ty
qHuzarA1iU4swqR+rnDPS8CFCg0lrIO8bSi1eZAwbwFfM/ao0hiaPteGZybd+sk0d4m8f+sb3GkJ
Tqro92WsmLwTtjrZnfUzB6lCPVmIEqmvdH3CX9FQbb/+/3FbOw0CSb5mgF0RfgUwf32i/vQ60oqd
kFho/W+Unro7QpjIsBf2nl6v3+4PAUt2+nQmTaA1Gkf2hyPrwYgw/WHtLaYvcmLEvKmQQ+I/3Wf2
P/yB2Iav8NZrUtNHFKnp9d7BkxygCOO1xgJetnm8MCHLaUJNKPz1D/Pd+ZuChh4OQsnizxqhYHaW
Tjrkl7MRJQT84RATsPRIqgr89n4zAD5A+0js3AWSGmySgUT10BxYQYFRYe63+/BYTUC9KVGOLMMN
Ozb+arE4+hsYFjrNW/3xE/k3Ry4egDaS9nxUS+l8plUdJlS29qEpRpLI+51hkAXXzc9qrruMhrS4
ZBSbAMhWRPw9iD7+NhZZBkwgJIO3OId8OcroUp9Cu8qIe9GeFGngnkYAL5LwVGhj8cXL8peNGguX
o5PgJlB9GuBSGNbE+I2tJsd/rsouBAWupOlE2ewwYcr3GlUUTw+9ldfS9Y5badU/dhmBvkwBj3Gj
aY2I+Yd7BX5RoSJIj5TxEM1lW2RxBPv1MKsSFrXWHFtXZUrABQLcEH67rN1zVrMCvH7XNkzQntaL
39H846RbArXgpe6CUSQsnAafcfLt6ZZgaufkyW3sw8E/zNexEJYB2yiQJuDqoQRKQn83XZqYIv3D
e9zsFPxt+hwB2FHTh2p7fn3CRUvwc6831BWxJ2zKJaIoIW3lyWL5aEU3iSAVxklBg3MH6WKkSztI
pe52063wYRZiL1qUyivGiEIfRrHMnsgJzJMeQ5OyhUyM+KYWvJomCIjVhjHoMr/PxK/Jp2N95d+G
0Ea547WvQjF4L8avgMEBmxR3/bBvCxkhY0tHjFaplwbdwFoZWIl/gC4iF6RtnU0k3Gvn2wMANvmh
VRJz5G7ICYnZ/SWj6I3XhoGzHbcrVNC/2Uv1YimrHk7RQb5Ltg4SHnjA5Vk38JxP5zZvvbzEMq+b
9QSZOj6y+y10pLFix296r04pIVKFJGj1swGdU273o75OY5aCULNREvvfyMWu23tUDb/d3F7E4Uwa
rivw+iM01bzsZ6bQpeMi6cAxi0niwM3wfsZPQKD3EeiALga8pmcUJ6EO7u5AkdHCMkaThUlDD14p
GFtm80AlrqHCx9uAyAew9MVEKdEFFHJNjgQ0B5qaBU9ILjGehVjbeWOoat30RbI1g7G8Z7bx+YgT
6CLFe8rZ73nLlWLK1+52EKuE0Zxz/x7jfneT92FWacbRCHnIpZvVGJTBKD65AfSE+O05TZFb3hXe
KoF7Z94CJ7R5VESQAsdm9DakFDgtx1rSuXLalvz9jinVLPtNY0tdS3N2UI6/Y3FIHGpu2s/PEgFU
mSB/soLaA7wJA6snbgKZdZxrUbq1nfwPmRQAT5qlIiYF0XhVvX6V0Xx6xqfLz8U6PCHIyab31/Ti
qQE9Tva/CkAeoHZZxTzP+iJ57scMA9zjNN2ykAXXhToxNYMJkxyFlP4Bj83NBHuztK8Kog6u53pZ
pT0tXPNm40ExXjcskVV74kS707RLbyPYg8NuJSEbMUN0vAX/PLIURDr9NRKPxyCWodtDupb/2EZj
J8qdU/ssqrWDdOLcNUViaNBs8xykeYWqsvAzXakQ2QLHIW/JwgPop96WbLWyJCPUOr1ZV1CkJLVt
tK4FLXhm3fVErgi7u/Zjm9favHQ+apqeVy/i60kwDx4iCwC+Aqo4OHQii3IMK14Dlh1w+FLWeJ0M
6lUI1c4InEzEYmoPu3qiRqgAKFmvuL2vz+Ev+rG/iROqhr+qIPUIzCZKHHpbpbyAFVHCTb19kCrq
LeeGR30d4UOjN3rHFnBn4UHsPfBD/2sh7643EPVS1DnOMBg5JsjpSFFqMm2to6rY55arUD3/5bTa
auwhoonbRZTFzPtJPDmdMwARChqFXFy2M6L+4rBDFVi4yOw7UqAc5MxapeULFJH+zA/Yng/TIR3D
b/wWSByzELNYgPfpotKl0J5zxq1vd1uC5qlQFKrE6+p1ALO+lSQ/uLEmzDNYdsSiiezGcTCH3TI/
+V3mbT1EAmpv0oRxChZpe+M+bQgVGqtOy+NpLD8O0u6hiulkcq5HsnDWMbg5K+bqdmkPpl77pLrN
8Zimf4kBbpSl4dXRXBBr+i4K0QDwgG3EbY/9m9yDhfuSaidM4AmSRmWQl5Ci5cZ9qiyFdzc+S0RF
atthhlHIxIsVBxPlJV3p5Fc6dncl+gCTi9SBhs4cFDvv8dSRzv0Y7m816ujSPe8ty8DNplh8F9dt
9aHfi2tpGxA2wt1Vcz/xdzehHVr9mBOUJrYXrXCPOhGTqI4oLOHKgS17GjvzEd1/e3BS9z2tQ6dD
imC/6Q6UIchu11fmTcGPdsTEXAdXNdAHnRJYFqwpiM3TrPB43Yn0tTCCnokoVCuZ8h53iXEM6Wzy
3TNAVQsdCniCKRKkMDomzh6CnfgQWEZs3F/j3g2swJ3zCHwd7elwSmETMIMQNybNfaBZjlBfXU3l
s1L8426l5FDBoBwllcU1KXoofXb1RobLfRYAo/QJclK39JmlwXDYQNBn8H4jxy881Qcnpt8cGLDP
5Ye98wM37dTrB5RCeL9fO0DqebsDJRT+Ne+b2a/w5NjnrBpltHiq+qWV2TQIOcRuFzx8SJppJ9Iy
8hjgP3AbQju2b1u2T/MqlYiJA0kiGlSXRkGIQMiKIPJUrsE9ABq/1YPXGqSM6H9VuGmCtBhhBSfu
iNcr6NsxMXXxZbhv6+jqk4kDtE39zvXUfA7Rq7W0nZbNM7wRjqmW6f7Yk3rS4o+XaEjjpaOEl+fI
W72brlkkrQoFXTgTbQiM5fav9YDW7CUSjjrs8RiH1rhfW+WlPxMwHG1AnTuSrQHCzq/jRTYr7Guc
UCpZEUyhQycgovxUv3kGSnRcc5n7Q52fPMn7k3ZFOsImDlbjSOtQoC1bHL1IXNG2VcAxOUvdQ6nl
veHnN2G2NgXZHyHs0OzfU3Ga03C6Ztnd53WYKP772n8tOTpLfYiVBWNCnF9z3Nb0j6VBEsOEOtir
HxP3mAcuY5DBacZcZrijBpVbEhVb0DbWIXAO2v5yQ822uUP/4roA7ohnfHT22mBXBMzz1nly4oYw
psdUOBrdK2lRXLQrrX7uFHhqmtOTBQHTa+3u9AB7/2j3/FyzcPr/6wL/fWtXsc1gSyv4TGOk6VPf
kPE1mlzpdRNm7Qt/sL9gRqi1Dio2sNISFosYV+1xfb6rnh9UYKiac9241TQJycLVxlGq1zu4n+Vn
h5v+F8SEedNngFdjGzplUAk7SRTsLADbVubDHm6E6+w5+UUl8eUEqvIoXpKGkztaQFxHY3oSH3cN
lg7tYu4cTkDT+a7TQnykzfgZQi8gZsitYYbhG/YCaXOjVrOSkL5DM1PGqWZHabqzUoWPysaPLdEn
LonbedpY8RbDqPju4sHNUyRTUVTK1zwqhayVbPiem6EaKjdf6fdsQ3l59E2LNOVqVpLMTsL3gsiQ
sJje0iWuZZnN10zPVttJcV0+tBY9Dlu8HVwtMokOuCDAT1zqEjBD/+pMzC4sgm0xoWmSDl9/igI3
8BcoO3vpvABMPOFaeMS3PawIbmJXDw5wDekHhz1Uz9v9IUAaSDIrQVV+zALpLPkuE/j5czobq0Jm
3HRD8FHM/Q4TkSQ485vL3BXjD49//jDIqzM45qc1tZJD3juSjpCGaLkbcO+YZJXpAzMsR78+lpQn
DhKWUeOSg/kmsfZmMkkWvnKR7TrCWenEBZxasHph2m85hjC+H3i1zKKNKFL79SXroQATF52i/bpU
9eNtYQavqItVQZVn0FvVKBQSQWRvuo8iL4IdaZ+2pp1U2QQBUiuts0Ny/XbSlCYJY5LVMncAQi5C
Ui8UZoeKmKOOUu4vw54FUEUgr77fkNs2MhaSifYzrURNjfoxU0Vt/dA1IED9Hvewi3iY/isv3QDc
nv4SOGlEQkPdFBXIrtXCVUTVezDFDNUkJyDEj7NTNrkSj/Ymor+k/aSsjdu/4BE7fs8kK3Zw21MQ
ilbi0druG32xrGARrzXnh8+dTdt71OXAKF3dBrF1Y4N9Jd21KLGq2+qczhU8ACUaBw+gAjkvQYMy
hMURHp8lvM/akmPdjAExLyZQtefWn2uOOxfkQ/XnnEukNG5yW34jnNrKzqdSU8VkE7SdYNrsvq+b
DOimZ5NVZmQAgbHgxdHs9+CnlNLn3DQ7tkz5J5k1k4/EK2MiXRrH6V2JaoPGZV+DvYX7cMnDiOpA
vGlVWOCfkZGOWXrDEghLTkBQ1lgzzc5E1LZMlga/ExAUygu9+z0YjM+YyjpGbu2SdVsuvASjKwtV
kPHsmBiXchJpT6rhc2ZF26DYm5KDUeyc9PNnQ9zFD/YceMPu2aNkcKS0sRpi8OxbgQZp7oIw121F
UgQaB5omwEr1iwIoF8mLKQ8lXak9qPFbSF8HMuXzVW+Lwr+XZzbYX8B2KV6Qq63XNNrIrQdxL0oJ
4rQOGLycHW+54lWvkTTTV3PpG441EJ3IJ6oSsZUYOSWvK4QuFHhWlC1xQY9naVTJE11wYKJVFoZD
Sa6bmLuWMbBtz2+vG2auuNMShyPdhfHlOSe4GBT4jT6SqKu8tQSHmMWagQQjAS/xxlyAJ6TQ77g2
kciGKQcTcc+Kgcp+JKIl8lOmEOoOQvttwbHfLqMJjj3ZYhROwVT34cvN0tmYmJE895poJMKFqyai
CIU92r4zDviePpHL65sxo0k4mQ1njZY5jkwkLw7pSD53pJAYAJqFAdV+ebMa5YKnMIv4Kc9odcvO
4BQOCOd2Hsh2KhE/PUFUzu/7QIYQ24ZgA2YM75pMr0wN61vBYXeA2oUWgVvto3t33D+DXcDE/VRs
lKLhsNs2QKZ6h0L4fP7SS2Cq6D8Z46XcAJNV56QF4uasjl3AfE5uKRo3RzH4Uq9BKTEdfBYVoQIp
K2curEoT2FTtLXN4Moxv/tgx10fx/wZQTBJ1eAr1QQuFM3b2pWhopMSkI1BZwvo8ctjIe2jrhnVB
BKvsEBRW9cDe54ljzJdS/AQ1FaU/gCmuyYtcwY3zg8LTQ8dZVffGPp2ss9aiDB+Mjn03pGdqnFuz
wkA14xI0o/R5JhUvVl30hcPHRLIPE1MwK+YjcXvWblpi9hrEyqRJPvRfl3tCbYX+TCqvLaJdiR/N
i1cK2cCTiH7xNHSTbsPPkmqGnAgZYVp2DoqzM1vtuS50HOTGfsOmERAzwH3sLGH11Nw/jZRcWCB8
uocAjTK+kZ8Had5WYtXtQaaFa+0ENdBWE7C+C/RX0RoCSEeALL6mmHyQbBGDH8ck57dDQtWwvJSF
SuM4Nioc75EQmqFrLqpI3DpmK9vSuL4Lgk4vdK03nAXyYoPHKnto+wC0JSHLeU34OyuEB9TvZ7yQ
nMw4jXQWtXJm8By1Q20OSGhKU9HgYRaVeaYJ4Cw+H9fs3y+cVbkilR1HwzOzsxzNpFZq0XfBDo8q
Uzk/7jle8XgzfN6vcfQ15XArOoX54O4rsAx1DwRyIINs+MYlMc0QgaYCAMQbGZg4i7PDw+NKIaF+
VE8xyi+6zSyd4+eSBhSktvZh9Ss3iqzJA63BKvIh69bX3r+7i7lGs9V+AIWM+3XmN4+uf6p3b9uM
LT06y4VmLv5gw1NvZvxMeS5wLuYuS4bRgzdbjqtFhZ8LWXCPqbX8dCAy0rXhcUG93NbD++vGSfk+
A8GRaKgELtZivoil3Spzlge5digIJMI2nJcSQ2JZhL6czip0rh+M5RW0DPAyaUOlfDghHEeY/erX
+Me8l6bxGCczslAreBkB/PuF5SK9bqACtVodFml+uqCKFRTbt5szbm3MB9CtkeROxD6amDt9zcxW
HN/+vvoX7LTf3DxRoek1HXAoWTrDoCKvB7A+vmRDccxRnkLUSkGc3IJc8RyP9kyOEn1IlX75x3wp
0j8EYXIR6eHCuGqqYdYzSTlXCOyTtcZhFSuOx3TyQzfhj9m0MJeJLzrQPrARK/AQnBSpLzYk0wxz
wmQiVt52S8Voh47K2wWOVfJ+csHMXH3dsUHTOenhJ9mGpRgNHcbaBVAYN/uRnJFin2RABMYxSvrz
GZW5TjTMzvfCx4d8VD6PA1lt9MeaKgh7Kjk0LT9BdCVDczu4QNoILO6Wt0gm/VNZ51JzNNKqqRb4
Hm84A0o+rV6C4ewt0mCmNQwnQz7W+12+uhHl36tyO6wH93J9+O+p2wXpMt9HQkxNr+iWZHMpq1l9
r+OcV3GuZCVS/zkkaNnSCGXHakAJkySGB92sgf+uxp4I2ezoHGdvseH9u1AdA5OrH1YLh8cGY96e
DTndLSTjr9XkU8GjowpLjZlQrxlMcJZYxVjXQDE2rzyKUrI32B1xJauthSMck62eywihISFRA2C4
NXyTHzvEXcwOKxphQcI1a+XLNUloZV8BKyrTiX0Uv/8JsnSZoHo2K3yH2gpBA0OnowUcgN5K41yO
cb9/kk1ygEqLzF4mvL/A2zkaFpyo49pHOEYh++Px7iuw2+/ifNmvaFlbWJaJ2fvJI9Mr6XMiYzmA
RtdKNmrE9Vw9z4VR+Vab7s15TxGCz2E2KEqPp+IbCyjydgcoquNG3nlvZGZNSe60X7Ev8xdVltEX
0wrFZs3UAlDNFzISqPtm6FwzSJMpdIHPh6Ty0DEStjZFGSSQAyBVvjJJEb7mNuUxMpff5ecBT/RI
dayKz1CWl/PGsFnBUBA75kWGvYhth7RxEiuc+EZnypo2U8NhuxAb+tLWgGOkq2sjl855KL1kgAsj
sofOUWsY7pJL0QMe8dVwNzBEzvQOYaj37L+aecvD38Bgovq4PlotgzyeX0qXMFRpgDkAtqwAAsXE
UfyTxgs5vCzGQocBCp9HDKkV0LDcPOQYW1pIHfRVkb3JYa9o8BpaPZcT9gClAa/TtblEpII9xqrY
lEJfz52m+8oq5oMtaaGkpHV8Y/Q8fh9HB8c4F11eIC2O2mBRvojKa9sVvCMkaDRh2tkYlsT92rfS
cqtBSYkBgr8br7bOAq1iOegHYgTk3kVLbW0ZjcagXmdSjzL/djsjX9Z9uUiPnVSRFusisPsvPWL5
N8CVGOdTE7O4R57Jrt+TvnQtJCDKOzVEdL4irD+T86Pv0lU3XhmQP5I7hbu0qITGXAb2qePvis4m
j9yUSrxKCuMHNyMKfVMzAiHbbiMW/NNk7XFkRIqJq4fcPq3VTTg29FrEXlmcHz/5E2vfnuJQpwT2
a0L9fZkn0wVIfGAnMBWvOwt7NAOCMHC/8S7a00hcC90NSPKZAxOUz2+sxrwwsm3hXYOyym99FgVV
w5WjyAJiSPUPasZt6YhNHJPSB4xvdZ2XSbBHlWPvRTHS0EPLanp3QXce1Zlp+woUFMLTuq29V+ic
lRPNKEZQ1D6YwQPLBKXC8nCEiBzz4NJ4inXrlADHIAk9jNj40UFpBYEBZU0OWHWw8JUVeLnYM998
GJSOnWhVcnP/LxW4i2bHaHnSToL2vKbjjnYHu8E95O/2MEhgYKitw1NS19lQhG7o5AHbsMw2g4YW
qHpDa54pTyrBTiXwOWZFifgDxu6063v7lqDzaRQkqfe17w4tETjHG3GvGyd9VU1l9MZOBfz43XrV
BSnaI0hozQW+aUWVEaZpyvBLKXnHTYl5XrNGPopQU7+jGWRZXmNx5ZAjpyD8tSfJRYLPLSNc4YDY
P2r4eOdHGqMEYZsmFSdsItKugdIe94nkHsENdwgk36tzw81p013Rv/52B7tvtjZulrizoPnAybgC
pItJGHoC1Bg4KOkY3BYcyypFYGxxvHySeJStzuUyZdkvC0TFV89hzwp+ux1WdQ+TNyH6b+aeQMrn
nAIBWdrTbljoCSsXVG5dBlzLqJpSjjDu1HGJM/KdEJHbUzaQ9jtUerdhtYqpI4Gut/3mFZcCR7Sb
82g6CTlQizcV6M/WonrFDCeZpHC9o81IIC1Tx0BuRui1QodPIqW2TDxv3rJHn0MUWPG0xTRAc/YO
mAyfZqQcQugzE+HJ3gcBNgHOYyoB3tEHhMM4UKtcqA86SUdxsjPUvJPICUG5QtEznRlPDigDqnOv
R6Knv8W2RrMPnT+Pqx13J2a8xSWSEtNnodzh7mcRwJpIorTCHnc0lMxXUytEE/zMinxPeN/sT0vg
P4PpBXEPdwdOA9lO/hz2RCRlKkMliwA5L77ntO460SyaSIDIILXQ75JA2GmDacGxRk/kkYU5O7d5
YnPj3o/jSr5u+7K+tqB3M7VCUdF+mMCaDUUhDuf3jic+Nww0Ds9lZv83EQ/i/WhRUhdAEP1csIEs
T2IZnbJhHnMytTeDyZHRNRAPTP21pm9zbbBqTnow+nN3/bZ74Hey8G3dW0UbU3wFei0nyJlxPhw2
RVXgh6QWv70KTqaSdeFe+2uoTjEb/PC+KuFpyk2ILv+rtnOHHLsIPRzvL2pB8eTWNVBohRiWGVK5
l2c05D+VtiDbCzmF991L3NadGSKwmBgUBqmJiIWue2/9VwPlly6xqHkTpxDusYGPif4dTFUvKIZy
Gva3NGU49Klcmto9Swhkx5P8IZFE2t+0zaKFZlSCM8DVNe8VidRjA+T6cEQkNmJ3ZKq6auC/G3dE
Wr9r9QCCI2sDW3m2he9QmV6UnGr+C0ooTgv4zAxZ4PJDY3uknjoRHCsOEkDPWBWEsCZj4X0nJ+bw
Tn0/1/6Ia2J1l9ik5azUmQiEgK058/BQHDR+6+cJuOCX6j0nN33PtUBqA9dLjRyug3toORL+WYHy
KNm6OGqogq3mzcPdYcFK3dbKeaaO3zWD6Z7HnoBVTo6Y5hQZDx64ftmTUU6QWp4tWUwYzz3kheFG
nPK+Sh9zeykp9bpFA07zzihNBr8CkhZdVVi7x9jAeRAXo5tA6Hp+JqmnzeIlrCcxIBdvwR2aeJXH
QUBz+o9u38k86JyfRzf8v/lTtXZed6qfl87thaoxNH+Up229kYkZkNuSTALDYMO89hhXV9E6JLbX
GWX+IZsY9V4N3ZDR2cLY9yaJ0/hRpDOg1981zRJ37Funyfr/h/lVAB4tWLRIpFQaXUi0rMG+zyoa
qtoAltC1f30IAHyHt6ghytrkR9lapVZRMzTKAPk+CS3EJTVETRJQiSL6W9Z044uKl9KcS0gc90ce
egblgsNCW5FjiZtZJaM3C2IqK+4ddr9H7hlyJr4UcjEVJLSTcKj7j6D4VdGafzF0Xw3UFtH0HAaB
EnFgWxJ4zDax+0JVwE9MyFhmodjBb0mdsUCqwsqbRbEJWC7gp0xc4cOMKLx/dVa0so3PIcoW/A4a
ubf0A6vkaeHBgwYQAnxPJyt/Oze3owPfztvQwh4nQkYPk+mB5BMJV0B3OPnICfMPRDzBBFyAcY0Y
JK7rmQ4nW6IcUCBksY3Lj2nZnyK+82Fm2iiw6JntXFjqpx5RG9/y0iJ36Frbo8WOZWHYfGdC5J2W
oydX0JtZ6uiET1TXmzXey1rMyAIaLWeyTUDb0sXTb0zw2LJO4Oc/1YW782J63VuZDUgZ56aU82yV
usDH83zNkVdUP/rVZZS/1+3HDmhWy2g6ZJGb58I8h+ZGvbrtD2ceNT2oHShZYsto0HDbjxLdt7UP
NBHtR/BnhhH/YpWMR32BeznB0hq3ADgkAzzQ2nNd4H3C3jTPsXiRvAJf7HF8e8ujuXslFFmgFWJM
2Y2wM56fh8gVhdS36OeyoVxS+VwFY/D4y7c4l2TxVQ/C/CwU7lddrCmw/GQAkjApxg9AblPTcLuY
rYS/g3TiC9aWU9VfZTZDSPmhh/Ae91E+3g6xFfCKLgR8OaElRtAjtsgnMKlM06TsReuclx0mbxT/
cIWJ1qR8gYBBcYT1tXizlTewv3OF/5eW0LGYMz528pE9MhwpMqwrpWCZKUaP7vA/gheNVF8OsXnd
vJGgA01PxXaKKyn2zczRY04bzbyqP55PkFq/EnkN8c2H5OwCpyj80QHYSa0iCH+TUvGt48MK522Y
ZWvDv7qOf0xtUfAgFE5rHXGi/7CEyBiqgLRHMqreuKRdkm2Ny31Mo5fYYVLdr+NtTJ8hG+9xhMTQ
KMEVq3roDmpcMTaih9kquPJyegGY1Qnf2Xros1QXuALr4dBrgz0KFg9GJnceg3afjSanja25wEsG
Zo2p7A3LQYDdjUN+4tzEarbpGUM9TDvQK9io7UydnfLsNJdb3Dncc6nI02Ggw981BkgHOCrBdL3D
D2s9rqYozBrcPFu8A7qpn9b7FiQy38uz9mT1g5t4Xq95L8B/uqsv8T+Gpn2YbTEc32RHmUy9lFgK
7s6wnpdxbFMKA/KDK4ES3zVO6wBWSLJOA89k7xlQY/gl6KuPPs70sy3B2Ia3PgYIVfhXhHe3dRDN
jn7qQ2GC28ROhRVNiXIDoYUAsTJ0f2HNgklyHg7GPnhUK5bHsO7kmHsb11ZuzF1EzkPwNH8Rm3Ow
Kv4UdJkLlvtDzbVwfFk8R3+egdJVdSOuB3q41NVE6YulrZPO14vy5zZcgxOajA0LtHGrOUWN+Y0E
Zraq8t/wDqmAZMZ+ooJHBrEsPO9qJulavCEj2tmhUayUwFwuLmNEtzn4JngHHIb3O6Odj8INvvwe
2/dxsOcXRZh7EPw13EvErIA7mvTR4SXFmSkAUCyLsBE4PZcv7BafAIT+5mPecvGm8hiN+l0IUiA3
KtdCCGTdXtovSp8XIIfuHHBrqrAPi4HGG8tRg08EYBxCIRmxj3F7AzI5D72cyVSKTs8GGY261oqQ
Lh3V5rOdnDEJEAGlXFO4/QPtr5XZF/SktPeYrUHIJRoSv2Bp9xk2AbfMSWjNg9oZtdqgT3qHFsb6
5vr2NRrklmwE4LoIlBE9fmdXVhJiDy2pf54SBBMLpGNL2E7ycaiBLtBoPBTxFMFD8eevonfa7XCs
qUREpFD4fT4Vs21yP/skDWm5omxChOnqbP0A+ey8Ircv5YHGN7JQdwI7Y7bIGDkTtOMEjI7Z40RK
72gWAMLH/De3ZBw5pBSTFKkvqCS0AMn+bZC6vQgA8554sHbdo1Y58eYdZxHdE2QFjwaWAQMS8c3k
u07Axodjq/Ldyn6ymfpfffdXnNHx0VUZoyrmrNw5DDhssXZk9OgNz2n0+HHZkehm7yMLoQMX3yDb
V6NYBY7lW9ZJW8BY4FiOKIEjQpD0LRYh8M5d85z71dPphg+iGan796xwad2VgzhVXBwrZhNmp8kH
+EsO0c26E3pKIedweANoRtleRAUXGbwbCvNW+dUpHX+LZFr2cXPgDdIi/2AQh3radvPvssP2D1dF
ZwrjOAg0ynvosGZrXzVFAI0iS2zdt8DSot+3avhev1UJiLaZ/k15uEdDoP8N1XxDOOPdRqPK96IC
8khsz7Is7aPRqTUXYYltvevUgPgfukO1V6YAjL0WP8yorAdx7yWXY5gx6n7Lv7Fpka6hn1g86tVy
MqvOqbV4o839h9YPQSO85xgpaLxesOOKkyOqE674KRsZ8Mfxdm8vbP1ar0QAbiidlJuKlL0KZfhT
/cw1hW4RcKJJeqDAFSNbLjNtRz0YnrVA01Kz3V/ldoNFbaw58FL97NBlq5qJIA9FuhSKr9S2gB2x
QXc0gXHHjoEWxrozXSmZf+vOqOi6f6Zif3g+LZQTTjnxPz80jqNc5qcqxW60Mciag+Nscpgjbhe7
dVZLDIXlp/iydxyI0/p6evk4iRkLDPltfLOmwwaORmyFsd8+W+rODGngcmmbNtmiwjo5KxrRPLll
pOiZMMEKmew5q5aye5szZyWxlVerYoH5S0teILL3Crz5SW7k95STqPhAiiGdFqqtipK29URDDWPf
t/V9QNsQq01TGq7R56LQmU8DmN44IzYRP/vwZr5WmgluzrcZ8/dGgOHTaPIVssEKAAQ9bbanTw8H
hfRs6Njrb7Pig3xFtUvWufebBVpN3iY0/AGUX4BwUlEeMjcTgVlLuBQiQ1EAyRHwoEhJBvl9nWVI
44FtlRUTq9+wVFyvPGpMCK/0ucwS5+5pixJ8F3lBoi931ew1GoxztRoLAylL2pqGdJbIJ1HDl123
IHav4+5TSIqh9rq+ea4arQlnbT/6UhwycNNCpBZJKg2ETYy65bnx8kKuYkXH3jUwtzFcZ/J6Jm89
6W+pOkrpS3Sbu02Ve5cy5tvy5k+lkzuvdcFrZFOwQv1c1KaQ6Rv2kMjLCFdl8T73fgDGh1Wwh/iz
uANWiQXOoW6jXy2/eVgHiuCpIlNwYPqo+imRE+VYJuliBVvyg9VIopA0hHU+z65D6BiZfZmaDW8A
jgqITnRz0U8Qts43MUhXi8U4oECjkubsrqteCLhgH/5I1gIqMYIv1JAa76ieO7uPpjA0Sf/EXKpM
kEgno9eVLreZLZPhCix9XKolQvCzkEVXG4ZtYlzn5Bl/HzClLl3O69HL+gEACpFSxCT4EkC4BY5U
ctwvQw+wSZ/xMDb1lLqJnxDxk3LVscBQUmiLAVBx1HiYMROmhxfANHrjndqN6UsrFRjSogD+a6nT
2tECR+qbwBWYn0efMNMA/I/AJktyHATdNPqU/XB0KclI+zWeFmSgQijOkfDk7eUCqyUtq9rSXTS4
3yvj9F/ixolq5X699b702LZOgx1Lrx1Ihvatb1PMgZhRjq3cqF/5EIZWHFMgHGqz1+Xhgm8qtBDo
envXInW2CukvYmoXkq0UGGZtfuAlM7ciw1EHetV3E3Fg6xaI1/PJFtjpDdc0dW/y7fW2zMugK2qR
iYajatGJCntdb4v9U7PB8/k+MeA6iiiCs0LpzmegXk5vSczPvnwUshB6WuD39S7r0tFjOtfMJbah
Ys2nuxnjB+FDupXHkB74d2T8dN/6TIPrg0SClsiBy0e6lynovv/txZCvDqmIPpRcHVa1WUNekJ6x
d4olKpvQ3IlUjrT5kA72LvXmPKT+93d9Zv7TkgmO/3v74/NjTMeTIPjzpVhFLlI3UWYLQXOenGb4
PpP5F+BUD2hov4clc4Spy1WcQC3lm5LzQIv9phO1yt7co4afzd6C47gVBLeWN1ABK8xhHK/sMNKQ
XgVMvIy+fTJseJlz2zvTZD1ODfzoTjdORzJw9JOlI5NIMQoUG/VbjkEoRQjUee+wlt8mmc6gEBq7
+Z7BXhV7Z4v3g1sg/tUE8g262NiRdJGfiKj1rGnIgkt4xnpiQ5f7kEn6VQFIvH9kyDE14BC44J+5
YIldXEOy1MT2TW3Tk4xzPUjw1FaiBbxcz9rFrFC1tROWBZaXHunrXCts6/GMuZFhZX2G6hTRYfsM
eGoRR4e8rs5rxjZ10kTC9EcAJwbD3X5voLdQL37iU7dKmr7S5VubyAhjtWtE+mhIIcncAWhqzT4s
JC/70/4glHjYVEZH4+0bf/16KyxBL9ptkNIMzEJhabYru3yPG1XR6sZ8p72o0wr2AbWgnv38Uepr
Eel45EXG4qU5EecY95wbZ/9y9K9dPoaKhN9Re8CV4vtif2Zj1A3hBRfX2yZu9gqHbqhJ6f4OmNPl
nyOWBzlvOJCG+2hRsfgMHLymKh2cwq8i92sLc/MASWUgIKRtG8lVj+w9BcO9oxFraJqb86PqVVBt
71tbBO+3mXINXLj0Uc0X/c1h0bCCVr9M+H1qKh3/doSve/AeclJtqKoQVnk5TC5rQSxWiKOf05oh
LuKf7/UqWRDvoire2Mh412hF+NOaq2iSyqNKrQCq65EeipONhqKyZLHeucp3N3Rp1SmzT0SrsZvT
RQTM4EMQLKfXwH4MQpeAuIJKrvx1gkH2QiGFrmg7DnCddDm0TVoP8Kvv+Ck4LjG2terg0sTurdrF
hQv7T8ausY91KfsAauRi22Nb9p6Ha82t+ZUQPjhqC0zjhT1KBjMwJ9CU4Gh8MUH3HKL+wCXr9pBV
lnqtPCsYylyq3rgn66aM0fWWCK6faaG1H4z+Rb3nuCJGUOVDY+ZvkVK103GSDExxVaHWEeZdX2iK
KH4wNiboMyLuP8K4F5n43S3QhI0O+9nTPGJ1JF76YQx+uTiswgFdAH5Q5Db5nHEH+UbSpFdHXJ8w
OwVqrlHTUe/9lbWa/sUCGIWfiiCaCUDVFiu/5LTPva8yugljaI+TtCKwcxvXjpsePT02VMwACopp
njLyCHKIVZ/3wzIpq87LOJP6hKYG1o4j05WBLpJyaFcpNNIAIAYb32URkSgA9GAZWpuuO8XTpplM
WEqnLJmDZcXWR+/E85XU3aqqdyJ5TrM6xgJQn78FXvjSKdsuWMZ/ppa7316aLK9DQm8kVe75oqdY
a+moqMiQwY/UbpG3yTBa6NWX3FBVooi0ajF0T3C5Us8QApwn8CUrAiwzwbVxnVZuGwLRZ3SgjyLj
QcrLUhKLUsenHsdFSnge+C6JCns7xXeegaC5gqxcanT11XkdVvYXoEJpFxhcmd2pOn+ntBXgSpXP
PuZU1Pjj5A4MpOnaale7YL7CkRmHXNNS1TP52Pt3ZC7MCs/I3g6oFHWGVbvVmsXXFZYXDoLuBjWp
8AndcQ7FW+Z6PtQ0cXJdn5Mfk8LpDSkdJLvsWneW3c25bxo9IOAXAzFruERC7eyQt5aMuRR/gJlD
SUni3iZnBQU8eFyzLbk8wM8jDds/C/ClCYWEuoREdSskwqlT4k2YM5e+89lg9iLUiIKtZ2QIlhJz
kZf1mAbwimBLxOKvn4Pxey1dUsNlo++HkKP0XTllwS52rSilabiKnWodSuLUGwxaylgbE1abKdIh
ZhCd7e+a31pC+ro86LdNxmxi66YCvDxtllXmfbCKFuGqxHeaI1+UCnlUdQ++MYedo6VA9T01X/D6
YY9r2cm/c/43IG0YcKoCYxQd7gMUKNB9Dw23RipYmifBfPxNL/gHG/RQ6GtE3S86aHy8AHbR3JwU
xRCm192d00/tTi6kC4VHy0QWlqWWfOX+4ySyzOwZofD5HVCmmUEfLoG/T02vpkm4A+eFjNesyVGJ
VLgZWouFCW2Y4LknIWqg7D9XCIwzYfd5OQlRbma1oTDnMiRNeYe9/OTP5rRcpdYKxMkwvjwjX7M+
o93PRdW8QDX49E1EA3sMtkJ4GzdCKYz6K5PVnr5jj5nNIceGerD6iqALpQUBRxozTphv4Z+rQVoc
a2/KFzqq+c0/tTw5p/BPALfjIGc2hOhJDcb7HxxumrK/ZJpuLeI1r62YfK6U5EfoNMnsTXUu2u0U
pT+xdoSMhrpGdU2Rb5twC8E4P21p9UPlL6bxeZqGUhilAjh4wQVX+8UNRHlC92tngm+WsicVP2un
Fy7c3yN8mL7wnRR5076c/WZCAKS1aEo/GLX20C5zu8yWkaJCd7GLRCni8XenuLJu2RqEEpgaFNWq
TZI9+/TphEHCRTAoXyHW81dglgSUwMOKIMaJzclFIW6lLJmbUr5VFm//CN3vn79W2vy87xVyMR6y
LD3H1OBIW1V9SAQhpwBvoz52a3znfb5m+V05EYqUzxM/jtqhQA4CNQBR6qI1qlskeSfoWL7rCmGr
uqXhH1H9lSlhcPez4+PxFnDus9myd0Y0jwUkJ/nJz6XN6Umg07penGlTN2I4aIBEPLh5fg9uD7Xn
SbHM8fflPPC2RDK2+Vc+U6611MBr85uiVU4kJaCsegS/bwAQNxsTnzebwTSXMUKxQkAT1uxr5u7S
TJvF8HTbcYf6MmH2Yse1lGsYKQYt8uoPTQcA2nnnJsd3oP7Bw8US6q/4DcckZBndRiULjVUykv80
xVGKSr6NMw9vyx26gBZtgfSOf7Z3l+sDNAn4iE8OJmo9LKPNQYQmWJkUzClH84NvZTEPRMhC6G6Y
cLqhCB9KGHoweS6s1MNec9Uu0gvti+Rz3C/wK+WdtRwNzFWtYVdiAB1+hGxbOQHG+uN6VgQuCPnp
cbRdXHtRnZf4q3tcrD49CXq/+Ydyo/QkuXX1daDsfBw5j2nYNnIHAS6VLMrLyQ+OOXBNH5xz/z3f
WxjvvJbuOtqF0tZS9BscGqPv9aeSbYmDRC6r5TtGo7CUBFiyB0GiRWdYx42rWLHSD8KvyUwm+DOs
FR/xJqyhxYVYj0n371b5yGf5/vzHEgUZT2auHSfh/ZryCOa588NjePbJGnxv9vf9+wFUcUSPONw2
52oUSKpphAv87SdLcWuRP8AwXfa7irVjKAZ3VX0SEfthax2vOYQcCPqdTc7P1VcI/dEVau7xrfLS
6aH+62409gMgyzmsgz7WyM8ONUgY12fU3uoRSXKOpOGGmToMC2cCs0fo0iGxsPLQ2spVHqWm0xq8
s7aJMcU39+HKKJjVM01/lIjE/KPpmAZy4F1c1HfvnFDflZBLxG4Pdxk3kgUYp2HO/6QkYgiUz+QQ
8ldmEPIDTavXTwOIQ0v31rBFOx86D5xHz9eq7qCeNnp8OJMIV7p4DjaQXK8QShxwUr/+m0ijsmwQ
1w0/WKf8dpt0EUXSmJjagiQIYZuYslFqNBXfff5KfO8Su8hxdkq+EWIDpJqdPICmT+Lxx69L8XYx
8VEgokhyv4nGEjm6/h0NAIE9eQUzMUh7z22sZrRQVBJB7RTMklGxCU9QqGYQ5la4wB3TIJhdnGtU
PztNZ3W7ZC01GRrBi7o1p2STYxgobnCVbvZHoXsfnVU3YOniVgcAPEfArBQRZeUJUUygIL1odut3
/4MC3wcoVYIPOK17M8cEUjlm1PmDHCLTiKTjl4PRBsu5uN0syHADbL3BQsceG4Mo4qNIB576l5ih
m2f8vGMEqWyLbMBR2cV45h36auD2eSSTaI6wO/WYNYLBaYHfGrSvL5bxxGBohCpaJZE/ogxzT3Pp
aMMiL2fvhLJUKeTHqKrBl8SjLL4Pw3VEpaH5dOegQ2SBTUPIkM9t1lSmrMwXl5wCQvQQdOrBx7lu
ohspA6wUpPUwyaFcgKmIB9SilfJtXZhdokkxI85r0VuTZEg29DipAHG7J7b07AYd98+/aqI54dAE
rOElyRKtl3mUbjOGoGFmu2Wf/TXh4KFYt74myD3qqH2oZ50FfQo3AJb0OSWx4+OKVa22O561J8IE
/Q8eYhPxwGPKNxAcpmXbZ92LdNNAr0vSOgYpjGDau7ObUCmV7JDdMLwftp7Zq4Ovrm02/OOyuDZy
dSFBddbOeP4IV9td0Vy7Zs1VJxH2D+S7EwAXlzkSE4seQJWhYDIja/uNgc60EgqLqH4SKnnAhxxd
Up9fUhwj5cNqxxMU5jGse2q5QgsyiEBgypBtuOGWJTn24C2UyIdJK69fF3ZibAazD1g2XAyZHB48
3IqOgKyKUp5M6P3IFYxWeocn8HPzSS9DP/jL1W1YX09QOUBig53zEj1cXwFfOoqtCsFRiWMAJdP4
iyy1MIVTqja118p6mODLkgRfUZqQ0ZBFUnSq9JNjfdz7IoiAZ2zndHYOGIBGtaBywjvpWaW9UO5b
X4T4h425pOQuJY9dzuWW07no+w8IbORbqU+jKnyZu5oFIrYlTaYGmGyE4taBs+OYYFi+Rk1hK/6K
jXGfH/SkjMD61iBzoxv0WrAbP4eSimWJjeabMnNJQrZHIp1Jx43FdHiFtDV1H6FLQsAo4x3I+VxZ
SxQ9xyGG3yMiZidhCQcNJ6DF0B4TujNbLRSnLOmUp79Y7E4YLktDgcjEHlF8BR6V2Qj+Dj4nyNX1
NGSrPL/IJuTT99NOMjlGPrjBMJtlpk4j7JD692ZR3kzXzjJDReLiq3ynpsH+etI3ePAP1ZsrF9cI
CyiTvxRzX9UIdYPdOJp9gtr7ky9g/5+Of5/py1SmGkl5Lk5YdCCmFQhrKLs4OZgCWcR/CzZEYpfc
2HAnxa9vWeNJpZm68ijQjPxZ3jw+j1WzhUJZxu9blNgl5mKM2cz1iStfs9k29H/bC6OaegwdaD4U
W0tDqh04wKPTybNL+LJOTN/mX8WQx1qJ2EoeTNqfjmjpxGgZeefIZwna/EBfW2hXpc5vTxyigb54
RXj//Zei
`protect end_protected

