

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
f+/ctYELc+/uhaDk9UPcPAJaXSQFIFZYBG60J8h0SeiQQmJRXrJaOeV3KVV/lgxJBX+Pi0uIoqsP
0dvvt0j0iw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ds8RnxyUdiC5UfagTnRdgf60gcPiiViW8hDU6PUQWVIFrIIkQkMyKnNB+w8Xr1qLiUBG5r4bOXXF
mErwm6JOoZIoBsQDC70o4vSL+APqLNFSv5xXApMJ8oplAbqfUWw9C8nrRU4CDut124eAXDPI5DeY
2JfMJZphm79HLBxzMU8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gRwcpx+s+b5LY0O8TRhmIjsPjqA3ufiQgXkVCZguAw8Z1suP9nPSCId7/spln53+f0/tJLCzfQ1D
fd2IUKNHJ4CCwxe5P3bfYOMwQGcGZYBnUI/rkBnbT4bLIULUKjdsdYIiFR4wj7A4r3rxdigXZASj
4bAQCWc/yTKuHPdOBkGm1xZsyE/cym0RYZGZH2+fxwCmec/mDDcJ/CpYhDoHMGEGbuBCGf8iBLWn
aeyZ9lCCeLqu6wdaCdWUNa54o6ZsntBpsV9wCPDRe9tE11ovPfBbXxn53PNK8XiwXSYMz8pn8OSy
qxbPTzZIACZ7R0Un42f8fBUIWh7tpxFHWyGs6w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nodK+3l/qqYipAuhJJUe0xOuCIN1x+TqZIbzLctg8etcdj4ns5ERwOiFTEWx4tFqSKSfiBrufhKt
yWt2sZ8CL8QG4oFnIznolrRNIehCN+4jyWbaGXKftDJd79ZqRspFhHLhD570bMSvSIgremGXk4v9
8wwP6uATc/QsO1FutHGO8KVpCzxvZd40lViRrR4PDuVgDCY+40pK6HkXuChY0nuCRXJET7H+tUta
9E+x1aTzVYUJ/1eoCVtOj+E7tu65BsmJ20dnWEHkyUeV1jA5W68X30ev0J7Hs51zJ9IR1Tc9k6oK
5cZGL67jAoPWt5mM6t5aS9518cZBqGf1oNIURA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
adHuDdS9NIcaGcdK+qIYLCeAIhoJ6/aK/3inFss/KwS901WcWdnwodtJYRl30WeSk1NA3ccYlgcP
qfRncDaW/cXj0qaABAOnK5VGPunMffN644DRlXhECkaoA/ySzb65JmiuN2S81Y++kCYraAnkSn1r
dHyKSUgx1u1NAyxKiVY=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sq/klSwJOJjlA17FRdYxJ+Jut2VAUuMuo7xqgzJ1RKtGf6HYfMcvDsg7H1p6GKxKsxGzQnDq+TV2
yvialaGKR25jq3m+YqEvu4alVvAND91JWodFLGOnQyQ4wOlFINcRBk9iV4KuRcCu6thl6yqz+fza
9lJ0zvBITt2ks0M8BRMww70MNqtNWaJF1CC3Ni9vAu/yQQYVeSwkcK5UOnSxVuhiH8z04bmGbmYX
GiHOmU3jVuxhp2YjqPgDzrKbdsoqJhjCq4T6U3d0hobbkU3Vp5CdZdl/0SDjWcHHzcK62so6sjkD
SzhKe/etWPbsSxqUReKLZSO5LheXEkpPy9MNTg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YH2g8ybH0nesNjg6E7y8jBJXn8tIKyyE0livQIx7Re10TDRlzMmCmwkIUN5tlGSOGWmhLVQbK0g+
rKcGQQ14ncV/D+goyDwXomf/CSg8QBf4hEnCO7AC7l/rY6T9MCzXDi91k32Y9rgSa8psw1rL2tRP
V4n7LZWwLzpfKD6nULSwfOxlRujBnhDthCpfLG4IyGF6xIvXwGHiPKj7eN88s6/dLLx+cbAaF19O
87YX29ndjw5p6GNVK2qmLkTN6PXDG344nzObIwO0uqqA+FVVCZMMjZTL8g4waFPmSoYkceS61wYA
ixxKVaGor3lvI/QtRPUF1CQLzsC2AYuPvMnzBQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jvCTnMZdPEi0pS6fvoWdHBB+8zNm548wh15gSC5pcwD7WN9Y9MGIT22qU2zoAQUCxDDh/cCPO1Yv
ADLZ0UhpYD2GjpeuWT5ghd4+qHg/CkzJFC+ZVH8ykfyN62KFE3xh/MluLBCWRsCStmZJ0WYGWgUf
Z9tmSszFQIuvHIcpusuomjakCYe158ViTxw5O5I+Q+Pr5RKTSyOK+KeUwbQzEyKFWzqyleebXZA7
oqsF9JxaiyEYCepL4kzaHuS0svOYXFReS//cViwJO3phQKvtD4kTD6UUO/VVfK4cTr/eE4lDEGtp
k+LKlNS6OtEasR8I92J44GiANgTY6Us6Bt15Cg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j5cGcfM8rqCCS6KkIv45MGGE7qR/xEFXp75tqUY+yuyLI98OR1gm3l5Igo0qt2LRcoEg4D1RNKOw
DnWeDNUo59EbHqHfiydR1fs4bfaSIqF6l3H1RQsLZBo4sI2WyMxSdByFFTGLb5Kt4TieIT75Psva
0GuLfhX8d2PRKhvO2rSVTOvN216IDzuy9UFfnJtMYeWnnhvRl/5WRu+Sz3OJbchfQVN3Cy4DX/Ni
ldwRLsO1e7pref4KcTGOk6rS1zTD9kPQmMdDuzqm7LeBRJWqvQm4c6gjU0r9BlEjqOi+Cgw4lVfF
uh1OgQ+uFd0WToDsc5z2+TxpMOrfyQgACWae6w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133280)
`protect data_block
DevXAZp3iOdVaYkccBS6vxHXrSQopJgPFPZVaC3zNfbGHPRmpU6obApAUDlE136rTstMNOCQ4SF7
LxhtI5lmRHouowxVca0IAeEw5zSVJkG8eEVq1b1YKgOAWOSF0FS0flN/i8b3Y+8JnMUuD6jgSbkU
oMUEGTv2DihLGdtr/LGQozI7Kcx6jta3QKNVSf+lweOLwtMvZGZ0ujhdi3oTBUzi7eAzUDXmY7Dy
gowGVwRTqJxfvqD9ULd+6VarWl0W8k00ZNCnIf1wlSonF5NDIkaWsSPJfN4xVO1zsTZEMQOALabS
SWkcEhSrwozTlgfBXfxNznqyb/GIQO8Vi/N2gLMsy3k9vabYadxTE7tS/0IQavFLICHXCb0TXe4J
YLvxJPkx7DnMhvdTeDL+K4uNjJeQSPR93uYz8qwJP9o5px6g4372hyo7jlmfcg8WkSo4MjD/KT8r
FnyLk+xysOMPcDfGnjC/WDjS5/ncMJr2+iR4mopkM+NjUPh/88YegnItNTnNFRGgmGL8Tg6qQa5K
+o/k2rMY0SWT1Rutx9s8uQHqWFH9aCjn7AfohLKVbaJq+uuwW8x6cPEpqMcVxlvPEx9dzyAtnLbO
uG6a+pAvMYEA57S6K34tjTmJmBo6GPNKUIyA1FHjZc1xphQnee4onXwKxZeVpIEkNNPIT+Sb94/1
NFg3hW1ynk70N/H05XYxhxrCJVkvGDEusZHpuJqXTS5OFO8tudFR2GwWp+DG78djpZKVVAnupZqj
B8eZtb3XAfUpk/DKBsd1LHEQSiXlKN4F4M4SE7mBZdUE9isGckk+C2k582tfbwJREd//DDoZ2QAE
ZsZR4fVcmq3pa86Uixf7vLcrY6RMrIYh7HGSeVRdA2mlTaYKW+UVwIffWri8m2Nyw5FdAm4Sm05n
AgbG9hCDE5amQAWHAU02dKIC6Gt/gmSWgtV4W3UZYXDM4d1dqalxyrfPRY+szZLZZs03F9uf1ddH
W28Sxh+mjhCTFXP69CjTAW3Sy4rAdW+WuR6BbN3PFgxmLcscBQ0Emr4+En+hwEVu38y57mWNrLXG
i9C3xo3TcYDWNQ2HkCVuaf98ZZZMYtNrsHTjq/ySaidq4Z+OovQun4M/L/8wPw8z7ZYHUppkaQjL
uNyRl/HwWvADsP6/CYGPbFOVlMCEcdG6FRZ9PgQZZXXaMNVLN+a3afCRUpYb/tS0feLOv9kkz6qM
dfquMDDPySnULtB8pwz6UN3UVutsnCkrEMwTUZseqagbp9V5GbOKDH72fv5CVheygBvpx3OrSG4S
Z45y5tsxe8h+uHfw1mZbsVymiSXwSd+4J7GJBtJel6lN3SaPsGoZquYk2ak2PHEhuLIOptCXf35N
jvaNzo/2VtlQJ06jtYKTztd8O0NESPbyibgMyzQrr6qdW0+BUoks4Qfb5hU3a27tE6t/JxcMSAwg
RXYIFNEP6ssqhJKtiik9bijfAHR0IvOEVNuxZUT5iHlenx4KmTV1Ui/RphnHak3eRD91nJJcrG79
SPq4FXObST23fT9klXOUby+FCS2lPnkumR6ZRs2TOu4e8ijg9bAU7OwA/aG9sJDqmknAlzlWRyUo
gyCVmmvI52jOoN60FYEfbMo4H/eIPAzDUbGv7ib25EHBzPHx5PjGksGwg6MY2FfgEjhyvlR4dhuU
25nZqDxdTPowXhYcqX7LV5ZyKKwDQyX+QiesyiCNiB601nnl0AcoY73Da5E/7zELyxR2LqbrmwWr
Adwpc+xQVa8I0FBh/qIHGDx3BaeIqw9hyAmALcukv6SM5XQ9ysv7jxjVvE4U1sf2kRQ2DoP1SutR
p493qbNXD7nn4yvzTELH3gKZ0qQv/0xsTcNiOYK0cYoErwl5Bz+ZYxBhoHiYnD3PhQFE3uIK6/np
IOjDyJB2/JHYQmiNWK5HWyeE/ERp9lU45lxAHhr7dY6OnsddxvpgbkpyH4GT0Gw2TEUdBv1wIynh
sJdSmT95BjDlNSnslO1vR4wco5YHKyGBoJFAFdHKSxav+RPsEMyWGOQ/ofVY2s4QF3FUwmij1S9X
6H1bwF6DlHvzmNpbrpMTCiqOu51j1CbXdixPqVRDF02X5sl3QpDL4TU6QPWnyPQscwh/XkY7gAgK
19KX0KCR/pEaAOyNNKKlFsvjL26FhnIMhaypwwRadmpM91kNonu0GCGs68ItshkuiKwlWaBqkT6A
LpbVTwXPpjp/tJI5IGQjSEKGLLwxBe2Hp/JcJijx90NIWTuMwNxpHafa4+ZEPNCfPTP+HFeqldpO
KMXxu3V3F1YfD5cYY/e5a/PADnOOmjUuxj6E9GwfEsZhVy40EvwN2NIkDaN5qh0abV3rPalAh3/c
pPBbPZYy0/IOFA+fuNsYIfdr6KGPYulvrYXdVlShWZymjQxcqmgObWSKp7v4pWANIs7PmRQTSD1W
U/uhIT9XlxFHYwH1w5ZbJCvsGTgrOIkzXHIXYJ+sRqTd1N+c1cGTrV8yLW3hi5CL0E8yzWmIIqdH
UHKa0IdZ2EfXGRdiDc30Y9eGjSxncet+RMHHWl9NQsFs5U73o+6qc+QinNeBqAPloxSPkUNyEib4
T6wY2CSO87Q//f1rDK+5FRLqxhfm38Y+H5zG9Va5iowDyBA/epSDoMKyhMmUOZ8erCuVUy3SeGmw
8VIXOglgdn8oL3z/kQ1LHRqvOoBrPl+DYZiOy83HKX22lfv9+h9KfmIJipJsfSajsXmTscLYKHjH
RtKAtksACusyyg/Tul+OXzDqLUtMd1WSI0I+9nwO99pzajfRbuLFNADd83NSWZ2jqzoH3gaW2utj
Bf2/nSpr10Obt5zu8NnNFhhrOsfUjwuuvL0Ubtc+uGQKvpGhSciwawcex0DhxWFNq+wIpgA0DWyU
CKQN7oFNLMZa0aaKg+iTYFBx9TwdlxUbE0xAyZxdT2copeLeNwVVjsBVVI9eTlSm8Ti+NFISC6TJ
TATHeiXS+rLTeI33uB3EMivamYyyvXl3OEG+SE2qlAPM5JjkLsqT8VyD46Bq07biINxgdlO32pFl
ygaVslEyfhXbYThhgoxYhXeFNUQzyFP783sS9/LocfQtRo/67ulyED5LM+rT2S09R8mulymGeSkY
N0LlFR/GooJW+BqSQuKMjvwGV9exa6Suhw5LeqbilfpjnnKwfpR9rTSLGk0UWt9hx5E87kV4bgbQ
v5ulL1Tagu+USWU2++HmVdeIsockPNJs5OlvN/FxXy9dNHhlkqu1IyC0Moo5u6PDnqTNxM/u9seo
8fqCzFGmsijwaYzVmZmKQT2vbxIjUS5BSV7ypBn2WDBoRxdfLlxIxaw5eMMwoSu8NRIWzny+c672
Jr4v2fuQOxBHw57+0nTll75mUc0E2AKG32vttjbkmtzSrxhnFkRYv5ExFSe3tf8+6zHekwFv8q2m
R16GqJSl09ATCCT/2pmb3iWjnoD97AJcNGJRDGrzV19D1T2zVBPkNrXbqP049KyNJG29xvxGZpnv
OmWiD3U8twepPKYJMsyAd/bEdAxPG1V35wjf8C1XD1ksmNN3VdPxMlWEus4OqVBplFIZyaxXWSTq
fKkyEk0u8/qBQLTRvo+VXXR33QSyo4+E/FnVGPlBPz5sClGhSD3ReQWFCrQ/YOuGsCj5WMtD0Rkd
3o+o76tF47V9xOYngwhsFFJiynog+CRpNqdath6WZUXZpaDEI435hP0olh4F1MarIl/EEr50t38Y
AwQy7GbBHzSv7m+E2i5CLS2yRLNQamiQCXbAcXcUC0kOX8M6gbb9H/53zPy7duVFk9nt1aJQAMrc
LpXPups924p8yeL3cEk8Zctxx36LZN8Xt1gPyY8Kq6u0tmG366/e6bBBPQR92sfci94nho3THVZN
mGv2kqGRI4fv6rl0J1hL3n8tw7fBgEs1KRTWaxyUKLcuuqfdR2wfOc1TM1oXP6t8aTO8JRxPbvFK
dbUMeNFLnogd/fMdzj1zCX4kQpnASGoSZCfufT+lCxpfS+moifu9feegJT+S195OhhMvyyTkXEEI
+Mcfb7LH4jU6Yb0hDC24MhpPBFOqJKs/YyWm0u3bb8toYXHLBVXyi+B1vXYyV1+ci/6azpYkV4+A
jsFFld7aNNZL/RqiCyh3PSByccEyAWlrHYiDGHQmZD+DGoqqVtroOadiDb+tdot6rxObsoo+nGW/
YG8qgfJc8rcl5h7jzibfYmqcueH9W4hn9eA2RG5H/RPpJ3qNPMOxubNvHrg+ERM3qLzdGyzM2czj
KVgcAfXnTBuHcKKJkd+O06t0kaljtWLSZCdw3GkxzPrMn6e40BVBvA3n9ygfkM3sN2FbaqFfEuyh
gcWfpxPk8JHt3U4m+8AaBQMmeqrD60gj5AfZvGtAug6s82J/TUa5tlIJ3ezGYpRWEh9hf16W59mL
DKjBaKt634XexuiQphCXsMGiEcVw4nj2V2ijyu/PjJuycDIJhshf5tvfmGOjR+OPSfTQ+6DtpuGM
UTsLr4wUke9gsFmC8P+CmoqOVC15t6KtXZQSm+busdnd/fNin6VRmhM6ofUB3BJcdNRRcyAJpUam
I4NFoN6HtTjt0Ehr3OUhdH4t0v9mfAKVBtpxGKCkcU80tgRN8ysRXMtgaDSugCqXBGciu7ceOUa+
NtZzhREs1MOoEd+TDejknmxCE5QiVlxjOuAB6q11hYSJbo3QXyNFrLvJmvjOR5mzTRcBgkP+8csd
cwblX8a/AvN/1iDmddLUwqssctygakgz6YUGcZcolgKGJEDjvXF5KbwgMEejw49Zz/a37p2TKRtP
2gxV0C1Git0aMHuwj2ddGnSUUS+14y6W9eEiccKYOQBIzdlVjDn2ErKU7D1JhVKork1Cp/+QDwtY
mGiVmNizFoYjGjyZHpX78yHyr7pJkZKk5J0qOv21iFqXxHAWXWvJqSGP1xR3my/SNbYNf9CCxkw8
H2KqLBHO+vh4CggxjtX0RaSmqkcDGzBV7Zzga0x5rjmJlLxxDDys3QNxobPjEQ3xWtOJJPxQhZKS
lWoBv/BSG6tpQPmSPnkxebSImloxBBem5AcjXcP17gCvFA4xBoLyZxLSzgDWlkPTtP4YIPGQtgmp
vL7JEzXiH0Q7nip7WQqcHLKVZAWPT8MiBLnAcnDB/LNtJkgRAnQmpVB0gwTa0yf8lkLfbwgBQwr5
3mR2Etjw5DqzS8x/XwcKj4ljNaNP0KdlrX+ieFfF5c0wa1bCI3CEL4P/LFJF0oHhuxnZqD0Ypdiv
dWPMXgzqWEk2FpLFXykurLT10mIM7e0EKhQ/xYeeiESHN8zgwvyiDGuy7TzdyYTME8JvxDLG1Fw5
EzgwH5GzqCjeyz2OkL9lfC+2Vw+6k3ql71jPwhEAw4ExHqiWXh8Us3p4OdR59hQuOsW7a8LwSBML
J/g8kJAiouGZDT4haJ2035nl8EP7h7gGMWjmJADndEihbC/8blZGA0bc2lwB9QG+OuGEozl0wCXn
QfdOWuDEkgvFsnyfv3+3d8FQrlLm/+0PphlDdBZHTmSIy9EmRyTJExlIVpnWi8A4HTdaDAhV43Du
Z9EwJYuOOmkEV0tE208rA+H2XUbhemQ6A9sVEKhzGALtfY1vL9WDugD/TawG2S2uwEfarx8UKBMn
B1zsoK/ILktgSn4FPPyNa6wsNZ5FPAo6Eux0I3jeChZLYatMsVhSUI1RRg69Bry+zJslZCHz9gnC
s6cZWhsTTKA12tnmc9c9MeP5XcsX+JS7ckkBrwXLg12ybksbZn7mVgLzA/hQu/GcmTFZ7u9k0tE9
vv29gk1VBiwgCb62mUjZhLkaEm9UAL1h0kijU+IAwN9sugiP34xHbOvFYm6hzuS+rLkWl3wiXfLV
sSNkDfuTqLwqqbSXJKx2bRGTJgdt1HBe5RkoJfCidIDILm8kLQLpD3OkRN7T8iPcCahXwL3liHJB
+X5XXeeBRfNtbXAQcxlReLUgRxoIdHHVE3NkOQ9S5sycxI5PrFTJjGJDSN5qVJxAQX+JMz5QMrKg
G3JaUlXd6NNcNbTJX/MiPtI4iJis8MarUKUtlXRJfcZCEJ4thY34UiLoLPj6I1Tqod4dfmEoVxnr
HpyoLp3epsGezpZIUxVrcgv6DdWdtBzVb1d9z6QxiHjWf2xMeRaMv9l0KMDWkptMJrzSOPcFikve
dD1o1jdHobvASr6ISKnYadEYI71N98Rl6QVSWXCzQMKWq51Pdawk6UhP64JR9Yzrv21C1EFjo8U4
D8uhTpdDudHydTHGnGqNMLeqGrY53zSdJtEcuu+3are5zVe2I5yrQMGra28oBHoimPZxaqnX7SbR
iyfBugY8JiFmmq7Qiaw/zuF7RlPyr8kVr1GJNByhtYJFADrfHf5kD0RwnSxAs2prfdtzmgN6W9PD
/LNlo7lHfAR9BnFYu7XPR4IF/1BXe4LVkAbM2kpbE58zpvzcK1RVdoqoG+NQQVqRHPcv5YBiRnWP
lnXHklP0ICO9zYpNgQ3tyVrb6uNzAsSVdX5O5XgoJ/bY4VGCA8Rx3LlSoiLoZiwpVgAulefzpzlc
Yv3FgDEIpe7ruwsV1CBuR+Jj/ZHrb4DLhIVSBQZmz98Mi5Y7m0hFSjdimUG2zES3KTNTLta+bAxN
x0h03DklTwt99rAcvrlncSM6VuNjY1mwidpZGL7ok6b9bNQP8Ax4jjD/+Bj86Sc9+pvV/3B7MjR8
WvEkYMz+jNZkERF73cclq+OlsaLCLw/5k5Io1ghXj6srGkbWyXJfenOt7utQfllNkbZpycRLDeEF
sxyb+u/LkDmhdMWvbAn4f3OPZpeVegRSZYf7Ajyn+k9VlhpTTxAl+rDagLA4mpH03BoDIpPNvSTW
E562S9mjhiLWv+5lJsH1WHmv8eogPMfvKd0OLTuUkGNOJB1l62030/8dQq1taqaWSekmiPfWfBzM
kPQJliWw8zYkCHxjW8W9DDRFujDiQYCIyzXoHRiTid8dmFkhrBqPUM1wRqTWPcPCYRBXhwXya6FE
G5c8e1n2INPuBioM0NhuifMhb/bRye5bDCetGXIts5LwinhkzVYb8w6rRsrb6LeiSyPqoxmwnhVh
+OY5D7dtPIonV4Q3Ec84vut1O8Lt2ayihkzsrNTfqa61fpEDcz9WZ3BCI9Jv6Cwp7S/U040eLBqd
7FC17rOhZTtlQyjESbu+f1HdDFXoTJu8qh3V18lnFWBb/YqsLwNw7e9b8X8TRwk13BFiizvpGOtD
E+TjmFBW4NaL7SACdD7Z4bz8Nb+IKBTZt6EkpKy5hk9to6+Qlze2tfebp33EflW0PGwgnc9kbJBj
dA6+EyhFfK9OSC4IdmsY03pVn0BRWi8tLBm/JrYwHGIOll7vNh0Jo7xRkbC+eKqI5ephPz9sUx97
UrEztmyR1hS6mYN1Mf+125gzwb9lo9CYXDmpCZ1w4B9yIUQm6LVLPC1oJHtytj4za+YJHCORHAXU
EsQKGdmuw3LQR55OM8OgyzaC4qCzGaIQcZrH6wAqJF7Ao9yKLtOnNwK80ElT2A60AeFANOWuo11z
Azm0igLLb6UEKSb39gVRPmf+GYX/D/TP3o2xxlGcAEzhuVe5239hdD9BR65Ioa8KGJ6fWO7K1jx4
6mLbirwu7/j5S03M0fTU9lmajktto9D0MIqSg0zvXw37BYjbWO+DVL1fSQOCV0FMEFYhYZYGR1gS
oa+DLa4uhQJPXcv9rbPawn59/5Yl11QCopKDXMuumN2/u4i6q+3QIx6RPllSLzrrxRdWo9wA0o6E
VEIsSs7zQYWZZ7m3JvoyDfYnkspJ8tHrexTguAoloyaq8UkBEhjM40rB+JXh9i+q3zduGGL5091b
RLwWDJD0N+OtaSiB0y/iQ+W4ysq/RSIpP2yOneW0SQc8jl0dvPsD7SHHQYAWueab4150mgd0dVLl
BMkTwVQAgse4DBoOUJ4sf1dtZx/oK/mFH0XF966EOhBWkBBDkAXeDyv25IvD8EJwK50rh9rnLvWU
2AJNBuqBZSzFNjwWXpXGBl/m0m32pqVGR43N0phOVSzQoRqXfULUcCb+CapLhSC/VvuYJGopEqxW
8FEOHvtRNbylSCSNZnXgpI3Rjcx080s5pNH2wr5U+k77oZMoxCXL2qyJoQdngN5tmSGa67cmRGQA
HmUOv3yE7wUN1YEGOFHqQxYGIqXSo0K34Lj5y7asHNbHZ+J7ZfON87qKEbvHV7AQcilAoVcDPAxW
OzNXhebwSKOBoMLJ/u425DnNoJzGXS1f8evristmwXW5HInvTYkIRJ7vvdzZtLOIp/Izy7iweVBT
7jZtS/tuc4mTUj0SC3SZAvOWJZTMRGi+/lnyWK1Wuq5/E9zPRkiuMb3rvu//ZyNyLpjYTATQNTig
wYa9glShHdFOEGX9nn7NwJl/dgSJVf/y3/ajJkxKJRlQqq94UnG9GW7gGc78vkF1yBz9m2YnkVTi
K7v14GwL2LIIdUzHkBdPqdcuIbtujnw83yN9ykd6k1ggwepAJmFzKMrc7VwEBOZ3d+FTya1bjIzE
9FaoC03oLOI8NQdcLrmUOK7pOxb+OQxdU6H/IQiFIeUglQsTx/RaLfKuH2WBK2nXrIFYzsBr5fXI
4GU4PXxGVtvlAGByIOisZoD3K8S/osd0rA1bcvEf+M1HEAtAoSiyMxxRQk010Gp2yaVCmzAJDQEK
y+LYVDbNhLEeZt4+I85zztAMusiu15SGMDCIVszRyw2v5fg9jWUU8w+sYheRRpdjemg+58lUIr7m
HWLy2lcm7jqxeBK0q1qJXxLpvFp2fBQQLoMhue3J/sqpWVujNIoJ1KecWFthS9H96+uFrVbNMftn
twfbulJo5rOkv2KQtEe38tMRhQ8y3Fov/O+z6i6HlFycGS/uXAvImXz0sU+kusFNfeXlG8VudTGM
sTcx4UNmR/X9So6z4zQHqmz8SPwaXECEP+Ag6THHibDqd91aojDkOrj39IP4ezWlOcr1WfUxCKnW
eczhbyyyVIkA9ZEvfziIG+wg1m3mSAtDxcjP8/9QK/5pYbR474glG83yE2HMTyURqO6Tjj96OAXB
PR4UoFz/Xt4O79yOukDbq/Rg2T2m07kEaVG6CYpwblvNOO4FQl5vPAfRL0u1JJVz/HlDZbTjdMwD
XUvS67IPD7BQPFkNOtPM/4MchVxp6IDV/qvCrzwioFG1uUdWL25vdajBsjVGeJkqmXCqakOCrqa0
CnPe+vra+tJjAzXu7gvz5JpHq+PrGQjpiCju+dpzn65aVF7LH+dgk6dbk48HY0uI1P9XzzV1uxFs
mAbRV8Uh3bBm6uLbmBTw5cjbxIF9cDG1VOOrq9x6Yi5dSzv9iDFBPNcntf1Qj4zBHBgtYHQbN/hO
yRuwIH6dTvay5vFysj6LFfjRLaPAtPgipzDgwdDde8O60SUCEQdi1A066yt5ZUPvRLNFQBgfn0Px
v+25l1V8k0Sh8ZgPQhO+LGjzG5Q94vxgIbKMIIEHMxv31N0raM1KizkVg5lFRRsBuRpCZaJvDqqk
0B95QhH4/ztDmhV5IhH02BCbZfD6Dd2vOwQZu+uM9SmvHUdjfGvhVEZBOChkLe3vHQNpErlNRmgY
HkfEROxBJH2TQakuE0ffUv9lBswkwQdIbU5ATeLtlLqrbQx4iLvaaLoo7pnNnjrbOETLTs0PWfod
RIR6G+LFI6u16BrjT/EKnBo0MET9RYnnTSFKVphiulATjQSEk3IXU0ibfg1mAq1sMa7W4K5AVe7h
Z+VSeVkwWX4SfeOZYXLYkKG4Hd8MqkVMUZ8QYTmrxEXK11O4FuDBz0noy8GBfdCCoyc5mbglyLru
P5uEC5JKu5lFeYpWNQqwTUPCj9jaMOnZfEqn+XHdxPp4lrL7Hs/C9b2HTMLw+n0hqizjLKI5N9HV
ghO0BALthqTpshdMbE5mpchdKqAQAiGaGi+q1IN5PfwEMDrpaQW+DbPTkb7+OUpp8OAS+WOrASRM
dWU8SYzJY3/odsNBA8lSmZA65Ps5Nqu5qmClKyVFDmxX8qjvBICVzh4iVXPEWXGS4qDG0813Rpyp
K693oNrkdB8C/vAwRU6QwHXaLT9ENWR8mkcaYwrpvPmSMICbef2qMeJJnEOVlDOgguPRPPhtItlM
hoMv6qxjDWyv/BHZxpLoDLTXLwDw7Tm6bg7TSWF6j0GmnASgmHmm3Mo/0cu4fFq5c1Vsu+gR9vaF
gSeYca+snofuLVLZWuiJo7KMML8On44oj0q1mU2JjygHl3smD7Vom4qwRRCkPhrlw63Z16LztiS7
msMHL1sfzr6WR1dXuhIouEoFBPsup8IPyDtodOXZK11+wA7Bvkl9cTrQPya7wivCwxC0bHY7spz3
aA2vbZh0J7c6ITroYbZRLREZuoPacACm67t86jEW/wVHzn4AVcgZhXgmww2zg3USibyk0sRDi0bI
ZgtHp4Bzp0/nKl0uMjXg4xtN/ev/gDHRR9fD8efAhyo0eOqsfkhuHJyh0fkZq9cquuWuYt57z+XL
s0g8GHylUQxw7DaoREoatJkOdXQE9kIU+JdcE30uaqYyG1BE8a4+brNH8ik9yTly4iIvPF4Jx02P
9OFvBNQUcasC3M6G86t/8vsec54oBs2Rkru+GlL6qhfSFNIELEVZjDLBgHgSFfa/TeiTEa+gTrCA
+xOD2U5ZQBosKIO61CyQSjLj5ND2vmlBhTaNINCtzCpxUMVpwH65WwOnk+bqzpskGvKIH2VL7noh
wZEEO+tnGwdKZgnKfSHaRol8vkST1+AWCW9xu+cSSFWucd573f2MqxEPTygeYPj3PQrBo6gSihRP
yVf+z5cjgJ0Sijs4xg9qwNWoWZEbfeeEN6oGIQMnmcAoBIWMKv0ql/kzhHxyEWPA3q5csXMrK7Tc
i4Sy83z5Xo4mU+t3RYvualY1CGtmQftmJO37JWM75ARezlDzphOB9o7mjcAgd5EcplJW6qbI3+Lh
vjDxmupbAVb0gnNHuea3RApkh3e8tA7WRJCCMaa/AkpXMvkIQ0d9146UxTVINQ33ofCef3xGxxiS
SENTtMtPBCI8PmYvFcV+AJ07m978Q9F1yU09PVL3e1qVdOLyRhHWZtsVG7ScLp3Bpa6wjdocUWK0
2JxKkNuK2xcHa3bWZls6T6QS7JVXo8pvK7eBida11wm5WHOT2lNnweTiOa+A3JxGrfcdh1jgvjE3
T961vTlEHiWQimPPSVK8HzzgWoLeKUZcxcHZtzBexhmIe79hXn0Hp9cOWf9HtYozML+CPUTU9twi
j7O0ugIfoHzzp36+PRUHFUvf6gj7uLu0GvnAJSPmjU1BHRxinjFkyBTCtm1FEHzV7H2yfDHGAqq9
yTaJQ2LSN8R6asfIux8sjD9bUKCKGpNGg1IJrmz8/LTFpUBFoF8k06rHwg/WHz/Pph3W/tEYz8L4
94me54bfNyRl4f4qADg8Qj8XWv3dSzO8nSeWfw6Bk9Q6QXxvJuZFSZAS+b4JX4M18vs816Lo3epB
7F0hUTm/AqX886Ts/lnFkJeAWhqiFK+XsTnKfJfHtWjpgwuYsJvIPjQbXQPJ1fdI8XMeDdI1XAq2
LE44WcOlHj9RuIBysT3gWHKg4itMRz4mmXQyarDfLYlB8Hx41ZAVzIUv0jjikanDk0A04eemM/fC
7T2tesvUnhC3eQSYDAfM/SFT34sXes7BmzWoRvKD4idmN7DA21t/15+h9Q4tmrg36b3E75tEl5tU
x7tt2BJNTzA/e5xx8qyoCHZYqlEwfEJnE3c6qs60K/34U1kqnm/hxqFs8eDqBEVqcTmKqlbI1H8u
GIIx6hnmDVeDvMAhFjIGy/YhaoDiWV9P1/MRrSTwAZQvH+N9mv+3rCVtVW3IhtCZAVy4OO6HqEbL
DkV+WqTzR9dfnGWzTSUVEjemqh4rz2we/b1cgKLm9xzD8exhf0EUHR53NDsr8hxtzsdeZv6A29v8
K+cLlHxWoisH0cCXXAWFZMcM6NsEaAQB1BqwBQEk8hjyUvIS/+48v1qs+sMj4SCwEEk2VpHfyo0G
bBB3uyXNfXYg3E9RAKA2WrwNyjELo7rOjDn14N53bqmYRnW+yOdCtbDMWT+BvfzrWlyBpzYG+UPz
IVNez+VqYB0QuHgdi8toA4Bp4lgVeIbaXUD7Wjt8v+T/zJ0MaxmsB0LOIPnMgF+KbRn4JLyAiUF7
y0mhzq1Buhr7FCzDPXVqiRE68hOqYyDygEloZi65+2y6xQvjXllP3HsoR8CujuGzzLQxmAB8nOf3
Fa/w84rVAOvLqoyVYAdOv84sSLPpP+AV3nTSsC/+Ny6vck648gKFF4rMzXyjfT7d5iR2WCTrkHPy
6pevtC6OysC81RllffPkhprcDnPR3Pp5EyDdTGYMgYzfzMcLUdBIxi6NT5yyjb5vNiqYELNG2kdS
Z6AZtNaW+YX8AAdiU1PjJwKjjpgcHnZbIkaaOydaa6OXGNzYQ+igmPNRRtuQBjSaSjpWkJ3hskP1
hYp19DoFHpR3R9i4cJZamXmp2ez6famWHd8we3nT6i3vlQF4DnYm2dGvwMejMUAcULItG2+474Yy
odRMo3vbDomLa4dByPTfE8Ye7oO/+DKymsi9YH6PrWl1d3Y2Zm88SI6Qzu+Gd0cC1c2dqFGi+ELa
XpuPdXjt9SDvq3EsSQO3/xG9IzYVQuEVVAeCcdrnnJB0XWCwHWvv/SFmroRJIeJon1qrVx/m4ocZ
gWBt+XOMEahRTNkjOpGtT09GuhpyzZA4qb7Bi+0RPL2FmJSwju2qF2JGJZD+YcKF/Gkfs0JWhN9q
PcO0uarGJNsqh+JQgjmqA1t5eA70Z40bYLIxoVY9FzA50PWKmD8809xvqG4dCJZcuHvdLW5Xv191
g1fUSAGFdzVyf40uVMnDBhBI8zTtIORFAimJ+hTVSkYHVHEWOId0MbkKiuq/fiBVO3/WL2h8nknr
yZppXz5QdC/Cnk0ufM7SPl2ESPuo2FXl3HSqE46ucLwq2dEP/5+SHH2TnYmUG7rKgBAE/Zze6R3g
M/Rmo3SA0XbOxtZ7AgHHmtxNw7r6PFinzAhojEW3lh8KvZtsZI/pd3q+gHUG3M1gvH4oITOJgCa8
atHkDUYZvZVCsURgW2Auu8I+auh8z6LhyHj2gLHmCQoKR1XiCsLwVrWw7RFvA/FybLYglDmvD20a
heWIQx0euTuYP4lHvRbe6vvxpbD2drmix9Fip4yCrHvT9ioBba80XlPZLqp89hXLssIxrzqEETh1
ZqnH9lmUcwxiE2lA7uaxZ/ZEQRPziMVzjDM3sX9hWWnTnBNTAkYcaObZ+X03YCLt2M3dygGDybI3
gmOKd69yAWL89ipdfNJMZbuUiwQMDrsqyHPfPH8S2QVM0ciMVeGZUaT5Y1Qh/ay5gircgCi+ECaI
YQH8hl6LJ4BfY8vfVXINDregU0I088WtGAva3/MnqM6JamwpX2UrHseSd5CEUhhLrfjl/+GUcF+V
ZxBGEKk0Ehtkol+d6zbefjumWuf03P3uvTV9fxd6J1eG88YIRYcCDPchCGw77u+TCXxelAi5OzTw
KweMrlpVUVV0BxQGNEyy7aRmGpSNpW9nsOYrY4QP8OboNdO3jv1roZikRXOaCfbkQHw93otqG8RC
oZ/Lbxeb1nXkTY5s0XpAqNMGYlcOVJBEfcs/13oqb5j3RTn87SQZqQaqeHIw9D7VffDKYtG+Qjma
zCXFHBnLA96h9c7GcYMvVyagXjhWwf5FfayfYUcIVYsuV5OnSbbSO2iZ1zzLqvUBw4Buoai47NSL
uA+9tD0q9BrGUqGTEu2rVFuxYbS3GD5hZyUgqQvsXVCtqE9ad+Z0rv7FWfkgWXk7VawtThw17QRd
OyM6Uo2kIPQpDVB8/T7gLrdPsq9xsud6QL0KeTw3zGEGYvfoOhmggkB9/JFYiKBbw3YjZlnlg8ax
uQ+LEmulp3kVOyqEUQCCClNymUPhj8gket6ht+jczgdF7gYxnvEIQ1+V0+5oePbc4ER0f/MeyIiN
osb3Z6bogoFb6ETPSsv7A/RNcMt8jDsufQv1w69KIw2wCuF47Gxc7vV2s16dE54j4dmqQCU87LL0
ArPWBBPd7SXvOCP5B5zPvkERh8vLlz+X3C6HI083H+YZ0mgSdDQYXkJ9/nA8gmaf9Pih5wVRFXzZ
TEQlF6dKocVpUO1dxecgMO+b7fkjBY9XuXKTElQdw9jgG5zuBLy4xy8IyvBcaN1xMufRaJiaM+KF
BEdyExVGVoQuAvNSg6vYEeVai7J24j6Pjve4rAVQNN1IttWGCErIvcTHSeV7ifiGWVMSqtXKUKRN
XLfvvGeJTs8efFVxO9lGUkDcPwxrb9Dbh+Vvr66TmTHLbWrPHqcsZiNQho6ju+AUjjwVdRZCMzYH
t2Wv3h21luNEngrhatQzKEYs2VYrfOK/G7C8bXIKhNOxAmrLLQQR4AbUntXQOYPk2BZLCnhGCJxy
1RgmAxQUcZPiNrc9eoyRBibulRGrkKr7tFBEZEmm99apUyPt7wIuB8UKAZFE4gmU9DOmerTcnV/M
HlLsEdtScM69fxvFt+bQg6/QZlARxNF0cePWz/066YtDDmcVu36O4WWEFEuAbXlYSGjNU3EwzW4O
zjGFbX+T3XFobTR4LzNvMhHPaZW9032LdwPeWdUyjg1iEP9e6b5BQXF8+QdGRo7W7xQAVkljPpj2
ktvFztmUny0PJjwOVdsivtJ16c/zULP9rdqtdu91StxlE5L3rWn82MHS94wGok5t2Cy8FyovikJK
sSjqyqZhL7xuJ0CrukF/tDhbMVX3Y7JihCuZkApHsuMox5yKgnfa69cUMfCdH7AIqtQq3YPM8TwG
UFLZwJooqn+IbrM91X7wgux8uTw8ghumecolpcpOhslSJdpQjW7dNhn5cI1HZ8IsXtssCdkl7d+5
sfnHC3NasHceUoj1cGi2zojadBPNsQsDZl3SBaU4kYHWmQcNQ7kPktwt3MyzRtvv5XS775eixit1
5tBcOydqbFpxo5JNpa5GG53duvVBSWJgdaPwEssCFGYvC9yngxn2w0B4xXJ5cF/NiCsC2KwyXoYK
9Af3VMYKSKS+rrabu6If10br7nUDpPDhRNBhWZiLZt42UoClUvXfdW6nq5Yc0GtIJ7dR8py+c8k7
XPTddYNLdG+99/LDJc+qhtviIpqr0yFbHKx+ZBKxzdlt0XyBCBRTCvXhFVBb0rZnbZ65yR+n1ApK
f7ESPES5wWRphgGDQeC6iOUvhrYzVjEjtHnuF53D8u3WLwJL50ggFwuoCLOBvIgvfvYeaM88If90
CEtPOaTXUTmHTpUuc7ErwFXiwf/uBAHeus/zedvGMCgVrTa6ju3ppnpG03TGBjOcfXnLwzexiDZe
3cfYT+qyzYJF2YPyDEIikekkce+u/eu4v2STjQdLOpcTeWSM4vLXsZxwYvCHj4QayJgL4X0qBxQt
lrH2fQS0dKMLaNIqoEvk2uINHTWEojT+Dxf1OSDEzMoJIWt/e17gfOTB+sFJuIvYYu2aGFYj2H3Q
hO4JNUEIeaJyS5L5Fp1WClvKSeMzsMfV6brM3YMuY5Ay+TTflnyLyssCS6kruFnDfbYjNVf4zm5V
5nKa0qiYyrQ6ETmiLQzTm2vyskjvrG5zYBJIVCSC3Spp55AhpQPQAcNrCczalt3NOoJuF10avBm0
IhZ3ZYcHCn4bmocmKeDYtQgMjNqs+TwvK2nTd/Exr4cFyE9u43Fe6hH3kX5Ik69Rbi3VXtDYNrXY
ya5v09qf2N9wDodfj+hprkf8f3xIimvBCO+2KOjAi7usouYUVhvTDYhHvVRmUPpBJVjFExztdvqz
vvd0IR0nS80bK36CCeAAS5Axvd33vPv5Rf9pHzMV+fIDK2irILq6bEYnh1E0quAHtgf4QebqlR9A
w7aIWmGuxVZApbOWWejXpr35uGP6tUSwasFl6i1ZjlCi5XaFpFiKFQqak7draP+XhPL8rkThvXiP
Jx+61OFS+ojnVnPIRh9WDoxAezhGfcKb9+8cw2uE2as7Qq+O1Eaa/MP+Q6G+TWBwfRnC02NGA7tt
zW8rKEJ9L+jY+XjUv4hfzlP1mZdS1pcwZh59AbtNWHOU1LpXreSLU/wVYQiaYaabKFGpagfg39uc
UkqmNwWTuPWPUpArBorGuHBZQp+/QfD9cQKLFIgcu9E6FCQORVProK93gPJL/rseTbwT/qmTXZCZ
UHf9CEk/EyL6L7owsUPS4y3vUBQxgu0/P3vnsdljLc1IOnSq9j6mxMkLlX2XxcvmbTAxE2udC7Np
Ugmm1tBSqXrUaCRms+Zdww1gwvuWsoYzU3y7Z3T2Sh1GzXJPstQs8NC+dhL9GxZI3MxfvbBJcJRS
JNm16AtamjjsuGPDAkwjaQYT1sCueFtgQ7vBqI2VIpGjDCHYCo3BqUTNLGGK89p90lEZlthsBU42
cGWimaEqOPk0Va3krUeA7kXhl3yVrhJyWknJm8gO5DO+1/XVEkYVkLekEQFvpev7rFYehBvorB3r
Sirtm9FYzkmin92liSf8Dh888ZkYUoYZHLSwX6Xd4wcEhfBP163GeTe+skbqJtJ0DsDIciVRuZjB
hi+USMTralZs513FXbFtUveP5kc3Tq/EWkk06DeEORQhRPSLzvsnqBzdzYEbkTfERgt6C+Tc1BxV
/px9S6zXWwYp4TpkwyrFA3Ehnf8wRzZ+5/myXM7yhrgdeWpasCTpRePfKvqnwTaBNYQuM0jpMk5D
xPYbTvm7jSFFr5wKIiokvroyD/JFELZdZqxs10KOQQY+sDrV4gcOghxWRKyYspr6mXJXbkMkPzAt
HkoAt5/Q/fsidUQdaOmRW2qgKwOM48FGssnhOKeo/IMjwolq0KYbR/UOTiFN3osia1Mc+NIisZu9
dzXG1Ao4JPgOr/Pe7SbrSbrYGCtl0KCj+D7EmM4F1QhKmGry9A+sHWnCaNgyqVAqURafl4SX2Uy8
XKot4VjwsyUjs1rHCxrVPStQwkfYTuDILYXy+qHOWWpendlh7ORSamQP6r6hSe2CgePFs+GhAd6Y
5uPPjCQILjcDSs9d6rxQxlcRV2Lu2+4fHrMNmK/+NIqCwjMiG7rlwi8iTLFASaem7Oy7NQi/LUp/
zV4EFkPbTYDVnvtdgGfW1b87QzUcjD1h2WKmsgP/5pGo2Hbu4QC7v3FZalk1GXq9z7IyWH2shULl
XXSK7cFcYrudHVmMlEQelnE8bYk27eozJ+MhDR10VrjIf/9G8gNiXVlnoOKcV9Mv2n3WGYambOnx
8vE9dk2g0JN0QRqGM9zoMW0P8uF9yOerslpz4ChtIdZtTMSDyOnG6Ay+UnPZScuZNSiaz/6SKUcq
OyUjKgOIBR/B692fhvC5kTYHbrYMBmbP8S0i2gnt1w7k1UumLlpZxNIQGozuonWguCi+NprXPtHH
6oBmFM9X2WSRPSdiubpUsDAgP0mT8Vj7NxIVo2Hy3j1bZavqaPBPOyrz5L9vCNIhP3G9gHJFcLrX
PLxEeNKq9Esk8qoFVCuWu60sRUG5Xp6sLvfDAN4AXXge2N6sZQWBeG+QAQWWBCm+eUrYCSU8NlVT
PjczBVsBP0zLTZguHD6Ee7P8npP8vYYfsz1k5Qre6a2ebAl2J5+ZdJngWe2iSho8JrK2+GcGHXzH
9i9sct+EA5mcEJx0/FEyf9WzjXfSnn4+N8xMlPfWaLROsVMsP4bKbAXlXev1w+9On/MowX3gceuV
ulTHz2mLgtuVEGc4UyqGqykeMn5Wzo2Z8N08LGr2dsMakitEMemaAEgveCcYMatBEBATavZqksc0
1LqEEHV8f69B7JnYN9vMRLtNbYL2p2f3W73L5UH3HaZPter9pKy6zrk39/0r5/a96VsHmJHXDYXZ
wBK+CcI8EOxk+kaBQsq8L/ggejfVM/k2HTr6hN/mX9yI4ec/EOjZ11FaG3gZy/12B5AcBve0R7vx
C+lqS+jqhON4YyIEWCi+W/TbVZLQd7+xXXZpwNlXwgYdLMYgh7DKTcmO5H65MIo6cD9xH3t5xSBR
LOAKmDveyn+fbilzldsi9hZRxfQJs19zMa/2stn/BWBiX9DwVSCAdMcq9s1A/t4SFgQJ9/RroApu
7u3bdM7Lfhmysg9wOdluucGGOtQHhNsoXNy9D3i2p9pFKrUmRVVSPffBrktRQ5qz1wfKVqyweiSf
XRzrdKlyB7LM8RiPwO9DXlMLzhGA4+274eJxKEPppBfIpgDjEGP1ytdy68tiQEhI3wh33kMMFZXU
7c5+ZqwNcdO5BtBoYua/mxvLncEv7Zux8HUh68xxvtnjEnPcWwXLto0Wpf7ZPgxTRxIGwuA8hRHf
l/KE8SvCqlqLwENA2/l33D8aHbrvQ0BmeNQXvgeyE99k/Xym1+tmSWhwx7q2eJaWkxBoiDJR+CAY
5oIYon65vT7dlN+sSA2OoO59n4v2yrW9UAltU569ZnBqbTlAQ35WMRTZHr0fe7SpgU1T7aKs3p04
BukmDCvKNsBXi7Ad5LRp9PIoTnPA09zbLikbgHOkp5NPItAv3oTbY5Q5Lt4zh+StrNS8Xw2RxLMu
wb/aJ6KBMgKZdiRz0Vc8GuN16yj8nPkIPLeRRFlrD6gWQTC7OSjOlcEYFTtc1Q6uEBbYgWRqK8hN
dlf1ma5vz7zaSabAWOeC1WCqDsNC6/ATxm6G2ruwLXFRpwQeX6jX1V5mhxXa8Djzr4pzlqzvxJ8O
AMcgprPCREHCJd9SC3EwP5p9dfGIAkeC6sOiESo01967bGF+6z5ev5VRKLdoIg6oPbqx5YDaoMZV
j7qTeyMpScExMGpiB4X6igCFkdImAnuuSRFBdAw96D09MTfmW7tBO8EJvZzVd8SjXjTZU+egbDh2
y+ekTrbdzcVg3hob8fJytIunJYZLc61UTxzqN1zhVyXRDXN1js9UKzNOzyIlyxajgSPLGoGztz1p
O6ClXAp4XBiZKAZJ/q7wzevsCmLPgWo96YhXisPOZbZZPIDMrKM1br8B7C7GJQ3LtMPR9cuTskxf
w7gxO70vl5swMEGhCgM/5e82GCDroQ8ikHU92H7/HFVLBP5y32ygtvCJmreGf8+BK+c6OVXVssM7
b8MK8JMY0jZdketNWo+YPK2GV/EB99oY7GS5kpue0I47TuitDMPKpjwGYluMASXWs+Vp8OraVbYY
QmMB8qtSk7w9+WYYIBSLQcIhRrepNfiriJYS1RU8TOgZocyrMQQZvXp49fkmqLTCOXS9TQm+VV1M
LplltoURe7IEk26VkWIl2QI9zTcIoYZ0wenb/tG8UriaNoBHsTEI02HfMUfNisbPqpzCQD02VoU+
kSyln92Nemu5KQ8L9zKG6Gwu4C/91En0JLGpWpuPWWFMvOSX2wTvIw9oH2QX3Ciz6ThzJCQKNsXZ
qMM8wgyyXPH2uTCJUTSBTR5Mp9wlMn5om47jHa/fG51ZUM8wceSIzBYUe5rXp90M6uZdacjnnS7D
mh6EeCOO1jNiN28sK8VI0w7pElM3xKr55WbyC7Rshdy9+IYHvGSZJkr0d9MIAiHoe2P1oJeSHa6l
wwn/IdOJSYBSRXkFR3fjQRqmkNSb00n3/HTye1mf+TTP6JDjt7hiUIocsQMcnHbZmXdQpFITcO19
SPJk2qC/DHS5eRUppWpswhx4d5wcH+rbnqhjmv2RuTfJtwRBw0IKlQFXnC2DvZCFbJNWhJIP+qgN
yXzl68yWe8DxghiYjfVc0FDQpI7RqbipYwuI/VuDgFJKFe+R/Oc9lnQCTGl6s2i8mSP7/Cs6unnB
1oUVg7EId6N/oeRBE/QXzIDvWv8XyE+M4LRkHVjAuEj0giGXbdMCFJU5Tp/M1aHh8r/uWnFhROKl
1jAJ4BQ51DlMCchqA8kFbDsZDZjeaeBdfRe2gZENQWU2Ks9xHa6RDRV+X3l6et48T6zuJ88tzZKa
biav/VKvHbjl9VR9dM+ak84ecVpr+BNnMICxfTcIQhnnmkYaupJH34zvCh0qDArFmA+53Ssjm0x6
Q6+1ZvmSM48rYJwaZAX5YnstgwMB7GIcBm9qAXzhvVP42+ADvA8tD/LCzZ1LZzCnhJPE1FyxtCIk
t+SmG7xBTVKuytipgQNWTNgIISjxyEFZV0mVdirxX8wzAOswxVQ94U5pbxoeSyJaaXoxLGerwFfN
8rD4Kze3VeP+SDgEJWedwKzMmngg4CDAUrprEymwbpsXh1puwhmnf4YF1uJ/AjZ/ZeYjbcA5dmrp
XkSUFvcghfaxbuvxBiSCQlRBp64T+caXjncje/VEQOx5qswFU2OZkfW1gLoevkb5pI06Nz9r7915
SiTdm2oVcdQ0MTocBAT7X+WGxTbVCCFBNDhdx38Pm5bM+a1gNpQgZMfh7Z/k/vx3nBZqS/UaLbfy
vDhD3q561tQJivk4ms/eO0GvWy5jkg/DwvdbjM08lESY8DOka7l/MjYqBRNsUFCiqIscYpI91QBR
ZwLCeSJYmS2RUFb9s02KRkxbmNQmj53Hid0KkxuW/rkJ0TKNe0f+vfbwtZl0UUD/vfoVsXVXXdUR
ozf/nbz4O7VBmagylPuCiQPIiCgaSOsEyvytL23rbqV/lj1O6wPG0dyqhEZ+MWklq3zSgzAyfo82
ZNn3YR2yQhyUpR6zm+DnncK7iHdAnVGNNm1X0kYjNLsXAMXZG47NrxSQL7cYczJnuc4aYszqyBhr
cOLsbFwZ6ZUsiJEJnB6xqaSw35Al8TZBXHPho/8W6rAGRRw6V+LV4vIicl/qQHdGiMkGnc0hQ2ia
pLxUnhtHEcV4KxhVAPu7epwYHx7yR2F6y7K2GpHHcogNE3t9kaZ/p15rBvXv00DpGpASuIvRFC24
/z7yq4PiBjT3JlNgI0eSZ9kwVj8fd59RG7oMah8fkz5S07VwpfVzQRNRPbxF/ttx7rUt71OdnX2/
jk9hlqfXFveQSTu9RrMwUTYsGp1VC5PiO1d6CyeOZfnYRMxuo9/Gq4dDcFsJfTkjDdPlcegzIEXZ
emZiCj+/geD5GmCLXz+Qzpsa56JE6KJ3ZGgwLM+wkMLqHE6VhoY0/dq2HPoEZCe2fb4yRbYxM9k8
wpQauYo1NGFkHzx9w7e1bPeuoVPTuuf4sgFFzRkeK0GC5qYaQpbNmKz/Gnep11T9kn/cDzTUiDPo
CXrjct6wYE6RGGjkyYN7jdL0E55Sl1qVRkWbgRcMDrHZpv59zSGirQmsFbwpQdnxXdKHboNquVGI
Sh13ztLAGNhdIGuFKrIXcZKZ9JQ6zf77gRothThlYtO9NinTLiGphaIYYW6KWvnpmsS1iQaErG17
uR402H5x4s4X5JDspiT2YlYx2Twchc8EAa7DrvhTSlI33tgcJ7O+c3k2hkIfjoF7wU2NKDWSZXC/
AENpuDqSD6+QLujLpRbyQxInTmb3x+53XR8XZDqch0lA4Y4mMJjtwklo5xFppyhcTCCXtjo0soqE
Ll8UJMxAFu5gQgCFk1McuLmNM4qwacXefTsA8QQp9blY4zDClXwkfqrFS/IVAoiQyuo8fus5vdx3
x8cDvsDUlT2fKJyq2UecUUNneImva8zifhRSJeubldFSX31mKCSYoGCXY460+UzKBz+/wBBb4h3o
WjxuOB+BvQTf+sqz2TYIjrxS+fTvGZ/h83oyOVJaT/0mZqQ8WAE4unIHV82TineLx+s5RGFRjlTB
AzfgRmLYjLUven7nR5zZn5AWRMhYTGkDvg0RSwXv1K5qYjUKWRLw2zWk/9Rt5WK79LhKeWhXRJe3
1k30vyTkQty6MOPNx5VHYKrZk5PoTFeFKw5gU85Yq9MKbjOavQNUmD/O1zeXpodVELtQWG6rR9pY
LbMxyGYoIwQckxFKIKha/bKoDHW/vbbQlVt2/Byx/b0xbWYT1N+s8pifHpO719ZE+HxWAGf7NDfs
doIGVZjDlFwhaWaO8gbFpoO0euluZCBmIgNV4NSk9KJ0PrOOodt3NKpmgmVny0b8oBflisT1Fdlr
Vb96Z+TBLxOG/gMvDzKLyoUaQOvpcuouu/vjHnQEFoyERMdqsdWInHrQKu69I7Vdl/uDpvET+NLx
eRtZvetpnRkr/eTZKInGpdRw+ByIMX/epkVZ3prdAoQoy0sV/DycX171P7nGEKW1wLKs0SYILzXg
ayjhDL136Wqp8o9G4G597rRkoWeIwpBy7RSqe5rti4SnCprWIOFS2M0TDBv/DA6uxkpx87MIGDh8
UzddLN/X5j/DGSEabvBkdDVeKClECupd5WvQGXT86Kzm5JhTulEjzJxjLho9riSJfdK15mEcGNd6
f1K5U9PitNJWIUjc6QcTTJ2XMx2dyeyWWWeJuY6IbeP09mAMXgFl15vAsmbQLLarRLOcA5IgQIpL
IdnAPe5oz6xxb9L4ni5ZBygMkixpAuXdUi69Z8Y9PstflDOsuftPyITrtMmIM8wUzKOCN72OYNRa
+O+/R3Gyp62hnaekRdYAcouj0CTBN5Wd2DPKLMjz1XYzCSyQGUhYe7PMcw9SnSTkqGWZuGGBeyuf
acdixHb2VWFERDKiakQ8dIYh7d1Z+4rHPzLWU9oGSWG95ItJWUiFVy9xh3ZiGR1VVIZ2nzOQIl8y
5ptSlmu8igu8g5K/25WmifPoGsXH/ajSTLFevDVgAGQgZEETMVFwfM7X+Z+8gxt17AO5TyyRSBc2
AGIt1NFO5NANeP35O43oFGuL79rlLvC0uA4K27GOLwrMXVWDgXzJz2O8v/ymWRbvenN8FxNEEhtP
peXaO3CpVJUA9ZqHsQh2joUfxqKVTMJGgmQJ5GXJdGkxoIn7IYQH66zW61E9tvfyqtEFTHqrIw5p
AgjzbBaTERfXIYBx3MBEeRE3keFWfcwCACZr3zEFNlHG9MDhN82F2md/lOAp3qxHyaiUcBHIJaWF
j4PAdQ+gw4luevgpTClCsMjngQ2TLlSsF6ty/hKh9A1Hp7nTyJelNeUFUzHbulroX2w/zDLtsU82
qcmffz0MfrauZOUwHJ8F8B9hPg74v/3KcCM6kjMM9AoAez56vatcHmPnZxxJsStv51959o7TLjhs
FGqfT+kOSJC9sasJR7d8a4DC7qacp4bie42o57/HcNaa8Ed7nc0RejRuo5N7ILIr5WipPnpMEnZc
g2Pl9ByMYFq+prWtClpjJYTc/lljtMyEvcynCjjE3GDoZJEo2u0MhOonu5V52NxrwbzCeoXFFfxb
QnPbe3OlK0oW19srtu5cCnYDXc+N+Ihledke/kgvEZJGL2oNn/B5uO1LxXcWKbWsCCUWd/xKneGp
S2BGmfXGbggYLV/GLYpKk8eLyxNrCGR7ONhIamv5ITJfGTxss7sv05nKudDKz2IrCIu1q/e5uewn
4SvGIuQm44g5QRIlVdevJCzYYWy+TJFjOhRdrPsVcqBpJlrzBlc1qRm/ObF4XUI9mpVU6jDu5czk
9FC1J0FMLsCk7btWCJ4Ra2dL6jme1sDqhXbI4XlNI79+0Qw1pOGkTJeINjZDoim7vNhuWHtxnkyP
9QxwhTII0Dct/+lg8QPgQ2W7uc/Q8zTFGfk5RLGKyDsOkYMusKsnJnm2ihqs9KWOsFJIjGIKM6XD
jv6SlLmYQsu9JCaDLkYN6/0timdrwSejyhQObOGVLSq5OXHeXcWvDdJ1pe6Gbdo2OpZZkjVOJ+F2
9CYne8pwOQEHQC8JNCv6QJG42BsNRikL6gs+zk8gmNfUKT2vnoOmlfpSVpGLzKNSkAz+ZL6e1H8Z
dJaT22vAvUIXTpo3Ph7dw0UpX5M/SwZNF913vrDpOOn6MNJBimbXUenTD3wjTjXNymKpQTAu7ool
xSnt7SdsgEvjQz9QJvflOwuhW8QR+bL4zA7DOKKqXwvfWDivOBrGygFua3247p4i62a6xQydfQoO
HIHi+YdqNqjiFs6Ucu+pMen9hVuJelJNcRU64hdpNpHueCRH6Bqi/LZwMkAmJpOZq0cGwdFfu5J7
zIpSWeXKXZJPazL815KsRLM6ptBHNJgKtYCnEEYa3wuBAHF7xYyygESpTWCBdH+74Fzn/gtCnov5
35gj8vhB7mbGtr3O9xtGYJY8C6NyEt8LDy8lIBUr4SNl6Nz5vu7BYqfAOmh5mzoKfk7MmQ6H2+hu
QiqqH7jkHduTEYziFJ3S+fJANiGmCzqkNJUnYTR7W4o6tDx8a5xr9ZL7D4FdNt0Vu+Tfi3qxkX7m
qCoQtWd4WPdX80MRuFyeIUoFCCxcEgWgPX1O3pUCs75FseiNEtNSUux6F7XbZD9urKR3Rbc4hqiB
Z8K3JjPTQhSUs9/rCWg1wPKMiRRji8YzmQjlG25jxeXMojewOd++r6k0jk+kfpFDjftV3J3pBGHL
1SGn8sWRqJ5cl6Q4fGrLUbiRj2HlTOlRx6PZHzitvMaU2vg5TiQgO/qpT9KtwSCDv41EK4CNSNDV
p0NqkSTflD/Z0O5N6HjRxIyCo9X2lJwnH6zzZg86OAaFyg+OTgLF1Ftudu46rByBE+fe8oSrfPP4
ohfSy+Jxtl2l9vvG71oQqFH8w6dd5WlS6f2Sk2TJL/6JS3mepefyJUpvH1heldVVZzYQ/fzF4JIe
b4q2smOGejJcd8XaA6TW7J9YyKyxUPYkRh/yK+hd6qC1Ot2UzRRGYuQshMqMZmoNyXDSXDl36lsQ
W0Z+k8VB44b0571fcqcWESGH/t+A9iD2RcNHD7BddANAd6NtZJodi6H1kC8eq9UxAGJy/bGpWONG
cunTYoNOO912DBuYU5gTu5l3pQmxh9Q4xJar/GSlRpAmANbk+H28qTquWdsmwC8KWieso/1kLpLx
e5AS3L1LiCq623d7lD/nyiadat/5WW1DlSl7EKxhA2KPWpOMOEMiLXpQo9Bk9WinVe3Sr+avlm3f
x+27BXhej5tbz6pZNytTP7BRybO/zCkXjeeFV5BIaxAsOrDoNQRidaX4cDcNpX8ocRPBtk85tK+w
mpT7kf4xXM30svsrtAT6k5uZebDvCB2I4F8xaa5/XTiy3CIxkUcbKxfkXvKxPATpWpNzKqp0UCnj
NhQDxx4178lsAq/E4N9kWbRT28ydXSrqdJJDiQuCe2+AaY8g4vY7F175TXRUfD41Yz4oNed6xTTs
7XqiChLVSL4qrRPQ3N/F1wChPYfeDNb7atvngS/PVhNaNggHYqe2GoNi1iyPIsgxvxMRvtw6Qq4J
eoIWtonsaS7Q3HKTyW9pz1Ctoje8GjEJJzzNqE6ADXV0Uh4ae1Ls5dVD+aKwp6K+i9F1higzM6LB
fMTpbx2tKb/+7y5GcOlfuPcQFx8qhFSdhTDpqladhExMAg6UoBj6ni/mio8R9x1+/BzmOsCbRgTi
ZWnuHB5CqP1OwRYpW/WmGfKRn/x4sT1rMJRRWpHNrZNoFPUH59B4VhnJIsw3G8fkmfun+BKPlcgi
YeCEGkjg1FSSPG2+Fd1bQJM+Yzh3yIEVZLdJ0CKHj5jrn3mNJsTffr5WfxcfMeKURrTPdf7l1jZ2
GxmTlhlRSXDknOT1Bqyzw7hBAC2+839fcrNvVjDq8AdKfIReBYWpL9yuhQ8ekgnreH1Hz2qSaVbI
KutTQO11vdxIasHq4Uw0b6gztncCoCorlyqSTQiBhVlRaAUWy3ZoC/JyM0UzbxnxfuKxqm9KeLWs
mdd9pwOPyCD+k55Zh0umVMYY0LItUJ/OBBOsKb4x3x8bK4VYwf4Z8Ks10Ju08yc3ubJP3NQHIKqN
zweOBDMYtnGVxQ30dtR856KkCAho56XSxTz3Hkl+OLSdgcr2/L8GzetUaBPlQ40Hlu9OhxXp+38u
ezNoVg+0bI7/dB/sE7HXHqjutHaI4oqk51rtVR1oOPqiYxM2R+85E4NHPl+K1gad67O1WenNq0iR
xLu2vLLKrNMFDOF8XetJnXHyYtgYOx2Oj8Md1/Aw9VEFU5CnyIAIjXToQgiNQgLJ+gykAZhiDfpN
Th2G6Pg+3mZw3rskIId8BgfiK/DU2i9FBGCZmW+L4z52GXZOfteuBUcUjKIGkPC5l4zQMJjbYjNv
AYEPWpp0aKVRgK7/LOTRgn7f0/GIFmiZW/2xUvGGvOEyebhoUfP/J4kUZRIZKikJqVFSUqe3q/Tt
P478jLg3C4N/rIIWH9YQWYxgl1XHZe0H7qEcm46eMeIJixe+jQFLNWrCsgc4n+oxgYzmR3JgTOFo
CQiVd0pQS6ACE7mOzp7hHhVt0cP72GKg8M8/WRtpDlKrpd77TcH7uNd5yfzI8T6GuFDq/jTHCDQB
u7M89tfrYdyXfyVbKgYdX7vv/SHDo+HN2i4I2rkDm5lSpPneqKLfNDRccyfy4XysiqlRFgRHNi9k
vlT90OnDEjCyS7LlDsb8FxWKFzMyhvE8OUAbjxzDuOJ4nTfkUlfxGifXzIRiK9VrFgXlHJZHwlFs
lRiL7yKTxjXicYHkMXinBqnLTARbcbJ2w7+i+3+4PRmmcQJ5llPE48AD4nf3KEytgrVKK1z+ZiNA
oXx2ugD0n79t4998HdDf5G+CxRjWlblQR7I/DKV+2IEzNJu810EZ3FehPzsnQWJ5hAa3AN40sXzq
9yOgbuleAe9VvFNmAbJjcPrOfbPcGzZIsDDG/zNMsI8S73h5wxSHlW4b7XR0dI5DQ7Z/LwDEF2W8
oVDAUBlObtjz2NTg0iXnBEDwNv3tucJh8Hd7iTTeMtPIXzQyS9SQq+uJgSe/Z44NK8OvdHB2Aajb
kFCE/BLRFRk8mvfUtRsWoyrjzsGDjWp9Qi06JnzpYymt0uVJ6WzUC38CeUfrIp7EaxKw2OW4GEe3
uMTpDhW/YUUoWIwX1AClnUwEZr0wPJGyPJ37EYFbl5bDwidazINnLK8syb3GChVr3CPREqgpws8A
1Lla71cEhFy5L4IF+LlFvOWCYSmiBueS/alROgPP0oXwS/Lyslxd5JowWzjBbxioEZxh/m6R3KWB
v54thq31D/F3zJsrbUnYOI6Jpss4/LFjUlmUDBg0jsQYgM8gMykdZbG1e+ZwB7EvaAFfTn2X9hCP
HOhSKpmHlyFAxVs/5uG48iQJkD9kd0sEe/V7MCeeDWDm3bvY4a4P7n4igU00Sadv75JFwBZx7ZaY
5c6S448jy8Ldn0+CPWl71+Er7FJiXKC0Nor2tJ3Qvy1Y4bc+WebSYcejE+IgLDhMy/cCdpuIMVw+
KRDUBTcKn0ilD1aRqlwR7Cbmc3FwYIFEldfrcLU6QfikFVQTBhTSEXJRD22uJU9fw3piZ3g6UEwW
RfadFWtVCkyOSC77bH4fJlkrF6GaTzt5EwMZrKIZ7jjFpJvrPilYcvP2dLcHMnCowCSKmpETLh3n
XHlqDnn7xKO3ZTFwbCYkDdhDswR9lhnsWLiSkRF9Ixs4DLTu5YHP5SgoHCBEj9QIcZriSYj/ndIi
qpHtVofc/UVLAqk0Oy7lbooI7kqNlfpf4qL4BiN2X5h5AuZACiG+K0OhliQJM65KCaSM1cAErRn9
H7+DF5Q2rkb7C+tPAY2d0DIByd04mB3FemDKxyUkh9wgLDfiC/515wA86Xw3rrY35/5RDEVk7WJ7
fWRBm5dlnJhkCQEVa2fynokdhGQJn7M5WP/GQHUX2UJ+9WqVpz7g3XpZwa1gzJ2SuK9ijZ5Y/u4Z
T5SxRnIR18/udORhlLg+Cox3nN948ZhC1ELORSOmoe09cFkarPInjEPoRwfSodY86i1mzdslEvTG
jUW5j/YmT05rQMCve8nXP9YQOV444hDR3+BNlceOZaokVkx3mNtM5DDABLb0JePW64idLN6ln1vn
zvEs8Wq+Lnm2ZNMKMrCQYsPA2YOULyIxD03FI8cDZC299kljrPUFVY+YH1MHpo7e2dguOqcnKNxc
hpeqeQz0CfHIGPHOc4ma8p7o1PsjYvFw7stSIRP6RlLIDpIWadABvLZsEHbnqQp/4MUzpIumgLb2
Ylft8FvHpRDftdxnw/7gTI5q3B0c7ShyH2zx0V4Z091V3BGYORqgFXd2Pts1cjNbmaQJRetbxW/z
EX9r9zesPW74LIMRyZ4tYWohdfC1QqxRTtg5UW6vqrMMFVkbKudIzjbOuVmFx1gD58hoCYpML+i/
vLqVDlNKbkxZJ1m88kYnYMcrXGaeTfVc8dfzKYTRs1CGGTU3+ronlZO9O66O4yLHh6CSy3GYVtNf
0/aukHX1QXnu3Io6Jg3JSrUF+vqYDStjkDzx5cvrctMHHJ7Bnz98zoKo6uw8go7JJLks99+wkIvY
Zw6OVS8Xnnm86Cz1VHhmc2wXz3SQ9eoHwGSiOJKkjs85c5vjlPuCQLclQTEFMsuwH9MYh6HFdsz0
Ibz/12JHPnTJPBQ7S8lMxObgXSpb9D/0StrH6PUdQ+XJ8AM5klZsJ48pQVeo1IP7eH0jYDMh0Cbj
Ea7V3gl9mQuVpWSyZnQ87Un+WchaW0a8DYy9JNf48Ee5TJqCUzRluoU04f3IhO8oJeKHVtsl+1WU
9zExh+PSJPaBBqWfbvo9vEs74WSvPDIBAnIYux4pQlxvZeAHK1DiPt4akbmXIvLIG41YpuTl/bi+
G/zQ49f+M5YdaJB9wgYHzfHhuFwbButyfUP0XHmG57rHqiJ9G36C2O9k52gcTYZVE5rUFTC2yFj3
uwxGA1YE6PJT6CLCGFcyVjEj572qIWQI6ciEOvO8Fcv9dv58po7IsO0gG001d+h4uDr1G3QD09eO
KQ1imQfDaG4xgAs4omlKxS1Km2Xus+e7PO0Lv+Y12k6e7b2nqSeghLOWFUx8yvHISrTHaTDAd+BB
JjYIA37DsNw6IaOprfl/ItPT7YvwiZ9PxRsLM5+aSAKoCppHO1vEHpgDK0EWvqJ3xQnfyO9h39s1
2cIb1Vl/JOoTqzius/pnd5jcleNgB79xobZJhk0onUyXZXzQBhdm1ssFeOruokNy7CfjMxXP5wy3
uFVLanDRA3CWlMalTqNx64NNl3N78r8tcnc8kUTiYtI3LFI4+kuqY+Wz26ygixO8vIA4Br7UfFxu
iz3x+FsdPnXm/tW/pCJHSPdYBfw3sXfaGkAb5FtUH1tSdaUyrvnqhdMd125UCDGRq36wWbE+xn2v
hkLr1jHuxPaI3XOdm/hxs7Sx2dHoO+QmMslZwNVQiHCxbQ9bjtVCpXIFLJjVLdKdcOE/mxk8y0hM
pq/ykUQ9AiHu9BChygYLD2mktP1TPny+5vrPYepjb5pDk8/o9PxD+0juCOjG6/dIhYRy3Q+1NdqB
LwZKXeUmysr2xckCRIg/LJiT9viQRIxC97auOnMi2yaoFgrhjlNBl183gkWdz3Zk0Gk/r8u9ckYQ
Y/StgOqBX67GldcMZ+UM6zYUPGXFzXG3yy4IU0cM6rGVs02d7yXXfQD8ZE30cyM/e8jJUH9SiFv1
KCLnOuzRf7YATYMAik1/FzmjzHInRNXapXufgvnwQdeHG8slQ40hQoUTGXJ7lKi+ucBdomNcM/um
Z0cfJIbMZR9Mn4Ob7jNVFaBOp7HWHQ4hwT468xgq+4Xu3l8/k3yEEFDYGQidIkisHx6xgw+X8ONN
xq54Y+dtMUiClSFynAhpH81mwZ9URU7NWqQoxwVNzf7MFraoC58E+Me6gnX0QhYceg6WlAMtbe1m
D3Fl7Tqou5Ax//iMYCI+Hx1xlGRc+hHa318TZawB8/xkeFATUIEKsqXZU2Vz3nqyFiLszB/6Upgt
sRDBWemSvF4fKFOPDfFiVF4UgDuZJv2QncQMj74frECLrN1CPudfeac/V2/eFuG9bvNiqc5h3tk5
kpf6bL8jXB44ZD4SrIv7bm5QRj1GTSDCBv7cfmHeLr2S0qwFf6ra8h++BAj6O/VcCmyaIbVV0yAr
+oPK/+6bZFVZptDy9ctAoC7EULwT5ilpafOMOEae/OCXTqqhz0HWrOQli9DhTqRoMmWBxxL4+aQs
lJe1+dibpqKnTFhGWHFH8Q1uSMSM8/7BmteH/KBpIcSR8PphGnrJBoWFJphrNGVoGTlR48XP9OZd
0zfF21VKBFf+kDGpKgYPVAv+LFFk7HZn/KK8mUW/r/U4U8tzNRONY/0uYGIRH7CvncQ7JHsIc956
ip4S6oBnqCy3AgHcO9GRpu9ERmeKKS38zaOnq7TNyepsx/yGlLGJnTdsfatjNjvXzZm4o02sKqoY
3uKhlPj/iAUYYJhfnwEez6xYwhIZxUAIK5O9CVkygl1msjO0OsPYbDraCCHhQK9qTluZA+sBAu3i
cuwLK3E7E3+RG5easW76ZjfG3fmK/BnhcaWdrUuZIiE59L5UNIiEu86gub9szLqU/PEf6VGiJXYn
S5RLiKTqnIAO3ykZYf3RYiXoQXZg/Cg5Vlf3totVY8pQmlG1t+h6zIfa1z/B6i7rrzoazXT7W/x6
7YjMfUZftZlN6ky3VykDhvuuqYNmno9sUjIje6OxSbPwvW2hwa1kL9EO2AK+SA+JfKQUYU4ANILI
DW/WSLi1/tYiBVJbtZCjzuXM+pW4pGmPjt0XqkYJzB0YHBkLAK9MDtbyl1Yx35UvVVK/2RxEnZCD
4WXE2EhuEHeT3CMn05f98oFvY/7fWwo0wkG2j22pCbaxpa+YQwkK7F6hGMkjGvgBrCo49oLKEo0B
X8QYf4am5f/IGRKLGh3TLzraVzJ0TWsYQ1UE7S7P9uEcGnZu0XbhfmkajgtPQNGP127Tl5KYF8ho
7ofg3w+lO5l2otZ8raP5s16m3vjOgVqIcX3mODmqV7knrGP59owntOQL9cgBFGNkZ9+1ENYqx0kP
tA5ekVm8jUWzxMs7PGeVcVgjq2gwpOwsuLs9UqxCEz5wNCvKlDlvv71ZIiRIzwIXElt6SejjwMiN
/DqsJrzrQtBgHWqQ9HH0+TsepI13JR+j2/aqnvENC0yXxdhgJvkempTxg2CaM+W34EJg9FpqGqGU
WfaOle3jqckVgs67/fQlDfdo8RcjU0h2izy+f1lBa9L0QQPbY1lcG6Eoh2RTMw+dcHi5mos/4Bm0
Rgrmr1N4iqb+VkzX9ZrdcWti9xNVyeYpwXm9TmrZAatKBtyWFqGFJJE8gaOHC77NrAkme2udG5OP
oiIM2bzs8EamMipxbKTBl1zsD0vZGOPMJjCL2uey9jOzq0qIS8X2zUfioddZaFsMDimOziY3SRJL
kEZJ0K8tE9p4C7+92ZoQrb4PVWErdF01V9BvaKnFexEMWQlgA6TMKtRl/0cNk9XpdMgnGBZk8B8M
3/6SUjGrHm+o+7hQ1MvrCkgXZ8rflR9Pvorf35LHiTU8UqU1etndnkN3Jdgg03LSDDx2Dzj100RW
lJFSxGk8nJ/teoCPuVN1FRLzRc5HKyetd9GxecQfo0fxLTBWSKywjLQOHZqCb0AIX6IEuSfi7MWP
t6cvSyb0Bb6RjVnFmzngVaPdodwmulBO63fM4i0kvMdcKSVAcgRDJSPyo+W2RpD2ERChDXsnMwio
MBINpobBfaTiZND4MQdjVDDvh5temgO0HMh/yPMWQYUyyI6AVxY1rciRQH2hQTKlikfm/kXytu/A
7DkK/Ms/4BZ85SaARnBLQjpNNvokTF2gUmRhcpBWBZC9rl/JoJZnA4Hn3OtsXgRif2TtII7AzU7I
XCarCc7z0zL0ng+O1F6zYkW3zLZAlGKG3zTlf2PXJ0uWyaWte1LPzH6ygKsBQGmz9UY8V/z1Rag0
knbx/kLlCLRM+Cth1CBfBbd3eW58ouGOBbbT178TR6eOUwwNY9ofARx81Cp5Abv3TVMJf4qFsLUw
GDGcSsY3zLzSrWiiZ/GYVXwZndmrMnHsdCJhZTsc8wCMsqMtkFOack6AQJW3nWf0c8l6vaShhkWD
nZ1O4OkI2PWia0R8eoaTDrnizbZg39+gQu9jVGwSt0u3kKxSOUerDfD/FkGw9D7FCbs5wZZOtvRL
UzAOxgI+quOQoJiumJWjCqB28pfyfA4e7/shOV5yH1bDSfyu7ccPUIWYHASQNqr792e4Cw5GK82/
c8u05NruN2uOgsAO1sMGmZYikC5BJ8WR0GspLQwGwHF/KhAC/B8pqKWvDMh4Z9YSlTAkANsGdCHa
4sYzuitx9D+f5nBFoUz6Gr8hW/YORb6RxEXRqgZiSAFg/gto0ASjCPVmTxiHngXSV54zqxjZOr6K
Tcs/Ge7alIdh3f9jGAySvlBEHnpk9cC1GeBodQuS6lIMvud43+TmbU+IuP5YOiqRhhzxOhUjRYOh
wjeqzFU970VIyq1Cn6IVb/UBI4vZRUP83bOLaIP5u/dGtUxuiQZCxuZOoFTYO4q4s5GWZ4JWCgN1
lbTcyU7hZHUyFhP/1bGa5qt5RXhSS0ZcKj26/gSvp6oPzje5mDCoVK1f3dkXYZHmMlI8X/Ap64k3
9j51dON6qgGws5GoHcuG4/rQqc2YgyXrNDZ5m6TDpTVN42NDAvP0kRhPXgDA612agcfnca8QjRg6
EtHQitY1FsJz0Gt+7HIKRM3meyK0+sVNXeNmhKET05LngIkfbHhmgBQVNTv4xwnD0CEav5g8ZPbq
1hSa3Rxmj4bz2YpwVNJsN8cgVWALmfIdvxKjlntRe7xaoufKsv3a/uKFqj5jzaqDyAXODkR/zW0T
JfFOUg5PQq59os3owyfUPdkZ6RijFYNoUNdKA9w85eHcLGls+HWozmZiZytBh71nu58gXnRJ7uew
YDGOuPADVkxYX6Z1GR6JHTms9MJXZ1NSastTjlzMqYPGlt9XyccYmo1xL8xocm9BTyiqd/CL/NB8
zv1EWa7STtzQKV1yARBrFLG+keaqGQ4DtfsOOIcXba4FANKkVocOkTwYewmv6pBy1/s+MxKNmm29
G3SdTIHQKaPAU4m8rAusAIiXmCnJ1ug0Ao0FH3HpynZFLjtueYfyCjJ2U+DgNWY2eKcIUpyTFD5W
DmJUQol9g7AOcqQANBs1AFc5fg8VKNAAZ0/GiMrazvdUYoSPCtpS8ZQwDJ0+TWosCol5qmUltPYh
rKTizxHXFT7FVQrI0gLUJXC5OpGffDFMsv8P7QI84sJIHmrj9LWnI1Ac6E18d9WJVRzAxRG8+dYs
+gHbScHKYuiJvmMViW7ISYB1a01rDhVElBDXO+lN1fEY5ERF/w52Q9f89FO7w6I3qn+hbpjDyLWz
EcrBT2Km/5+O58EuMQaIp3j0lBiG6hjeTCAXgeAtHlC0x0ztSZm4PIyBkIAx0EsTDXw7Oc3Xvk7x
5FuNLgpV1VmGcIIerjCWsQ0N+JXmThTlmu9TDcEUXcKxqT2OyEWzzwYyOsqeS1xF5MftOAQQmr0y
h4lrgIYfg+Uc7suwkDhN+8LKU57GuM+XWIx9xaVRs9vOjenJ4R5DK9xrypjc8YqIZA/UuYATh6zy
ZeruCCtxkm1QNYCas7ZNQgcmrMRfG8Hcco2E7lP2fXOt9iptBXAudK3JobvYCXS4IScWVPSuTbX+
ozRYf0wE9y8I+1F/Edz81z9HUNwJUMEDrBf4cYiArttssOeY22O+LT60KTvReOXJNpGvSbWRFQIJ
0ZZCEptFMU0DdiTX0zk/w/wDOyJ6qaCwcJTJJ8UnHcKXdTViLn4Uu2H2SJPXommX1Hel3KjZ8dCc
QbzyGbsdN6l3OL0N8Fjh2jPbt9mc6VDgehjbKjCIsV8CfUeOWWXIqjeQz8xbJCB5/3KT7CUjBanM
P81vysWmU9Wr4OnfiLcC72JRdyYvdOUmgkkIObsUU0H/3gzb+qX2DVSrXordsIxddF5T2CjayOoY
oSiIahk0CDXeYObfB3Hw5gs7MMmA2q3hKrRy2Sq3gV2DbPFOJpLgRHWf2KuDYO8Nm9ihZVcDeJRe
ZnnIu3ORvNw4au7PnUX36NUiEgZHnRz9npiq67AgLfnLvrCLXbI5GY91pv+cucNbDg6KqegfPP/O
Vagh2ttfhbl0hKSTa8ZHrOPjogGcsgJPTzsO26shF49FIHqXUbY58xiQIbKNmHiMnA9FcK4egfVv
gg/xFIzHutRZvWQedTehQHg7Q+8Ob+OmmtmT+Xx/NqgkpWJlP9wBETbiaAnBHKMrorD7eH34DR58
g76amKzqRuTf1w4xdOhopi6U3QD47Cfj3lRRx87i9sBC7rJMa4d0Pa/EWvkknpkj5y+dfEVWc99g
gLPvQJNJYiBKYktiCrD9RmooXUoG+vhtaI690LKsblIMgadURgviXf8vU9Iw20J5Cys5f7N1bRt2
FAccmQe3tRpOUHt1CHQULberFqrF9Q0JDtEy7iB182/QKpY/aOGXXqxPcH5rQNRFMbI1/J30RVrl
FCwxTfw+eE6NZh+cS2qwGMiG88g7w4+cPFmC2HtiL/b/r52qdFIv1KEfkB9OO60etnn4L9a985Tj
bBqBagpvLuaKYkElKAU7X1LHtvVJ5EHDYW6RtBCb6PhSGlquRiUnvRiHmVXFkEz32xL8QULXWfQT
3k5MdjAfkpYXDyTdvl+pDS02olbe5A0Rl8krihLOjxCZKy/VFJKs0Xei322sWvqODI70bI0iBlV+
5sXj8+EZTjLhozZw/cFj/S0h6P+bofRwh0AnAcU09hLuLvko5ga1mJvX3SOZO5q8VOjqmVFVObi5
EO4fhuSS/HN2IJP+Ypv9Ev8soxWwWlT2UQT4J+WVS4bzimESB2600MCXRDXM+YSFYGwZxNAAeX6V
5WQr6ZmUbc3HQSYOqIg92uvSKf0+lCCj1EuQ/uMzoFSqyseYhOXpZjyHI18YNmXiorzsp7Vk3LCw
IkU6asQq4vw8qLm58axLLG9BqDIQx1jzTKab0F5CGTXFjY7Pm8L35GezBGtYp6gZqYoYdY4CIDzi
s6FjuitzKpZwL1SGxSpLpZy6nFOfUpNpqNaO6IVjcTE5Kn0QQ86VbN04VS5+3na3y2ciTniR+UfF
HAiM9+HwinDZCEGqNaSTD1U++BWw9Mc6zoH0cksrEUo7JB0T7t5Ms9D5JC10BH8V9ia1SxiLjE0Q
28B9K+ZIY3LKgk2OYN2mxJJXUHr5No4T31jdZ8zizORtUZ7/Dm4V3hxXTFeEnfZsmsKC4Gk37GXE
lXenhNAUmrxO+BJPA/w+m4C4wRwHx3TqRnvq+44HbI041WzwQ7noUeMgOylMCiDrqMERItnKMv29
s8OKJnVOaNd9Ir2/2eO08eqT5I51eGAP3E1gItgqZB5xouH14eVyRisqwd6ir9DXzITNjr4c8xok
/2zXXz4kWMeI8xtQ0DHPO9kg8hw4a3HSK18Zd9ydicuONb0MAI/rEokUrakObrTjUYAwScjL8vrS
mZxO0dP7FFkJ1FoKFt7bgWOX/S96owkPmwGH9SrkwSauHWPySd/Y/spXAG4DXfWjZ9rL85BKYQ90
h/hjF7ExpsrpViXz60GaPjvN0SUO/eHiP8cwGXuKorngVLfczqN/8mEat6AivSo5XFK3lknAOz8N
iISQaQyuBOOv/JAsnqKoHX1QLM0o/qRw+tvr+iL/imz6uycIVg+SQR84LikscXj5Seer6ddpLDcD
B5aViXSqpmIyQiDgngh6w/aoNJkQOBm0uOdhzLJP24TBjBDf90atm1a3hPrE7Dg9MUJ+j7mI7qDR
2vic0CgfSdXgXue7Sx0zJYQbRcwtsBq/bxTaqsk7TRGzmGscnHOyv/dGZo9SOOFMDd5CVJ1JslOS
SmF7HIrRmnXvi8tW96zkeesDBYd2LAYbCtGUiWASSPCHmDjW1MXBr5+L+EwOVjKe0gUHgMm+0Car
xp6ft68gCI/IPrxgs5HXXDz6pJPnwIIKfgy3qeMMA/fb3A8U8IOPkvhryH1A3EHDFCNdEHkHhcju
Lplqbtn6yczl6HQCNrndStXesxjEmgPG373/8dZPA8haL2RjWJPKw8AE6koSz8yJ1AaNYneQXEnP
I7+S/7dNy0hEAoY57O48WuX8rziikK6KE/5FtLhsZI6MiubwbPoy0/cBjjqn9KA1lUFCZMjFp7fb
eU3FogQhS08md+gBumT+5E4MCLqYPlOvn/XPORTYCYUUDQBeuX1Gnkrj5Ld2zl69UE1yfMrgJm9C
KJIhz8llD7lM21aLETDDS0lYBa2/cn777mlDRhhIkT92bjUBu2a07iLEcnEEoLtPmIE6de1Y/QQJ
d9Bl5gZlb4dttKrIlyBFSd64EaG10A235PG40tXlex1e+6Fwd99WP3v/p9Qn3Ow9d/QDzUF2CnSk
S0PUhRKry/kRMCLwMM17MXrGjArwt0pnYC9Wij5q779ptee0x/b+Hr2UEfQo55iGewmihGFaXpVl
aeHyh/COy/Ir7SoHZCJ5QiLqaadMTF9duDIH73L5UqbtKfMqUdElu5UaK5UbMyCXf69qxXZto6IE
KK3/PwohCjHfXHubtFfu31rzeN1GVvZodB17uIyuDciJs61Ak69zmqBs12NpkxbRMvtJWy7RFP9B
1ENNWjU1AhQ++lN8TY9dVI6QrGjB+xH6hNENXDWudipAgIRtEyj1gCE5Jldh4UvZN1PzAjVfOdH5
MtP1bI9ZPkp/8akvjlBVf9M33Z25P0hAhBTvCN/mZbwxwFVaPB0usZkwa0aFjmtUmwvUSGxiarCt
+skRiUHFWbJQE8IdFVGIWtlgt2upRPT4FOp5PhVaqruri3e1NK/HklJqMIuWfrljZdfdjDaU1oA7
G3C/Zm2oibpiPebzJRGSBm34V3oHjIDV8rV9oxpQ1IbI13bHfv9SCBK2QjslcMVch1utxrp8l7mB
1C5TZNUoQSKjP03HlZJdPa9crbHUeFpGgsaQSD7xB7Dt4o1KdhF6jrHPxpu2h/MbXKqDfcGiZF0N
2sJRH5Z5R5e081SBREfydocJATgnjmwi4/MqJVaO5ixPVUtc0bjXKKHdGPU31kt2LRbxEKW7+fmO
J2uGTczI6fEiLo5OKTzoRcXeb1pV0n/xVHbdbeLTqxbOwZIF/vV8no9dnRIYpFsnrYqwx3Sqb2Wu
vpeJ9tcensU2NMQ39lzix2B9aRIw93TLYqZrHfDWB1pkXFcfcjYnBJemwO9LHF1XaBt7FkVOzLKt
DegA8jwKDRnhDLt8AzP0AilFSDcbh82n25wFkikUUNGhb3bIaVIEsk7a06BIeour5/9OMDIH9OOv
JBTxGK3agWoNsfCyD5zWwdvH+L+r70bZaOiQ+PfWrbyeuRay3n5UvbXUrnVzVTFiTy9MDxrzqUVe
7VbjTSTPDftYPOqw+62HLGNUgWKZt88yriJutudrfXuuAV3d00Nolu0FqT28eZWFqqKuyt3kA0nD
0o6xojJqZngNh7gzcUzvGJtW1U+29yPw8B49TUTIgwwtabojjwv0jM4NLaZplwcof1nClfn37Z3B
FBwL/fb8/HgH8gT6hIeipeLfPbkLYJqbVVZoNgVyysXeUP1J6hODPRDKtk4m07r1BtvtcZLdtlqk
uTVghhc3sg/xqGLV/kIN4B/OfpxmbdTSswbD/BDelnGoKzSkb/mlviRJCiNdHA2Zj2Oq+awBqffI
PlZjVODhz+hPN5xCGJee80ixM6VvMRynpDAW22So+n0I9tjE5gJPImzoTL11Zfj6MQvdYnXxGQ3l
cYG2iavnZ8gBI3FhD5Oqq5ipFP6L/GId37ufp8R6RrGsAgvrI5riRObXneGIFBhkHrNjXq4nkTSV
TGdPzn9tXwnJiJRBDxqu3ua094gUff8dJK35K5AbA0BfLarV1CJ4smRIfW9Qkcomxyi/ChxP+kcR
uz10k9UqLNt1hZ4nidOo6t618KPZ+N9z+mKEW7Qcxlwu5Eimcct3VOrcn8UvTVOq60naDvkwDOH8
XcjTPEXLkWUhgwR9qTHBaqwBW/BxYPJXFeXqbeVftUJ7/pMB9jzHwLk1nKFoclzefAtXGWDltEUj
OJNkYAD/8/+1gWgwD9LHaUIMGj4mpy14bU8Hmt/SxX/I1prSZafThm1z5hUQ+8ajAFxw3qFc96E9
e+QKKaOnphoVEMD+zkieCTLldTPISx9uSTGof4moJnPaY7pLLqhXAa+Ij899QQZ2vChs0q40y1IS
TuK3M2avqlmBAiHm2pBL3oZYuY5oQKBHUGcQgAYPiBfliBEvwpAJibAk+Imu0bwGYBVWTpjcbOuS
9Pnc53WF6Xb78WxbcGX/gMjpGvPP6SWLFP70CMvrdlFs1WiUca9n6Ba/a+HBJGsZQzgYwtxx1o0o
mUKK1L4wqDRI0sKFQBma/jS11vjPkFc1CQJGX4z1qI06ATgFufCA8OTVGlLNqtXAg1A+e59+tSsZ
2lgx+pUlOKWDjsjhZlWIgE0QQrK919SzmChhdNrEe/PSF8kd23dvlEff4lEOKG8btnrij7jJKNMo
JW7Ik+tPVMFRYNzOdHas+G17D+Rv4moKarjI0EueM71HaIzxim1vZB1r9LHKU0Kk9TFZIY/J600G
ae9/GO6GFuJqWk95WVbt7pZ1DVWG3hxagBUfp91A+gFQlp7xxRGb9TvrMa0fiy9+v3eIwIw6xWzH
+lMmmvwf+8D2SVSE3dAjQ2st+yegc9+0OPzWcWQX0j3jlIYYUSp/eyafbdmTRfGD6z/ZHqDluSYW
cWarsoZ0kayMlvWj8zB6sTZhxwsX77eRZRfamZZVZYlfIC2lxpYh5gjrTef1K3AbaWyv55X3WTdK
T2Eqv6eJ5zFES8tMBi5q3xm3J2xXn5ohMUtiyR37zSt836uNczLeU6Q421tATWyJdG3iOyA7EbWh
/yzSq0kNO2Pc0Xz74LnIqKl84n204B2BpFBwquzdBkGF5GSBmXxk/PkxKaJ/TjWmwfeSNqfkB+JV
yo2kQlJ+/csTrONM5GsCqLzsVZ7QzW5a2Y0XbDFQo6c+xtG0SHx945c28xeTAZdgMsf9+cKeV9Pf
ExVsKotBLYyoRPulSpYWft01WK7eBzLz/Mj1trOBaFwZxA8WhTdWZTN1cJzbd8r3bBDFFGKJdcWx
Yh03TKTYU/zI4xk8atmZsSlUzRpop+RpDZqnUDbo15OfXetAb2TFg0Vee3e6L4RRFE00pdqLmWiA
BXgE/bNKlGuVHqAcI4GZwLx5rd41YOOjQu1QKdLrxErUHJAchUMpln3mPFE8t1Rd/ncujGx6i11D
mIih9gG+CdcS8i6vmV3DQyyiP817fMQvbyUzBKaF97n7+5DI3die2gJJH5a9vVpRD3R4tGWNUgAV
61xvEYcNZfJAxvl6tvV9doeqwBufM15drI5ASmppG7uU1iOCoWLLlKxEr+FV/K0pEmbuNp5zVIlr
GyPoCFdtts71LZeqAqxV/ZJgmrQb9Jz/aCSWx0GM/s2FT9lFPwNJ/XWGulKto6rsfkU1u/Lw8BUe
QGqOtx/TXjdLopbxsAhPSLE+NFYLNUbmPZTX3FufLa+MAuXfmWkyKH1pmN0V0PlTaADiN4m5KKsk
SnZqY0tAbFQt2RqjEBubHTvYBEMiJv6HWc1M3gSmKQVk01BgyTMqbPOUjgSSivkMb8+8T0vNxOha
Il51ftJ+itSjZvu8w8d6aQ1zWutiuTGhlhIYgUX/YDU5+egctx5pto4QZzq9SVBZN6Dfb1jLEhiq
AZwUo+a+jRyfjU0LZ/cXEdDdajwthdxPUIagMFStCfTanwoplXf1JhpLyzKQkNGUE8jyEraiKiCo
Xn7L7I92nCtZQdrxapX5DL9WvWUDPVC3fqTooFXjV7O5BxufqyOylg8nzbtF/HwSV2w2RBL+BghL
hi3kXbmNjE9vXF7AsIvT+Wt/vgnzsGXwzACbp1EYCN66arOTtA2AILYDc2jYRNt8fHNHiUnKFNE/
YnbmVgDLrTc9nhmg7y/W0BDdD0Kh4vB0Cefm9MQB78ipViPwvXuBbyptL9lCwDmNz0kofbA1iksA
JkXvhg7qrUznRi8nvHI3QsuxVt0sMPSFSYlNmJ0rbIhpv+4DNqqIgzqQnovWhgbI3I7GJ4QYxfFo
5uoi2ss33EvnGH9OXu89akVdUrI37F/fqh/HCnVe8iPP2m13UMkxPdU545a8PghK+F5Knep9iZp5
e0sReKac/SqjkStizU2DXUf8337E2ixIldNXk12lpWSRv0Z/hP7m/MeDS94beAiJh4VY1QQBUk02
bgeqiIGXSTvF8rgzzZQtyDNGOWkSUyLQeOyJu5lSLf1LiJ/4P85G5E0xPkGX+g/tJkgRh4vhW3mT
lJktU3MOEtSsamJH3oaThnWNzGWvT3szBXUfJlflrp9cpq8iGAaecDjHT4gYLq1PRcpHOmjuF57b
HRaBCMAj/DZ+aKZP5nSrVMV0kSd7bdhXYtKaV1y4rPzWeltSbyywvpGNQMWmD5Fme3VF1G0TBHN1
CrXtiCJwpKfo5HWExuotzPybB/37EZ5O5rOorVhmAslN0L7sNt1V6yl3VlE8qcDUdECX6o/utIeJ
nAWzhpxcLN/zKthzfRuW8M4etdOvc7fff95qJzOJLtzXgRl9a+VoKCj+KCBHCqaKNRhNsOOIXm9g
+wJEEqtus9K9A/Tq7Erz6XEJfdBNFMjJEIKX9FDGF+x/NBHowNSvGTrjPS3LyTFZm/ow772LmE2x
wSpsDmiMQp6fLdr+OAd4JvSWcHhHmAAoBLfbV6NpCQrAPZHjMGzGP1DnQ0AoY51+NAxNUPFUz8v6
t7wAkbxhFEFWE4pXtYosLiX2b8ywfvfYy4e21ZiN8VpjDSMAa7DeMilpA8RhTa3fVE7o0aM8q4ZM
S96JfCSK1AF5WA7Dzjvw2athTkjjto9H3z6CWt0wi23kgED2r+boAwsRALO6i9LKwrXyMG55Vf4j
DerUligDWBzozPMmfzHWPys6Y8ZYuj9H7oNyiGPmTrY3Pe8DQPcaKlKFzUTjRE6iiHx/F3DY8NQF
00ptnjmeQJCUqafSSQ1jhBcrzDSOurXlehJ/N1ZaLAkGI5NVfaGg4VUzROV2BMPpbxtpVDCs3mkX
vnmvgFdxPb3uyGDC1fT/9GOnWbiZ1Vf98Snf4ciMN7+eht3mXmxqrNGEeZPouwuViXwZUt3vp6WI
sSZnXYgcIarXz71+ZIT8zij20LEAUc/vcKWJUcrGiwKFmptnUnjezgIyF92809ZUsXdkm3yX1JSC
TTJprorlETQOiC44fBXgMWB5n/Xg08Mt1eThBbWIn2uJB+N7kwsyIjmrh5sPqSUXfWK77LzRcRyY
iSz/XVsu6Cfr+ZenYe0VmQXVlqnNQFIIA6PuqAALcyemLodv9JFKQs7hS3ZTctzAvEU0GtFIOPeg
Ptew0DLk1iG+bpdJYjHwahPURWQ9uDjpFMTgbHyVqMNKy72IvQpvZNKgfq5TRZwhVqIV3lk1mxxp
YI/9rtqf7Ug0G3G3GI2sacuWMQQR6oNm/muodAzSeiDbfhTNfGN/5kFcwLq/FBbeo4DUscJ164mL
pX0H18RU9rGho99bAqPXEyJ75p4KtkfHcMBFWcO4in0G5ID8MUQ8HIhDxWIuXaKkqEcQUKAGimkS
S2bDrYmdPGF+zoiVwlAmhoQwdLEdUMN2p4cpAxw6GmSR+4rB5VdxESI6BXalC6eJTGgeUyvNDobe
F7r6TraNh0jCziEQ9eEKBcALPxXIqW8n0wtlZPlxXyEF0hmK7V179jZa69kobVoGP7Qd8ZKWFt2D
UWcra/s9lHihxKsrCl1NcFTAKGJ7j0Sony27BkDwYPK3OMAlHB/AmlZlTYC/XX8C1QKgP1VrCFtg
w9kQK6pInvMt7DjYIcyAQ+FDdJo75pu03TU0WwJ0igyhd0e9Bt4Saotn3SoZlxca5dQWCvEIZZCD
flnlMwWjBAupuxqaLU7a9srXf9xpkfJeSy5XajLXYMd2QBmfUvJntPOBMS8YG1ybmmiK/zgHEf0/
piJOQqpR4rrfNEHJAu+4PLQdK5JEdkIVWSOUlNsFJG1OqI5TC+ZKl5JWWEeAtusWLX481+yc6Sed
VhpQ45Eg0Ci7Ru9DFNDOKD7RBZTgeOunN3qbshExNbJXHz07iO0FuiQ87BziDHfZUkQV7uYTH04v
z5j0EvXgdeb00dwu1hLt2/8EXxT4l22KR9n8yVb+RRtgqaq2uiPIpOay0two0mNuzBExnAIM6VAy
pxDo3hQDoGo/0Qq4u7C4RUyVKItimAbXtjDEMRa4MFTU+qE0iuO+IvAepYtZiOg26b9PRHTMtzo5
g0CzdyC1/GdFu6jgUjHfS3QYamiTqsGQPe9+ipQ2WjDgv9Ii4x0cQcqavi/Ppwog6mO1rqZIUes7
taPVc8zwWX9eij32BeiX871eQYv/rMx/lxJTfu1+orS7m3rkvadQgaKwvxjglsKh/Yl9fkT4xcJR
FM1WG3ZrhibCsnc1gQybxtG8UN1qxME4If+zqO+nqrOsU+jUi9+cMzmd25TfB3jct/m/SgefWhs+
3x43aDs1buYugXUDnJNSiCuCtlspwFph7SqSMA+lfBD+ALEJtcQsAXD5QoDMRktBIx2ZFJOmHgHz
+iF3PkRKJG+IUT1MIAIBqAInJM8zGQBcRLCFs0ScHZcBr/vHyfnMnjgqAURz2VpxQRkX1jIHrMuf
8iFEJM1VVeAI5t3Mvlai/7clq77BvfW7JKgsp6+X1tpb+d/8u6PbxPLx1/bs0jbWM5Qi8S6w9knd
hxHcLF6NDv1yMVbC3POJRc+cjEgM0qE8f2IoyOw5QrApt0FbVpuo2GhfOdRMoBcAD5JZjnVCO5U2
BgSQGSfYKuG8LY0r0tJErY3+hD7WmbU4UcUjOFGX9JfIihw/iU/3WxxBjoylj0SzH5nj7gbe60Ar
0hBPDsNdevi1lqvn0OWVlP2sAArztQ8PaSsAr+Xtz/D9+GyaD45b5FlwFHwxZit8gtqLwWOSWtcb
+8bt/8j1Iax7L/vNJeDSMdXPvMAAQkVAJMc81Eaue477wlAIclp33O6iZ60ghxMCq8yQ+54fh4I7
VsmTQTOwPoA+bJAs/FFkn4k2Tr9nCrBc8oM9JMOJZEKdrfuCsfLQOdcG1jGt1HhD02PL8BmtCCtN
Xjr2cFYDDVt8Vr/vwFnuLnzBWjxSKcyJ1UtBCHYLu0XI75q03UZ5JQtEbhRxDP/Qfa0Tu5Fxs5SX
IzeUyqHZ+JJvqj+bmPlNWSac+++q/6EV4+WWTjdAlBtR7uPUwOKEvHIAMDPhoVTl+opFQyzlR5xd
9fkGcyKhX5JkUnOxh7nMIBYuW9HMwACGjFqnCaR24l0DIgTq+hv7eHhvz9gywl2nw9ZdLKMyQR7t
JkGPEwj+hgQiIMxvl1Vm67naELIGkbPAZicOe1Q/MnVnJIvWlkoNdquIb3Yt6ga9jLgWm/afxFQM
8FAILHbKZt1on0IO57kXFrF09FYKkzEysgK0Cf1nrkJVZebtIwoJI6xdDuaYEhaTJcqAltg1RPW/
frRdxlgMOAAGKVYi98rFdZRFN5jrApxC4tmAYCtKcBG3e4zc2Krr7KqAzFrvILVbWlvsaEeHHsPX
cm+G4ysNFstce1x0VxeZCc06SmusJliDO0QGhlS5ipYsT6DPYCDZEfYGQDvg52F1aGsD2mO1Out0
+9+vfLzngdPKknWwJtPD9PovTu95U3AKcxkcRNwCG+LinZWLOa9UsX/t1awF1S7cgSSCqRD8OpGH
c4x7vuhN0T7kdSGTfFkoyDXiskz9s80MXhXW8NZHgVbKT+yGBa2DmcjCjXvHshDATwQMePMhHs/R
9hFEUulefsF5N3OmaN6ZiVd2Q5vMqMdcQRyi2OfVEUf+SJ9zOPdeEGD16iPtaD18nXZM7q896rzN
TgC9PCULYvBGU3KTlnArHZiTEgh5RwWGurZuDrMAjUW5sRiE2m5jOxMwRqwOd/WeHT96PCVN5K8i
CkaFks5E63jnTk73RPX8QacWvY15hAlAcJMosc9Z16qDk4M/Une7QH9eJbMeeuxSqY0bqacK+kSx
Ryigz2ZtuFqu4q9GWDc6EAYSJmVI462ghimTgd9kedzFfh5RMubtgSP10jixvBcnhnC1qfrSVZAL
p3Rh5k2Eoy+imDue3LxIL9ppNZ4WXDwmORGv2jOMFodWAXWyrXTFlLuEiF9t5RPEYTR2xkdu90Dn
nmR7mMML4IcRG0zmVn15y2gc5aoMSgTloRvW5cQ714nDlFaDiBuYGKYOAfzGJM8o9g6ibyOTX3kz
Xe8lh2wUY7vsRxpP559y76IBC04NMRvWn+QUf4jtIlRrr52DTM58FFVFLIwHhfWI5SXWVWBi81s7
M/MPUklVdWJDCFKeLyOxel1enWiZskPzG3uKvPK8VFDNqUqQTtBLinIjeAtK/BIOdU3PwNhLEA2W
Bw9J8Hht5Pq/oBnfAF1Etmxb8idI3QvpKxY1PYqVfSSn+vW/hZNVcWZ8PsJweZnU1hKOLVbQIdNX
FJdx1oqV3rVS+arbOxMYzLiiXeHJyNkyI3eZB7mF6PD+K9fTKOnSYdPDBK4P8qgSM1tZ5E0kNxEU
F5yemUrTcpaTU1h1WyOMybX0kMPwjo1AxaQ3felwYL0W2icCJKhzY++G0EWDR6PK82yqnTyN3l0h
QAVl3GS3X9wsGtUhVX/ZmlZTUSmD3I5m3RtUQ5k89BGV52DjhOsSjUMYpOqwb0qW3Y20zXLsxX9p
NmkQfxoxDBhBvdiyz+X0X+N3IsYGik1T1+EjnPX4aPMB9g/g+EPVwlpjx+Fs41BeUgql8+2gWXOz
iJiv4PH/w7xlkwFX49REfS9dSRS6+/xp7/rakIY2tKepbq17b4cMZsYTodq28uyQdBvE6SPgioyl
fXCUb3qIKZLx/xOWhXky9BChPI4Vfsxw/Ur22iyDyBIjWQWuXFsu0b7yjG9ct2xaZyewoN6SZnnl
5oTlFOuk2yYsUtkOmrHEVeWQa+I5407NnlXrSmE3gYIhZIo/Xs83XpB84mK3QrBQFrLIRPJGO5f8
/RS/EfrKMko2hpk2GXHRjmWcPye6e38+cLRSZdYk/L2CtGSJymmLfWWxtACezFURXGapdT/rdsgg
FGNR5aoRSeA1nOMlUkFeAuDa16hrIpF2nR+FLm9yFIIlCiqvyu/HnR3Xk3D39Eu6Wdqmm97Lq97g
YFfO6NBHq+nKnxzGeqL+wS7HIXv9wt/J3UWROAld5alO8xV1dcdd6wG2aU4nUADc3DqyFfdtI4CE
K+7PsXHavgJRAWKtireeMH8fD4tOfnYvgSHUqh5hCDSd2cDcpg4hrXHtuXLGjMlLPVKa/HqaDWNd
p2eVXp0ilp/qfU5owZDpA5ol9guSeE1jZeroetNfu2NAAEeUbQBkpq3TjL1gR8+/b/C+qFuDDIuQ
fwl78Qi5IZB6csjZcPyXP4icc1rsKiao/R8ojOeAoP3mm/yd37p4zfDqn4XDrRROwkJXAR0UhzDH
SPkxj3eTLgLPEXXKs6DEpuj6iPHqmYBOEpwD3EBOkmGx8r6honu0BQzdtCXfh7PXZdg8BpBoPi97
2kdGMK563I+wTLSi0rJC4Scg3mNxEMHh5U/fMEkRbVeLYJEt2mkSZbrAp85AvB+NX9zBjORUhn3Z
IKQMF9XYbF+Rao1jieCCd1+70JU6KgAGxYIQHJogQTyTDTi9U4pco7+Iu2b5u7CrM8RCjjSBE5Hl
cusknIRC9ayj+kJqnTZg5qLGTb6pzr/NBJ+NtUeYtAdixBN3PC2ml/PCcxmGL5NK55yWi3+Pa1mu
wz7xl8NX1EMlsbgmbV53ze607Hszz52I4sYHTQYl8h03o7NMFlzdH3kYGo5ET9oC9Z8c6PGQPkik
m0wRSRmqnf04gtZZqf4ZH/kb6E+o7gmS3G1Lv1EhxnmqYiUapcRI2tT34PbhLS46DmpjyKTmssxh
NFvX57dQJXl3G4wgI7/HZ2QjK5+lRD7cBIASeMZjirt7lfHq0tyoBWmTux3JDLgEPdB3hKDQpxQ5
mb5ISSYe95Rd2OWA01OlolJ8vR2nelFQWoqMlhg7GLPdQkPlOUq8a/jZI0BweLC0Dveo8nEnvElC
Am63qIJyIfmdEBQ6Q4VKGyYMtn1j1tVJdN4adHWWup4QkPK04mAc1zlY3Yk3yXcnWC5ggLPGTfcP
MoKVvEPFaMqcVEtFd2dLGB3RSzRJpowU3o47MS+tx3AHrhTl+NCOaR8CJCTGZEcjCD7Gz0Z40nql
lVIxtr0qDDbfBdNgoa44RxRYAf1GdYlXwyD9nYNAD2qmSvDAEUybTfab+CwU7h4UuF+IM3Xvqjkx
tmM9qV05XAFWwpY0EfP9Mxab4ces1Uxk/KD5i5H4jHzTNADU3MhiavdDwkAjTsZHdA5ChhCR1oAK
zIk2ywhfCmp8sgQVxRpdmlCa2ywZWGXDistfTTbazIjSQ4w/D1Fqj1vJNLUDMnhnptLEGntj2F8Q
04uJHCmgw5dy+OUMW4CkuZO29ItR0J8HjcNCgfSaL5HR8EKWvyJXZk7Rl5aPRpFHzuT7ulZlAnil
oy3AgxX0hAVDldMrhykFKwqtZPZL/bxhNV/rFLso9Hv45Y18B3jGRUZGRD2+5OLH7qN5iZ5ZcnZz
n7NYJnBXVquTHzavufVWypaHrA8kSvUTgklhAlCVoFvo3fMixSGosH2izXJgtNtGXcQbxMtb4Fav
JTwk7WE5Nej/GBdLA8B85tLnKhWnRdttdSi2z5IugEa43um23l1M1GI3uj8M2XPboI6hqXEaLQiz
Bkfx/jAGMOZRA9wk7QQ/LIhgl1jn8zy0y377FMPYxi7+RVRNzVJCWys5hblLydXYSdVCrQWfMvyZ
mrqxr6B8/LGbUW7zOx0z7RelK5THt2HygdZlqIPS/nCa6vxv35I/CqmcGzD/cynm4ovc5aw6SspE
Hw7sFKtAGNKmV6m/xwLuoJnERf+QhT5iRUNoRG/FDre6opR7bt9Q1MeAoWuSnK2geC+fCKciUcNr
vWO2pcEMwHrSdWFifuLx3qBkB7ESffvMnWdL3JSjqMqkN9Zz6z0lbyE+dlhMkK44pq8blLCL2VnU
BqRDiMHOZYvha6L5YWlm+EwhP0qF7Bg4qQkuK97TYcBjvxbFCCArAvkf62iCJcWPznqRER3xIQ8f
vcKH6pqlXL/Dd/4PVjOClf4tO8JAG+cp+3M+DZltqssUFmmaDX23msJKehAXqXfa834jcNUdzv61
yHKTm4eSh+DUq6bSXueoCl7p480YOVhSVsG2Z6h9UVJ2pmVITS+2mVyjpEFwRQYw2vCTgxn5eI2U
fiKwcycoKaAVnmMFE+Ic8ze4tbzCjijf/LvxnTQe/W6KV7UUmUHlyyBvCZIKSUw4QjJjrKx3ueUC
sc5XLqcRB9x7r182Cf+NWMidl1aIz4f171/EXXpgBprGFBJFJdXCIQ+QdnRHiYir/VHM1NyYWT6E
nBbWjDMOkRxje4FIk1/DgiMNp1moPxw8MF375zT7xVzwel0du/S+a9QS3Uz4d7elZD32dEkMMxDa
MOiw3HALMTI1Sm99CkauYa5/gHb5T/rMLHRmQzG1WRQagUM56u7UdYqeDc29RzWoo28LKLNCDs9A
z0eBq/Y8rtrRZX/LbC8JApv+Kb+JEpt670OgGbFkgoX1GiGlOqIqxS/LMPPiatRZiLOB2DB07wEL
2rviAA4ALJu2ztDJbV3fUY/P7vpBNfxkzIrS864UygBIF4k5WsnYwyBKfdqTiNAHoDGxsuZlJpAk
2Kk2BbcLKVbHL9xSd8hyyJPbcO9UCn3+7Xb/qNHNwNdwNYUzj3cYKLHiIodMs0bWaTIXM0gVTf5f
/5WjW+MT4iKNUfajtLfK0g+eDQEDZKXsgLJyJRv/CYAnDPLlhwI1PzuiX5cE2IcJXwi8cZFeKqGq
SUwKnT4/ovTCr98BeDLedHeJjFSFY/YuP9rfsEe1nGcPWlozaN/dbG2MzKal9Jjqkm+sTDTMOm5y
XciLRtxERIPGAXUSXztPzooQWfEBGbYyg7IVsvWq1HNdwJ7cDpEMv+QhcRw85ahD+CE9lu+kkC9y
Gz1XYju8kQWr+Q592W+Z86HmrAxjZ0O8dXarDQw61E5mBilnLLyzCu+nT4o0rllem3RJGy1Co9WH
Ug5ORVD/b50h205kGE/3sPehTWLTSIDquWjXLzfnw8WZAUHBESMhomfxDjMVuvJQSFEYjTeVlwsh
Co22tL6fH8xX5OJB2bPTIdrT/Gc4oGR17gorzVWpigbHOY/yhYFrldNHa1z35Quay0dA95c0BBCq
bwGZ9MPRBRb7Xt3fmrV5CuKckwxiw97GZgRbjES3rqjFUcBTXfNTnjcK9TXeW6ivhBFQiw3tIU1B
pbGlHhdoKDqCmlNjUU2H6Ad1wB8rdw8PC1BEWrXPf2M/lTpAV2mXJHEASayZJTrgHfTUuC3NSoZe
5htSidzbdmp7VNblANeXKTSJDXuW9KcBV1qQrvN55DE5rJyoNJrznV80BuQRnO7HEHf7C7M/CIzd
4uODq0M21Bhu+X5GWf2+PbzUQO1gOJ80HBab/waWw9wj7bEjiIasvMFF/OsbQ6TldE6MZLqKGle7
a2p0xZjQz142f7/Rq2aN2EzClR+QWogXruX+WOKAzXX3OveDbMd19noLi6JJX6pW+Bqik/A7Soju
tsVeFIsXZb9EaPVTHWc0ksAEPocAjxXd3wj8Fv0vrXRbOVeGeBXWykzX5yH2aiAcZTHq+itKO59l
xAGYhbNqM4aUyk2nLqf2V/gYwe11A8RZE+o5KQRv5WFUnaTJJ4Z2UunQylYGxEmHooIOfDJZj7+x
oBN4FAexQxEmwTW4f8RNolcM/E8kC11wxTJzBNLeLRsm3g1rpKw/beFOLFab1SZlYHYZ4oaBsWY2
VFVqJA68rZyVdWAg6z4tpIqkECrZftog7dUul2Q1mn47q5cj+Nlcmqdo9TikftlrhI8V2/YiRKay
9UGYkEIxQmH4hYYeyZ8T47nBvNYRrk3S7eA/lN91vSK20sbCVtS6qR/zyTSLpuNvhRRVn33Afg3a
xU1YITY1BCwYLx4lhbV0npgmRSWH8QRG7OOePozl5QCVh+cEzFsasdW+M9IfXkAgwrdhK3mVvh1h
Sa6S5ROBcgJI6OPRoJJOEwSWUjOeqrjk267YQ0SYAOTLUkDwmp1aE8APcNUjoSJMtmYkoFTOBf0G
8IkH5/UcvMFeac0dI4VgW5a5VEoJ0eUez54GZv+xz2ZCUcXjnqyHSz+ZuHzY4eYPrn8qgJn8L7LD
/YZOGPwUIWab2JzzTvyvmQAhdA3L/aK+yyQ++RWYYbEXHuQ1BtJxpc0KNWX5QpMZlo92BAN4Zr5S
FcFa+EaVgQIRsRnGExlATV8mlFRNJiNZMMJTnwCMtNy+gxc+Wlb7vYlzgRiHDIAPaAkXEBrA1oon
K4huMyKTMzyF1ENTdpzt/UsolzyvJrEts/UHiQ0jVNn+b4p/f6AhkX3xvhgJggItImhZ4ak4ksf8
3M4yi2UesYPw1W8Bx0//ncjxkCER134RBkMfxlNfQKs8rS6G37XeyQUWSEFlSI4Gt/MSiX1XDzdA
trTOX37u7G2PLwSbVwIVDj5Nfef2JQpf/vt/3d9XTNtXpbVHSFsme2L7lEzLlehy7LXR3eL0zhIz
zPgOt0BwcnZImT3NZ8SuRjtZmKfraEUKJxohJUp5xP+LwjUweB5SObg0Z4Y4KK0XAjDt4MAeo6OD
7jYSmrqroofJR8p/jXdi2O7F5zwAe0FIyeupbYuPIhkgb1LW27yAd57Nqx2OUfZu6HmfAw69FLhZ
PRCrGsrf4zQDt1fzH6LippyDV8FMUis4rCfyBh309eXkqWDA+3NdH3GHg4GNWp1AclJ3rDWJBvLm
lUR//CCN6VAYqm7e4GjfT9Vsq+Qta7EovoCw/QxytLd39YXN6MBhCgv88ArZxD+dsQLD5drUDwQ6
Ms1uRtdN9EAf24e4ky6xnX1ZrV4wrQkd4Lb/8RmVhjVGqQbJnXRUKOPwKwmcpPw3UYfbiwCOZOaz
AQiw1pLd461CugZnAVbTe9H9OfNBjq0Z4DlWQla25+RMef9fImzvj45hQWmdBjJHDO2yXG1uxdCB
e13UGy2+muq1p+YUQxgo3DyOXMxWnCQRgDUhLzxvMHOMHChQxNZ179dNlbCnrzO6nGdKzgArB04w
cCVbpYxdTHhjU0OT1FJPmLegMeefFvEGZWXL1EoK6hySCUBI7MU2fUx3mB6Y2HHdAYbHDjEid1HU
FKdHoHpPYdH/W5WAus3IQY1LuX0FqMx8Ea6p9VHXbijN+F/X9sIsjbGkrSrxNSh8dwX4p4cuRxwR
k3V6BMUxS/fagf3HEXCkfomESFkkwyVT9/jTRhVO7bbb8OGB1vRCT6gznl7lqffyiwyAJvsr7NnG
KhwPCaFIZqYPT4DkNLT53uAnKUsQ2Xh2eIlpwFeJ8tQauX6a44gQzzuiBh4j4WjGjATia5sWjv8J
o/fQ3lT6BQJe48lBUWIJwIgMbzInJl89IqI+3jWs9lqL/f7GhPURj06KgXtN60qDrPqX/NhugTAl
7sj9sr0Ncv0CfVc92up3bMg2TBCVWmKYJtAokH5iGMcu+B/arXg6kdy7LHNKMMzZ4SrVG74SpYZO
HmcrzTY+JzJtfTBy7q3xqXt02rcUAK53RXR+IWjpGoR0fgvPqzQRqUBU9+ZKc/N58gXNpPh4E5l7
t/gd3LmUWcJiltcPt1xVcLJTWHBZCUx16rShk0NVvzjLAwvGmO/qwS14H6gC5HtoEOVRHy6TNaJX
vTyRgwN2bnw+4P6A0v9dO9RK1TjQ0nxforld8aWKkq1DCAC65jaGOWwVuijPUb3p/FmU65FoRKji
VDP4skLj8XmikPO/Ir5pndviYgm6lZZrTBkbT8L5S06dRkK/0qW/Hfk4HNp1Z3o+bQB2xLUMxJyQ
Jip6a4CQY2cVonlFeNeihCEhobC53UWglxyubVHOWAobMjsNBnetFf3uAjl5crl38bcqWKtwPnuT
XgJiApvNt84tquYTEon79fE/klodkWVHLcVv9N3rkHzhLXUevnQmlcHFN8pz1CVwySdK4sJo2tAM
Gt/OD5Jc0yYOVDVtckNwjyKlSD8Gnfu4l4q/aQchfkT0VW7VnbLG0lmAHKO/wA4uP1nquHwtuuLY
qa0cAKFPlnm8JxsoUsLabcJx6KFS4Mv/GVAnOzkg3FXpioNJ+e/DUAeY9wtQtJ0IdremzX+w3I9j
4KcuiklolWqFoeCecBw1Q1tMM7+ZpvsX1/vV12jyAkzcnXW+R/ql2VWoKx+zDnRBBzRpKTiBQWd/
HY9sSCeO4bEIbzfH1V+L9BjEy5RDZxUdtBUjzTjreZbfvjDalkH5+E85awcCHNpRBUNVahJ6p6/N
vQmWkKeGmeK0yNiZKPY3GF4R6EHI5GPWT6iCXtzLGthoiLem7PTXWQoaMEKqDclaODc0iNMtwtHT
1qX1gzTgwee9SUN9OYYv34WJW6JAA1kpfzIA9MYhFBvMqpB0ui3s4uAknRoU9JjCIwZd6EuXALxg
3vk4JKT35l6LoIEi5zqCSMVOxaHTX/QLtLZ+WKS8nDdACPxhUkyEuxMB4spL7B3poOu4ehu6Z6if
Z8JUo1M1ouDWoV7xSSprBdKtalukq+FtZ2Z4zdkpX+lNgJ42cyj0apNMva91Dftl9kRNtEVQwkUo
ErDXwYPevEFLzgZoF550aFl75aSSRq55JiADar+dNV1SPz5Q7XfqXGDbIY6Iv9DMJRp9dlTOJKst
QeDLat3LCUHJHcJS9dEgxgVZ2K75DDKV3GfXRHpUY9mp6tRVs+Wk1edQxeQBZ47VMxtmVe1Pm1o2
IRL5GCuD1nNuSBis/NoLBjY/MXttfoY4oNgWqA7s4H5JMACBZf0uGaFAiHpQrJzefXX17vxt8/Od
U2NeIi90nqSQ0NaIpDFvmJY6Whz0BWBKisackL46U4fG4m9c5fMkOtiZrO37lprBqajGSgnKRqLy
rzK49XXK45aF2RcPwOUy0sejJZWD3KHBMjm3A0HG5s8f1l/dyBbbB4TsIiCfTO7hkA1IcXEzrzoF
gv7eJ+ky6XiDdiUFajo0kb1e15B0K5aaXAdkGunOJFdDdYal3iNi18fwlMisZSPF9LRUcdlpgi/j
nWGwqgH/0ulSLfqnJeBxswPero7HtPlug4gZmoZn7QbJyN4b45s3yP4WBV0bpv/gyz7x7PRE6zTi
hsVhr7jyb7ItxhU70h4gfSMXB6lr52bpVmDJ5xsBsPDEoL7MDCk0GmZIULQL1NOGeXZ1jvlbn/J1
m/15RupVc7WOTx5Ds95OWqgRbgLofc+kux7TBntc6Rf60C4PJV3PXCKqQW9JWkhxXqvcCa0homJQ
u5WjJsvWe3v39zcMMHkdvrxiI1NwnyUvaKPXlQK2oYJDoi7U9ZrImIoja0wT3ljPAdTsZp5SJ12s
jXnXTIxux7hOc3d/VIkgqxJnWmXoCo6vHRB4xEVd2rpSr6kD8kfAB8O+3ebOguI7VRwyglJDNziS
Vp+x+b7dtq7A8qb49cxzeYjPfVANsO73qp+fY7HZlQPaiod3f4qM40+68fjQp20wDTXv4KAeTvF5
wKnRT9MAtC7HR0ZX+v5f8oly/Fxraqk1Isz68kB+zRtuWvn3l4fzQOq+Jx7M3rd+vAa4ehM5zvwv
5FzAf37yQ3lQxjxB3hDhz4zqZi52dUtx02EVurbrToQs8xTjStWF9a/K3qYTUENTxz8sr5T5B+Sx
RqiIopXnU7Is9qwErd2Y1LPQ06kNf3xl4BTqpJ376FVGgCf/U/ugy9HYg47JuQXkcB3k5e+09WZg
+k7Te/jWidyA5ZtFEtin2i3G4RjYam2wcKmRyIILmi5Bagn0301sJ5KM6cy6NCI8OduXlzd4OaKL
rVPATYS60Hw7ZfK5IZPYPO/oy+uEpZfDsVzUev6ZrEor0GBvoK01LP7IGx2XtLSNEzM/rJXU8x1x
Mc+zjpkdZa8WIg6Wp+owvcQuZTk6ZuuM11RYruqNpbRD3BFYK3xEQnoc8nENSwLf6NFlzeUcYRbV
p4Ofxj9XqM+JMDSQk/Pf83YQlXknsCBB6UdX5CnpEUOitXUqSPk+hg/10BR6ofVhJCt8tZT7dvNG
7sFvM41i2D859yGyixB71jCAHFxHxomtl7ZBJT6ZjhVG70RtlEoc8RU+8tCyQT3agivV9gAuL3mQ
ZmGMmi0vgWKF7KaafRu56LYR5mvWWyNQpdP5FH1sJTv1TH8NBXFhUj2fWHdRzMCkcOKOVdy7r7pq
nkmk4NaHY84/Fx0eOMe5siEZj6hLEs9n1bo/lRm1fPjJNT4z4MQAM+wLSon/Y3yYuOhbMBnQ4xL1
7GppDUCNz4hOXl/jXuua2gYBOOARlLXVJKiAtIDx12VNBZQ18p5bpO0oPQ7ZqyncSsqptHmfu3Nq
2LiVjGPM9tvnv94Q4IgYztpov5KMzXbxd4Iu8bZ3L1t2O7StU5Ntz0VaSoOk3cgtDcY9RRULzadW
6WaKlDcVFuzzm+YkuiNQwY69tvUEmfwocQPxu4ukCG78tvqCw3SifOsq82tR5XKlcFE14yKAgFBV
vdO2XlU6rTr6rmT4FcbvHxkGv1icAghe2/Qj4jmTJqoiEySTYHd8zKs5uuYK/RH6AngVOWT0tUZ8
mF3VRq7AiFzEcvft1mlbcWEghA/uIdlukxdL58vr7qchZ3YdDyM+p91hoQnBLFEqSdGVFgGcLWLw
YUh9r40BD64kAziMiHM2U5B/al31BMfAW867JqnK5/Eh1sAojncEHgBDBnoTs1gm4332Q6lfflFq
DKyrOFkn9Uuzv/JvfWt5a/4zh6yNXHQa+EZYrdtPDIblcKhoFsfybCw2jh2qJF/v/43cA6BYKkUW
Wzp9kDjdN0lFKIX8GumA6D9maKWf1btWf6Tbf3SinhdS7Yil3VYPF63yP2VGwlXdiqPUDHndCLQI
IZ3/Ac1a83YBuM8ahOOkYLshIWwSopOFrgXD4A6N7Z0ug8nZLsRiYsoP+7Izdm+aPUqIbDmh3ZKl
jnZsJuAUH8pGIKeIycDslJtykRoKuKuljtwq3iyQBRaKQhUCyrsIb4kabsK9BexVmiWZIUVDq3ty
z14gYSPs8GuOljwTmuc/KA5STevS0tyuTpznKl/4UlUAlYnrJUO1IFp7x9tsqR5QzD98DwckliKp
3bL7S/qHHvMiYKEatI+nkiG795K4ZQ9ic2tmo6Gz91cwF9wFBcMm7aZ/TOLiCEmodre4KDLzkJK/
Byd8DoZTivtp6Q9qLYMCC9Aen1v7FW38RF9uFac4o83tLYZ6DEX4QlW5EXQzzW2C2ahISf1kWW2r
svhfD2WVzEA9+14EuAWl1n56Kot86ExQRZ0+o6ju9va5mJhTMF2+4yz5cbDnu53iLdEw+P1pjff/
jltokXIYrtlNdDA050WqJ25o5QJDdd7fOO+NN+R4y1kvZMauJTUTAU6YC4WRXEI7W5uBaBxDfapZ
ez4BbIWZ+1hU0R4pw/z5qPMDKh+/nOvfaYwgrHBBkvwr4wvhUIiawioEY6o8CZe/rKMtV09B5W8g
lqz9iosT0CQNNl7hBcERYQtC2Bv+1nBZJV8/54kYfgMhvmdvUuhdDdW8NOo5cXk1V4ruNdU960IL
lUMEczHCFWTB8cqW8tw9Qkf5c2V6rLQtBqaVWPvIhrUFB41lm+eDYxq00a/oNRBvWsfAfAa5ojdd
RC8jRWIEG5sTpN9husU1jLSEhXF5tFu4CwwH2dgCBLq+VzJPmoYpXH66sARkoA+d+xZGXZzQLbvr
pz85p0gkyWhxxJMTxQZYEoe/gLkrPc5DILs/ldwZEnZJszJb1fav8BkKejrl+C3K1vUUXUFRlOot
nBZ++Q3ddomiydtdiF+7YB2eU3Asc4nHCJmjCRlCB9n4BHfexcGJqT9iXN4DwSWFa0C14Z6Q8+oI
SgGKK9U/sEojsEMemX/u627M+NCSHyU1wHLGK/hM7ZrVHmvDruCJ2msnvQGCLhx4dAQc70v3orLB
+cgHigI6JhV6XPUcLJu8mwtLvt3VkHnaaBAhWwVw58WqpCIxjo4KawpYKytxRB3fsHP5+AF9tM4/
rILfGFbl8UtKxqOMDSl+DbxGe5lkAmp2nkeMzxSKUx9GzkshLGWqa3BowpYSi/9uaOBUmhGq6KJy
ucUdJscgxid9jIP56/Z6xukkobMwNBn87IyVcZyd4WTCAVtaaK3MlItsWOyrelCukuNgA1JzNeab
Gs/8NfhRwxGwCPmbmG8Mc9xXxEW0Xz8WlUkGvClh5ZnZPvPsUP4BwpGlwsOC2m6zx+u8371qqtRN
mR4UuIgllDblUXs7FpcZ7yKvfWUSZSwfovlMZcPy2hjaj58EW28mx07SoM6sDuxpj0KSxUT31ivJ
0Znghxmfb4MPLB+YVBmd9rNIiQgYsw95gNuPJxlbyda+QRPBXX3wvgfPfTQuX9BLvEsEAQBpgI1Y
alcr9NDOAB/DBE4M0qZk2SB6t6PM33Z9sSBaxxwXxYi1Fo9P9042bv73p5Cn52l4alKxh2wtWnMc
Hml0HJRximLQJ/A6OA14utfUAfkrErrNeyK7MZbiKdzk7cYbKNxmwtaEnenVTcnejAnCbYDMI6Yc
szJk9vUk6766wctc8XRJcCSYbCJ9azNzDxxjlMjidOkh9/AbWnRzIqgkvlogjBuDjqQnePV4ZCz0
pvE8C01ZsHirRR5TOTgYAPShEEPkOSNW7NbowFXQIMxqLu90yIBROz2WigyCpGxnnkjIqwoVo0ca
YKP39+HZti/hXHO6Wly2bfAiI1tNiUnnKYPVMVjD3d3TSs5M9AKqLV4CVkCWgh9vlZ7TuG1KyceJ
UvFne7wWGOmoQVndptn/y+tGH5Z8pKwJDt6NyNgX494uSLNsqh+MAkUIOHCEhkbFJChiorTorIny
RHcrGOPdgLFPVJg/c2a4BwxKkvsUZEipKYQwa1YGHJAv0hPl4OrnTolgxXzyr+492rfFUGolY0MT
+vAdeEr8ZJwXv9Cy/Q9r9iytIEwA7Pvu18hbnu0tXOHyQ7YIAEMq1MbU3s595I1lMC8rYz/cuDje
l33r7S9h1tOooz7oXvKf2doOWWeqCwOuaCo8QlC7KMwOHo7WZpFfWqwE7svpF2gSlhBGVME4y0vF
z0xIyWrMaWtRzisEWTH+C7JEFNGvCPJG+fmUNbU9VIoi/2EDhjw21rR/4oiQV+VmJLYmAwvqYqa4
DSp3VwvYDCnGJpTUASuVzNVlwbdPzLmCqmhZD9fxw4S5IX90gkQO8cX0PfSBNsSFRdI8NgfvXgDS
43XMVlZzz0x32by6/s3Ovf2j99ZwQtCzv7C/ys0jLwgSKmyhcvpROMMeIngV6sFSvW1y2DhJcAZC
Dhizs5JZZVokjfTwIgYHusKlBYAus2USY6SuY35liENqR7EwIAQ7/9+3sv7KGVZ+l6MsbpT9Al2S
p8c5ubOqocBvtv7doLOQPRgEqDZWK3E+/tXf/sGYBnbepwBvG4bRKEkDyPuqknzi9vVDI9H0s6B8
saRIGMH1+QnLWUyxaLwKnQo7kZjCFqYzlflfKSgGzq1YZm95YW4Yh/YNihceje7J/xYMF29IXhHo
Y1LiM9WHrie96QXlvRvh4bVhcGtdKKzrXx+0Sx+mG09L4jPFL7q30NM+fxQI9cPDlk63t8pvOqba
7um1/5665+jlwGaP3w7y492fvcPwksTWJ+piLJTqqxp0tYyQXyYDUgRZF45bA8EMKJIA6E3NcBYF
gdGWPTHbbfcNEpRXaiVFl7sJKzt7gM1MlwtAsjBvmnc/Zfv6zMfnM/55pHL5BaCJZGkRj0VFU1Zx
+0rmwfUIcSNI4lW08IFlQ905sGMgqxXkTR9bl7Vbcng43Y+0b20TQA5ceCJVA3uRfbJh84tIXkXQ
o8GAC7cb4Rf2o0UtFabeqOim78bLBCFE2tQZ/D3OjnNB0pnNgWFdDFRlGf25Fpp5EjDaLfqgKAlv
X7Vk2bMevR2dkyINPREhmiFFvq5t+zit2dpUlp6G+rnMplcn2g0G1ErIPNJRALHlwF8xTt9MhpgO
cFZO6CpAuH3d++ZRhgLjMeHTAREJ/OJNshNc4r/vQdvRH0ujBotDS/lq930r9X2m7razkGztGqS5
4vSZyYZC2xsG8WT0oiSh4sE6aHWCEyFuj1F/wJF//40a7oFpJ8R4D6oFkKs6tK72KYHiomnBJBQa
J+zrsHQs+8lBornSl/CQsK9OD6g1NhYVzwLLlPTZr6dFhyxdOL+ARA6mAAnGe4puevm2zEFR4aa5
Dnm6svRQ20vfKCUEfLRnk0rH/zfqOh8PKXP/cgFTtj3QcU5j0yFgPmjriLaFji8Ub8RbDGckQzcl
qBWoc7sx2RJHsFyDDioIiWNRIBUWiky6zCGrGmSaWcgevI5fSHLGCWs7e7XmHqDSu2Jj6XOQoCbE
HgJrJSizruxkZ4m46CZR3B5hONMSP6dnEM3f9WjinWHOdb8RCjPWRRxFMdXqobDSScytui2MKoST
BuSK7Fztkk5LquhJWB0+Ex14+X0Gi8AsAOvPyqNUsLXY6jyVvIhpq+G9Sr4JjXL8WaGd2iKbtFzS
EBgYbErEEpY+jdE3IiC7xVJ/BcLaI9JDu8D793YLHtFpRPdfxhoQp7UyUTjhnBCSMDIY1FALY5Xu
JMXLcVo+bqY/nG9LwI8oqr3VdGwQU4P2CueqI+sW/uEASFm5p1gN8TpaQx7ElVyeZi5XzJG0lP9z
s8hzeAhuNWxCTtXfrrqkGhf87/Kc2IqUQQFCkWfA2KzJq+yMQWuraYcjKRmRW+LMe9KhlTBEnW2c
T0mAaH16LC9aKVP+cujEYn7NhD5e9nj8lRx8am/wn1kaKEfZ73+2yZn0sAek9TyuGh/nsfu7bMIC
ZEtQsNgIqQD5b9GhdAKVybgEPsqSifiTfFvu2KvKnVnG3UW0SBsXmCYaZy2pyfQaWziCajBf/sTA
YbO3zsUjlKH26ZSQFEJarLvqH9hfeHb+uC9hqS6n4m8yZwZ/yUjoJq5sjGVysK1pVcO0IayaPVbo
88iQdGGNZBhZqteTmNvUZk17lv4Z6N/JI8MmgM9a0hkhqQd0p6QhALeGpZCTQuLSPRgqPR08XHba
VXGrcSjsla8B9DbnlSorQZ2IvYDMPg8WdOOBD7b8VlivpXL0me3n1bnypQlI48wizztO4rUmfV82
PkrhvDuPUL8wtgFPTWFKU8mQ0oSQzY+p1ye7QBccaL2kDQewcIHY9UhOMFDmVUSfOkBmHh3Om98J
mR2N97hbW+6i27kaWO7TbE6g8Zasp8S8pwKbN0ZAtmDtVigYbcvQqoa+T+v6r3Cct+a3d8eA3gkf
Ckm8CyItX1gWhGVCEEg/27S5SFvWV66zxrxRl9MVpi9UBQzVd0XvESlE1ERyUwrw/1UFwuXhfeZs
9LFbZXDZdTzENmNLaLgWQAc7/sslLYHyfb5G1aSEKyTIUHIpyJfBoo/uPYtFILSso2J12n8RgyWQ
P82wUz2xoLgAchJrynZHWC5uw9TfOWtkAK+LktnhH7UaHgokVRe/b6I8bmRNCxMSfX/CYcbLZKI7
AjRLXuceBV23WhgafhbHYdRxhCVc94giu7MG0903i2Nf382KXulRZqSHdFWFlNn/r2jpcDBBprwF
XJtZNQVtX2CqNHRsPJCmh0JXrPZR0UesmMwwJAOtZEYb6+Paxdjl6MEMDFsY2SjlaCBgQeKvnuMs
YXL2UcGzRAS8rg+BBPjnyxFrxOjueZzzyrfYP2w3a8CfKLrY7hRxxUaoZlRG/fF3VJQbrrTQhiUD
7cNgVjGtmnRPB06aMgHINaF0ypFvesn/MpffcXBOiAVJ2GMaUHxO05I25TT3xBxNL1NehXgpsTvK
qHWAShtf4D9kAXZKHwKuISoIaqyAtO8csQTgqtd9BbknmFN1r1Swrm2rLUP333c8S0QImLreTXtN
UHs6j3xgA2H2wJQjAWh5xMVCgrn9LgxuhXnQoCs+U+ONKcpodonOYvtJgCu+SyuWi+2UTQnHsi1e
uCRqkUoigbeza/rSiP1Ccs2PtglFUeGLiqDNJhItqlwrP+lk2HxNxW0ujUBd4XdSrDMQ630OFRYG
ht3ynJC4DSFFOxalW2o2PMr6x32qpFIQNZZ6PC2gWTT/TmZZ4TKEfVKASCYF0VX2dH7Jlyhfu3sy
DyrlPEBnBj1TGyovTnj/nG4/j/dX9p8AC/x4yFZJqqhB1qmMn3Vv3KU/lroHHAhrHWhBo63WT49m
SaXaLtdEjwQ4fvIxff9R1Tn1aFr9N1YEr5nW03+9aHeVk0QXWrF78LILlFfEQ6ay68Y2PCHfjfc2
deL4pjPMp+VRovko2FIV8KcdGRe2un2k+F2NsSfBLDQigCYlnnZptIYha/DyRbNsgxppJtulDwpz
bgxkj8QChI6n4Ih0CTkqz8ouLEwHR/jUTutLasPgwXQNvicCSRUAlse7pA5lpmpED9cqRi5yjjF4
Kj8LxQF4l+fL1hjX0BPiOmMv2NiGDIBJxdhGnvwcJx0N5MLbcmZSQZMh9sIZfpTC6J4HH+1Onsen
qrPc/bhsELGd/9U+IYv9nHB5lUnCejZfEbZBf9M39hCPVhKIFbvKoXar9k3T/ErL9lXCoh7Sz5vw
mucfYmqkvxSnrtPuiaZ9JUyryn+GldpsN/bCRXcyyN3UCEsmT+rSj34K/WIgK9UV81aBystwfrQN
6VdX+noJn3PJIH7CF6gjwuc90NeUXKIzpm0+Ql1frSff8nBcuLBdp9p2cZeH1erls6l/2lYktsJn
/Yl7c2OGaG/q+ag7H9SLnaifzKEq34fLXp+XaQms10NuPGZMYql2DqbhC9gwPqWQbI2bqkIAMkuH
VD6LCHY+CFkf9SdP4ML8K1Xzm8Vwcaw8Yx6ga9EXNcrn7suwhkevNVDt6r4QnX7J+j3qlvHXSTi/
j/qXsPPJJzsKhCiBoGoDI6RJWUmgmdIoOO1W6xg+YGHvKU/MfmT2imhKuNTh6Bg0RuOY1pYbVXqR
26r3eC11Tk+HpDTRac75S8LCs0oJda+zZzfCQBZ/Yzassa/b4i0m3XHe/6Nsc7hIGWAM1VTEB25D
nhP0w4N7Dz3tNDTno5DgYlNwtGwJ1cuWnQ/vi95UM3Cbvc/z1SXNp3r0uXZ9Q71+gKDMmHVdVEsr
lXc4lnyUBD84KBPswbOQhFlJYvkU6mL6Lyj39toW5UDL4o3GTJ1pRa2Q6S8Fo/zFJuiB1Jn6CtFp
mnJ5mPWZRh+Oyzyrl7RLibHa5fS/Oac/Xt775WYTl30+Xc4/sqbufiWN42jI2mYopr4TWimoBzyY
jwM2rnnkObHr1y3FR/oUQpgU6MdmRVDVxmpfnRdFUzXQi6pUgSheKiiIchxzsWNnK+hH5tRel5BY
UtfoOs+yztn2HGh/WeyNnf8Ng1KAk5LzEZknZAuijPRhWbPXWbWWTieh7P2efzHORJ5r/pjQMw4W
mYhR2hi3q1N2/3z51QMCwG/HfWbkDm7KKMetU+lNgvd5kjYWM0WF3zc7Q4wfbtRsoo3t7l49poIT
G9BnWVHe0fA/W9+Yro3htJhmlxFdU1OaeeKFYCL+KpE8qoBmoB/ILZdVsXzFsK1PcZvpYq707Qnp
FSI3ySHW9h7KgjBtJ/7H+/pRZToOJxmG4SDHLvkSr20sDEsL8IE47LqIjc+hu2eqKJn0le3PJEgT
VlL/nzCfpXKnx07bJHDJ1WHP72koznir3nEpeM043TujYziCkk4XYtquq8Ufr3m8kQ/uu2Gf79U0
4xAj6BOkJ6PHtqVXaTSCf0cpwVSxqxlRfMID7AYBlYANMQVv2H844gluAVL6GEdXBDPTt1NbCZM4
YtfivinEQsNRWrb/f/gIkDkW8+n9ckG3QsDsObd8wKv7KUUiYIiXaNPeDSBjNU0mwem+3aJopmc9
o7RifMLk3kRTqM2JWnjC5iQEvg/KtsGAMZUdWAmktex4wPKakpcP7JwgfKW7Bi/XsvDPtawKLdge
HhsWJTpR9peUBM72JdLz/ucOSQIEzlNVR9VubvloeLeGxpDZc8MTK6+v6PPwQNRwzaU+C2OTZg2Q
O9oJnArpQiMPBW3wk+iVRqwM7+HuVWfJJNywqAOzq5z2c3oWAdHRgH4/gfN9W6jBm3Ym0r2mDywp
a1xyv3/FGZeu1GZynRxSvLKT9MYvZXAqiBKFRDWZFDkExdLfL2XYIoAz7u80uJENkiil2FZohE/V
Co23ptQO8oKI4l+ZJ2hbIyg8TL3UHdeML638NCo5J3szoEwnv923hg3wJppvtHVJlgvAUvbIPzMc
b4Yy6Cvfjb5VrJNAEu/CQyi02Mgi0/UVh4Usrfhgo4/Haj/Uz/MvAgJ9aEm9g1c28YkgxHHJeSgv
czwBLxdiTR77e1EyXMYC0SIO1F8eZEGm474Mpiq9ncCKkjGMalwUWLTyYkZh3okR82u4ltZrERSj
g8ysLAYoC+sxg58SueTFC/FIrc5gFLfmc6sU429efVP6dsVK33iQsFI+LDc49LMNwvWU/gBFEwBY
Iplldz/KkSt8gVbjm0sbGQahU2Gvlhc80op6DE/tZxhbg9cCjlQZV0vvY8kXJDeGc9+3t8V4DJtg
jvQYyXmdduC/Ir4jePVdeMkr8kjNmRZ/qqu5kCQ3wsQ++KRPiu/4lGvdnytrRDX+QTNoFZYs8Mal
7UsB+4X4dz34zLR/jFxbtIW2gXZww+HxZJ/+2FjTR/L5YXTh67FtMNYkDHd8NfTqnh0ZV6JIMjgM
fUzqOC0GPFUpFMOM0l6Er2xk0DON9XAtlaOPUic7te9TW8fMj7nAIHSqVzNfiPzkqwjl5uTUd9m2
iKFQUBEd1DAuI3euGkkEgC5t14/eH/gzy0Y6rMMVSZJCNSgy64Ul9KjylpWnbzmFKX9ue4j/UfEu
gC72TH7HvDO8TdI3hCiKroZ212q1Jw6xF58rBq4T1MChdu8Ob8qIAkFsS2UIHSmK+6utnzlozFHl
pgcMCc/mjW8bD1xj90fRX4kOKobLUHNP4NkI6rM5dT3USV//VuhewMJaXKv38e/2eq+YveXgrZ8o
YeHpDhSOHILpJ/4naxeg49Jaqha45D+UIvgn22jvp67zSiZvPYxo+EXnTR7tscRuEzUeq8AWXPaz
4LIhiJ9zdaibIguuFLOKL5y/8U+eY/8LPnkxCwnpMq0NxAc5sC9arTxnsAqGELv7vlCr85yOEEZg
RKUG0P7yxK4FOfY2Ge3wfbNJHRHOkosPgvfZ2IoxO+GHxvoXtAJtVOw7DAfsJwiWml+D8vAPY3Pw
80V1vKjcg/1RGXCDJS6g/SPt2D2JXuT6OUX4AtvH6nEOhvvEwivgGv3HaiyVzRFybuP9TOcyp2pO
hXmo/cNwB8c69cidJw5gdFAwT41gxjuKVOGJO1WS6YyHvn2BeTQh6lBxn0Dm+5UdOzaXocGGbkJs
mh+csFQ8bTmNxkMsrJfN6dTCuzrI3ifQ8KlM0KrR84Bi4O9VYyV77eS2u1/f63nUbrwYqMLd0UYP
9F0JyNlveDkMFCRPYGTHjfD9ZbWhni5MmEUE3v5bHf4D8Zw1sjALfXLW3suraWJxjchnRLxqZ1WF
TdwWqF+1qvYROgSud/X25S0G9O4z1OylVAbUmtrV8r0sDYycgTLVoh4LsBnmSec7HjapI5k2BK40
5ZYDRVtS4Kn+BL602AAMhxphFFyB5q8vzxhDWs7753Ui5AeX3bdj4Fg5gGld08IzlYlksNR+kg6K
KQFBYvTxF32ANLnajYkCmHF9j/wua5vvpdo7IOFMxKKIwQVop6kPTnjK6W8ncy9KVxfc2dNbMFvG
bhxKubV4XDUjjyVG+hsoF6dES6cqr4hZfL5G+YCJ+RPcbRZBSbFXg6xkxrS9G52Pe5/VaeQ44Bv1
zUREBGqNYO7GcbbxMagroYpFWl5z8lCI0Hra67t/02qguWfDOJ6wDnOW0OAlXTOHP2w8o5bQpFQd
14G/9D/rebYyROuRtl5a0eLzmkStko9kOOT1HAboQPRAXs/ofvY5F/evqyOrVOyFd2eS8Ji6K4C8
6K7gSt5F4mGwzv+YwYony5cbd5lAi0fSs1AemhaOHErwEdgy2Xhv81aXtlzopsq3sfCAF13IfuPL
TqaRVCmI2ItlXtv42F3sldqMwc/Lfz/bD7J2r4x2jV6zyb0cSJx5iqflJ2/7VMbrWc0N1hqHIy5N
6R+aY430CrRNZp/oY3iQjHbUtUf1aHFih3SkJTeu8j4Fy/Bcu+Igni2trJ+bMgHr5avHoHNhfgmS
v+5etr2yufCTJMPJPTp7yLCN366Ai/qiOYPioE3DPUnz2MrkgTbyvX9y3U35QjBMfsXdYb9eGMDG
8r/Dqr54G4r6azcKdisUOHl72fLxxmlFaqxKKH+p7E/SoHs+l2BLEr773+Q6uBXpvhBg9eJRkBFq
uT6EqXaxH9001wtYvhIr89bQNQrspRcD3dSIzKHmdY6jR7peAKcrwsjhnlVn2z9bajKpr6liHPI2
XN8KIIIJKVWFlQvWBDgGq/oVG9FxvTUuffSYzvthG3gJm6KcNkvORj9APiqgLHA5znaTAaG3gtm9
FFpuyHNdiNu5+siMHxI3UxW6wX0AFztj1afGVIwhBvA4gLTh/QMCTg5WUlddd+/tfbWajgLpuSnh
1HU4CQQa5rMgjlrq4UCJ4i5XdhE38zmlqQCxEEugxm5ytDUd17iHT00dLo5PD4Ib18xJTQYZa2WO
n6Ry+gNCXH1t2sStnEGB0kNTK+fGT1WamMWIrazHqy84bMwGashmv+F4hcmnDLk9dSlXzlLXM8GH
C9f2eYRQQ66ahnvIHQBhdROiut82zfMbx4zh9HF4JmQNABJOXJQzirlEThcUKBQNRZ9gzdkvLiBx
iQ6/1XFdcaeEDw6knDVdHS37frpnrgDcaZm0AAWWVkRn5M1T9UXny4u4pvM1scxbtjEKvYvpUT8f
Lxnei45vksFCpM98P573FsuJp50WPAux7g7q55jkWecIPShFUxDJTncspuG1RGWAxJ4oousGcn9c
DjRsNOjVDaRe0K+pwpmI5ymezKU0o95sp1JxNeO7agYcn9XMtBR1+mo8nfvzCyTG2rKoT4dOfOHf
dbJX8YQ/N6Sl2NekTwq/aR994V9RuDkE7/Q4QAuSC8sxb28hL5e+bcikZ4rF2uaRXeYWWVvBXqU2
3jbybjEJBigJ/UyxwJuPfrU/9HX1ZYamIqj1bUfoHXv+bCWr+6LVOcfD7EiMgA7Qu6kQAqSYMK/a
INKR/Rg1EUH2slakK81C257pNjz2xFjRqzzWLXqq7L68Owga2nxHyPNOHMfq9H3CLdUj2aQwYhgD
++htYQ7sl9DCYJBYC479fKkdyxqz1+Spo9ew1njrXquRxqX4fCYxQbzDh+Tnc8NmqAAZ5FAT2mf1
Z9+Th4DebICD8ZaF8Qz3wmAJCB29/q7dE5XyfCroZ8g7oBG7TQH6LnKqAhG1OWK8uYd2zyVvyzUo
0Zg2pf18RUSnn0El5rsb3uFrIs3lmUpyZnpT2uBOL/6XnZQ641NJ5j4+gne3wUDNwbEN8G+FE4rg
A8jm7lGZ2loIWZIT81YjgdyBzZov3MvomtlRg0twDZbtQO+baIl4nB/LfT9j6h9XQ2TlOH6l68pm
mVjH9H2qtCAAGsXpylZgVX2cMikqZnXd3xkp1qPJ2nIN0NO8zhi5xZXrfSjjPf6kGtaS/02hfSch
oq8B7d29D8iWQfRZgmcKXuGpzS615rhrOkoLWwEiUG6wz0qcASdmrHOo7AWrn4wFtVebTmsQsxN7
8zntnkxilylVc+rjuyisv0+wao6T0R40DtDfeDQDefczpGHqmpr/mpgliUTNV0/E67ePukFDZpFi
Awl0gS/5dLXSYomRcO5LbkHLfUYhmX5BgbwUWfas0Q2VA6A3bxcJvtOX6k50P1h++4R1fagy7BEC
J3dVLj6u5Gjy9osKoYZcm2NuMEuGxlD1XIod8mDeBpWkOzlcxynyKM2xh0a7qr3LOS1we5GexejP
naDUET7uF6U2qfZrezWOBv5Wcp/eigvySMcVCF7LhsTF9EhSp/ykidh0CqwiNyejCqHtyOE7TLZ8
r0ubCe4YaINXUIM8luIVqd8pOxJyCWBSMPqVfw0/nIJrZKXkjhTgjvWGMyDkujCWNt9tIvGvftYz
R0TtTSIHcp0ugbWGp5oPDWmpNcjF11n8YRIpWiew190AVADaTW1APWD9Fj1KevACpeuZn6BFRWV4
s33PpVUtqOeT87HRJWCXhKGAZ4wngTOuNx2v6hzgUzU3GvqGGRqOZDFAcHKcfk/4evat4fW0Yu9n
OdcmPKgwC5jjRyLQgKNURcYUA3kTmvxXJ/a7nW60/JtZBZmhhhP1rzpxKbsttX5tUZ8DsDfLa7wl
MbO9cg4y8HIw1UiC9/EopfhMPxAINg300Hd2G8FfM4ktCXZUHiEcLfr1uU0GElNTsuNCnJMlooSY
PvYYx+7fgK6XLF4v6wQ4eNShKXXiTJqyUCH/s+c2OP8wdGSGrbq59L8Va8djIBJ7bwuvS7Q8Ywce
cjL1HTD4Q3eD1mqX/8fbA22zZT/Bp6dSsZ8yFkdD98XQToh4bW8SC6q3KbEARTMbt39jWpKyds8x
TQkDFC63CY+RLNsLFg4wGoQnaS6CKFJjVqubAOKZEHvBLXV5YgDuBoYBg1vXqeRV9J0P1INiZe/l
AqA5iZQY+ajHyAsZFGK2y9fF8zW6LrFw/f+yzk4hYLpNKKTzCrtrJ0cQbnV4k1iOvbHWgG0qTD6p
ktESpwfj0IPxMNHv+1xOnRHcv9RaIP+48e2f2dWQxk5iRe9dehHwffFttNU0L27WIoGSWbd6Cgg0
SlIqFVI3YJNNsRHUACVoySy77ptrJxQg5T8E1JtdcrP+274eWo+q5PV0Xs9ErCaMKEh4Awen/Imo
NN3OigZAuZsAC7r5kBPQXRbRvP3PBk8ACJuzCu7cInBHnT+CPLQ86UFMqhr4+C74EYHGbOtxX9O7
RqoMv6HKPQbJwp3S7tSFCPsuiNxugJOEBaqEnnr0tqSaAkFAogu0FCQHILjZsDZsn0gzY+jDzTpV
BincYfrZ9qGGikW2mjMrZju0NVqTOv4Tveo/Q23hW1cM5O2FtQEbKlTT6Pua4EIDXJLMdLu0jb8V
igRkSF47MYIRKo1teDqhs1tHF/IrMXCgCZLNj/eUVr5xyVK98GWyM4mfycjicEU5o+4ZTNpR5KZ3
2H8R6qNE3JRKsykNYr3TI7MnDCgBMEsXC6iBumpQLXgkmNW8FjpshtVxATdXhh6CZLwVinIbhGmZ
Lr5l64tjrRC5YzejEwh63WdQ088l4R2icFtXRla90UYgJ+8hHKcjtZ1j/Dpyzw9bkAa07emEb6ac
2qqrqvnhqjZzxh3/5YUcVUO49CSJoIMcNa8Tu9u3NP88o1ELgNdDs4NZj6Fx7wCrqfsgcR5e9T99
UQx61NH/Bqy8ZJauhiqrmZfqY5RwuUeaRUth6LBRrNSx4iv7MgaDjA7JgM3q6L/JDlJzXBrJRdSA
GyMM0lqaM1f4JToMz9RyR8GrgE6kds+TZJiFX/4dD/dHRsQaIcEdx4C+mOvlLUfgonmU2ycbWXQM
Kj/VAh4a7GMizPfT1jMKjY716IhPcxHsze/kIbtYpC/wPBNDCxuPrzER3bzGRvnGV6g4lbiAvgD4
M2VaGyZS7SLeCRcLMIxNrs7bKecg2M4y1cSIcuToc6eYA4tE24fCwV+dcCOn9c4qJYK1Q98ezUEu
tbvS5v2zvpIJj5Wou/Fp4YuMbtWeiZx0CIP0DoC+kXwl3a1EHWpbXidA0wf9PkxBf5CQeOXOnEni
R/Vmp1hDlccqAHJHKfgmi9GkWhgn1RA/hadXEweW5JG/F6musIrZOGHQU6i5C1GJtrBqnrSBuDUo
pcFX34i4NcDxoOow+WL939KMZ21GfIFdbqaESttkadhJV27hhjSPVrDDrhiwH3LW0UlfSWal8+hV
q4VP339T1+nmhiXLmxs3FkhrXzishUCzvmkw9opKjct0jcM4tgilUr2KSoG6A7FmkhBDISBlsJgN
rkWfEG18c2HEdMWcI/FM3JKmWT0/3PuRt7utyn0AMFrKUvYd1J7fWMApXrp3PpiEdrm8bbokDuLZ
IAIaoZy7irAZFjHkT96i8Tqy26aOxkymjdWg1PZ5DzIQYduUgrR+GvjRFHFV82RyTuPF/z4SeC5E
e3OHFiUNXtw3DS7aCegatWfzxmwQ22I3PPPRvaHoF851wphadyyViTIo7gf8v9XA0a3TK00JIq16
YkgWuqtjNR8SKw6c0dkXgTqI1EWVnYn0tHQTnXL5ZckLfMpPGztnqrYbLBnAuVNJq+N/vSuNOgNb
FbwqrIu5gSHnuItWrnFO3vgdyuoUj+49B+xxtlv4p/PjAhUxRztHDxSI+odDMdiQrjZCOYf5V9DL
n+ft+0bPfy5vzv39+lKHcJ9taFi6ceem+4C/kBXGr+eD5sxM0LjDkRVCXfosebeKjjQdbRhY8M8M
BXPTwq2kPcjchzgISO4XaOTQsHv9lr+e3kDL7feUaleDGDNwynqPUw32M737RdPSB/RHtrB/AS9P
H4GMXu58dVhn8ENikwiAToP3VrKDH6tEgK06m2hhOsIObVcxF1GDnrlLdaxFl2Ve/ljXG8V4mz+4
fzmU5/rk3y0M21jWwZznlIICemcwkbm/N8fxs0rJIUO1oTwewBbOXAu9ETzgUxcLzn6vYJsKofw0
NQ4iHJgbp2KbXXegAgvIe8mFv5yQZedb4T+c+OS7bvjJnNk1P/hz9Sf1XY9pVTW0z7gtsyyJMNg3
1id0RWZP45t36M18JRyGY52+bnuB/KPaiUrDL4shoi85CuP0FNdhQcsiwJn66QDijSuZny7xAAbs
utKogbTnmioerai9uSuzZKw6edsTBiu1Ef8wmnsfJs0fqNe7IpKevfVse4svSB/Q3zZw3KO2lI87
B0V6Hx/uVDP9cTweVIDlaLthVPmOLtbY9eIPiRXLw0V2qhW7XSK781vGzt+z5dFzTVTnU+bQGH8m
Wmkrzv4s0mF9eG3kpTKqb0OK2fxoH3W9Nse4ZseAoh6/5j1Na6eNqghhHYZO6el2dJPUau1TXrpJ
AGBBQJB7L1y24H+bhA9TPz72kVZav77YlFFvnfe58HrKaRtTn0iozDwwOoeINfGUxwqPlJn51aH4
dymR1rdvklJbmgEuU68Rf8rIKYEG9BZWo7yXBOdZ9Zw7sovErdlpHvndW5ywPJhcg8p9sU1OjIHx
hFPtCKyNWGTatR33MFI72EO4x9g37p0ZDG8bSOV/JZwtL129YwvuifyW9krxxQOjieQ7xfjqh1jO
4HABXm8vjFY9lQ60l/Fm6Sxy4nFBuO7dhbrc0xonKkSOwhqjfzSSnQsyo38fS2eqLCsmbvElghdV
AKl/s/5dMNZxMa722jugmiffO2W6me3mCX6rGhGw1DNyGA9KP5/yu2QUar1icRTrjqOhurTrXkLt
zZ7WsbmkxKiOhVI5yCanhqcvYyiXMxSGlpb0HQmids3kw3Xzdro1cReQbcoZsYolm52OQ6FwxAyx
Wbf+cugkU2u9X3qnJHN7j7/gaqr5MLcNmNuaoIjEWAA/cQOz4jX28yCa5BI122emtW146gOyxgSs
msJ5xRLV6fmC4RrQgQU/fNf9H73eJFdu26GS/+TDjeulGG9RpCR8lY+wuRhgf88DwEsSqUMKf4Ef
tn8ViLYodw9ixljam2Ds9Ghv6lFdj0xu4dAJLYMX8Hb98mHF+K5Lmg86L01h/8ulL/w90qH4Vo/P
yYJTlrBaItcoi1KqfHgSxbf7O6bdu7Pz2BN1szx/kJtpBEOYxgZDI5TRLKl0ZK9+we/YTAUJ9wDT
mrCtnjzDlE7bUZOT1AW+03kPWATVtRN92OYMVMvk6DO60ON+FbOKNBrDXveWfFzsqCMYm34KUkxU
iJBzjbJRK1QWsHm/KxDgTI1cI7aYIVZyX1jrc+XNGhDKJZTLUgfGjUeUaeUHci+zjxauo8pJB/ed
7FIqIfuiiJYS5QfOXqdZdcolpmcjX+Ydl7GCWwW5/yKfzGzAIIJOs24Kp6A+SyC5cfN5nGRsCuZB
nM4InH7ukzQqjeg4mSsftK+mifeUkq+sHe4hJj00tIGiJgiEItYLAOTjOPlg4T39h9IV+uMWThv4
/ymPOPeOb/MSIy9mFQoLXmKLeNs9qkmLifYwXxF3vuwoyVcVl5qej0iE1tflxiszwfW1E/KY4JLa
dGM9iT+IE8r4KD45PB9HuV+doHpTgoIbABl1NF6Rw0YwLW3goNyDCJExiT7yfbSKC6Acxc/2cWup
xwTxINsCLD8GXJ6T4K0Or0SDIiPnwP9g5rLb6cY+Wr5V5b3wetJ85kpAgFt27ud6iNPWmmDtXRPS
tP+51UsLi4fxys7CD93IKVp2e9tNx1EdXevu6eSkK/2MxXNYbm9Th6prmFYD1Zery0OiBNw71yVV
SPK1o5m1vUcMSezOIbvC/r+rm0frSSYfIInBIAOoifDQX3NHxGon5T4DXAvl1zTmPqO23kIPSwfY
jcvPZtkEzheqfcQf+0CmHgMOEly4znamzrf5NVMBbVz9+8cMN7vleInuDGef9iAY2oiFaLRtT1Ex
ByU4JLicxqA5dLDDtPhIygh1x+clKRVaf6n9jUKLuCciUsyCZr8GoiN08p5mANsCsx21bOAlKzFz
nmos7tfSJemCsgVspsgZlRF6migyEydO59U1rGbEXQHr6zAenKCTIH6PKNCpJlg7mdMw1qpxNZcn
hdtMUgFRRLrA8k6G2K5PAkBXZYgHUFwJTaY6R/GndeEv1dHXJVzgbyAqctfLBCEhJAB5ELxyvHru
zG+STRDBYszvWRxyYCI3K38VlaGG5HMrkfIxRPPs6HptMZXnW6BHz65bb9L2re5DHtRXv2h/Eygs
UPwUsPCgGd4mnNOJqtUetAJc+MTut6HVC2UjZ+tvS5CUQ/0kWETXPwNtwnLnHyY30A6zR3kv69bK
QzIQTq1Io2YhxpjjGWfyPITDms6kgyhZh+KwwUfgFWGbFmqUR6R/vXGKzp2UAf2O/XE1efH1/ZPj
WfG5wmCC2WMtdTbhGraiY+0DiTUhFkwA/ZG6MiTQknSErzOgBaBJ8W9WpwfxUl698Lm0QBLyyLMe
WDVLj++XY7zuW2oUV6slDmFIkOtbHEYDTF0ToyhoNW3fQ9Z3CJO9t34ZbEYci4v4XX1pCwHq41nF
J15QfJ48lBYQiCEcUzuapmLFUu70srIQ8h1sA64s8Xl3/IrosRGaqIx7naj2HONk4Q9re4d+7Yb3
atoNwu2YRL6vUWLqaGd3B94djnmleK4+F5lTvxTteT14wX8H7dcxH6c2n2qyCYmluIe2iQOJSUGQ
DHxpT6gkMAyCc6PHShftF95MF00BCSTB6eZPYGH4zRYpibuDr0xKUPCBX6L2E/LYDfIuFktoagCu
ejHnww02ZObEQb1xETdHwuQbsKB1hz34ZltyVN7ljtQfKLpjnfmMi4OxvzNt0LK7cNoyzDrVIU0Y
7YujBAx8nB4pXuOTLLVRmTjlMPkV0X6C7gzTmrzfwaTRt0OXD8BZN8V4NufnFSNINE1juyFlFt0m
oCP/UQXocAn1LMjr8/8tPn0e5ufAnYPGxGRpLsc+Czi5QKEa+rcGdResphQPqFws9QNodm9NSzQz
hQ2Wuw2VBBhQy1BOC0lckFqjhGVW0EcvgMQT/jlVVMIzohSL/HvdvPpm903655t6OWxj0GOX++Ga
PaBPr3LT/nLWnVQK06DFx8StR0buY+0MPfhyShcieHCbDNn9hAEsavqqmH5DPID+rpUe9zZdx4u9
MR/SKl4YvyW1Jy6LDGjvs+kiseFSjKmrVUY/oxrbtfCgBe8aKnrSVlc8kRLqK9v2dqVABswsbxHK
ffWu0jEdBdHymgWL3XYnKLnooe21/AcvKjQU+kDOJcrxT4mIIaYsoy5d30BIk+bkj8NPoVfjN0Yr
65FX15rN8YmIUMbc5ZrCpSsfaq3gYYpE5TjcJt/gz2iK1BM/2Nw4C/ZO9A9t2e2Ut6n5F1WA/dZi
7BisrW9SNxvn28JlV2B6DCpPrWpeJlJR3rcQptOJ+B6By5pG362i7fSohi+t6O3HRUXXbk4cS7cC
d5yLtISClLkgu8Dy3SWdLOy2gYlxSRqNrgoGyvERVerGhvYD51D4P4KJo7dpSRMH8hvF/Rczlde3
/5LOLHdQM2TiYlOUgvEyk6NWaYaOCPVDcwngefrD9G9KQRAmtjfP10BPIQGJIoPPW5IAlUtkwMTa
Zo5F5vCA2apwef0DGzDGveZwAhKszMzGS0qbTDeu90eb1dd+0oThiWtp0mSZdNAgJmlHAKd7gWkp
E26X0AAaeRurwJwEeNnSQaoF4u5kQ3sYGdecpDwAAtnVy6OOo1YH+k1Kg/jm1dZjy9INevVl0X47
fdehFA83LEmUzgieSzjgVQkYCMkf7bvUr3SwniyY82a41q1mA5+o1XPlrrc0a06T1eRDMe7KA4B/
e1C3SvUqJdR9nkSqhf34780C8jWHFfEGsKJqm0JojOer2lCVVhs6md6iA6AnUsC8VlP+pg1714hO
01XccL9UohmO8/k0rFL2aBEuZJbBRT206lCUAXLegssEc6ulU05LRSL1TpLQdhdGE25QLOZx4+r+
FATJu00qU0oNEcxeLNRIAWDoe7hA2k3OMMWraPtWU/h4s1ygf6fIRXvEiNJ2pSTDKHK5YO+0M61X
HP25RJRDMxyCIbRFVaJNSwjDAkZ0Xo3Hh8CAZXJ8+AOBjYi4PXwUq77l3nYaVcVyXhjp8lleY3s8
IA0aJbwgrssI47UuLuyzJKmUVWDhLz2UEqMjN4vBFg9QuOzvrJdIiPB/3Mm4GqZ5KHUU39MFm7Q9
9AxWj5FTwuZJvNWjR94FXtrBmFMkHVroEP+X4iIrqUWcwxGN/xMtP8CEjcViYWNjqIgzbaz7Kh5v
0R9RTG6r1+gRlB1mEjMq3K+6G+m9ahXFIVpUU7WPG2+7XJ4aSYdx2e4IfLwa7Mc4DTWzvorXcxZ+
ZyzU/n1jE5tYzQSQewFyD7MIJ2bGY387BxuOuLGMNYAgwjKFyKS9xTFaj6KaH1s8SlljM0KYREgO
t0tG738StrY3dWzC0SKItuHkhWxJtAm43jNfE4OV8VwWGGlOjrSM/eIg2zuWdK2NpAiyrYsl9A2k
RID+Vvo7sKn3oYcFeX3sQQck/riayJiB0w77bWfYK/hODLX1iHOUf0pCbGveQuR7C8zH+fvAWJnI
wPAqsP+uLIx+iki7RQtOdZ+tgDsH+Xb6jq8JqUTf5rNE0DQfErFeLxv5yQFe8wYJ7S/dfebok8mD
TaDG62KpEeQoGrSdk9HnB+EK/stqvwMG+YEHJUjPvJWyDttAd4kkE9Nn8aCXfFnSUq2p3gn5DBiF
2jli60bi6gEDQMoCmXnleLNNEQCYpz8we/KeQxtsEpmRlm7O0oxNdCwvviVrkXpZKnfACejKyVoC
ueyixYL8byhRzsV909wUdfR+y/ebkKf0PGaD4j9JtHHL0HS+prsrJi73j663+6E5yMyHNPtC/04U
AanJ7XPkgvQTxal2B8Q0+s0V3MoXJVzYxI69t4d5eGqQud/3Fwz2uR7bA7XOXMAM/R/IciW9Hw9P
P3xSkiigZi+X5l5meCKw0MN9a/yLMfNSUzonGTdWM8voKoXmSjYFgi9Fu4L9L9AZBnaTnPOripSI
RuRIl8QDWA2GdWqqSZCIjfZSg+QJsA31nk1GT8awWmBBB7DBEnkvLdRgf5flVCCcE7XRtT9pVJQ2
sTkPRHCzV+f/YqQA/h9W4hRHgwn0zl+5EgtkgHRab+YpLEAA4/EHu1W3MhlEUB/kAdJFfjhdVBLr
rM/HSzmLpD2+ZeZYi5ernbm2LIHemxvEFrUA1smJxG5gw1fq7oSVRk1+cKx1Kz+cmCYNVWSWys5P
erWNKsJWN0vWxwz3B5yLuMrbGtIXegJlULqdh7IJ7FWd7J8D1g8BPtZEKzi4Tu57JdRXe4QyWKe4
bdpHo8OwCQVuUogHrCHAyYMxFf9XD54pf91GL2wQz/v0f0y0SbF96VyYTW3MUTYNBexRxbESJ5pf
9sBrUgpKVsfkwhi7yFs2VKu5a1xWGIeNYJxhuoz9S5uH0YoDS4t49fAqPzLLsVM7uVTsr8VdHFky
10qyp2PHok3veq4T9UE8MRY2rp8g1/V5lrzhhD/bhIH+uc9lNHc4gsJS1ISU1FsBQt0Xk7xCbKvT
hRrErghGUqtxlsjxkJVwc9EJZoUz9+os3VAe1P3FYWn8iqfCqbsI0J1fEbDLh71oD8v3rdZ3UxF8
jW5UyV2syzZR6s4SLjayDze5QO7W0WSJm1PphU1ianht9csdDcjyJCrhRl1GepQjMhqfKzLPL2Aw
TKkOtCngOANqiDswSHhK3mpRbZgPqO/C+We2YsjK5QXBUo8nYEQNWI2xmZI6pBq72LWJgwwHMh0I
i5q/HJtRLh/eofpm+Q5LSHdQnTtRKOtYNyvrjJ2tidlFrWBMf9MCPPqqEsu5gbu0RI3GAYeVHcSs
Bc3CrkPS+hBnhjOJKo2lCe/gZGFMMkAZjAn1x+GmwEjSUQGIzn7MT+EIKHcY6NOEmrnTfVqAuAk0
uTHnLIJzpze20mYwW7Z1uIivrI8UuAgPyUM/brpn1EWxay/YT06jUkDd11S2Uwz8IEWNnDQH/yES
lqDUosVOAQdtwq1tNwpaSJOe8tSsYcEzA7ZuGa3umuMAIcur66nb6fBYDSSBgn5Hl60qI6j1+CSN
A+UG3Zy7UXSMfp6NWdjdIxFxEaTi/DYXlgmyUrX78bpPQQYFqztNdFkkCK8yAbGGddQN7VoIb63o
EwKTDhjHow5XlAi5XQJXq0pkQzddjJfF3oMh48413zDRlKTJ4r+uRz1oCnDJp+hAqNCQ68qATUG6
GIFRPaixhgNINcQZrdL0LpM11ftVtlosXBXRlwy6+hDM/prS7tEBP5deO7Iu/O1nSystUpSwNMdh
V3PJ+Uq03hUvHKfh7pnxdJfxCaJXaWMv/p6lF6eeqJFfZlOtT+HkIVBu0o/Su4fTduRwn0lvVhOi
XptGh6i7DYPuxrZJgSp5jA/3/FNWcPDtZCcASjfpLnXcX270VXVs6NeHtv7iTQabl/hYhsYxPvjO
EKeRYPjxw2Ozufiv1x+S8xG54+NWfPxRxQpMYJwkg1C3zBHlqqrDJzbTDeTg4yT9jr6mcOhAp74+
Ci3pilS3Rub7Pu+dVKo8WjFI0F4EpS5VtGZKHr72Cd77kslUBxK9ROO4YbOTzkiPlznBOyYJEhKw
UQ1TNdpSWNWDcz9G4+qfq8KUIvqDs43hQK0FKlYRrMuEFSXBVIFBxfPdlsjW5I8CyfEPtjfuHlKk
ZmI+HJOFGlZ8vMGfhz1xQHGMcOMJMo91gmG45hp/P8dv48CjyqKJKSEadCezuK5LWMxiVtOjxg5W
XsFOcU33M7yBxCObhIgFNR7lEUFOxMFzBDR9LsJLWbCcaaCaIMb9M3kMWptPFtDY0IAfwy3wFkCt
+VbjymIFPBXHQ9RUPBkjLUQ/VsBj45GU6yxHhXcH+f5KxNk1dVhkujbfpCtYqLQIvNv0v4hzrr4U
97I7XCcv2Q2h2ZZVt9A7ZnLiiR5r/wCwwc5pWCsokfQDYeswnSfYQqIs6zjog1XusNJZLZ7zx6FB
mfuILOs3noFA2fMzx0G6dkry7nYjYYNpQDi3uEEMQxlGhWe3zU/obUjb72AHdRrrBtyQSRs1E0pl
6wC3a7y2rjyZ9NeAfmaOfbIJvrUtBlz0QW/MNhTvrVbzc453D2ylL3gAT2eB8dkIskktQnxUnR2g
I0MIbZhfokwVhg3oOq+M7nc9GQHXdo7Sq0q4RmALX6IG5DM4jH8+trtjMAK1Y8wzv1tAdK0Zpm57
ApZDUMdnzOnMNXClMIKvC6Ef3McQotZWN6GMstqT/5UIsBNft9qPwrmZ9oQlfy1W5Plx1CFqkJRb
BaLOiuartqQxfrtw+191RvLBHblYDEPFuhk5hwzFNGMMxGpwcce/f7ksPtFTiXDn9YVbixrmL5U4
PapQ0ZTEBN/+C2lg+EE0ybOH0M3FUD3L2Yl64j2waQWpXtqYyZD3gBeCaFJap7sEIZBbkBKTeiiF
oD5pA9YDVGzWxvQidHJUPPpi+QJrcNdJ26D9jVFfxtuHk37fnG27R6YVLWOrVW07omTcsEu+nv8j
CU2OHCTqBdBl6VxCIrI+PaiLVqjMU1uAPMLBGpjE9Pggfb7NBeraNdiR7V9aXwNFshQyYYUT0A19
iiL0WwLR74Nz1rscViJ9dm8P0l9x1frtEohkgdGbd5U74oljrzwDJlgLJuHBcY/GPArtVN+h/Ji1
0aY1wRrX0rOO+LPjiYm8iB4LuvechmW83LwAkCUWDi4w5YSqlSZVnhxicwJd5m0bT5vTwP+V6oGe
8XlHK9FVFJT7c5YWRUBlpURJtqI2nqk4ck7Z9yTx56WHYMDLGHXN7ZrD76b/kFH2aICwgaLBD1sQ
WmpF+IlCIs7DaTGoqD3n8ZylgN5mwlakprJZqSkTNYKdQo7hVC8eErmYsV9xHQ18X0+ZGiNWVzG0
i7grFfZr2leGLp45IzqbTgFlqRXu+ncAhLCrI8HWgEF1oFQigWHptg92w1rst7GHcIxH8ZiuK0iX
byAZZJjn7PPvfMcyKpPmo9Fmja2RcuQ9NH/hoNUZoHI1USs9GQ7OJv9071gZiqh2EiZXSR25WFWY
W8sM+o9AoGRYuFgmHfu55E/HWqb9Za72nsAufDRnIpaCsphUfkV/HiYowqRyHJeqfPVVUuK2RG0U
hZfDIvEjxI0p8QEm71jspR5n3fpYK8QyX3pc1riOCZJSH5s9E4cpTSO+fFNlHVgugKcRIjc9lql0
8rNq/Ozy4dJCazuIwWJRl0duOb5ME0NZPeMUb5m1rJ8MJ/ULDjVswtLthp/Zi23db56eDnDZcXC2
ydTv4yTFmRW8PmKqMbBW60joY1f2/wNTbpETWvhpUAjBZFh2bkAEApKLChlhKKkYzHx0mOuhtvsg
qKGPO76l2BWGL9F3ewwUA+ECIPAWJG7HptFYtaE4Umicj9gMpSBIzD+LtglxIPVLfwiSbB36Mg8o
GTk5FrW1J6dw8D3TZUxVNBd7hR8xiKcRFsqWHyncht52zxast3yTNT/QGJiKrK6wvjBOBArvwUEK
LXiKJiSKSOdwbJ/G3pAoTC2zhAINXjTdLSYDTvctDy/g07udWNVD3J+hs7PeDuvC83o4KAFX8/2i
AbZPmIwPcBRq570/FkPixl0l2JjqeaQYMR4yqzcYv9YKAqY5ltypwPHJ+UlrEAtRboDyn7j1TWsq
rTwOr5cvQ5sm7ybL0rXscw6R9M2m53y6aUhAbcXhESaXuzb1e/nacaXK+iBNp/ObpH/60uMqVo06
zCRmBuBnjHGyVvFF5fok1Vzah0KppclnNz2TgA0BBdu7mddPkSZZsN1iGLx/e5yb9F+TOCqI1sCO
s7LI//zPEvZhFemJw8jkqet3Ni03Y1/7a6SlNIw47ByvnABTRrFBlDPxhIHPl0416qTl2sti8pwB
3exLLvHt7A6gxHklQuGsSMideYSUKF/QFstpXmnP5JTXhMVlnJLGkbQxMKk1ldYJOUlMZNy+aSrd
mtbs3G2baJmm36i/8a102UquTsCzCZUKc93pYKpsAnL7RwrLQMcqEndS/eC9DZRgDRr7eRO7AVUy
xU8lDHtDlzFO1VVUGLlB9TkMJNVgZGTOOVXliY0ABZMn6D3yUCR8HuwEA93fRLJOiWfNmZukSejl
r4QAqLWT/+hkzkCKGe9HBmmzeDvPI7nQw13/V+/Cr998NE3fwJRCulPX8D2bOePYVF4Z5y3hIrot
tdvhFRONxtrXhx0MH1HBmrx7R8jBGYJs2gCTinEX3mWdkh1ESGqLJuXE2E0rwEt9KCly1IXz76s3
U71L0SbsqmRmL9p7+weBd7l6NOBeeJJofkH5K+CmI8RCgrOCByAUeVVxiNO6n3lIVzR274fE0zt+
cQclPKL0NoVykGhetkwdSwGdSow7dBSk4gpDCD4KZ6HrasshOtUM4gZkKW3ZMpd39H/KXM9ND9fW
t8/OWPj++MR+Z1iTq5w8NMzfYbt1sHSZy7GhHB5tH1PRV6DlPqhaCfLDXOkaXNDXarCtOVOcPlrm
jSpkXXLeIMqYeVwviieLbZhUDEol9/qv53HI8jMMvPkF5EW0EjHO4ja3QmYn/AV5HKqaa5vT52RH
MqofpQ1TCgCoFIuWyBuKm9AlPWUiN1FNQZHsFBhay8M9EjLncngS6MDrfANevth+ZRT2M8+wXdSe
yndcZwkFmBRJ9K8wXX+SpGG9uquFaj0FvDbHEagxBDtUXG/9Vt48vbI0zosk187Na7w2ary8R+mc
b8Z5QrzYAU1jy5+byzUo/OSmBBzjEzmplpCSwYeGEh2sn5Bu5LyGmHcqpdb/x4s75nwkORe6HbLt
bJSgjsEYcI/l6bXSh9zUXMrI79/a3IiMPJ6kcjnl2gM9AmufdTID8G0L0XHcXCL792WN/yk/NTH5
uilOm94uKgm2gbKdKvv0JuSdDRO1St+ZZv1kWmX4OWSkaVfMQushBVLkzSpFshhnR21uout8siSK
eRfmIWfnRkynhL742X3DgnLi63cqU6vGEnIamQw2bT7BlOBih3PrJV/adFE69b9NYm/pr06uqcHh
K9BMgVI2rsmi0XzmnGYpmVCBrEaPCvtV2k/YzI03MsvZclOkfhTT7CsaJWNuU6ddZummBp3UoPIf
TX2qKYSShbz0y3IKEIqA7YRbCt6ulB2CJpgURjjPhU6HXMXkC0nFWfIfIqGv7csC1oq/fRtDPE36
VtARWOg8b4XkKxYwI1dQB18tDdF9ePt7SlAfwqESxYwbBtpOrB1e3DPm52EDbhCI/TLxd5T3c437
c2NeqZQAbDZV4jztk8RCqzMtoix4R1gH+qeTgVv00Thv2pLE+y9Uw+UrHcROWKYPnDosSkFVic31
J0wWpFeP2f8mftB4v3REp1IykN3j+xPaf7wYBPGdSXov0yjUgQEah7RPl6lIuC3GMStoOM0I1Qki
un0DmcMJ9tmZqYXf/yuGF3sNJFNSmOAaYrh8zEgwwsCpsYXnT2KcYnvZBdkrKK1TsgWgJbFlzzDs
5DZfxOtRnSCZGJ+oA9/AsOMkuXp7zLhbYnSZHKCcWRWIqAykQNZUdFP+3FMTJyUgpF8ApvXjJ81m
/T+lDA2KQ5441LJnQhg+Wgkw33Pc3F6Km8GjRdhE1R2nLmkl9QMmIoYANvrep9k2ck45/bn0Cl4U
xtEr+cn37rBOqGFjczSHdEl/X8KYa1yj75sBOJB48yCeW2590+tdZSX6/32pc5+z1F1HuslG6mC2
heKqdMyggg6lKyNvzJ4oPMvFW8DuqAtiXMYTuvuPxhvaGSi5NAQ89Kl6Mua4M+bF0mGlfl8xl+Om
PmKGFlAjCHcVeJL5Gz8QY67xm0lKfzyuHKfCZsUvMQWKKUy1O7oHI+qN76P+xeeLJUkJ1sxrMJ0e
ZMQAFRky4tc8mhYMulj0Mk0Hdb4iQ5FbnsYGi0V3PyO4LsGAaJ13Vqrd/Xro5bkP93Xxs42elYcC
s1xXNPWBLfrmBcKfQyinP6jUH0C9+Wi4ntmhU4SQznKaZDlfZI/F3kduIJF7miOtLCp2viYgM1bM
+lJWl2s6ICQnz1Hxv6XThfAhMnB+YCIMKcAvIKxSN8pc9v3VblRYoj6uhuDmXdHosra1L2r1P9w9
g3uIvkSoLozClKsqC292cauGAC/Vzicm0CHfukYHCPniu7ugyQmJUEV6mFh5dks98MvhpRBHF9Bu
4fjNgXC7yS+er79ShAUvVjaVBv7e2yFf4TtOr4N9gzBSjCpET2XFbGDBqZibU8shuJv5WPZciRet
snuJeiSj5oHQzTZdIenduuX8Cm8UgzhM4KHnVTJRL/P4c66TztqnKa5eQzw0SJhdpWp+8HfNXCiN
/nLs+QQdsZWzt24qx1gutu4nY6W0ivjoF7OsrZAfmWQ7VuSh9y1Lx0gpfSgD7xf5+ELN4f/8/s+G
MFiFPi0OAXutMSCXvzUWmeXENMi8jKBgO6ztU745cLEGUTq2wFFJNxEVdaheT/JXb1p1OqAdHuAz
UlCW5XoxI/xMdEekIsccz3RT4uNsXn4MN5Z8itL1xyo7xlsCXg3QMIuWsnSqo1xrmrlVOH0KhTeJ
+wrBCWdI/N1oiGT0Fdsx6H1FJ7SP0vWXfdkYHDolplQ3BfM4PWglFGCbFWhD7Tkkxc0BdmPZHUwq
LvZ5rjWsbYUZLw9vZ1LZm0FEptwo1wDzTMamC/1nhEmnRqVHLOqQ34gVgu1JVimFaz4abjkXCsJk
WgnF1R9n8kwBLDGvrSWGtJWaJ4gpf4ZXmgWWLzwifl9Fi8VribkBEry4CeB+wYyfpumBQlxWIWUl
DNWhMUzr7qX3jrCiRCLHb2vOMZeNYdrZeYLKfmHompNP7x+kIckiedpJREQ+Hm19YMmuV4ca3WBH
sIRq/si4H4SH5z+SEX+L55juGm5OY23kAmD305kLhxXe6/1CKsPE5UtI+wLq6uvn4yX43H91QE8s
RWhUAAgelmb/zva4gBZhLe452a0yaLRUec8dem6MHSADFp6q+UG+ems3PQcsrMY/Z2s2amEo+zGZ
p37TL2Hvgwh5jDnxWZ8anoQ7u3k6yT/cH/8HQwA5vwU7cYJGnEtCG1RFZG/yFZkgVg9pVf6CAgVb
xAapKoNwQfNzCdoKdH9Bs8RVhMk/yvZA919HXK8xOHXOZoMT5BtV/PIQ5JK3cg27TrMZmR7iSIug
+w7co6mudFUC9Vu9mBGbsIVSBQ63GeppOtfL1mn3Iaa0rJJNIAqGrnuzQ46LnmE9tgkfMbXnUx4N
6Ypwo01FOkbfJqHNYAHbzQmNUuQ/GT3IvIrH42tAOuBsIyTNHU4+3EzFzvDwTE19WAY0zH/ZpJAk
kAVBneCd0isoxaSbRYvpqm+NaVXyt0HTQr040/uOKl1U9kdNGJ4jVV2BpbKKkrhfUAJpThqaa3Dv
SVEnGDMXQ9XkfzH+zJkucqdfjv1OMmmfLkZqekrlZtB+CXgsC71V9qZhCPX8WLp/4e6Dz8osmxqd
rfZFxQKh+Dcc4Z0TMVsekyaS8nVhRdSho4bUCKF/xP5/8p8MtW9uFu8pUZ8357TY/59EXwE9rNgo
0bLm+RbKmdHgW8g+9JXEeb5Oxzo7VHcUMed4VVhi0kh0mbLpwQxuUShiavHiag5dz3ob8pVBs/oj
qEiod2IWRUDorwFI8vvFJwlDeipGFhV2Rjaq0o5N8WzECWdkBIP7tde73lnB1BTef1X9PbVVt8yr
pex2HvY1g2qWtHg3WZ8wQCE129PQqkV+Xkcx0ZPKO5JHUejSzwRx+Zceu23lbR1LweDIIkZ4f8TR
tI5lz0fxc6O9tFB/6FEIXgC5Lr8838Y1mXDrO63Y7AshW9kdiCPHOz5xr6CUWy1WYCNzC8cpWj3C
ymKEOW4ftcXbpgOIpQ/CfhR9jMdHypOZineEnaD6d/WQ0+HRx88+/jLwnso1FwmfKzayycYmi+Dt
XIAppoLulcAMlAT/yML1qgPZrTHVoNhci5PI/RGGM971dCZQ7FDxEC8CkAjfDJjRxceRjNH9uJYH
JA1rqZ1nMoy4mbR0OKInY8q1QQku0a0Nax1jsmbFpZV5vAIEaaSUE181ACzvtoBhaBBDbpwq5FkS
U7M2mPH71xCqTbjUcB2wmP1KK4MvKHyyOpIA6/sZTByvRxy0lRaT/X7G3afFeWdF1pWbiYD17y+/
0R0bi09rxfhCFJnBatGxFdQGapvfOkFYRE3sRVPBmYovjJBHDqaYSv9ufuGm3rXWGhnRm+D6AQxd
Jdx/dHNMMoj5fkOOHWGljMpoJlUiJPBB2jOmDMvisVx+R2+BjplTNyw9WvVhPqvHIYx2j6pVvKHH
etquC9BF2UNpm84/o3ZfQ7lNHE0M2hoXIhGh3g9opT+k6abbL7AhGyLBd706QcXHhivDHRqW1zvh
TKBf3Js4wCL79iXA/N+ntQYpDAOKdmRiM71+0k4VJnBt9MghBC9LCs7lvP9IN5qV7hIvS0SLv6c1
5u+L8NS18i8w0fW5eJi97W3SbOtgoMzRxp9h+/BMGBAGod2r83an8cijNvfQ72ozVehVJnFL5rOR
m5Q+ybtOypnZ2kLs08KYwU/0g+mhocuERa0vnn7h2a2GndfyEwlD8gcf2dwsgQw/l2L1HnUSx3d8
u8sZtily2ufSNP0xbeBDdmKV4oKiy796gWlEFFzoDbb3dsY1U7vXQQqE8W7gFXXtTVhYSWa1Mweg
VJKArmO9i7TeYt2BsE06B7V77wRkybBUibv8Dy5id3qE9s6l9Y2Z0Nv6w5NI8Rt+pb4BxGOC+oYg
A9/KDjokZidBoShszcPe1mSOB/x0QSfyGetjJmg6AfQbUCGzggSvnFFhdco0+NV3/4+qAnd2c70M
2DNlVzDrzj8rfyXyGzL+uFXZ0I4EYABDmmF/t8ssrkpbOxmuqnnrJrhWBY3g0tQa2bGg69YXPz+a
QR6+KSgheRN2e/mQS0m19cc8+UNQrAT9Vs9lj1kO8fkxu9bON9Bweh20otHUkvtabEHvM8907qv+
IlKfxWeTPcQSJbl9H5JMKdZy1quB2b76Yqe0dcUQaszZZWzvMB2le1l+rHI1NqFtaosY9R0aG1MV
P8IcBrDaA9RBRE8Ewi/S52W0P6T/q80xXKSYrrhzLN2iyA5fzgfabAIFI9FYUK6lBLW9Q88PdIEj
GYUqvWDF53Y7I1Uf5G7gqO/eYCQFlururC0lU1wLQxV+DmLiw9Bvx/jYKZqMQrMMB0CuqBl3Y6kF
Q6gi8z7EySQW8WwRx08nbKAaeCwPHFgEcKYIlmPEJV8cXg/Oq2xwbrcWzQV6s3PjBWL5YmbczT0w
8QnRJ31U599UgEJTtFtuhT153rlqVuEigGrKEIsCj9yODBfxslyCois+AQYTNYppNCqgfRG1YfhG
vRodngALXvbfY6jYU6NWH4PlQgEjg1EMdqoK8rXo6XW4TKISMIWV1RqyJQPuHK9s5cQu2IzX86sL
rcdcznRHYeHda5w3FcVWRz3lSMFfhNAHM7tZ6A4a6lR1yMYY2LPxD8Tu0i3xjon19GRQPM1kvTVK
IqwcKc4foaqLObGVV/rtgjDzHcj49+nLxeZ+QwOYcd6HabI/78AGkbmxeNy2qvc00Cc85cUZHz2h
Ryne71NEbz5YoCF6/55wmxgdOrUaLtkPTZJ9JNQ4ajMJcFtPvA8EY3rpy8DNUrTO3x+TLrddlpKK
z+FEO+VU3KhjYOTmUvcvwGLlw8v2JSdEPpw4z9YCIMSk0yQFjporL3JscUHp5kG1YArOsA6lRwP/
/XettgatEK1ctfpwHTy6l1IcSCkVHmFTRgCvKb4cNYXaxWZztZavO8j9HeZPYydbIedMSs4hjuHL
W03tywaSCqlzgX/wC9jgEyQ4U120bcMUMu92s9IQMIveWWb063OMiA+l6tOTNyQfCwHsQS/yUT/6
6iDBsJHAh6W8FMjwitWSOHiaALZ5aIMJjlgKJkvzEyIecmf6JM0K5NriqBzLLiELEMwIq9f9lNVj
vWHnGZQVm/yJ+egEJPN5kaDTvI9PUcrOleY5TXPA6nG65FvRy4NCEp5YsQkBBRkDWeIsutP03OQB
tWs+sv+9W+ZwEgFv2oc8GwGVdVdeVwsmx3br4s5trKjN4i+LWfmgqUsS5HGdBdjNJSDMRMkuTtlF
vrW+cuLPPkTzE4RwpwH2X7jZYwgFZm6BSThbAon2uG3geN2de2OvIWm7jrNtPL63EKJaZyT/S+d2
5ty1rD1EkgNCLlvMyWIIDCDg4H/7y+91oEmiSfvlzggzcD+CWmSMATn4o+e7AciQ2SRcVd5/Ldu0
iAmDWI6qjgY6OWwzBXayVxO6NaqaY+GquEJTmXAb2hKMzplbSJ0EOpYCnXS3KhmsIFDrTHfv4xk0
JGbedHzJUWUYRKUs+qe9P0ug0HrgDm7Fw7NFlgx+fXXAnXbtgIlXAUTM7trxJzb6kUUDmoxTf7oa
8JD8+yR/gLE1cxH9VNv9GtqV4PqYoxc0GO+UKtvZU5v6i4uH3aN5tj7W73dvKsRndNUgusrR2Gu/
xozt254/HhflhHG2FeCV0pYp8G7IvITW6j0dCvVy4IyS2TOJuZBzNulJcn9GmDZTJh2ODoSFyPd4
6cKgi8UFqIu3fqdFjvR96RVOx0ELKwtiLTLRoGxZaVcN4iupJP4y+dW6zlpJcJ79ck8YlHJB/Px9
QVXazv1q9wI41ceg8w1WYixsZIsuLgu0YoJ7YAN2ompIzWjBUomsjm/9/mj65BRT1FAlm9wNdIZS
jXbskDLE4tCDlzmzFHP2j25Yj0LtClZckfbVDhiSY/pd+zZtSglSpTpQyEjj3bfY5JXpwGIhVeBB
p46Y6AO1FH/X3NW/BBViHaOtBcQxVyywc6w9lhSgm6gH/vQ6H528j4VXw3Y+KPCVaYGVuALiGjes
NH8BCmwS1nrVWt7E19pxwOrqIIXQdP4Sg0tUNpzu/iDA45AfksdE4Br+CNehUXJAs23YNSaijHgs
w60dP3GqICrV5ucJwM1BgtkxsTEIVsaTZm1mpU8otcgUFFvgmb03HhZ4YEZ08Bu6KmbuaYpa1bsb
JhuD07QKAVIMBhalmjTkSzxuawBkTujce5zVUncqfYdxV0HvY8HpXb4+cnnr+qAJZ1b6h9m8sOfp
ojevs4gYiu37wEp5PaxhzZjbf5KNRYX/dMZS5P6ljn/kMXrbsxzAGMk/p1tEsTYGsGbC/iLp13DI
pfYkp3MLwkdsGAzIcUIno+jc5aYJ7+19F+gKqPP/8W3h95rfzIBfMKyXsStU9Gm8dHf2kPOOewrk
gjjhZWh7N5RikapKWFQREcL/Qmjl/+0MBWXPH0GnwNG89cZRJOLkcRTHI1i6yC1ZNjbFqRFj5MUx
aU1aX+n6aAAYaf6n11MRl67Oe+J5EwcsVg4iUfhiaK75ucc1LVmEvgUwMH0c7MEYK6RQjuYXBIrJ
ndpYroSktfYHeCkaraQqRd2lrLob2FpJ6UO7makOU+6n8Y1LYnH2+rHYxdB/vM3Kp77MqGLkQ+r1
+WV3zxlqy/cinAx1co5APUQkeBTAsQhCTSS0j1g3YUGRdwZ5aKCiOOEw0veKBjc4A8uKg7ys4AO4
6yhZwUc4NGZU4iW5da8ZNz/IkPppIzGoBM1Otfgxcf5+CKvmKiet4hhokA2yYKnIC9MvNOLuQpVQ
WZr+RDfy7mYiZN3EV96sg3qKDiLf9weWvaUowPKRCl9a1zqVFGDqywfEN+Ui7iPvH/s5r+i6Ky5D
XokszgcQ4aNKjHWDzvAVNSr29vMQfA/MUHX2fEM7Jfz0ALIhath7XXH5m4aUiF5dU1Fah0faMvg4
yEW3r6dEqMUTc1yj6S1Kzx7G3aKwPBm3cZT9MnzlxZpKTvNZmw9q+tff5f7ZmCzat3pY0MzllWmw
smlaEMHuXcl7QHgRK9xqIwKnDfzY5ylEQiCpApywIb8/+gnbrbC19CKz3Q9wEz1hel1ojX3pzS+z
rxSCBB8VcfrdFL4KrDNOMMUdxvt3OT9Oh68QcDpUB5aLH15KJHc8Jqsz/Dm0pC7G+D/n1qGtpUs0
KVUO3qU2rXSne2Qp/rc73I9JiwI/yiU6m+0Dr0QSQmwvzNEoxwYY7JcQm2qFHe6bqTmKtrltIVvg
PZbneEFNaOy1VcoGm8G+V2DbKY2+BMVZ/pokMEMrCcZGtHutxIXrrNi+SjyRHuWgaz1ZtEhWT9hf
XJiVAV4H66/YEkyf/Pkb5aCJbz+28+B+5xZ2TjiV0yL+1K/hNGyaBr/walN811tTKhs7C0qiCinf
OFFkS5R2CXtks794M4QvFVu4PvH5v3q9w1Pidq8sFu7Hk82wnSyXf9kNdhq7rI71j2zI6gnoJMMN
c80TYyP+bqvyCYdmYAJRATHgpJAxRIrNXpSZtbKecHCVm7q4rQe4e2e0BUjqD2FiQXQwsDnUSDUW
kIN0G7ouDV1uwV76QEV9RDkzfAgPmhWY312briALPgitr/jxnryplJb4pRqfaPLaVjmBO5jrPQOO
zywL/cY1EhRTNWUMtFNGomlXEvvK4+CjIkTnF+kHngJK3KogVnHbWpCXksAY7RHWudHdQZ+RpUVP
BLy4K84CBbDRJfi1j0oeWRHM5bl8l7ADE+HeO6K4rU386ky3IzUYPMsr9PnvbVlO/IJYWv0I6Y5P
AHnI60PKXHInElFhRNay8XzsdH8mFix6y0gc6Hu2oyIUA23z951eei1wZBE3hsaBIbkhcm1ZNiAs
wEqTIZ2kT16oK1EjXGfazL5QPIjeThPnUENjf/obbtcE5W3HbhxqFcla85pdc6IKhw/1+jImm25d
sbockVTnnOl62JewkXuy6ZWwAZP8Cxw8l8LUntJfdbrYFGH7qPnbcTjPlln5Z5xJcu3mEz5qrxuh
dQyUw/y4a/X8AsH8ZchnafB8dhCZgsnsc54RpaC64Tj8wRXgpfoX0fSO7PcHI65oNaipw9dUpNJy
3GOMSvwUtKTB7AgocwurWcPqGpyb+5nbGf2gGo6Ovommgww80MVkicG7gixQBrZGOx7qSOuzEXpE
WFa0cVxzmmB77TKGXAgLXBkX+WkOsaeaPpKU2NMBx0YN5ZxX2jvCg1lSo6uIqiGdMGqM3lhVStcn
4yHWQ3GIARToIAQH3M8X1TC5ZN4/F9EesJqOGNndn0LOgCKRCY4UEKNJwvdZ6RrHsd2078h9b4ap
OG+BtcoQMcsvb+buXku3QJT6Hk2dlI/bfLoPpe5jCjGmRuAFMb5Dz9wECeg0YJHdvRgPB8dTXfcP
2svu8Xuy25Q8g3491XTPerkYvFPjzHd5wdPWj7yW3cZwkZu6ul3/lfvFUblLyPYFL20HeObB1PoZ
0U0PXooFuK1Z+vH3qbfLBARFa4Z/KUPSxcYLhyfwaoVvN4CSe8JYJhPHUuttpncipGVshDpAN4Rf
cgyOcaUIGuWDf3QMVqNPWQT5oQiIf3ZjPpyJXiKRFibY0PKM6dg4yLtrI9QvOr/7+6DyIHNhIkKd
UyBRa2xr8JEQfprFNn6MAk4Pise9nFVsuzdY/7XGWdvrwQU8sSK0vN9H3V1Iq+R4x1K/EWiQr8XB
+P9SXm8SvO9RpK/DQFATvbRF05GI0LBY3T3X8AoZcta35iodb4EXD8btsvnhIF/nWEzFU0m5hF7Q
PQIXFRASvUKIQncn/BEWaoM24yjstsdLfDSPCN+16NE0VPGDRojh/vgLEAkjj9tCDs64SoNHKNfq
9kGolxQrzeNrHqtsygQ626c/60VaLPqDPpI5O0CghvnwMZ3zvpyyNTEJZUp2mCgbelOdPo1E19+B
Bo83fIO3JSKP0yCx1BUKBLiIUbWkOjyLCMJu+BG0rt3fkOYoMEq3vSDh0GZWBVwOxUQZ/YXWce2d
mlNDDamMw0UQCNp9Mj8rBIRcFd5tad0yTQcKUXlZUb7VUa6Z/GXSTgGi8IYIZY8nL6SannpAErMh
hrHRIeD4kJ2GBnE1SICaJ4KMnKoAnByUU04UWwD8jj8M8Egg1mvyi37QUmkvG5j9ZOpEQbJ5lwG8
ERh8jdDhroOu368nGRAa9UWTgHXlxG/D9WeVXcTpYlBGuGs2ACxSAyJh9DxJ21qbqEQ6/lQuKwwv
kHlq7jEAaAX/xPbzBYGGkBkD55xa6qHoOXaRa6SCvYJGhCm4V1GZiYluw6iK2uGUOpLnobmbwiiB
FNfQdT0cYueH8y5A4xvXCOQV5rsK+frk1qmg1eLrrZngdalATQGO2rGp4gmKWse9WLTdy+XqTcBY
oLcEu7xCEZ1f2IjJL3/ZWrEiadWxoX0FwiD9gXU4X/LQ0b17pTRMMIq4dfwFhFAOBqI3Y5SHESQ6
ZkM2Xqyp8A/5WmeJ/YPdBMGBAW/FiEH+S5JEg4PrdcX/6yw4AzXRRWk3WZeexOF4+FYNj3hUau93
gWIbG42vMlxdC6jptQrr19c1aKA2tJ9xoe7mIszbs5kUiq8+2eybOuQKw+1EV8jT5SdnDCsJh18d
HHFhEfg/y1pTyel55BufW3HioBUlSi+C7ff1UGaAotpBpDZMtDYkOPhF3SGsOeWhROpkTDSCk4OA
yJ1K6CEjD3sc59sBOda3nyaWUDyQOG6y62uFiqytoCOomAagU2sU5dUPIhz6Ect7j6+VQyuNG4Qy
XZ95tU1ChlIF2vT0eogmrYuWbXRppCIQK9JgRgtXP5+nUNCDyDdREutYK4+sfKIUamU2Zda1n5If
GPD+2fGwHQRI6jS6WdgPmZVabmYFFzQgT6Y9kAmlBmPnfIuIgozMgONYIEugoX2xfADkblcU8avw
Ouxi/RSPMEaXs/NF1jde6DsRiY4f4dBurCmfRVeCfinXZpBi6V7S2ctIszOGAQegYz+8UFeCWq3Z
NTbVINzjpg4FjrGOxS6K0/P+WDHsjuZ94Feq3YZvXlUPcZQTMSeNGGiKZ9oiZIt0PiIjkKJGAeuY
1AwhBAiGYLuGf+mmXvqrPOhlyUzom2XwC2ft3nEZlq3Pl7RYO0ByQXp7/IfiMEl1DDNrYzhNyHCD
rq/sKyOtgL6St9mXU8Q3jfXku342B9wbSAcbRiKQYZFofDTf4UgSkPtlzL43NCodC7RoDlw8wDrL
0l6NcsszgXSuzsPsAnNJQcgXcpeFZ3/MbiyMWTGwsqIOSUJroeuKCO/7VIcnLVcyKIVRP4YGOlXH
y4XHEVGaR6afYvizuB9DyjSHrtkhQSGT2jtdBj9Ff8aMh/6aI8yy/rRLRmFyQlurXYAqJEvrb0qY
B5e92YKoxs8xM1rRroyr65TUiZhLbc+FeloWszi7S3dUFzDtwS9pdvXQq4hrWooOUu6flhlpLZlu
VfwLkMalQbfo20VCkTwetCdm4yNhx6wpK/8qW4udUi3PiwT6E6uDXAyPFMWwaUH14xFkfj8FweV1
oTGj+68uJcvcDooToavZYshhMvCqf1F7oALqiUKCL7qyuV+xEc3JWAwtu2ugg0Sd8zzCX3wxKvoQ
vOzUXz14aCO9aDfbnIXNe8LBvJ5SzMUCmZ4FPkTCMSAaMCzUhTnab6ZIpnGGJcDTcpO1MazWz26Q
rL85j4EGZSqX5crT2BjXB/pPg+AlqMD+EWqcPm4Wvqlg9RukqcYal7zvwi1VWoHuOcs3bX4rfc/b
zG36yP+B3uyYT937T7+Crj2tkt1uRcWKRKsSOg4VkBntncZPNto/UIlzBLdRv96FJgnyHSCdywnT
vrI9VsYsPpjO3GeNq13NjUOxdUtiylRHg2uFIbyxaPi1gZjkUOk9rC9rVe4N5UFpnctwzOei2CXi
3HMY3CB/yfH/Qg3pJFBWktesz6funhegr1CEaWxdOFdZljaMBjlT3mACRrVumDYMqRee6Q6mCh+t
nJggkcu7NLfV41/QWD7l+GNBiBSKgGnAXTO/Vh6bfWi0C8rUbgOsyY3dBDZSA7rUrRDBlSZf2ygr
KjHkq++jvnYfZPfz+hpKSCEPfNTSGbKgv1r8L9qLp2tyeuLgGDo0ZHnK9IBJUb1/y0tK+E47qpbb
f5Jojd+5CAOFQZwQ+FifCNd1x4zRZrAzQ0rCPcqDRRtfIgSwX4hONqmcNucyDttYwVVeeBJ8+flf
Yc9WnXw12ckmJhdUiPxzteY5Si6QKBU1n6w51Iv5xd2C+Pvi5aZ/ZSfz1JWGRIE+2xMC+fIr1F35
M8JsD+Bty6sjo+qDqOTFFAxbbXx9IJzzMkhmR3E/negfVzP7iLhumI4dD8GxQLIVpXfIUkPDe5ja
OklDheoVrwHqMivnYCeWwoK00w1gk9L9qJnYt5AJYN4cp0mMA5AqsBZTbpSMBppHqNiudE2D0y/n
XILuj8ZS4eXVlnzyaBw84Kscpyt1CscbWUrITsKeZ3C4mpc6IuoaBx1KxOtV/Gdv+Oncj5fIiCSu
Q60auLt3iJTTBuizPPoCtQn7GP+4cAwImgyp4vhg/ktlJJMQ82vxeGIvvZdifVVjjLgv388Q0dXF
kdF72oS525rK1d15+QSNOHsTag/qlIIQcncefkWtFXhg5CPFeKp3DukV0frgvMIb6jhWVs4vfXxh
nUNTrHi1hEjEeXUq5QhjYhZgMp9WqwNNSGylsyvtVxWXJ11iKS6nJMxNYIc/wmKf08v7GpBf4Dgz
fqhhKmOUqj4lJctsKy8uHwfh1w3pj9PU5ejQ63WX7eA5U9Ad5EPNlB8Ys1NnK15vruvLEXiJmmZC
cBlrfO86g1bz2JAPl5cWdnbxK9IaoTLg9o6ksoUBLR4oh9UMEIHltz67TA+rfHWiLBOOvPB3C9v6
64s0D1PFLIRxepIRz2eXBCJf7PIzUG2u/xmxnMhinxtbTPTc73zxONmMx+Uvl6BvBfH2PEC+e4xg
CzVSLnsvlXHl4bcWVI4MxraZ/GqHy/VGC/2iAKsYQGvhQA+o31Os/l9Ddn8ugAmn8s/ApPzCO0Ou
XFB1UlzwEjP01KMjxd1Xt8ZChTIE1DLEDWFxiRiWp0++FivLCTXxTUOGv/D0C7xyMAvnjrL0khRU
vvfLAw3bErJQWwy3x1ytSgIE0piAME7H2JdOtwZE3NmStcySxxtBgLWnKHY5CsCPmd1RfqUg7z03
ICnXxaHb9yi8+2sAVLgGFgyA9O1vD0JZqtEMQpek0QogpM9aEZvIiZmwvDW0EZQsLq/LSXyIIj27
8ROkusFhxnxKHKz7ZFZ56/eud/1Ut9rynvRjy3HPj/iindFZDYPaNUqANtNbxTPHhyQzc7HP9oRg
iRTniC3dwJ9btLF6nIlDw25Dn10MG5n0p0dy2RUaUed45yDNXReRpjuoQHus1BjfprdTX9pksqFv
YYEd5F6zWD9YNO858/bRtWp3TyMb35AkUbfeifhkC8PrbhxRh6DwZw/kpEJq21QibUhGx4KTznjf
ZFEsoVvZqIWhhiYRRq91fW2O95QHVWPdVgNPBz/xF7f6OkkQzVqK9Lc555NIXyXE9YXGE7agwD49
iJGPrpLQFJp+CctShjxoDUhVK+N6XJgXW+p3cm4nksz2WWy4Yrd6Ut3Tq4+aobBKRNqqRfumFLIz
B5GCYLEbPbM7ShOqEbNYMEIsyOH08EVBcjwz0nKbxKxtII6mwfY0/6daNWUac83bHMY25y2wUW9M
WXI9AmwdDtXNYTFKpsg7mrnJ9+uywjuRhpIaxmpeo2dyk0+n9EjCvZyubknMi1lqmyxWZHjCNV3Q
NVXl43sXdAgdh1cjMAZ9lMMVgLn7x2N4A3+kRqrxI/2IB84MOCLEFFWngKT1ge2xGrDbGiYOJLRu
8yc4XuWhb2sxr3ck7airbKWQYiHWRrmS8/wcPJvSFTzz8ZuqjGKqldnzMnaLXmPzkJjiwzCQL+xN
il2nFgU2IV2+Qd2frK5+vDDCX/IKUBSiTdrP87Y3dLOGiW56yzkLPk51IGRWvD8YuE++Tuk+kEJl
XmnGFEUs5F3T6be1vbGxG4NrXl8JLYE2Yvc4ENJrmRHX1Jco9PJS3X928kfVx90z97rHsP7T+eSE
jl/bpfTBghObvkB3uYcPzjlBgDU/xcCCoHmXccn5/NqXZyUsTTiV8pweurnFGsaDXAIbzb16305l
RrM7fKw9cqTPyZO/B6pTxqOGFL/bjBlT5eYrxpJAqZBQROJNYuMMLe93Ij2n5Ss1euGABxAAPEsu
i/D8HUiEs30xXp5QIJctxdx+/AZM4obB5hxtroCAHhhyl8lF0QTGI+6nafykItxLaw82Y2JSMHde
tFbSylrQP5clBwhz9pqszbpg4Q3MKclz/adhohjw7tc+eTc1m6TagbY2Xhmyrwv2pHri9+g3H7sB
v5Tx+BAoVsNq59fR0F0PKafzw/1WxCc59mUGs9mY0HK6RRPttq8ZSPKAiycX0JbB8psp7uQO1YLx
qCX61bxO51PoaiFVU0JncUmbjQLUMC/4XvtPP6RvSn/ZR1IKi0PA8O26jNp4DGPnGU1Oa0vUNJzd
cFeD1Q2rtd0rMJWSmCONm0vLBMewXffBGe8pAHWqU9b/lEBl6Edp9Zj/gcRVTwhX93inTrztWjjG
rzyJIIjDLPIGFhi5K7Tim+WMvvQ8DFbD8ohhxzEiOY/B790SSDZ5qJx+yh0aN4HK/rzV8Ihwb4rs
u4tZQCehXTziAmDD4VrPktO0P98zCD+tFl9Eq+3VQ5/cGTqRrXSi/8zHDqBAlT+HSsXuE9uTrDz9
oScd0q68AmzyDRRC9JTL/2qahK7DPPy+35nfWBtqwSUQZH8Yrqoa/fx0XbeQSh6VSiZMbQ5tj8Gv
me7vbbklgtpIYunWQHPMQgmNukFG/o8KjAp7o2I93OO9mbsOgwZY+B7dCpCg7Y6BqlUJzNdg6hu5
r5wuYNYwXC/CkWKlHM9loG/7HEY0NeRHJOydeiB+296e+2o7bV5zrWqh+Us7hrqIduZqI5nTFYYF
f6aG8TylxW6k1/wvECrlpAPPo9mFXAFiFEhdE3lz3ethA52RcqhElOUbwitwh9LNmzDGOJj2d6V0
4492/zYbLKiLfFDP0MpR2yC1yQo05j1JIusoViQb7ppxD4gvL0j8EyakJsj2qLpUwJsaxTHPwNBY
XQL3a9Aqy/mvS+KYFOnHpirh/1NGq9/6IJsGjUbgEv4R/lm1crfLYr4kyJSVhqBKB+VvMvESrxS8
iokCaRh9HfLXSPfTSfgP785q4YEVyUaOsrtXCwDwAfWVu552mSzrKmX6PNinMjsvMU2rafCf0ins
6B99/ODNBYH6K4397eQj3/eTpLgDlX/WpA/jcWxtx3uxGns/WL7olmoky2yK+kZ6aMMvrWNltW27
3+c7/uMFnLgN1KHBnComT3QGOVMUrRoP4Ukttj2z/bwbIUocfGVW5r4NciYTGUEPjikEDI1/cYoj
nHim7dyeUwJqxnUXHrw/YVSOjoGtMtLWlJ3LRsSN8vyjN2ZhC+jboGk1pUS4spXl5CgD/bEoUuak
IwlQntDPIfk8zGlh/o1K0xJcxqIbSjZwr3Gh1C3yRo1oO2Wd9KOztuD7rttmr3Fp13N236TOsGMz
NalO0dd7G3Ssftp8xNp3PvqxEQwZR71RM976p9hVs1bUUhFRxbXfJgWNOcs/SBozF8aQ530JOuez
/hkIbNgaJLtptKspDXaOxPCHjUqaHpaK3IsvdoyBF0uUgcduVoNTm3Qm/zxLIgsXS5FK4Ir46RdB
tDe/fKUij6G+BWRrJS7BAi27GDYN0TLvfEEw8BoehaDtLZqIgiWHHdOlQERbKM28DBUmpYBnyMXA
SEi3f+BuJUOXYED0woZ/Rbi4yzFuG4jBgd5PuRuM4wrQh5o/2i4htxo9yXBw/0TaxXdo8MaJ5nPL
goMDzCWge4K4dg9gq6gY3qxHejFzuf3ustdHikfNe4fiaHof3HmlAnF6kGdWOsdOJtXQN4vspqsI
3flBjPfzcWIa1RUk+0OuO8KTAOgTLIByLKO3MDL27TfjhomaPR3e82p4QpBYZ8vezdNXdRKt3ave
cDLkTuU8scVclZzYX+sPYBa0QvwXf6now9X/nd9JudwJNskpw9hZF4PTW0tfRmiWBNUbJ2Aa4Sd1
Z7f0N0DM1OqnK8OeLInq4jBPOxWkJ4jj6t6RCCEkuVLJ/ORRxVY0m861vfBdSp5rFngiLRKl42PI
fT82OJ4Vp56o8/wnKeXLlYxCLLfcbikTmrPB9l2duWAoQoM4Ek8JQ7tl3qLbAqBFHfk3AKA5uuEa
VVGctFVKgGvBTvUIp5Fxy7gOzaH01QkXpyrnc7OmwxYr0KtGu4qs3FJms6drSlk3UctLRk1Nvy4x
HPUs5mhCnhSJ2cpTOsYeZLORSDYWl/n2+uGdJEIBVYUDSNDx8fqks/vMCkY0BrcsHwYRxIY8nRxJ
FbH1QHMkDzqJqSNIhNjIA+e88PAi4FfgpMqHnm839F57u8AhpBS6jq9RpYL6S8uqIzQJyzGQbQrM
WhWonrcvf4HLxBwahImxuLelvYB1s2b40wnNUOmbfsW6gR3TAHNnVUOnnsMlGQU1T2bIHzAOTFdQ
dNXBLYs/1CqKs20vPFQAy26yCwzWP/RdC6ra3Bwv+c1D176uoFRjkPppWhNxetA/7JFq9tXfp+Q1
KqYjnQJq2aBQkY0a3Ax99y5T/f/g9fsWit6FJhAJwAUEDJhggOPyRM8jzL3ECOh64dTsm56sBBBI
LUjyD15GEBKofyiLtq38cAyqA1RebLWu7v+Xqran+XPlpcAHZV0BN7rahpy3p4Pb1TNvgi6b1ke9
It45ii7XEJ8hAjomb19TtpM8J/RiRgoL+MszMZih2bR4+0tuEPi8XLLbgxvWwdBJgLIUtCbGFgh4
4dyS5d+1Wd0hGaN+t0/Jmbxkj7U3U0oJ8MzdWamzm/xQBt0CkbXdvqITZZmue2gCLvwzVJ7+Ar4i
FPxkeq54sbmINeOn2yhNxep/DIfVdPQrAPK8WjjBr1/B4fPXEbiiY6fehQuYcdsP2/3B9Kx3jLFl
In4yOd/w21WWtpSK8N6TNmSgj8qjewm8C8NJONZ+1wbAWLrvQnrVu7hmftgnGkIwtqMBrpiYo3b9
oJQyHa6fxkRcz/tPdOZUXgYgtWGRa+7spJf+DtJYkl6bqLB5Eb31QD+FsaLS7Yb2n6Rgt9TMtbKk
4t/qyV2Ybqnp0zsNbDdnbY++c+NsthBTphTfFnNg/DLkyT2Wo0fROUwzztzWebkA4KSWKYHOIufz
pXMgaDpKCG+XwSXsqnSyQf+WA9kKN9PRiaaKS9ARQY17pUv++I4/Lqp9dMh8PNh3cvwcIOcxYAWb
BCkPDDsyTuuuT9MbwTvCwN+aSAWO8tiSiGfhi2tb0RqknYTseE0v5TYh+Bs758lvGV3iD2wB4VoQ
+B3fonBrS/2QdwCmL43q4dvvUrqC872SNQlky1hGpdwSSu6wzsTKlLw7upX0aXTpoO7e/JaIotO2
s+JoX/dMpWqtYZq1hStWojJMdpJTTl9rVUwsUqTIAsV5eyjQZI2ev/CJ7J3T9FKEvj7YmtPTk9cl
NiI19jPsovyv2hqdWMjF/6Y2Iea59uOiU2yxyGulxDtpg1dBTITLnClByIp087kZX/+vpOHjBnSE
pDQ6jm8yUTVDJYzx4/n4raU6BSpIZD3voUmk8/5mgxDVL+z+3srN8DL3WaDFjm2rKKOuUwkHUF9r
T5UB/eiYsZzAuufptCFhy7pxdOI0URh6lkdMeCwKc8cEhjFYJ4SeSfG2YIKwWiGADcycOAz6hkqU
jENiGbqyO96U1I/lu2BFk1tWjhANbUj6l408kE5OYZTbnMm1Rk7KDpIqqw3zMHeP+E3paeff0it8
nb7fW60gliMOUxo34osG7H1TvEjwTiNvCSaaUJtQ8RhelXJS1r/8BFndkV7XhQcvtuGixqsTnw3i
zMow3B1hjGBw8PDuTkCIvFYKDyemptOYAK3mOlrZtSWtryeNheVPx9hazAhw4ENKirsALlwn5dav
37/XVkV0UgAx6W/cppxEIVdqj00h+EHKQVrswf52tGIsLxcR/TaqqfURa2nMN/VbMgbe4MqCAVNR
ZADt4OiCLhfa3LMHzgee+MlbNo/7LvdG7W4TI647xYPsXbuPZHAXDgrs0jSB1tgFDK9nDaFNjhx7
ZfytrtUSFgc4Abtjtkfp4yzJVRWEoa3+Pmvq7LbfjvKSp4rVhG6SFRpJcRiDHm9JC2nA8uLHCBxk
LnnDSQbMtm7k3+qlWcCamUGBo/Q9hFbgNlL5X2WOOSqndKnKIgfZJ/e50QVFzcQlMelOjnU7axyp
Ubd5Ml0Jv+34rT/raWc1Atzb2R6x+MZ3MpunKQ3QgcM73v5IuDqj98cSZaSq46/8nHce8zZn7Y1X
a6+JUaRVbE5lWdshAGaXpL6k03hM0j+c9HDM8kHzoU5Y8h/Ym0Hl+zmZaIhlmK7CfP2fAvXXU/eT
wziSX6QCZSqKSB1EsGnplxK6yx9TeMizNPGh53dXvjJbvHCxr1KNm4vXs7j6zOdu6gfDDdRYCSzG
mDJtk6hJeWtE5MxpmW55brl9IGYDCLu6tMyT/2LKJCSWprkUOzi0t4hRkobE+3jtCbgu+H2ctfyG
yQ8xtWYacXlfwGAcFKjdLYMMmLGIaHvF8cSqDqGIecRQb7uzgLE9qfzcoDN13tD+kd5bA/153jTg
ji/zZSiZhLXxhbzofO9ie5+WKTz/pDJ+R1i1/BjOWeaKYSED6nBJyk8lHjCi0ErrTZNS9c9vQkGZ
BJXZgOmvb0/ITInzA3HeuyO8Kf/zRbHEedQE43N/s6yH91/h+TSzUvMQn4U2eIE+9ZtFzU6KhfRX
fs4nXDJD9SWk0yOIoLt3JJxVQlScCZ9TYWFtvhj2Yu1cfQ0zTw724nC0LukNZanq3a5qRxEAjzSx
GekYpJzaUB8Bld0lc92BrnuCZS7cUJ4vYPOt+/MtxdV+HARF3+TE+CK52LG2gxydla3UZ/T5r61h
iCNWO1Oku/McIS+e620ijDmmgDz2WSU3j8W/bziZoOBFvZM6jn6MmzUBhFaQR4biVvBYNCl7KACw
T6cqubMcfyCAEdEzLrKVXvdlfQ2UBTktbTavfA3pFPx5EA83+O7F8Sk+uSvNHMbW6Bdrnke42jYU
Dz9gcdwcsv7YW+ngrcnfvZxpoq2/AHohmHS3TBMZht4BS0y3yGva5wxFFiNgls6PX2S1YD4lQ95Z
paW4cw2a4kXBxuAE/njb/ebHMUN8FpTCUXXqXpb6t9XTdlAN6ir/i6IMNgR4YKfIfmI0azbI4E6C
3l2GiKdgABpBM9+EmY/Soe/gOl3CP9NR2YeYCO7lloNnvUWz/U5P7T5s2zcDvrIAstk8dP1PJj73
WcbNuAcLeRfknyvfFy3VK72REUWMK48BzZI1O9ZgD3h82BMMhtALbHbwwFtYNZUbRE6ffb8QAEJw
WjwhsmkDQDw59JeDn6Cvp25MC99zxR5vw2w+lQWdvFh+Wrkz6Hy7G/DtigeYRk9CZ2C/o1Ryysqr
QiNMC/9neTzAjB/+pr81EY8YdDniMwuiqAwEX7XMCmwOlXS1higu1WTRN8jUXO3awTIODXz8rJzT
W7DmVcJFoMUDQ6sDw5/37hJE74fUcfcgmSU0okifVM9Yi0msODR1AEoQpIac4mq8yDAnU8ilNAp1
Mxp1faoFOsDhiE3UYe4IAP4qGkxNvugCditGG8ZRNI2mB7Y5vnlmGRNXGCxlb/OYBc4RsK73SZN6
nKIMgOKZ4SAL9k3Q0ZYede2XGwFtngWBxCc5GakSaIa3QY/plR9dKy7Wctj76z9LRz4x5pHBkWB2
SSizI1FHcVZ/P5rAY9kc2A+J+gr8hIArgjUi+9L89kuJz+rgxPv7s95YQGggcqSIussSbF9MeiT2
F/ypEuwxd9f4QyiYzOhEOn4kpTEUFyZQd7DiiyKgkVIh0sUTUYyrIcY1xzKiH50rz0tC5lOJ2L99
Eel7i59D67hcfEA6KNy4x4zaT95gRi9gUuBThRNKSS6AkpYQzM85SN81jBqhtF/BMUnHOyAaYezd
l7sDhq33BdZ/XVs0p3GuPDpJTuTJgMa8OZ52IPawJYqw2Z3j0R9jct/xeucXgSFgcRfFy4U3bNEc
ObM9rmteDGRiMx9d1eCCZSJ5eP4LNxWaavG7tQR6PrKHyscnhc51Z7oM1zHC3ZSM231C9Nwbg/C/
LjbjuKBA/29ntZfT6zOp4IRvtzaC6zLNC8nMDYERmqhE//ay2hLf2DGr6nKRGa3maMmBF37Qd+If
RzoTt/E3Y7DBNoKWUP6Yi2YYLcL5b1STbLpR4XzFDbALHKZlwi/2UCwwGisRKECV2AydvZJKKcNQ
kMVuKXI8egzGKAHk7UBf4USPK1NKgWjiGPkDUM8f6BfepqyrzwRpSPLBkOcWtZcZ9JBvFjnI9xgk
G1enG6P+PJ/eea1BDjc+od4VZLvGSLiIT4yPPulH6Af1vs4MpmiPW5lzN3m7Eo7loPL6DT7pXRSd
RykRdEmN80yqpsDeh61URqzNovLTL2049sZLg8hjdCc3uiSdbcRV+jW992LQ0Li/+PQV9K64VKkV
XLRDWLaORziuFDfAbcUKCvSkYiZ76ZtkB0wjedY6MMDB2Hszh4Fg2ayBDy1OmAfJNgs7e/7DpStB
0M8NNT54nda65r4DOEiTZpf8EW5huE3pAlnsDgFNmxf/UOlaV0vLA7nwXR1Fp41gIJOTkrSk3ohK
6YjT/BkuN3EoTY6jHEw71TyV1xmAHnfTI8D0y9Pb4ZeQ2ZvxET8rYb33G0db+f+rfuTWaUrvayRq
99ARdZsniCj3HLXUvG5MOGZ1+o4GhODWUrvbcSPJ50IUyXLE0Ysq0LUOcoAKJ7oHGzS0h4Xxr8RH
I3OZRwxH0uYE2UgCZyMyWiazqfGhllq7S4uBIRmUv/BHskzTyXaIszCKakLE21l10JbqxCW7GBCC
y/YYCQBGmYn27BzimTd2Qucj/QBW9olAdUXRL9ZLZTlsqF646xoBkhYd8iwr6FDVKpMrDh6ZLMCy
LfkeXx6mpNp4dNCismyASyVn0O2OylQI/nRLUM1pzHmBxM26dSD4xC6qVXe0V8fUWI+S1OV24aJM
2lcpY+7ux97a8WuqJUPr5uP0MlZEXjUCvWgKhjN+TvIT5AumKLaTvN0310qc0gyYOXxExWXadewk
XSR9gdEdVipIKyKqTSFU4MWSGg2257f9kFjJC0zie1qvXPoNyIPrqCIhDxg+KjqIbgyznQ5DhO0X
3M1WbypCzzkuNVI+oWoTqmotvckBjWA0aTxEANqSzoDOZvOIgl6+pkc0yJqDv8OzpDgePezhaicf
rhAJp0/0Q3UKmFB5DXXVnkEC/2PS92soxs+2t44Jt0toel2tvqG37O1MPDWXoXVqXXMnAlPp+vpx
hfrzmtBQWUtucuAI1Otmuqc1sNOTPrzNPAjDUAohJOunHRiwUp3UWrDC1mb6z8Pn6xuGavW8zNEo
C8egQS1FjinbbpCqXh2LSlbC5ZYz/6AaLQXqkYxFbvntmzlckqCUQM/V88spduUT3K0Jl7nRgfEg
9YxHk0yh8lKwJgHK0jS1X0dStCCJfhYEzDG+mplDO3zkUCrJU8FR+CXLBNSOMjQBBLH9kOjzrvWW
nZMzBMXkXZDUxL/KLnafPRivk4fMTKMSp8AwFbCd5kzWfIH1yHxNsZmm2cMDLsK+Ysz3t6c2GoCD
pNK5ANnas/RfWQoOKy4x+zyyoKiIWWPpYlbiU6SeO//gJWYTpsmCfVGOKq2Fvv0Eg1pENiiOUrI0
4oSDGpMdnW6yu2t0HH2akmpAzzD/2O85GpDMU+ag2ISocfq+yliq4pZLglyrkpwV7vzO/tY1VQvH
dAwEtbsFEstB9Kbs5MwZ7RRGCHWIpj2szUE4XBYK/OTCR88pkYisPxyWHDEm/bDRK97Ug3lytIPo
jOQSUS6RWT16NbEssnRu5VxkmZ7ZuLMO73EbFmFGi5hb9C06F9GFKxL7WAcfeDjnoTbyLjXnpyGn
kb9pRig3COgxJvTdrkJ167IyHUAl7f5Hx+m8/zUoxQLS83Gd9zLW17RPKDg/MNQKwGxvQ5I7ltqQ
3+aJmE4yu+ClsOBD2uoLKox92oaggnV8S6UMe9TCcSl5U0dE4p9120rJENjHfdYuYjvmsxl+0vUl
Hu6huLQoaw918rN/Un0PJjK4hFIV3AJKwsb2rJLRFUm26qXnr1dTyVxQ91FZ3zQttRwJ4G5cIXKb
IgpZ46UJZ0LbHZknSODNV9D0tL5CjYK9zFfnoh4kFGiBQ53JukMOVZsFpSAaTDTGsEOQmOzpijGz
4JCRksqb05DeXaGosqkP5EmIb72zvHAEUzvwrPoDOEnH43kYbcTLPB9dQik/3riU9iTEG3wExru4
4TxHqmvxOEPVLQiudeht2kJOJo3POKgLA+k7qYZsJWWFB05zTQL1cYt5Im1EMWjURhUbxEV3fTV0
iRPSnNw8sJckXRUC/4dpHx8dk57Y3nJ9lcDvThRVqoy0Y53pjneH9bIFLbId3lHazScXoRkWW/BF
SZhbQujd/iW7C07d7P7tYK0EKB1dwB3plQhR/q+ACloyvyWPuDUvn5auZGcjpDqPZAXpZRDvCSwH
YhpNM2yox65SZ320Q94bhDORPq0dDH2+m9UdEjCTmSJzMgGykes/7CVpCSz5Hz2YhCtj0naDRrcG
hGjLPv2KZB1fXJBTKoH0xgFqX5v6SzYWfpCzKjAfpSe/E1+ZbsawDzIfb2oWBn1kB7z6tka6xpq5
kKgPGLWYPHAhC5ljb02W2UWepbgwePfg+FosbO2nRwLtHmQ5O+rnDswxSSm4NTn5MToK2n8qcSGY
7aB9YJGe8oMle8PsKqJ7ISEWX1vYqeaUteSiONLsRPfUePdWhMnbFX+mkzxa3kMtvLNsfsM66bcW
KCjnLKYZvAjjAlgDt44bYu5SE32Ar6bXx8D9wJSPstexSokS4eCyzEtHHem6ML6HiE5wg6f/hssi
XqfApsUY0TZsPDhthNruSZg2yvchzeQB6+yY2z7Iw6nIqn0dvf5bYz84iHuORFfXTQBQoZMpbbeU
5+pnJVOSo+SYSygMeZBvhHbzAQSSEF06MGF+0bRVb2VDoJqC4g2vVU36VXQCWkt9LWsPcRA/B2U0
inH62bsogS2EOiL6it25x9C+eLsJqPWFjxKFTnOiyxcGcUmOqNQ0yBhuldQ60eM44Xh1IzOCbUTF
el3K60KZQtlJSMuJvXtuzFcPE7350F/+eT5QkRPO/pRQpg3WcG3iuJBSO61aRYRpkuI/YjFDtQ7n
wMDPOb2ywnBubxM1As7w6DJT/NtZ1cxndRRXUdMUedWL4vh+w9/egPrz1QbHYlze7T1A7xp/xSJg
wXf/9U18w3hPJvlHjEYzVpLak1S7FZfFWg2FBj8gMAXdO0l1Y/WcBBpjJ+mYoUQ+uleuFsxKEhEU
cLCb6BzShmhFI0paKbh2GqgHTkWGx+IxMTQJOYmGYJB0MYjghNO64w5mm00cAk+QY0m34pGtKYFk
LUt4vq38KehcdoU7X6nAkWkXgADuaOMNxPZ2IMHI6Ejh8g3dJz8xq68MPnvpCmTkLF1vmSSLSXXE
PUGUSn7o56oXJDNnczhNC235bhT8BTHnD8pTAnAgQrVeG0kqOv/0WJYZrXT9XNnY4UaEYR7NZw/9
3fFtdL94iArdrqoz/gYolP/LLm3lruWZHX3NtPXsUvUmqFf2vIBKkaaeZ7QMlfEkfA2z2d5nLrVf
jmpELiRNUXed75LICPAuhakQpmvBT5wfXIKrkzFupb16U3X03N0ZV1Q45TqVKTt7z75314JMcBTi
6XMA3zfxCU4AuNadUFBKnOfD1Stz7+bh79D0RV7ln6AEgtXKY+N6mQMy9sazhFB3wHBpBZ/zIIEY
5x41xENYYRRmF46uaCIKVC0jsQ3QRBb7BYvGt4q8Ih5U33rA/NPSov0bgLnAawD+uVogkr/w1ILa
ogBHTMihDl/VFntDB3rPyOx7VVjz8c0U0Pg8fZnEyZd57JEW83WVpKempFNSixqVLGo7+W0EAiQQ
Dz8/OoCSsFxErSlu1W4EiRO4oneJ9ZmUQixq3yN3HcD5CibOQZuLYbUG8NG44VhU5E59C63KEYeL
URgfPKdzU+hs6YT/hRnYkZ31SDd9c1qDe/UVxdNq1i9esOwjrua7bwwW86AuDQS1xsf1Ehmg7vwE
dgR/eazHIChtSoGi4CLYGNbHAUjNkGbmKs40a3R2sFVsu2fLIEA2vtW1dWim82gB8z6BGB5tTozT
r+G1takSCTOfJsIyo1Cn5CbBXAZ+VdAruZSoFulPjFLaR3sxUQtLJkZ91McJoR+f+FK0NCrml3Lo
IeIJdGWhvTfLvi4oMKweyYDZ4eqvhMjXxIY7heTlptPxyWRF2w/1WKenC43L6ud9tYOYdSR45Co/
v+9/ZpvffQaT+DJVZTn6Tn289xkzBBZj9K6wv7179FnORRJNyVZ1Z3IpOjgtyGY0Fh8AetiQKwDe
6QjKbJVX+HX2WHgIPfzfa1H940X5eRP+46/GgSxmUM7hakB3DurL4K46XEWgs1IVB3E+hCXp4S76
vcUm5jhdRFg4cF4ugnCDfBJCHUI3FLwkS7e9/FuxqPvc79B9/h8g79rXfOHTiTA/r2ZtPJui0xGf
HIa1lqYO+EvNiSZL0NNIyy6ghJBApMSv7D+/zFGm2WvlKIWilEbZ3zDF0a8W6x/T6rD+Kb0Kug1B
trjzaZMTLM284d6zWjQfMO5oD7FfS1Rma7hE7zHTHG/jWYBYjJN5TK64nlNahsikkpMTdKNxIGkz
p/fL0ARyCOd0T7u7KtIGcGDAD5DSRsD77ZaqGxEWXHoMq00JobMOt0xk2JV9jhPp54dFGoiQjd1V
4U3tMe2xeNTvZWFR7EpFjyjq7tTOGoN4pdqk6HMS92sDY6Vd0YlKgiUsFE2DCFqXwx1lgz+sh0z0
ErXLFyJF0qnZ8I5+nqaRGoUukTmhJbN9cIJDs9Yg0k2Ba8QRANM79y4CtilVWaA8Y4EDJ2Cox1Jc
nHsMi0pUY98iGkEaJI77LpXM97WaznuqgoP57bjHNceUdLvj5ZTfrYP6u3vf7vc7hGJHlS3fN2R3
1s2IwID3C76YUR5QuMA45WJUO5D08Gfc9qgxI1MOgHVu+dh3RQw13OsflkxV73QB4CsBJ0gcOuOs
U22o+JQfG21ovceCDWXQ01FNVpmKs1i5HQFc65E48Lz+gG9mhZfxKJuFR0g4kpT6Cv+oZwY9zhnR
DYYz6mGtxq//rTBLha28tqL9LD4Y0EfYBLYCMOQfxoOC6QQ5u3W9sG8NL87UqhN4lhdE02uWd1Xz
tS2omSOyri1FDSu9JUplbhTZuCVnVWz13u9Q+CmYVZlKsGFEWTsw71+eJ7fU9fFVfHzFogdvAJ1v
MnPsniaBkYMZef6YL/BK963spO4D+cAnEilhr+B6D/ZfvDpEK83WJthxcqXwLTXNOVML37pxkTkX
pIspH/QwV4DyShAI/Nxd1yzH8CgWnSBMj45nruO/9gAtcivPzeZbG8a/BVCkYxu+vyNQzOMmDcyH
bY4PREtiN/TbL0EF1ydHzVX634puv7+765KyzpNVw3gl/wraWK2rnpuD7LJTYgApfy9F43Qp623r
bRrhJt9I9EIfS+Fyqfpe/u7zMQLs2UwVJpWcVf3hjhcpglqp6ofC/0zpkp53SRRFsvoT9AU1nhf7
euC+qei0XodU7PzZDeyZXsbIgZDeZIPoy9GNCVyJQGd1jeP/zbEuJYj4Lv6tUGg/KfRd2fBCt/KG
Lc69Of1dFMz6wK7mY3WfwnRaBHb1ps2Nu893V4IMqvoM63K0wMh5ONorDKLqJQM3pb7gJw59n/yM
2XOR+7RbB9jknU3Dbq4hBiefND0ECbTMbV3OH2rhIF/cVFszbQorW6FumVV3GptdWnGc3YXJQUGJ
+tM2dars3AgrBjk3AjYTnhMngv1Dq0WlsGCQ0dIAUG/KRdhqrGMkZXrR9vy7FMrrD3PDUZekWkc/
3JjkGHRuIWdcFPwkqNMs7fKvjHvoRNWJK/8or9cGiqlVVT8yXeb1LtklImw4Vkgsihaa/40or523
4GzcZ5yi19sqUVUtdmJiDXGWjdGpWFmWZVBHly5UEUNZqQCe9uZZ/X0zCvM9O2aNXARu1tTPo8Xv
vqL4A6YP4EQjGhsFnDCQTmeyos1QzOianUfXpf6XuPUeooXiddyyPxUOFtHSYjwUaMFMjUfsAnvP
wseXwL2/tBbJCRsXzmXP5BC21tvucq4uj5ht9alKvRzXXRQ1A7u2tbvxrT6qp+9evS/rvqPf1goP
LigZWkLsjqMFfvWPIchnZhiDlSSUYoD/Cf40jbBmLJfxXuJDoT0TDdVzfXJLM8nEgt0gWb/Om5GN
TffvHi7G2yhGwk/8DW0m3XNA98fWKxavGtBMms4Hg8jnTIogag2rRTKjyz1CkGJamtsWZTEtYtZM
N1LBlGsJEE+Cym4Th87rZXuBWC6L8ROpnnI2H3MFC47YX8WDK4JbkRhrnR7rHNeN9JvriFm9gXxC
SB2qLduZceyhDBPmofINkmiOsWfR+6R7uPhlvAg3UWXym33ZuHqH+S2CHmpjjLrck92/8s2zCNzb
2xUPtJ+Q3gMtpUGK2vCZ7aHPeM1Ly1bdv9U7134VdRQjLERHNfGFK17eWS/Nyj+OaWKi/zut3aJE
QXJ60LZ/fOGMEqQJdpeO1BY287NF3yTtqQh/56VGXDMJ84i3y2H6c8tfgrbnvDX4jj//7dOGSTfh
3UzP2cA2707k19v6fMgt3E/mJmF4Oo9wYMf/veJSvio/qhhYT2OSQT6XUUJB9xhhAo3YPqL+OQmC
DWlLbEOsBbhFROExyay0HkYWNKNTH6PKjotmH7ZfF2eDk7LH8k5NmKZRHWPbG/khzGaM6ggGyLeA
PgCnVdN5v89TMMg/UbA9EHFWZMViN0TAtryc2zBPMFhJpsGXYJtFDh45f9em3ttXXLbzHi2vETjo
5FKnvngCKyqZWXLsV+jd+FlgPj+3lxp8yCk7D5L+z+wcoxVITFjRxWh52ZAQtqRMbSbEke4Zx8eb
8a8Em9CPTauOLgP0jfsa0ZziOM+DzXwB4inWY9MqbKLysZ1R1YyTi4O2Lqx5QJx8iBX0m7XpUyI/
kOcLRHn+q8vtx3XZLURvHzQdA1c1G4tR+JJkci8vIBls6zyue7+Sm+wV/n2j4ZU8eFkUx9WbSM1C
SN+MisJUeKcfiRYsyNw5cJLes1DuKDLMXHueDWkeaCom8Z+VmMFXE/T6L8S6oT6HyuDdrUerRoiO
RyrkG68AMknDFxGLdS9D8u+LfcuJZ7KdBJ5EDE/zwFzgx+N82EyxQQvzo07p7bzpxzIf89VfK1Tq
dlzObhwBvOx0NRjOQULme3HuwFBXjaRQB16Lm8eiaTPKpNdiVT8+XWYbp8TVW+LgHsVzw9XaowRS
+sKKDeSPfW437eUE3is2uTGFFTCmLNTBJv3TOBTchai8iQh9VCYaFFlgSTABhJ27b4C6SkvUN0go
PdkubT9CQyxTqCkt2FgoQKEXOZ8MWTGWhyOQuYx1r42YEfrc8rDGME22Dgx400SxHQ7CAGlxYrHY
C7+T9seVgDOR7WKSH85Xr7CIkaQv5Yn9QgxiItcFIqDU4M0AIlLbaL/0lnFDtgL52rwZpLKzs1oP
BasVUTKL7wV90lineFMFZPSEPehinwDCXr6EKwD+q6stfnQqKq2+Ms/J7Ho55q7GOuqHLU6BW0XG
Z8rEaqcS/nu9CUUOY32PqoyiESt0T02QxEGMJwG5p6bIjUwIPuUB1/ZdwKGfO9+ReUu0zwHnwjG7
Xv9tX90Te3fiPH6xCX+vM2m0mphpJJV62UrZMtJBO/llRpziR78Ji/j82yNlOeMBJQzW4EXhuNe5
vCgz8wKDFOjdU6Vtg6l3karqjgGZvVxCxuxhJWFuplaS7DbqauSgFyfXz738LFSLJLn7Daa02MTU
yC/yPl/PSGt3NSD1b5z3ekNKO3oe8LCtlCIDzSb0GSgZ9Wi6wHN1iLwHBowWAJ/YGGNpXE6V452w
bCp0snBsTdex7gG3NEp0ArPTqiYCASa+e8ANd7Fwo4YCt/+MP8OaAIa66/llI5gpUnqB6+RJn2dY
0Oe25wK0BZKP7Z/xYa6FM8hyRr07z9xoTbo7IN2kfBNnivjPiHYxobx0Y1G38LoBrZi/3wCDVsBn
m2Ocv50N6We+bow07gq8GjJpGQDEqVydUDW+Jck0OmU8kW1MIWSH8DmhBSSkFzpSteZQO8AKFAEM
ACz9MgUFlu4CQ/Xtm0+IidawdNLnf1/RR0cql9KxtOvoSPSb1TdRQ+F4kY5/4XVoD2S6n7dft63+
VZCWlhbK0vdBr1kWozX8AlAZZCBzIymsMlyu9YYReUsWG5YxPmKYvvX2CFf6PfNC6FdJruYchQ1l
AW6YTUfTGkyxKPzeRLLywVlqXp0FkgINi909UzK3GDkN3K/Ft0HDvHFybykrzVQwTbtp5FBCa8Q2
hdWxNDfDGblSprvKIZcebHlIWGDggtiZP3dVZbEvqlmrbX9kAczTxhTh3P1eY3mmzKb/9OSiYAxb
U7nWFJoEqcv6hfbRawDc0zB86tk5AgmVZqyVOwtrzqzmyDyp5RRhIojcOZYHoVVw9P3zGcZlDy6G
ClF3Acm4QhpgTj9o3cuJjRtJFHUbpOV9Az+qC8hMeRte0DD+RItH0MKq4ri2Iv4yK3gOxOSD2GZc
rdXlgBnGayc4oI9iTecH4Q94TuN0JEXfTPQamndW5UooBMg/V33oyCRDoNPYBBymTnnYMw8ZlH0t
PquLSMbYz3IIjPkIoCXImwkeTeDDtplW63PxojUPDRCi+KNVJV7um9nf7qw+AZNMEC6ZvM+a4CpM
AvWGiIZ4VFGWlyZSWOf3bZlKQ7AfHhIbv03mXd3STu47chncan4BitXl77JbbF0l4K0TCFveHEO+
9uW2sRgzuzO0HERdUFCKchjZw3LYqtjGYvXA7oGuxECbShvSKgl6zdxdU7FcZX/J5FJvbgzFF501
XpUayPvWCr9lBihNVpq65koPUPGwqo8LA7tzWLJeserVRxmw/YL5rU7C7snlX0fXgl9gKdXc+QYM
fqm1+rTUySUvGYEsHUDaDkCFb76E8f68gY7SqVUkBwYlTm5LEra6zRcPYWIgNWaQGo2SwffXekSm
Gc3pnjrnmtEF8XOzmWPhFt81GWUMcqetTkQjUPG4VVvgxlpwsIgC9DWSKCojDpx4SYnwJf2mCWTy
B9qarECtmBBUQBeoIsnVaG7iYWIp3dJ4z4O9ePMNd61Im6HVzsS+grKID/2zaG7h+R3drx6VEb/W
pf6TpJv6cUo/AGVGt4bzendi5wnp/fV/NFk5lMZGMwx4NqDhPyq19IrV+l6gu+5ZQ7FP9xuw0KvH
oTtjGikRMXp9h72IVPk7JtiVLW0dTgjQG0DjapmIxVXQoNzjZy+yxkVMkyt7EXoTzw7WCKcGNssG
DKupCABPdbvNADH2q45V1TdDDuCLS9rfcVWuJWRW1N8vd84RfsgJAy3vPHUhZyGt/OnWVmRSlzHc
7vWUieHaxcCQjEbRj5LTJD/K6gXRElWkUZVJ+A008UxLtPhG+Asfh0AfJF7PFZwJPd9RPkNPsxo6
81f2RfdwIUVVhJffErfI+xAyrWZ7AfVHreRwW08hxM2rGDQNA3fpvg9lEcUpfjDO67I/lJN97rKA
KiLB9G+eaqhLSscGO0KKmPwZL/Wi218Dl73ecrbNLLxtSC5L50ixhArGWMMi7R3eO/vek/pqLKOQ
XMXGTrFzAF0DoiO595yv09ZrJGn+BpGePhsnpsBqwfHwZUJlC/ycZtERDOxHKq+gomOgWqN22elA
3bKz/jLcy7RydM9vXkcyTpzluHq6lEQANrbGMwP+woPZGdAWSi7OBKFnp7nuDJvtapH2cnW1L5FW
Dw1ANDXhZ9kJTn7ZdMmvZOzKji6kmpeq+9Hy1ZMZcPQqd3pF2K5RDCKdJ/+pgweyLIuTmcDntnaw
5ekoeY4ooxeyVvFW++WyLeJCR4jWrDgq9/msD4lqmrhRD9PNAp1DPckhKS1pskx395XY3ixO696Y
R9ZRAL3xBGLbz8XjrKiwzWZKEnqBsdT9SRZ2nAXHYjorynbtVA44kMle9klYG0eJXYEcC56UO4EC
M/FsfhIMPPuD2i+Y/kiKuwdxRg5BpZY25RmlrlpK+KetMlXPMhVOiqzn/jYs0jn/RCxAFkG1J7yy
AzVqBmLpWaqis4nRF2IYpPAQn4dg5DsFoasxyD3+CrOfbkZsVpcb3MXmt0v6bWQEe8JydxT35p6z
3BJc3c3KFXORgYUt4QFZGIJXSeQ676P7mflRmNE9UaRwWNDak6e8uA7+5lPVDWTJ78ZSF+urAXrd
KWI6m13afKoYMCuCRdOD01Q2hxK0Nq2E8tHa0HmN3QbmMbwm+Na055YELkvn3rDVQY3bRL2nkyHi
/BjuCLdGqEpjRXqF2M9n0Z7SX4NVpQhNplIFAT421RMHd7OrAxue2Y48Zyc8SriOp7Jw+0msUw4k
eODwHFOjzrX/yl34gyArXA8oOwG7+v9uFXBYsE7BqgFIVcK/OV/7hwZz1/kGMpftDF8ma9gaTO2T
j2P+mLM7m3eOGK4nWkvS8GuEXNxeZ/QwfEtCXbRNCkZnBXzepVt+ZJkjPxsYZhMTSs8x5VR6ry5h
b80P2FxZi3NynLMhsbkAlwR+3WvgjJQ8Lp0L1+xR4DGha6CPw/L0GrMVwcRYpYmQ/kcJHB8a4Xss
rcoZnn/Kuevno/WHqq3i5E905R0VPsbMT96JAQUouFBfQxGkCCfIKpnw0TWs2CvhO1HLxmRZXBEC
h0PP0SdUa1VDqvvf08tnLhLwVzt+QXUhPQ0J5AXXAQNkobcMmRkOJNM5rDZ6FP5f9cAwQUI8ah8Q
PkS88yYUmL4uYJpOO+CoJhGeGmbGDbAfapji0iFKJJbRtqSe34QLSk8h6cfg7shj7F6N0djlpLnr
K7CGyan/AqgK2rSaJUqc8nspXVDmvtehX9zIMUdWVF78CkDUDlGNCxsWW1IAgl+SBgHVlY8QEQov
kp3DMji4GOCVb/9cJR3aqq4E3LxnCjnWIqPpJA5cd21eQWWAltUVW4WxCYkbMmSpVLTm1Jf6y4so
FOI3tQWEzGrFAnl8QQslie5w0Tj1HQi6uOwpxTWVJzhRxEC2wR9vgdeZyDIhvKTAvtj85N23r2qa
ZMLwFsPep/UzHV+cf8B81zVxBWqafzuIWajyK+Mqqw3W8XztDfBegom5J/QH/3pThAPB9Rql48lV
kaxE5Vy4reDX/9GvrfFcDInzfUGMe8ViCEECYz3LDhHXUajx/NuqUx93HrvtKOmQ0VPgTm1pJ9Iu
4EmpaVsrbSsXPiUvwWX7kPMknia0W+XcHxu5h9NIBU2gnrEu6W8MX6LPSY9TPJS/NvWic2Io49ZR
2X6Gw/nVy0zc7MEq26Y5Jfp+YsIDebrO0lBB4oDEQU2cRSlxawHPTV8QISmiiAhI1WI0CV6Olmf2
9952mHqPU31foDTstC+pfmpuVP0zfiWgYbrWFYkaJ80jgXAIwAHJvknpjR87QeJV1/Uxj9JvP9yh
7XNqW40pYTHVpNzHWDCc9abpKUkMp6MlfDsaLuF3fj7NHtK4a0o+61h8R4v4GIEN/JH8+vFCux+5
ro8q0Dsgl5KotQF3yItDnekN+mjaBh7hLQWrTnxHn3OjeL8r1BkKPsOMtaje1j3tTmgy0D2Vq8td
/XcTO35Pmc4qM8npTOvtut2OTbPc5cwZFkFOhq8cfMumUGgP/lpj8/2SQAnUIjCQCs6cgWMmnXr8
Jf1SrcTB3yNN9cZ23dK8wvbaIViapbPGgHSIz+yGGeehjIUFMJIxIEliwY/hkWCYDrBTZDYVr+Ri
O3zQS1/297ejjNeCdZNZb1atUjVzfz48NuCd64WrRSr0d2g79hry/gox3Z6+9hZmFLW3Jad8pxH6
GXoPddiOZjNTfN8Acjo3zOWl5O6oHRXKVRydnV59yavUupluswfCEyeS+ZLb76F/tDh+v1TQa6YJ
H/OBvQqCr953Wme4Hx3Fr+WJQZxoh0mJsb/NNlC65JFjRDajnQ3QNyDx98TUtydBW5lMB/KJ6Ec2
4hOuy6YIZYSrbzUKTxs77aabIedLrZa2G7ME7DK38bulPvI4EbQBsTsAuZwpbx2hdlkfZ+ZCgWuM
K1Q1fDQT2oypavo5s3/+B18smV28bEFcqPSrizgDicbmMIcFmE5ZHcK2CCPxdtMP/81YaacccPFB
VyowMd929M8vMSNF1Pt3xz+r8v+tY8yv0NtU08x+Ov4KWf4uoKj6U2v0is1AtoUly7Dhfs+ZFcj0
8udT8eShRvQ0WMdT8N5CduvJR8QN4oJzOIJrMciHpn8wISJrhFs1HL8vS7ax1NjBwANbz9IzIT7K
pmnoGfG3KFsXvwxbZTWLfdppAyNIhDWmkvA4/lFrIZwefsP0Ar5Rz+vBdCDrjqbtZwOEwVxTcSCM
ijhR87qepmmevh2p9GML/7kaIucm5AUjqwAVaZPmLmNkFe2BGqtJ3NMVvjpJKBdnIKaiDwiLvCnI
OPQ+YUWiJQgITqqhqDwWRfzmGXeh8EjLx+Y2mjOqE7DFzkhD1x17bjCf1Zs2260eOsesp8jAELRx
4u6jynkKz4mzAFcnzDYD1rjf/hSnEGQ49DhR2TVz0vE1zU2t4NSgPT1cUfsvf/zG2MhkeiBy1fw8
oFbl7Q4mpmwnMXDlW2e0oF5MKNktc8k1CNROg5VHlZ5X9gQYy6Qp+hIvv0XyxGV9zuWGW76IELIW
r4t7wzHr8WX7CoU/iV8FPrdo8URob1K5MlISdp7yNAah6nyEZWxuL6RH2a/4oe0ySi+4bqFma0Tm
uABlDby05p7VZr3NVG4m6P4RXBhKQSZ0jCHdwgG04K14gSlu362KyMBCiXaoA1FxB4U9c/7X+GIk
W3/GcC7yyqejFcScn/7Ym2VO9Qmy+bFBRmYaL1blk8dmVCEPssy31Cd2sbS5Odz3XRdfDVk2exuL
/VaDGQfIFs7K7yGQwi6bECl2FCD3sYA31lps/vrw4yp9KnjOuqeudnX4iQLSIFXOlL73gSnyqtZW
Ksv4wumakMYQbJ89Hi+9N8uZOUS+asHCFKUhZjCKMh8p+dmcporXppJHjvaLte6C/A09UXE9cb4j
FULktDeRb5qqTHqHJLOZI9zrfXUhTUyo76FWg21yqV4Dn2CFHRFdHZYwcJZdq7+St2m0d2m3ypb8
ijR+a5f02pZgdCWlsdULgLH0Wa5v3wuBvTGUTGhIV8/uh/nrgcRCYFOnw1lPxxLGm/APkE2uLUWY
m12D9Jie3G0v7+qjLNvUxTLap/cQdxtI46fExcrkZKa2Uz7/x+aeq4zkEHRk7EiUkhI7fBblAkG7
BEjvAUeBUo717b4mV+66CBTctdDF8ju9Q7+hE56Nnxw2t6jcxNef7kTKZtAwy0X7gmGH5g7MNmjt
kCJZxru6WrO+4NrmybkeDNuoqcCTMl3s6xdF4yn9nuPbjfszy0IFcJqNwqjcISTZWSyP8482z46O
P3stwPAtepKXMsfjlWCFIcpFL8wzV1Bs9yCPJ62Un5v+Q7QFiT2IC/+/kdmehUFjltyHtNUczqKq
X5OBEqRFLsBw5uVPCbjOhy3G7auMhW4STas/76Tjwmyj4SEWofRt/CLszernpDkEvCFRcnWsbxzn
7SnbmZz06kPwE0OI9nvjeoTB+88OIBgpMXQ95BijUTOEGKUw6IysJCG1YUEI09NmY+klElIwhkWQ
WV4P3WK8KmpJQx5LsZcLFv0kUPPoBQT5IskrnzY1iTcq/vICtUerELLKj/3KfkLBIQ/JMIaukcgk
1tW0lyupywEIlTiVamLpCVkEKOcXLZ9qySJo1/46gl0vYSlNkcjf3RkdXx0YwU7hUa0C7YvbRZdA
PpI7x/Mwxn1WF4lbvQQithC0JgtmQT/gsUS3VL/2uH8lfL2t3YnEi0yWsffXLwoCbDNrSeoP8RAO
8zLzfvDeSdhszFRHA9/BfV5qgqdv8cl2PN55VHd1dnWtNEn/iMaL6VJFXGo4DhUeA7meu6KnRgRW
zchULCrOM4fGXWdUoNGddd62ennexY0G58RvnyCKqBR6CDJV0YdTMMKAkM3/5HtBzF+KEQzWHLhd
OyI01lj3u2nBuwxuRAqHvRJOqqbnS6sEpDIb2LXz3agc5XWaZONW/fecWf9ngaLrJxf1CteC44Vj
wMoEowx9qU8sFaWiP6gDp4Q/fNL06Fss7O8fEmDuVOxQJnp4EMjcU8/q91bUfvIBUajatwqjRsxO
kmGIk1bVIiICGjtC5tEDS5DjXUETFdBD2kg2b0aQUUEqmLt7tWU815+JsutnnjBrln3y84gd9X31
k2UrSqmpNmyy7wpcNaK0dryU3sEvSbMQqc9ZTg6fmEKpO887CaH37N7jsq3rsDtizk7je0rzPpop
jdsZYhQtaI0Uj3VEkk58NFiUBB08YdMi4hrEVXfPOD6p6Day6qvI0NJ2ylxqlt8xDo0l4B9BwO72
4rKGPaErXgjrCETqemfR1ikkTsgU1MJS25/PDg4ix5pR8BUYhnGgKzr8kxUzldV3MX9a/o6CXbb+
THrFYxzCAGOl3R3Md7JQpitT/rr7AS0kMPnKCLVOCthYzxf38+D553FbhK6XKYDZvRr+4e6uE9cJ
WVNJPi3TrKBlL1Dco8Jz/GgQ5IKmR92lRPmPzC3Mf11lXnKXcWbCWnx4IupQFudMAuqM7FQT9m+2
eq8+dP7o9C6lczFXAoIGSZ9Z2LyfzbU5r4ngweZIJc6OqQ9qLdaOLM2mRIah7Sv+dVnP4EZNY3gk
Yv0OVTNYWGAWWNNJJiDSL6N6BK8VywJ8f+UVCyuWWiRQEOgfoVStIinSBTwENuPFsF7xgP74Wgd1
a+h/7O9PJAX1yTkiPpyzlMdH9MvqyDoEvOf9QbMwAOobMyceKA3uy3SIxzlX/TwktzV1HFArIC3F
iC9Vmhlzq1yi1g9ToPGtwD0g7RTj4zVXqmx8GcjZhbC1EX3cfBm8q07C39UKIuOJ6LOyT+20azps
GKFEOlGqYPt9QFhn3NOG2hbD6zjUjNRGFf5rZ6lFj7VGTqVYQjJxJrohjYMbCL9kIMn/bYRWdxYa
4luDZ00zjJHAuvBMEtOMBWHjyLayyeoPR84bFHGsFmFdGj8IB5ULcImbRICfo28eRvG3mTx8Nn3F
rgXgG5+lqd7gXxqtcekgqA72eNHwDqUNhjJixWL8MV9/Q+w/hhLx+wGZsvQGaF+Tf06gGEIZd9AQ
HYwHvQS/lzWpPBhu6PZ0t/zckplqcncDAmqUITLTUEN41vau1fkBfI5XW4kPlD9ruKP1dUDATFCU
kyohMUj0zzQ6+fTRPmcmyS9x+58UQElGwBbiHj1okY+KpdBxKGkGzkLAZaf8gyJFRwSEHtl8ih17
RC+beEjdvsEgauK2IAiPfXdi/lKcOA/AUdU3SuirysD8c7EA1gt1KUhkCLdBBkI3tQM/xbh90Vk+
rOaTPIH8fv8eBwYO0JiBSaxchyUoyPlPFQMdK842sVRYtJZdUKF09D8fYsxFL9FQ65ctEvMAKu1s
y1stSSDDrl92MV5sshVlIXD+sXq15wLC3J1X5SHl9agbrM4rMCGiWPInn0VCxOhRs76QMarm12Dd
8A2mPlSnDGsjWeFSMGiM/jRBRhq7TaeUuM/w9mw79iP6V13Nq2XvuUSbfX3S6DC5M7dZsquZBe/q
DycniBT2LgbfPDE/yKHEppt4w32yiwm3i5ewHkoUxw7EIaSsikdC2rdGVY5LR3k7z5wUqQSQ6cBH
MhYBGrv3+M6G6LJaeWLKHFFah4ZMHqgkNX6jAd/1DsySB+OevApgu6KujPhYCB69fClEOsabe5Ar
dNjHSlJvLw8mmKUDg4/r4ukuA3Ag3QSM91hBp54+45gC/+HILJwdre3QeoZWTkgVm8BKVK4piTmo
abq6ymRL9MXGCtwnpa7qTT5am3smYeMYKMLUeEc8e/i4bSMubdtK4fC8e40HEcSZIe5Q4LjuWCVC
bhNvCc4XS/IGZLZEeX7A1XChAC3jsg+3+yt/0zXDw4y4nnOH0FoFbkbktcvSrnvG7RytkISskEWs
hILTjhbaVKaNI1veCx0R8oBzE3cTjJnPMbTHQKVs+Lcs1CKRjkBwJ4W9l/muPH5Kn/FMKHdeZ5ZH
rLj0xOK75m9fQTH1GJzpum7iwbmZflHLqw4to3ML7esu324wAm6mzTqU/T4aMvGGwjqM/b4w7/Wn
52dosJhqkmmntIPU+48uDWlmLOZjIPbkmr4UM0U3joVTOufiW1wxPdwLsMFW7NQIrGustecoi7cm
kxAP8RxCXqgkPxojG5hbFSLq1gYcNz0IiOF93twiSU+nuwv5H58K9zpdir9UCJu93cXntHukOlkK
yzriQ6T8xsqokO+ukC1J0aV4KCgkw058c2BMc9hvZKNd2MGpgMXUUlCvZDjVO6/YwqTZN4YuG4Yz
H2IYsnllAFtXbJ1ksvQCvp69nuWdqvb1+jqP4IeIbkBl8COIE2AFnXuqXWAczNLMVal/MdbXd16m
TFRYRytLNLqJIq/M5zpz0S0w2RAEZNGjnL5XDZjwcQVPaOEYeubP1VnQVmNFyuOioDvyc2b55ckw
mNNOS5ZOoUeCFwKafAJDK2pNvbDgje7EsW6z8e271rhoEacQ8Qw5jj/k5lxkaHCxLP3qAQUyq0s9
SlWCIxBN0X9uywGQvS1N+5XNU0pAwTKOhx2HxbCIKEKY6jIYGMEnPYFMvmjHaJdsAfLWX9dwTumG
8XSfqJI97o8P0NVFx8GsnwF15v8s1R7DTAqjyAdLHckyT9K+tTIYRRmQ6ZI2c3BYbjh86TRDSags
S/8VC/OWRt0YzZ+glKDpTJUqPoZhaNx1QAN8/RLeMgHvE0KKwfqGMdBrBC4uoA7KF3CT+NuFxjrq
PMNmiavqWHtTVR4DlqxfBAtkShgyNjmFMqSvzBP/6F20POuRs6szCWAnOiQMKrRUTjtt6yG8CV7M
jJoFfNTidfKwxJv1rT22kmlroqjNERJvu5/so6QZse7H9Q4hsA5YfnOi7ElzvdKojeAdCWLbVucO
Kr2pYyt8Ph3iPz9ORmlEGlYj/51Qfn0iR/pBc+Xp0fqT6XRSoyV23ELI8V1SIS+FWw3lkoXjedKp
SKsvbyh/iNw1GQXpbTOikQqimyEvy++iUeXkcmP40ErnskU7CHjYj98OJOLUBTyQTbxvs5tc4zJG
a13dfwinmyBAKkl/jJZtoBKWYmjnp4CBFb6gUEZHZtGFnVukLXmK6fv6z3m9sEW/ThpvE5OhEyp/
tIf896z8EMREhJjQuadnYlWTA0m5gdGlxizeDpQRCRUq+1WTeCYeBKWVKu/edn6dx5ufH4cXRqMB
0EvPjJCi7tO4smJdqM3NSXQ2PXwY/E//zCN9e5Ar+VBaMIo0NWSo9tpOC4a8jAhKhsfDEjA1LrVp
nL9d+pVfH/TTA0VIqcPE6usGShAt3A3HY00pUwGq1lgxx93XlYRfMnUtZNxxjAjn5wY76AHWg2p0
l0Yj9Cin+kzK/N+6an2xIK0scw5EvjXJsnIhUoNFLt9x9AgA0WGddnRmzGDnandTmRX0IMaKxt4D
hX9eLRj9jSNGetsBZ++GfWHw7it3kNMcvAfhMCPcedM7IAZT3jpSzWHWcrsJ/kDWASUIJ0HYYVlO
VmiG9Zwm1LgaSdQwMOc9Ma6iIXJeD4bKQFlVsEJUZmbJkguc1CeiWo/NuT+FzatsfnkiMVXhIbJ3
inrK5+jdZr2BOiMQGgK4+Wh6j33x0kMHh/1syI3T8zAW64vXiuYc2mDGImeJNv+wmN1xpYK1xA7C
moYFeCNj8wAfYe7S7qqFcfyDPvKHOc/Tnpr1MmANA6Obdr7BIbRFr5xI0XrrOWy9pfkIwZjuLhaR
lC1lR11vjvSP0jI4aMPkSK8HX2POMrj8Bv7IrYl91Nsitg4npdX13RBAumm32/9Yq06+e1j79owx
AMfVX0N0epK90O30VDSZsTvOP8dDYPDvxtHWNdP6E+y/7neJFA/AOKjB/Ob7KVZeCKGpQ2P56rq8
d3mdbL7JFPnE0HHaxlij9zm3WUF6ZdjP/Wqj4MHiMgek18wKUDIt7xoF8bMj5XjlX2W5dtLz1AZ3
1SEErRd4MuYJ73ubSyORAxPbcdywt7igpdHHe8oyLFEAl9Le8qh0iyG1zlVBLqfawMASsiOEBY8O
LQy0KtFS9o1ws+YBb74Es+jVedvY13xgtZ2xzZ3SxSM34p+MVmZlDu6k7WBsz7qhYaeoTfMYOsBS
uyebkxAVAtUSkN0WQ1AbmoFfNY3vY48qv7sDHcu8Q+7pMr/JrwziO4LsOVzQzBqNtUhW0lUOzC1d
QbiRI/fEoQgTxZ9XkOwxiQNRdai+Y5TI5K2E5u03Rmiu4SmJwfaQXVvKpqEXLWW6lLsWayxwbelv
t485VPcb5zagBXdScwYi5uphsc/cjwuYfV1i47YNazT/nGul4o5CKZBkpjkdAHChEmcM3WDNL7nM
bWZjdJuDUT+zjaE3/od686l4Xtp8QdaQge5n6y/4FLVwt1Ef4Seb+zSaZP/6rQeIudCGMwPX7Yec
2ywjKSL4wCRAsgj7umsFcQ5VQpjUY07XiyyA6HDq3beUBIieqF9WMKxX7GzbykNZqrI9c4u8SNiB
9JvdkV+uEnZ20ouCGNEHAsJ1Z8kwyS4xvoRUBXMOXje1GMebkzdXJ9b9hYveyHSLO7IC0mAoHn7b
nyBrj5Sx0CK/+e+J9ArVnHfjSw+wYv6CsWXZa45mZmmmVq3BV9tedC2eaonaWp0mgI5qMsoYJDHq
CYvKRDeQOnoEQygNdPcv5x+fiPju8IvMrng0annKEagNJwrg2Aw2GK5M4HrXi4UReJtlRCkkWCwv
IDpNymHVm4+Hpm1ftK7J9isSwImWUlczZ9gmBW08b8WAJBR2eaO3/sXlhUiF0lS/LS1NBi51rqub
igty62xh8d0rCrXtW9Kdol3MzG2QXcAsAEoBwJDLm7jt6Lh/CFIYYGRdfMsgZhIWwM6KB6IRFSRI
tyNz69QuoJv06lBRWM2JwyZofD1jg+oC9Hg158e+CvBUzLOh2/9YJLxYF+EWma5qWPIlCSWA0cGQ
GkFn+Jlz+PkLNrExaikCTkoIGa5C6G5vqa2y0kCNZ3t+T/WrSCg0PVK3tut/MDh7Hlc7lDgNn0ec
LPFztWNqxwCG6TpWpIThTesgY5VFSu0D5LPc4V4J9NlfcNn1vw2ud034vzFTWAzDpQ9wp/MLtZiZ
flz5yGQg5B7iFXxYgxaFFFmzI43uSjF+NVizzJWG9M2NRVt3v1v5Rkf18U/L5q6iyFtl6prjP4r3
w6U/UCEGfAFZ8HvHzjTbb0XqbszMkZdKtA4KrE46+Z/l7L4EDj3lJ1r3kF0Zo1N8UMc7RN2N45cb
RYzs98QpxkHDoydYAQ766HD4q5E/mVK7Qu8BtMaqPWiXmTT4SY/xNDRyUnZ0U+ZsgodAgIKghHOc
ZgP3z6Yaq6XIyo9mEjS8fwi13MODC5NzCHk6k7krQ6K4ztggAFenX7WCipRwwsXrURbJvkXbPGkg
CtO9y3mDzk9zslAZjyKGPbTOJuXFlsHs+CpSO71453OOuW3n8fNN8fgpbH4g+a49hvLDS5T7qf6J
DJSSvLBqvypz+WfPJcYYKHViivFFsLBshPNegO881z7YoMDYAYieht3eFEtEwzDKpMP3U8mjR0yz
90dmf5wYlNtz9FF8dC13JYJSxlSE2e3fuHqM5HvJe5Gic7GIeruaFD8LVeEd/TQNOOXLU0ILmntc
LMGr4Dt/CNsyPXZMxmPA72UFbs8bBXptBIUFt+Hjfkesaho464pUS+W0SyptEhrKVO/bxn34WNe2
BB6zY0V83MRsSXwWdEJEHzMuX/1Y2ArDzwaQoin1MJaocs0cWRp7h8IEOXfVpQmXUoL9QwvAL1U6
GaiX4hLzSWzpUnpe41aR8dhkBcgEAlASt8RTdODSWPubkhvEjKDUdFUd/+/6z75mkWR35y443rUr
25qbd7xDxyPqFWBQ1+odhhaWi5DzUUft1yciFeCCu/HN/lQFz2egGumzJkAS3+iwaGwUw2spysZ6
zS4hDKefNeiH3dLhxzYStgpArvP+10AhYn5itLmU+sNbtVTiRGlmnM1xLPoULxaIvKZIrKlJqLb7
DE1En9MDcd4YKsyKoIDdQoUDuoILiSxYuu2tEWTvXy0TpjZ89xpfvEbVgn9Mt1umoJqZQc8EdOua
wUh1WayhtVeOjD6iubrdswiV9IjgBf+uNOfl354ZAoI6hDCnVt1yOrM7v9xA0FhjI3rzJFLDwvLR
ILqpwb2DnR0cgA8eAH2u0+cLwzwd0iPi9sFkCfO9ZlYqeRjfIlfbmtxawkji3JXljSFypQjqY8n9
IlHdt7Ufdc/DWJ6qwA0Sv0ZMHhINlQ11hvWx7g4RC0/r4Z03lBCMDyKGsuDzb9fIgwq3Fuy+o8Os
OGpAAvk4eGQ81mbUwk7WDeGGgREEFYS9t+xC98xZ0wiTGBgxDadY5jzaAVnkQa/hq7W0xhN5rHFk
bWCj6IyqER202fEHu3cXiXt5piitS4OJjNJ++lP9wBY6BJ44/C8lCcVAof9xlDXbpIqfgUdVnwLl
EtG3T3nGegFqHtXYKFJO/OdXOA+rJO9aXXPCvYTabUJdIZ7QirAGRjVBepJRVtv0HtKfkTdYvJN5
l3ZGTLmd9CwYIk734lrE9IJ29LfUEtSc8bT6axefABGPOdDXaGA/IPwHOSBJMfB6SX1Kp/AZH111
kS7zwcMbzJB8MbRnQRK5BO0/zxhMBSnLCTSurZ9/187fl372A6By+EHMKsrxAXyPpVs0ccPR+oax
sjJbQSYTVMsEgu054s92jJ2AQ+XeyzRdikPOMzFo+1EN9aXowegnap6kxE1Hj32UY2ew7taDlPk7
2EEm5PbeLB/sMu7fI0nLJDskcRz7yMOZ9kXQwPByOGLG03otiV7eqa/bHtIzG6yrOZieWyqEmewc
nczISegh5oo7oos3Ft4xEyMUBHjr9vW8ZtEcD9df4Yhoagv7PYWSDbwU+tQ9lrRcv7RshmmVYAZw
g1cXWB8i4+ZTLIt7r8Q2EakVm5OoY6n/AinPljHv55oMWAEhY9f9vXgyBEFJnywnx1wAh+q7I8N5
C+Oi2uOXmjcFtIqjGfOp6mdWId8n27BmgBQ7gbszgpH3jFoG/uK7a6Gj4F3qJRxXi+Y0kSwmc91b
M9jXhF0ktSkOOIyGHqX9zHL39ut+uL4XcxdETq+mrPlo6gSKsDNv1FQ8K5V4fEAf4xu4nK5FuSgr
mioe0QywnUnOr4zHW+4E/YWJrdtct7vsjI7M78g/ytwPeFo++0+kGuuXbgUT0GvN9QZWM4EUyjbs
O8dOVDsNAixw2G+3UzZt79di3rM7ymsw2pbE+bEeYSBeJWaKrMybbQO8OEL2nXa22SgQP2nt0j71
YGBSep6PV51w3QEkKrznyZMbifoWDcmhNygiV8C3fIeaLLnVeAL7vxGxyd1abHXI5Q4E5/SSNh2O
fACSbLSet6D8PBUT8lR01d0eeHm0UU/gBgg/fvCaDC+SlYMlq9flXBXpGlQDnEKrvQCRmiMBWyCH
cpLMc6/lpB12bsC50EiDLLeSyisMnKga1BX4h0PQhAL9FhGvt3oQB1HMofXiijREMv+wxJ9REGdD
OupUqC4lFusbCqaoWv/nPXqHYCJXKxMOQN92e20XlXHgQjsSyqk0t2+qk7YCDs6QEehmJiR3GNL/
LkPD7K+GzAnCyI4YQJkze1IsU5U2maREmXPTVbTOiVlUsZ0elp6raPb9lpa8u+WnK8/A4Zf4lxT+
7qVqb2rKfxY2RIQkgkk8lo44t1SHgRRyk7O99zT1iC1ujJTHccFXpgxJcxKyU7YPm9aXGu+N67fU
CQ3j/Rya+wEyn3hV8JIUEp08+DXVd9s5/uhFvoOr7gBWyQIcaeMFAaN7vsgxJO17pAvsQJWyc0Vw
n+c31i1FnXuF+JcB7UPH4kaRbcHl4NlLNVFD2GWmgqGWybAmkIFskli5lbG4JQqCPW93m1JCmpcL
OV/btyk5alD7mgtdESBa1s/mr3c6SHajG2K9F8HVyquxGLNrmnGxvoj4NeiorK2v0diB5h9r9LdY
jWGUD0NEGACvC3YgDs5uaT5sFBb3S3vy2mWby1paCUmitihmHRcgl/2Zb5JIbUBuVfc9cEy+dvPr
Ur8B7L0d2XpEuIkr4OtrVdZJaYgsrABMU8TFelfl4KY/0Z+z+hKA4ZIU6WZ6xyHbzBHV2VmyQdC9
DojzBmEosjB62LJ10eCn5R+ZsdEaQV82u5CRermeRrTa722ADb6QHYBvUFvH0dTOr/cxXMGH/TTw
2g6cyXkHAs3EiacQGEA1clcniIuQoX7x1fDKIqskV71/RF6H4pHSLRCN4PL6TYz1ZI0bBCRqFWhV
BFcWLM2Z2typGOORdj/mImVH/PfHuwnZrG03VTPNQfqXj8FzSHKupOx/517SjiQUetFifpOU7ty9
+r8Slqr4+y0jSwVlRnUhalSoeBXnXbhEwo/fG9dbOSuDt6+czyeUDR9P2tamhYZuPjm+jhpWmucM
CPv9pFxz2psLklT3HcuU0aI9+kc1649hyugLnvf3VsjY79UW3GNLwzZkkjFMeTXP2zX0iZ6fuR4S
pWwjVIeY7X8UKxMTjZCcarm7R61Pf9fS7Zhrp3SyAxao1r+WVT7LR2P8k2QY6yi10m2xQTgTVuJl
rk4d3e8ooNpQaCYKnBn0iVXf9OQuYNNNWt9JYLgN0Li55loL90NxOupNQh65c9BKvjvz+j7nWFkf
Z3oxdWwawKkzokRJZ2W0BU3+NRUCX2I6gFWf2jxymdb8LMHe8rEZ4xEgpQONxb8ViSw3xsk6M5o8
DDpJ0lZM0kQqRQ08e1hRm/EecQF9T89da6TTHS/okESYRheqyekGg/HBGzqBKpzaIXwp3xspusRY
EQX+nKh1m1rpEXXhJ9hf6IU8VZK3+J5viHyrpbyCPK8e65brgVG4oTZlBbQIsnt/Dzny9/+v9buW
b6x85ZuaxsIEs+afv6GvkzMcX++wHxqBr/qcuaIBPLyLJDnkNCLQyeBrrfE29craETE2XV4M2qeH
It8lP90dKmAPkegiPOknvLsOgIRSs/clE2gVkXnvXiw4EALiCdnOhz/9SjqXRA3DXOe5dhod+Oce
HgmOlBQW2htLpqCSzUHYrups7AOkrHlLI30TowePTlJUPSgBVhwaQ/6A4z+raiiTJ+bLAU6SU5Lo
Uf0eGvfsFes2BQgNEuevHsCTtccqccdOrrhsgn/sXKqK3UfsLByip2AapCVosNAgqcj2Vx3ff2IE
mn0GL28ZSwENFt/ZGqtE6UR/7KxT4Mk46VzEG5VgHSMgK7GqtQlWUlLmZCcYySuhxCpF6GCUbnSW
hHumBRu7kTSEwOf0u7DG2gG2CKpq4SVswZGbB7NkRGNb8Gp7C7/aP1qXlsRE7kEwMV+Q22z62kjG
+19xjT4sKZneZJMoFzA6/Mzp55zrBntETaaY3mvJhy9tFuR+ueB8e7RPGl8qkaDKJSBOXVn4UrEL
NJxC8lJg1wZnsot+hLWolbOhmCr4vZtBnJY1xtaMX39VJw/zgBR4PvHYdLx8S6U5XWG3ppLVzBrX
SGpWZIuZA574n3SyawR/erUrXEnzrzMTjTdUSeoQYYpXykXWp1TTXgq2mXCn2qv1eMvmQuydZiM6
wSRInR3jBe33I2kNMCx21ANhQbJlaAVgoB/LMUVL/iokluPSjZ7ouRmv9+mQ+HoeC5prjHMTj4eA
CIdZxV4yl9/krpbeAmt//KJnsAlfLbD7yB0c8TTicOvkl6mcNb1um0HQEyukdLHawBruSQuZlfkB
jh+2XxTFeAqfzFusoecvI8Ge7glybrAfNTLIJ1s4sb01+6m6eqVn9lhXs9OVNNcwsKBCFkCWnTLm
8BEqKcHrwJE4ZEqSF51/+d3GScVMUtare9/voSE3CUSLjsCQjn55hnpUtkOAwDalGzgyvMbOWenS
jz+L9hJKHiLnEC4c6Hev8uYwbIQh6zVxb+bHrDnLgFvMhlYjKNjG5r8UbMNEdhRT/kBKqvRLDdA1
epoWtySTuaDLt7h7vDjKaDzvdqBGAoMwmxPxQBxl4VQ6CeNrLI9ufI2x3ToCdBiudsGxQf1+kX3U
OIh18B5Tcs7KvctqpOXkO6AIk0/dxxY4CpjURxIfSAbf0C3+pRFyp2eTcLVzXI68NZc4ml06QMmk
S9oUGNEELuk7GQRsf9d7hWD7npWzzLcWIzsrYeG2zBoImKfUroe43cfAkJIF/s2BD/IHUdfPC3mN
kPafVSUJxKUI0ucsskmOd/I6dooXeNdCn9td54Vj19H9AgtoIYNimksfqILV28wxMQdqT21gZ0ds
ygvM6Gegt2ElCVH5CCmdZWtV+uTMRw1GLeOkQm4A9w1x9FB5Xmb+aMkF3ojiL6amiBHZL3rtWx8N
3pL/oa/KZ40nUa8T6UjudTv08KDjQyMj+NbnjN3l/IlIT2kEYy8M3PKCHLwH9a3lCIPI/8xpSc+4
cjpQSye0GmeBXKtuAmBCe54wx04UvCgZOllG/5j6Erj0Q6C2krdkAOIDaBZgqOQl4QUtHFXx93L6
A8o3sKSfPXk77ZWJt96cIJM/TRF0evQYhSnf++0EAOXIRl4oBaRnYqkymuuOolFTopdRrJAxxmsB
iCHpygS3CaGV17ePU8ajoj4gj9HU/1hZJjmPFfwweKbwWECrxILzbQHPmSKiL810bb8pe1iDB4m1
XI2YkCaSoOVkPeAbwBpbbcl8N4tONHTCRcghrgXVFgpJgdqs+ZU6cDbvasWWmZNuAEQf93cwsN/1
LM3FIO+zc3ECmSSnz6q9MWg+di+AFC4I1gTN6ueXPIJ6bPEEtSXFP1a9FApdabqtqtjknb9gq8/X
o/zz/v+EYLUKkwEUF7braKjSTKNMFAadx4shS4OARrz1pfRHu29JgETnxbrcXfv33GN2piOs06XR
XiOzOM9oFv8eXZX1jusHh3lKemv7kBX1GiSBtkyJrFShDSdrhS4s/965JxPSzIMAT6eJPeWYv4aA
0X7SA65aezyP7CqLLp0QbozVUTeU3iaZzCdfTjn11ynNzCOjHTt5zzbbeTt3ArEQF25XQGs/4phH
ITS8BsJQFjORoxN0++qD+C1WSBbvl8UI4ocCRF218QB5W95GMtMHtDi5O22DeFzo4qCv3QqZ/pKA
iYeITm2+PVjPaGUwhf6wvIagVQm8x5VdO28qKED3Lh8Ks99fqob9jo9c3V/OEL5An/rlb+Ym2I49
6Az5NQ+um8Da9RSQ8u1fa1QuAgU9d0B3fGrBN7h+V2jbbnNcNWRanfYgnMBMr+j6HDUJ8MRjbZHR
c6c7lSZsTQJbOfpAol2UITW9bTAz7z/yCVqPLKSSO+O+ofu+V84mjeFcTJxxqTKZfc91vZR6c8sf
ovWxAqwcJgZ2fhQwwGOmvcHWVx3aD7y3fAB+fMzpmRBEy/FCYPk6dCEWeK4PJazR6eyg/Xpy6ELO
k8XcVSkPG2pzBQuQJxfOUkaozDoVRZ0mi/a41UV9rPjBblNVhP3ZalqDGqbJRzVTn1Vhc7YMpwG6
DocvdaZ6U4v5pGvMQ85atJCHbAGchzdrKMN/lyaqPgGa9kYNaDaN6tk0eJ5351rE/7/vv4eL0Q/u
UmQwIzl47C97XlZOXTTMvrhVP7H5fU8VdK8/WbZAp3JN1lF3+ZMLVTvEW+vog2jh6wNH3aIOS8ju
+V14E3uYk8sC1XyKMLfzIBwsaXsQjd1+I97srKCh1b2s5puwwPTWXdThnTX+I/BtKf5+rDFNiG0z
hxdv0y4X+ImVwYIVjZMVGyakMyxhLDvvZYyOlhyOJOxV9mCKTtVIWxNNu4I6wOYWUpQkLUhwXjmW
C8uzE9rkHjxTvYPC2yXrDgYbXOCfit6C4vJTFR6NmrLGk2W/xMmV4KL28hXF8ytwVcXFdJiFWgST
MPk986Yjp9G4EfUdqvJrnOQk80KvdybFuiqsBA4RKrjckXFNNjIckheSuxc/97EI9ZXYBLJeJwor
2w1jaMm5tVKQxdf9OFSVMfv3dvj3M2hl1nloHqElazFLw02WsCBFjPUbc3Bu73eW+zzlOYFtQnS+
mlYD3jYI+xL+z7rJOP0OcBooVcVyKwGOS0vMUordVblR7Y6Lp5bIkkfO+NE9I/WyfZrF3pyf64XV
3wMZIQEO5kDyjnjzUZMPiULbO0dvsZ/ItUsT/qCITus1hwJ0tMeTjz2e9vd5D2NKoaTIbOqRtb/d
HrpcYZ0DGJTW8BeLvMvEpD1JuiLHTK1AacXRhKFL9g9bDXwflnWJdjauVxpoZAYHdZFZUkMV2M8l
mkIOgSHogX/mg77BrEKRY0KLjkJzDqkghU2fvgJzbtFS5GRSVUx8Kln2qENqID+wfWSzUWKnbN2m
9hDZJBJpYVBHX4o7eRNEJ6cIqd6+5FNiCgrn5deLFpsgSigIV/siJWMOa2nTy22IvUv6KpsH+mq+
48bC0JxIe3cqciYPQpMbLHyn11rxGRUA3FJVdS0CuIAzcIu51fWuc8nonvbtppzkV2EL0M9vSzIl
+5rwOpMH8mYv163NrIZUTjyeC85gs3CTHo8Kc7IZZN3CrAJ/R3DLxkrj7Qnr80Xv2xPmWzlOP7gS
+t3Izk6dhH13LKYo6iY/lSGFMFFfaIAmV20bWQFmLYgPPNP/ha93b/zFTUEVvaUTHoQes3jEN4Di
fBDC+xTEbxDi/NlphiWLCR0NAX/cXQ1jF5+hqAPi4XwKO1tb/asuyVCBR3EInEKrIVuPo29VTwhS
rIRQdyceCpKOitvL5PzRxa59ABjac/wmjf0IPVOgwZFoO2PYiyMucp25UxDR5U8K+ZdkxdwWsE0d
dUl4U3CJNNFNlJw2lmZwRa6pKdprdwcu9bYRArnyan5l6xvge+g2Jiq8dapM4tFsrjRLzeNznPGQ
jOk0m1IrZJAult6+ysE/dLD8qV01wx7+/pFWk6jkXxs+J4kfoqfiB3VLiCS6zN3fxyDHNgjwFVGx
pXMwQPnBsrCdz2ntTgKGPpxZOOQb83aoWUKVrqiYeqcZLQ2cUHX/uCGo/LE8es0JHiWW+/dfX3jy
VHDIJzm0/zXeY76RrQHLwmWWFc/sdZju+veJvlG1z24Y+IHAyW+7XtT39IvRA5PNTsdjD4XZJaqa
QcOsAZGbDZyPJG6fCSThugf6jpcuWuBves5CZZptu70c1OhVWKjUWaA48ha+IRd4GnmIQDRhlg4K
xj51q6aQfOeSarqBL8EhJi54/6UJfiSjxBaoljgj1Tlbly3YfL+aWH3e0suV1KQsKnVnnOU6zC4q
BHf7kmcWzXxRJO5BLGdmcyF4f7RSZoPDwADR3pToDSBK0Naar4i+oHrRbPQtL5yIL2laUhyfbpfa
REErbTsjqRlWK5Oo9SHu8FIfSAVo0kfdvntdCsBCab8UWecAYeqEmDYUbl5/DwXHDnzs8O+DWcEq
NZ9P0cgOPjH8Ej3j9zxnaST1q7tfPYFU64QgQoWBP+0rXhi2RynBY8nwcMhf6WvDQzyUgK/A8+P6
BRzUOOLTpUDYXhyuUgXtul6L5UEM1XOFuciL9vLT/Tp9H46gjeOg3BvJnPBt3bFFH5DZj7DH6xfq
Gv9yii0/hsORfo2OMBrqcUpBGLu5pXONqy+rCFZv5eeKOzXUUgBIXnwSTIGdq9fEBJoJA62DlyUN
5BlB4vVyoL9WJawL1vUKNN8Cim6xIB8Vdj4Thno3EXA2i2fLHP8x3s2EsWobbhry1E4XT/QHgyMu
uiTS6DAcndAOx2xVqX77erRZLyiiw+J0wRjU+eY/7PFm6Zf+GPTZ6C4oJyYQgeuf5Cd6BikVLQJV
Ewni5bDCKxuzvMR6ZcKIcg2HyWllGCGM4K7Rj6Zy1sSjLOyMK2lvBPpHQGFt6TCZiJBYvq203Vzj
MX2rCoKLKQ6CPPpEb8bfv5uxXMsNy1+MFCpkfzgK80Y3Nduy0MyDXWOi97v2M7ATXzJ5i0J097PG
xxya+7fPyVLY2bfcTsC1VJgvpYwPFflf9MFIJH5dxTQ7Y3w4HgFJWAURONBZB/P9rRss77d5achC
p70CyLQKuos44Ujw7tjXT7ZnaNIS+mjJUn4b30IhXq3YTnPL9C75PoUMciy9Q/K0eeEygkDBxlz1
Zaa0sxf6phXGsBz87pQSBtg0D4KEO5Wv8PB3I+2XeJ7S2v4v1nwyly+Q4KkhMJxMY6qixgbDCOQI
523Vor6cdsPOpFfTguJsjwpyjCinbNa4CyST+j9cDTiuFNikjm7drPbCgUdOj4o1eD+Ws+X5e524
eNy26IKuD/CBzuwhba8RND6s1OLNzLXLjZQvCI3cVzwxMWfVk0IG2M8eRQmpqMc+tUF8QeIAG75G
LlSALMfGLXsw+QxKiGFRWXQ9mc9FdQCSN/AbaAWrSO9O+jjtNjmjgOTrkR23pJf8mSiTD31jsD1H
HBNVjnlyy2r4m4lgVC5bsuxp/cH70HsM9RiPfap62SmB2OcqNmkWp0h0LJig6Kv132emgmGi4oeS
VfdjbTx5mBXxpw6BMJ6hRrE5R4dxH3zYj59p6Rbv2pJ5afiSUSW7dv+1E2tT3/IppIbZ1VY3IgVh
ah8Uu3BWYM2yn7UOL1p5ed84GgRq7b2SGjtLCHOO+FQQdcHPIhqLC4/PGciycA9UoqFyXbgpvf2M
1cko8UhON91Ck/9bKs9/sDNYYXSPXBeA6sSzoTaK1MQ+fCgmcGPJAwz1jfyt7OBcdzLfdtemvgO9
HL2PK2h7KG0P0ut2nzP/ZX/3nQ9RqLvwJmyaF+t45LGwLWbl7RHT4KMg+BiFviLWLwmb0TrKUkYt
gb6eQAL6OuAc3iYSueOaeZa8xML586TlVF9JO/V4Z/uUbq7A6EUy6/fXWYcp+6/fweeIRh4JG5rX
fh5yiQfjc1Ag+ZpF5a+fORRIG23DCSPFqbw3YlfBlH+9GMb7EcNUPvBQ8YxcbL78+3FA8SiHSGwV
PNEP4gX+P39M4cc3aNyZA6fvXgQuLvVkY+h89HRtqfFefJhKzYEfNQ3iF54uSuVHpjWx3ApEaSZ5
LmTavwnl+GTLmQWJhmk+FmW2Zvo8f3QY/fmBfCOqJQdn8Bz2hrmOe3T39LO/AWOaHFHjiea9VHCF
MiM9IKlPUq7BeSv417tde7kLLrgaG64cZcc+50OZ7FytYcm2XRnSS2r7h6OJl6kamcNfEoxmKea4
COOvimeq3B+K7rxfJg6/D+Kbm378E3qEDdPtxCyQp/q2ZfMEUmTe6zAfKB47OFZqsL+gWTLCayec
6+npFoi2x6WtwiVZThWAT8Yo3wadQHBd7FhbjB8NlXJE4lp31JjEDTnmMNw4EibxBuWw7z4voJTf
5KEvRf5gNAtV4Uh/vlEI/trDyLoAHExji2BxSZ/sIgJXQnAKiMO8n4syRi9Z+3ZXyEr5VfxvNbYF
qS3IcVSkzYXhtACtmkicG6j96FRUhe24cbU/mug3VagcJYddLxQLDgd5lDqI0o5N/myyehTSzyhr
ipV85HWM2/ya58F3YFylG6xNd7qDgG2i1KQmLWlAlr62Qd8eQRUYUA4xqXNz7oYJ5mjkHFuhguJD
Qv9a+ZhT7GNbmaSaHNrRs9mkR8vdCAhN3/xpyJhcZ4X9utTt36gVMufT8ThD4JXRAfXQtAMdDver
+4oBbXX7LbuRrk4wjouUBcVIR7L4aOCZFCOCz4O46CiXIaJ5Qw4SQOJCqXi2IiPGX2kmr5pB6Uje
oPnSQPlUogcTsMoneax0903ucmkILU3e2cF1AfnRo2rjVsBq9Oi/RNuFvrnJ8qsfP1TySkIqM+ii
XlX4W+bqtPvVlW5+jocVg6kDF/Fo8W9cgfp2Aym9jWOalo2OnvxL87WR6mTZjVnEJ8q3720XM8h+
ufrIPlOgJLBvSKQZ+baIhtm8TURzCM8mqVu5d+SxWXlWqr9NclA910f0e0En6MfsIgYUqHKN09jO
F9oW+lS3CJHRxp9tmF60L+/oQ6tDGkxAs/fZt8EFmX0tOX1WWanH5eTbOUKoqS/SpiIoXDg5wNLr
8tOWwLwLEynmOKhF70de31M0H/M5qVklV8grqhGtEzYaieYhz3fU3/lPef6BC3ZFdv67zWOR8Pq/
5Hg5CmeRfKnestMhq8Cdw3WAORI/qz16YBOFMChUjgPkHYLQYvn3QMtwQFjXvYzp2HjaoTxiEMmk
sDGXHmlnh7c7OYCIAai1xyaLFLc5bjkdEwGOf5vLvYug76PI2oH4TG45gvhTYrh3KW+AgrySLWNt
DppdVJpKTaqEGoWWU8mrmS5pEZj9cpFURWremjIYTm/DW/SZmGb20IZQ0Dn54edgV8DQ67EcvZOd
lXBTLfPQUk23zs5V565Twa3869I9vGxfPtes1TAi//Hl9LZsRRK7zaEq/cqZdUr44HXLxOqREYEP
n4d1hBH++/bmB/9YZYJPFQ88+r1x5ft4sgQc7op+nbbvFquJSLMT71YhnpQU1NQqbVGSbG/13YoC
XBxaBjTI40LFMt64tSK89yztBMov4waGQfr+ZFwVNhrhEx8CY3wddDY8OMPlObYOaq6tJTBqCeZe
ivcMBeAAeSLOaMPZ5/523VYyI+5lc++0pIKFgas0rjPKJUZjbHQ1ebAGJujgfk2gRtfKE+QeDH+b
LGDcDzJpuKcEsEAHjnDANKVQWaT6THWvRZW36Oiq6dtKNNpi1Du0Q5o/P9cK9nfBI57bwNfGuExb
4AhvVwjJu62YgxwBADM1xAdEdpUj1dkgP4nnfbNCTJhEVMfJKUyPR2eZIP6NUfMcSn143/uT9k0L
vPFgCN1k2Nmy0vielM8K7y9XgeK4NZCbCO8roRahJd13KF6ZWTCXYNiyZYqxv6iwciNrJMuWNDgS
xvVWGov4/GYCiEETQ8CR+qUSM/jUwYXdpPj8+6ErUK3DiAa6rMbQfY3P+Th3YcZKFCQO1Vlln86n
guSjYuRkmQ++ZWyaKgjtTv+dT+h+piJOOwLfe8R3iAnKN05XN9A4uGPfgj+Cna0hjnmUAQRojS16
qMvv0mljZtvTdTauNDhRnD2q7q4VwMxG3hYSyWpZ+eba+5QCpugB2e6l0AUBnEArc4/9ZcecTJ8o
9WNI7CQLLyQytLd+4ZxzOwrPN1gshQ3p+J8SMzdyhFt2NYHcA68SOeTsccjptHkGcNwp2YWas1hk
jCdvPDVKY5Axs0utgn8oAyxmrIX0hxFdzBbLMYFIiQvL9ej2kMsGznv9ZPR/Er0Mtf4XTIz5XKcS
XrRA+bNA+wNgcPOz/+J6kn9yMrEmhRlHXpoJLyiEPHcKn30JK2KzF/57XaEhYZ4IflpMzrfG67Nt
2R79b6c7s22pQYiDXux2AkoesPTZMj/NDqag1tMFhK4TX7s0r0zvKKmWSyoccudjm8IzLnRQ/pI6
EefgzIKcm6xSJARFw2x6HjC2ZoCObnwbPWri5LHL6pqXVWamxQ4AN2s+WUYQ0J/hR4pXyGn61eKp
/ACBGkP+jOdhd/trT/lzORDtjAmUDSjbP3dEOnU1E2STw92CqiRxoKcFYowrHlCrLUeWnAHmMqQX
p1g0F4IR5EqNonRdyLS7oeiWNGe9ZQRciIy1p9iIMxfjTgb3PNF2pn5/x2BIAlKi6azOOYqqJfGZ
q8YBB0QmtKwFbNJSu8rEDBpGpxhEF5nTZe1Uw2DW6i9a477UrsyDDLUR55pEHpAqvu7SRVvJV8gJ
qz2goPOgBu/ysXSIExIEQFb47UmQhhBV2LKOx28dAGPfac3nCbSVOmbLNZmSgZo/TZ6GdqShRqbB
+rRKiuM3ggHemxZrHhNRNLYtkw2aqiatRoq0M9ad3MoyYsBn60/m4T3pxWsY2unZJ9tmLoo773Np
PpPO72OIqOgvbnOkUees69unx/du8Y5xHt78b353wPZc7QP+5FKQ7zTNCpBI7noXS7aYi2x+JXvZ
/455kPtw+f1DTVbdd2QLKAgwMmHQsVjgO4DPFaXTEAnx10qOLnksjQ2mGiThCoaKiSzzroED5DMt
Ky8WTtHQKDyE1aonwmiRcVKe77sGFclvtlci7wmoB518DmoV8azMGVXOjMMyFqWkuovepELJncV9
8LVBlDgS3c0urm+THQX23jBW8JWuMQd9m9AULCpPrhQYt8K1ND0IyNKrwpHVGCxQ2JCaRBmLU5ra
V+k7D55QedsCEkKwHjoovRSiv5Gk8iNzhH2h/+G1iyPwSDkgI6WG9LH1xAGB+kWkDlMoxR5LryVC
mY7CaEgWLyQi9lC0bOS0VVgO0fhA4tQwe9Mx66Ld7X/07NkggoF+y35An7EimJksMQBWpJPETfaX
CMF7F40jB4YIXAQom/PkzK88POv70KlVCtRId8pj3g7EnFAMkT50eU30gzSbwCPF4XXmazWiMbK7
78R+E/mjS7OS9WnBB4qgTf23Lwr8VA+zvIADaei5JGNXum3oUWt+a7jvoGtYUGCwEc0CI+NEc6Dn
xUy+IJa8i5ksuLYLtchYolKrzXzs+u33AiXFoDi/DdzCt+G4caOoIFBiadTO30xOfqI2aWqErGqc
1zgGrEXGCELNYiWsa7IUQJwetDbzMVTBVQFJuMMGZlnIoqyLX4dvhmoPBHGbntNCwKeu5rab58Np
9pNmKNtkz99bJwh/kqO0aRzbnUy1CK1oPDDNfFkRBkuYCnktCMQJLOlKgh00rLBe1HtOK5zaXyPq
DEHN3x6LehdOUNIpJDmh6fkf1rAakmgkIKpVhrTs6CRyxuI5YTAbiQe9W4KErEsQI+mQkdfMzXqr
vYcbstzh1Byd966kHo0O8/qZmwaiUo1VEcTqMGCvSCKEo/rpThHQgILGVIrEEUDel2/sQlgalYHp
t3Fp+XaCt6BqnB9WY5rtnA6pE54jo7ctvuk5jnv++thSs2I7dFuTeMcKq4XBdJBhYavcg665D/bg
AX0aoiBQi3TS2N7CI81kpSRrCuZYRJQSDZ9YGPp2JASxlDjqecDCtX1Z2EaysrSwpK36SZliXYkn
mQJf98C0RVaDFIkjdhIcDUJbryIdkpFFmAiX4l61WXUApG/UK3tWMjpoHf3UO6YrxavBjodZW4/s
9K/e7rxfdnDW5mFYGpUtBcWVlZolp74JN6bM+XtYyWvdY3owah3LK1isbRamcT4o6T/dJ8eivQsv
qwM8ZZpDd+bQU+L0s3R0PcFXwwEYx0LJzM19KhJsWAHxpduwGftjEdxDdhzXK9qOySifvjbB4pwV
wXCuA4muMtcFxdgRwmrcuXXyKe+H6aIcNR7af0fsBoXEKhrhNxrMZoqhhmddz5RsKXJf0QMODz1d
0WI5qZkU7ID1P95RsMWcrYH8w9KsrosJPe1eSKEecyVbw4Xzmg4E5ECKDBGs2zLn5v/7NaoVgMWE
Cdpr9r1U9AdyG3k6meYuNJLNoe0oAy8NUh0nfoHaO4+y3be5g1wC5IgfaghKfQffzrwYFxPStjny
4x4Ge5QcmfwyOukBzbOUEtt0O5nrYgg+Rk6IGas+X9O8jrOYrIBX+xgZs2Ikq8D7kw1KK+vfaIeh
LEKpoZxJla/Imxg7WH7IXRiSD8oWoBS6bqEsp/n1UL61frZ914S9BAVTCz3iHyNhLfQJaLV8VcpF
p9qKWwPX8NETzaes0AhulUElLVv9gea8T7tL4Loshfar2q/e6d9xtuPoQvuh4cg3pwoF9zHT90g9
lICAXJ4rrtffK2Vr7icmseOTayYRAhQIlAi4AGVkYmZM9/GGOIXqCNtRlIjkZPawJtpe37HPtKSY
QyYP+wLTXgaetDpfAV2hWF6ozDfA1Th/18nCgMIOPzz1zd9VXgjylGawzNmSn2rC0rXqhh7THFih
n9FTbl1N/M1t1mJpHwh5SJEgy9+UMsErZwVn5/gyq8JXJlhB7oHcJSgYFwhLW3eCYD2s84e7JFH3
z9pupQ7K0kZmrDSEYCUqwekd7Fa+47napGPk0nzEPKVQAJoQWV+wpYXD2rE52fWPJr9QMO3CyrvO
92MmF1H5TQ8HUw5WSAhlnWTUE3np3XU1XNC9ivkeHgIet/TGUdW+oeC3vQZyJOC5oZtVTCzVeZ6i
G0cmQXChQMjUFXPtmNQ6WWTG6z+JYqU1IcVkxG6wFVU9zDLF7iDqRv5KLsGzu1rrNlzotg1YovBE
0liS2domlHk2y3kJg+8XpUolN6uBd9jA0C4n+IgXwEUNw1hFWyuw3PAZQRwqwlEZ4JkQy42Hnoi+
t/ogWOmCJthPMqHLw2xsVPIfr9ZCQh7NmS8rz1Pa5IVR47Kk4TREc8WbBv83t3VCQ4gqPO+b4Tta
CwVoYlFVZO1aHrVLryJMnMDtQOisUmLsj8dlzO7fYuBiEOq38JMB8uREjkUKPQKwHitt09qTLA+u
aFdDJPV4llADem+63iNpnjIlzpC++oZMbCZYR/sWfQSrBXR5ypabH0fdzzVtiBTRgICy7jJFYhcQ
4WRp1lJ+0bK13kAYnt8N5eYic+1Nh5T6JSvp8XOpS/Bx7mS9w48r3JRkdZrlILnnWHrwHbr7ui1F
IRGQ20yi01ShZVWcgAByOOCx4P6VzabcD0cmw06+MpcF0VVAXsAd6gbfPDICQJRdSl4xeIXRK3q8
OGfnZmfWpjzpJX0MVlLrQZDczfDVGv5/Y++WmXCV3zstqQoehNAZZXRjASOcfBxpbfHPEKWZiint
Z4K1/uLsL+4oaxqtiqFVt1k6JG5Sgaq0nL46yB91qENJdg0LSbczkjzlFn6gFTbmPT3yuwRnRhE4
aL6fHOurTMdkGb4fD4KhCHsHZBAVQeWULvtyAxfgURJVHH9ZcmfAF0IQcRxUyKSgpSjbU8AFwKmV
ZX6V9MqxJl7PreSohuvu5tXiZqLhhhJtBr7qNEFUHFPam5IYGB7tO7RA4lwZhraf6sDQkUOXePI7
D2T4EdqMROfOQ+eiKL8ZKouROcfgSZ+UVxthwF0r0ncsDWOauaVrHJlZKwfTGOXusbjMpR/KlZYL
SEsAb9kFJTbixWBz2CVA5jwiSmd3pqw4nOkSmhcZI6DK2Eyx4prz1DDTudtmv6sqp5n47kCKNG4W
/v/ow/N3+MwIAmLEtrVWrzY23TAspAUQ+Ouk+e2DoJDVBR0RLPE/momKfhOobzhVxb2o6jihwcK9
WW+YoSnTtpWSZq9AfUzGd+VKd5UPcG8hFsMuusQDZV+69UrXweh4PG5hbyNB+Gc7fAqteLkwjFDH
zfooudtoIj5jGc3WkpWNSz1USLCToMVzxlkmTbx/TTgeBS+zj+5fzIwBJe0xhn34BW4Pn+3w3HSX
ctUJ/uit9/L0ZZW6cOQ8Z3X8PK6bf2kn0pOlIh21GqrluJA77EVsR/W4QLcELn1z5cvj63+r7Flg
0UHNzhcgYCIjaUX01Et5RQ5o9dt39RAQz/1RbVm7eOiximInFIhycF3y/31XywmA+SASdW6D6pW1
kGY8ARSZnSRysQ4vKOEIK2PNl70aDWpJg8CZJ4BLaZkH+t/vdyTaCGuG7SJube822wtsJMKBy8vA
5EK5OhJGQ7m632TgXh1Li4Chje8gOskeDstOFB4S7sqKC1iOuELqsrHRnXCfN3JWLXKY3LjOiCmq
A87iYC8vR4/n9TI7tAEEkDpVP5YLvDTv2mqEahJcYSgs5dhEuN6cxlHe3qh/lKPFlaMfHefG7pbG
Zl+PNSKfMNzupYhDYnIFAsTkNaGGh4eaXU3UgqyEAb8xalxftj6j+kF6W/o8bRM+rnzVq0JIIkhm
6aEoxAJJlvrhWlO2KIDqsaHYKl3sGNA4K2OBaS8HTlL6CrrWxz5ARmfqIKhnh6JDr7D1nSeNYahs
5aRW99bJbriRogLVK3TQCH99WjhK9hOPvEcIjriyOsimGKzOp65Z1iHdcASARm3ZVMjrnJK60zTR
YI+Qc9pQlDidiHtdS9lLAqVSACPh+tvduGNY+8eYNS7HUuQ3DmoVpwvv05vBN3060zyZ5onnUD6J
OYyx707rEWKbqQr+oMFgw+FP8DzzqvxtXxgkoUAX1tbbPeB2uOYQ7w6Ovvv8pxWbqPzq0ZV0jnET
picYSKTDrD6t/odqWZEYofIcmRAIs2WRlWBBVy11dRf4gwRdUCqt7i/CZqC8d3A4dIC+DH4e08pE
KW+l8m3GJ5QVWs6F2whZAvhhLNVBjjqCAz69nfY6gTUWK84Bc3oTVFx2jqXyRBMMWLYfqWYp4AhR
r1bxS/Jpfaai6aQb7rVOKvU45oKx7HFXLjIZz06sWpXdCEiQafAWSD3gjptr/wBytOO2OkKGY8Nk
jdL1jdunGg935TxRj76it7t6wVoa5CWWPKmziYHZnnS1sqCKXryjPoUPZP74PETSPisvHHpB1vck
eMfL0/HuTIIf53d4NU3g+Dt2O5gdw/gX2A0lMlcJC5y/3Giy3t74wj04/Cbfes6eqV7M77b35iBi
5RFus6U+X8pykgbcceZg5d3CM60lSSovPXkvJr+3czPAiRLPJBzfFi24O0p/hAUO+4ogU0RX49+D
r5Cc47WLxE1j1fuxWL+LehN4WXXTyTg0y/ykacxy06alxge3wagNcL7lxcaysSgm2otllpK2TyOC
m3VtXdafFLKdzWjwaKB18c3eHwDvV4ol2LHz43hL8X/p0YX4grx7BmhMEDauX98Vc92LbhyOgEAz
ouTDAquhM9PJ0WC1eKbeW4QQxaYQQR2+KhX2A6vWlP6IWfgt6WAhBLBZAdF/22sSAVSDwUSW3QQE
ui4SMPNNM4NvBqwIhrSoLTRUxwnbvybYy0RuJwmcqPz0kha/Ch6xCBqlyRTcLH5rtNXSlPDPnge2
RLUpIzb57Q2W7nxUg9UTrJtqbQYERBU+F20dlUwYUfvfUL0Z8+VikM/EO3DzgwmtHR9XBDeqU/xl
94uU80nF95DZA19FHDMqcEcNoXtk42+fK0fv4rVfE4gAxOED157Jpupa/WHlopzDzipi82lorz73
lbsu/ExuRpo+4bAN0kFUSx/kGQN1K0SpnIc7XJNhTaaGmu0NIuEPON+NmDd7zXDn9/kTmpMYce2C
QJuSsczyUF82jzsVgl+42VjE6IVV5eCw7KYC/AGqCh8HHG9DnT7+itA9vt8j2SvIsCCltcjohAt/
7WJuu+Xqmu7PVT5KU8fNk2J2U3Da5Jv1or8qiORHk7ncKLr1UruUCzhdqDonStx7h6Fviz98hGeh
M8/Ct7skd02KReH3V/WyWiRvkquqis4BIQo4M7v3loZoX7pTEMILV8k0c/DBWLxZabbTOqsmEv1Z
egJXk8iVp9igJnvUgBF9HYWmvSm/hgqRbSjGxdSCE3I/m/pSmlFMKmNQIbIxDbHiddXzw1zJS1iF
6Ou0UKEkVlESdOzfejN8qYhFe9HEnaJYR8GQBRM4iVtOkjnCUU0be9rOFkMq2yf02HbQcTpZsG2k
NU4A/m5GhTS0vPcYPDuPPDP/1x7jr+/XEUmHWvgA8foYVgQoEChWqvAM0A7UFv0YAa7c57g8GoO9
OokDJ//wSelUtqKHElMMfY78f0wRJ8ewGuxQoUGOk5mj2vU1/maNTxxdos8nIQbMP5TRpa4xUae2
BjZj0tuZh7JCHJQ4xPtksEXb/btBfhGkDtDauFHo/TB57V6z5FvyPr1hwdAYL9Yh+PBSMvw+NKdz
zJyFcVsz7BBf5/nWUMCPMvp4S7mq90AxLYjy+wogCVwCy31gJpQTozCHbSjzIgT419+k6Mt015FA
q8RG8TXD1vdrA/gpZcuVzmKP7U/OTK/jqXW2Qi7k0PlbrAlyx5j1IN0112qzVF/ow/HAHwwMX+32
br0A2bmB6ObLpyNUBnIdV4Ag89ZCuH5WjTyL/G2h4cRqfz7uIO567Z3CW5oWtrsH72BoaTNhi/6k
5qw6sLv7eYDtxpqlDQGiON0+a1oT6LaNpVF6m+JM9Qk+xJsob0mYOmtoA8q+6q9PcCi/dzfea7xH
uD3LYBPC3xUrJmxhgZspOOXkxzey+ZObbv1bxXFGe5vjOOKky2eMqTlGeNvNYJkoVkeRn+tAOZuW
aRuyxVpEaAvt/LXjB3Neos9qYTHpp+BQNYKxaJXMm4NmFe6DYmmobIQaXp7D0YwP4swjdAWx/5XR
t6FcMNpr95JCJs3ijSpWVh47xq2lgfyltBl6kjxzCdHiwBAv5a0hYPYHu3fOagNyKMytHMr1le9c
p57BMWnA8VNCbUtS1grJW8D013AhiGW+hoOlly5mldV0o2Wai2sxSTOcvvSzDO9RbCeZjRAhj38P
hH4zU0VheYw4Phy6OaqCnR/bPsucmorVvYDi5HEdyy82gozurIxrApFQyANXds6hJURZpHwRMMPz
2PLZ3h3mjL+sKzJ1A7Ae0ZosXNzgLh37TMKPpgAradXDmwDzFiVqPBIkBdUKFxWzANRbPIuWQlo5
1q/1/SsJn5pu/PtGD5GAsQOwxcRkWfjW75b9i0JAUTIHiSQRHe+04+PnSVy/RAFRwITKf5hLBArf
qwfWuc99LSdDXYSnM/Kpb4AigZtNud57b9GyMzer0DO2hkxGvJZyhSaOnPL65xg2vsa9K0FPIygm
U7vytELFzXwburyp6m0I/J3qttbp5wq0f9Ep5LKj0XSbsFkVh6TEB2jQ5peh/DLXb/AjKeRTYB2z
UqOsgwhQ5IV1WH6+IcLa+QTH/zKWftN33QGFwsLdf7DXnb5KY2L1pRzD8ec6R2pM5IfAWw9fiV0I
/Mxh6vl4s0Q1apJUp2PwuIMdRJUHBDrj76w5hXTTBREQpc686+iV/vRc/Y8T2x7TfkiSSdw1OFZK
rnnSHNIZaXDknPI4YcDWSBj1eCTun2OpwH4W3+/8nCHnmQPsm3j5bxuSFJBKnihWSyusaKQYtda/
llHTsOWLYbDsKTw1UHWVzA5nN9ek9+3H9Q4pP2dD6JNMsM0QK6G+MlV62xEcNl4xBjVK5UoU5ozX
df4LXogDIyt5+w0g3ACpnVPd3JzjLCRD/aYvuMKn4QAusYLyBVNYAmVclBD0dPbj6JPxNb23Zp8G
xEsMN2TsN8XARyDNa/ccMoD9EN9wfyMC91mZFPKh97yquML6a15Mc+r2VdGhFDdsgnXmKLen7SSM
sIHjskp5KYQ0lO9Yov5fxJFg7+/28JDVYZAlFgYgOBH6RP2vMb6lZVSA2PHWYGOOll/ZuNse0xUG
q8GSpIllaD7uZDK5yrgIDqJmkVoeTftuuMmNWBjN0lCg7/Ct9xODfKGIrXjBWxuKXQ8YPB1pzap4
83nExKUNgaSZLlpSnZQg18QvyTj3FE/TnAoV9p7BOjy7sK0eoWwx91xwzmBuydXFrDvpSQELX4l5
EqVpldazdcNJDHSycBR4yl05NUsC7oOKgZO0JeWpvrcr7VXlHFllWxz7uEUBtCyr17krWFzpZpN0
muGBWgMKOyxb1fq28AtN2IxA6doGbz8cbM70fcm8KJLdsBfUztRADeLuUDG9Xi05dfVbYuti2YuK
Egg2wk6LB0HUatZSeFcINCYn7oWT5WSpNyHgNkb0Wpu3f0/ZTg/GPV+n+3TgB8SX48o23BCCX8zK
PHlH3BBqgyrFvEAA2ruGIEYBoJ3LgC6LsaPN2HAh4agFj3s8cItfFBHpKjcfjzrOI1lBE9IJ24xH
3ZfBJMpSzhZXbKHMSs3ecGhiFwu8nxg+gsxXrMJUJDa00JgHqaLOXekBBPw/VA5GpbUnnyU+/esI
jlN+M1EckupnoZx0m7wZjWNe4/0y1twaFVybLEO9R1Ag0+ZZu8NYUrkI2E/DNryyV/W2K3X5qNVC
glTuOpDDn9QDrbij40ohOU0sCWXcO1tP4oCFSQj+aueW/93rAU5s+wfVB0SEpXcTmzYisw6PFhks
bA04vSu8xelxiJ/iVnfEr8lTwe+F0MXINQs3IGje+BZsaFKGsMGuLvNNdzGIT7ltHT7rcMdtgOOu
ZiwSPVfgCLzJUp45lIo8rllbnbqXrd2pUnkLyVBu5OBfMVYPRuzVppmWx2qygO5dFhfpd2nvBF/t
pzFcEsqDJFsYHQKK4F2ymFmr/d+ONcgxwJmRdUXhf/KURHh1XVCwsUA2DyE+YNms+My7obJbxQk4
G1oTOiBB+hL5t9uONYbZJcsz23Mf+o3QSt1k94uF9hSgemt7rCEX7IwIpR74rB1RbIPhpp7eNwDE
KeXM5uCRZ2are/d4jhydtVwaP56yAkgyOZ8mLPxuxj7mG2O93z3Nb9JNhte/Jcebsg/HkF98DsG4
pvtOE2zDrWb/7WoKyn1GCldiAgANuNtDo5DYZODajpMkexcIcpl2ew9tNwleFsXMRbXxw69tLmhz
90+Sro6hLmN1jHZPodSGVtJv65KLXr9isimwJV0ht3hQ+EYMD6vNErMTOMVfOck63cEXKXmtkHbW
3XlzqnyN6oA9qfteKtjnJdiG8QJAiOch3OLpsvEiMcx6yByc1vjx1Or9MarhnYy7VnQeJiH+2SQn
US5/ooqVlqR20fYsEOAGTwBvfg7CWyEmMBM9aU9zXh1V/ryhANuyyIAt87OBYUW9UArkdBgxcJ79
z4BawTQogHCmlBNRouA/qaggJqDtePK0ovu4vEcLPM+gPBexdYPLwgGmMufPisEgAIENorsiy6PT
+dTLoaj+hZmn6Muk2M1mPsTDsO52CWTXQGCc1n+QHsBNCYLigyFEL1cM2gwk6ZDSgqcyvvCP5xC2
CI2wYab3vRIZHiCY1+Ffge0rKJWTiL0bC/CQdCn8LGHzLCdUp6oje8NKHhjlDvcp/bqnWdsg7Udk
mzK1N4oWWKNiSo5wMI5yYAoAF++xYYRzJdn5pbQZUG/BDpALMWiRPb1e0Q9TGFym8vgWnG3cZzhE
zMgx9olhdqhgaph5mpzAfNdgaL6k5fwVcJeRib10uw5OVCv4zDg5VzOYSOIY3iU9KlE/Nb5UBd/c
X0pNU8DxpOi612QE71OwVAt/WX0CKmJH8wD9+M+cCWMpv29zlrkQDpquu5nSk2cdVoZu79spYA+G
u8hLhKuPPVTU9zwuBlQJ8Nf+s3cvph1c6V55TB2gy3Z+Pt7LSg2LZkFkM5zittrQHUq3WGm8w2GM
CCAeNc+zw4+V+rEeYGktsD5JH08NdLdi8NzyL72fJn3wA7DFIyXJjsFBLKtaGJuKNe+fyskflIXU
wC4dlf+XwaRL5zPMnw5ByhsEIjUXO8hyzIiYdYkWgwCQfVJAr7YPaaGEbsitJ331yHOkkuNSL48B
QoXNZ66DEqgm+kWywPmOf17VFAMHr4aps8OVNsSQZZsCyuly+9CBLLSx+B/M1EeTpkTd5tw2TDKO
luV3gz6w9SEPRBa2dvk1DksQ00KhNw7os9B3BpqeSgsP5oOWQ6C6bXyGmEWzmo2k/LaVOFYzIO/2
DQ123p4A1YmUNEvFSF00oHpijZDn9U+LvfaG+yYWf0VKZvKS5oi8/CwOnWhJ+MxGOCKY4ZfIY/z4
r26WX1iF/TMUunlEgBRgl7TaIJHNKgMRbJxs7TojIsfj4DvdU4e9qXwPUWVOM+5qP/+8v6kRiqB9
ulsV0HYuueoYwa2j+3C4QfO4ctMa+7XvPe7wTKCaDFBgkSVQbjwRokc0d/CSOjxoKAww+5z6cL+5
DO8SJvwZg//PxNX6J+QdvlQCYkN8+XuYq+dbKYSUwcT2uNQNia3c3GRk90nGB6u2g/HAZNTWgUpY
rFh+ydHU+GXn17iUXtLNqD8UPv3Dt+vWytDwXHRWdDgswgYh024FqnZWLABpuiZMv2csra+J39s0
9HwchuUBmfCrYrID1kw8IQsODUDr1TWDNgVwixJMY5ebLWgxB4N5jqjgSM65ePStJZUYtH8MdUEd
S0jOxjz1WoPq1UPGaqR4EGJf3Kj+Id01CgwdcqHYoFLUFF/nBfqYcc8oevo5yaihZk/TeVNSOCXV
EHysnPVQL36O65tnMTUQQpsVNZInVrwUiejZ/JWnigzde5Kj7WX7h4e4XQhAu4EvyDJrAooD0jp0
MXuuaTdVxvq9W7QXWAYpcS1TT9JA+mwLLVS/fZNPWBPIxab+U59wc2jXHv38y4SkEhBr55y7vweF
KH4AtdlKLK4sJxQv3ph9mg58h0tFXWE+v3BiI6oev89/7PHtiXM51WPO23mUfsIlng6/hA8GdOJF
c98vuOHPpMO/y+DsVxj0+Apm9FOICu6xatpMrmFYdjsiv8aMgW2shP0LQy9ocAIw8Cr9NT8F6hxe
0SMwnEEjy6myu7SsYnAgZE/CFGsGntU1QwUaM7/vHbAdbG8eH10nDcPCX8p86Ppf/49M+g0y5TAG
AlZEflPXuycPw1t2yzbKoNTAIrm5waOFqh1I5kqGzw4pkYTVw9EpnOO1hJcFXh70q6FHlH3Zk4QC
tqA/7chOEq2mnGh4+WaN9MZMR2qm9GXH8OcwLPaO+tkXv5YWaFjZmRDDr/GKlPYrsM6huse91PFk
4U95jsfsYSfDgOIxcreg/xpoyHXjbTzx9lFbKT6C8GPq9cjVNkWZcKsmhRcAu+6pqDA5KGqyay+9
KjroCqw9jmcd6NJGgBlRtwDV2KPLDkZ9oVf3INDPWR8SlY86G94Ogortjt/Te20KMvAmHUYtgehL
kl/CuUlDYhusbhwumeT2JbGaUstUFRiZrMzjdoizX3E48Ii2w4S5H4vBBuXHx+gmANaEJ/diCiy9
kxE/bjmQCTiQYVaS6bqoW8GDGKd6m2g4JQ80ficzkt9BoaQGlxWbrdbQY7qQGsrGg6DAgV77wjuv
bZZCh+a8WPi0kHpxI6BPTyuDI+xLmUWOmerMRtBf2tta/9PlVizjZ91XQncGz+vX9wyxs08V7aA3
1CGdwme8lZLMiQa/pnE4yEbnp73MOKP9a8aQ8cd6NCEmRxLmQsX18XvSTnS/fBLSLKj/42i/Lbmu
b7g7xvlMOcOMbcIgTRIgTJnDGok3uDEAcgm1NtfuoeOSJMIQimjdK1hF4R0s9EVHCl0WWmpLujSf
Z/kas89ZK2U3QOpM/ciJoV8UjsewxbEcASEYoBJ4OTQBQAzHgjsqw3VisFS1VjhFv3zxqHG5glnB
E7dDijxx9k2aNozgQ7beS1v8qw+vCvVJz3BAErhH+N4ttnVa1tlkZFGuJK/CSA7Pf2oLiykZXNav
UROKk0EYIqurV8UgN3V1F+yMe2Pf5OQ23FhmGpB2iYo433jrIT0zHlD7Vn4grIEjsLri2kZtOFoi
wOYq/dtHI85QuL4jlZVQ8Bo6vTYpx124ALIBTgi1ZVx1hXA2f03ynAVROB+lfhheJCk10CbaEl9B
4Hsn1mCmK8l52wR//V5TJG0XgspzPfcwQj7gFhPjPs6L2PMadxxbIf+TeVO1rhPWsuSPdZdrcZIP
X9kZsI+ZROvafUy2Hdch6TtvFVv1LAoPpSLhbPvLqLNiF8z1KZ0j3h67bloLfLjWzpgLOE9c7BsX
pLI3VlF2VMyUYfxM18QkGF17rlcEaz8Oueu+gHyyL/ubfJlGeB3Ex0pBzXKz20SjBkhMSoXu55+X
zOnuqXRo/ZzuYKdiJe7JL+8ou1RkwonOt2TgaUhwgX1VIsHzVD7zQ7/iay43lUBwMkBCd8an8czQ
HNm9WcyTbGavBEzdr4zTbMneLQ1ow+UIJTiNtOzX1So0nud8ptypkBfJz1jltMmp88NKWMggS8vY
LayAa6MZ43sIe+xkfJRYp2zv6/2Axr2g/x33G/UnbRIasyd/Zh6S6ckPWDQ/Gv1GLSfi7BBFtCG+
0Bh7asHhO/oNY/1PMiquR3epvLT6gHOePDTOw5dzFHzjNAPENsjzCqyUtzjQGzF7k/CzpBX/TcQ6
0p4dh82crc3LKeqzM9TzrEKFpPf5YOM5Ov60y9hVKU+4nj0NAogWhyw2ldtkkSR9xkwf44yZHkA+
r4KLygdHgklvC66bI9v2mPTfk3SV4MGZr98S24YvfwzLAP6bOekEPu1vqUYqwdwlEZ6wcWUGUFRe
NHYdzkO2s81v5Un5CwmNv0v28seROwqFFrcYKvX7p2BbAqIT2qC3EVFtDTU6QUQQJw4dRRxslnus
EuBEZDVFZzKAi6uMeOIBRxRNqB5++ISP5OMCflgX6BQ3ozT1D6FyrtH7ciyxIcUROL7malLnbfed
M6WI4ysj06hQPwDZ3rB2/lIIj/3UjWZlw/nb+teISx7Q8LP/to0rl7/d0+UMHgrduwRHVw+XiNYZ
n32NPHA6ykGpNCh7i5Esc88vp0JA/k3/BA+Ip36weIklLE4yZmQS9SmGuejjFxvwiETt756vf4m9
B5HEcRbo9aTQZWftbKgWvbbixIvDMDY0h/xSkd6zxz2CCQ1owl/rtsr4k9CDkZ+9Q1YUmrxvGdNg
Bxd+NF/6aEuymGCTA/AKHVhS3W/s7TU9CjGuIJQE9oeTRqHP2Ibd2oFM12Ba3rUt+ZJlDH2y97Wu
OpVQYWD10EbsXxyla+WJaeAwiUjin+7T0aTKRwnHNEkR4lLQaIt1Kg5g/eCmxRB1XEGUOE2IjyET
42uARsISEK6WWCV0ENJ6tE+TCGdV9InWA/X2W4RSijfEa/BXNOOBpPgNFfBkmQUeO6uZ2xlCoFV/
qmwfQcuyxbKz5j/uEjRDIESTVkh1p9vygmyOi+VbXlSQV4ZH9eD97bhjcSLD8ulOcybbgZ5RRviZ
mDhNRa1k0CBBxf7rVXN7vXBZu+YxxgYhmKsBmjCvbcXZIP2ZvnUPlQ4bcepbrr/C0+OqQTmE57wY
YgJGIdk9Nyte3QdRCn6CfZSe47xc6ibwl0521rawmUDrVHTmuyKch8hv33OFgAmwag6U0j5En20X
+5e/ksivUJ2cfrtDCa52c/LLA0fVMTiuYIyIY244mZL15hr9256ORdkoLwekQlwCyv5hATI0q8yu
SfBDN6P8Pzk5r3cmze+7vok60SAIsYSraT0rdPjKud2NORvXz2Pgt9stnenp/mtMJdjTmmHHvBB/
LFCptyITKr1BK23JESKZ9Ul62x1Hlq+uvAQEafJKmi8hH6bMx0rpNmAoBcufL+pv30afm/qFKbfG
oWQ+3TEQpjuGjLIu/p3x3jy0ESfMqim7jB0PSnUCINA4zAYLhFXgvTTkq15zzZXkI0UtXckCeKQv
3xF+nBCyhPcQIN3ZVCaRExGbZcVLXZMpejyHpLsUhazAU9rkImhw+0WusXlI0OT9fSLnffsjC/qc
7bbLy+PJbGah9uo6SZsuKTYVIEeib34cce8MYCvSphIsSHFZSYnQ7Ru8+llflInCVID1EdQA1D00
lJ5pCEPswQsa9r9nHer3GK32a7s32xlbZCp6217zAT6a+xkGBZzdlawcuj5stElMcM4hLrgNpkU5
vZNyZQ7BLt3L+dUQElpjX0+YQJ6DllrifK1Ch49TAjnERfm4Q03hqS2ECuROgz4DkWJxQY+nhZR8
G5eNuI40aBqNjh2BvPRyG/7uVXRQj/a3KeIWsg9NNYApOnfcjR2H+GjbcFKElhM9imaetO6mvlXg
mC6l75wECyrDXbbChSzyJWiWisiXbCP1hu7M/k7VLwfTTBNpJCD9jtct9VyWXujzmmkcIrO9Xjyp
DAHAiw+vMg71o/45u1XXwKCk8ZSr3mt1YIUWrJroOkviLt3RmJ560+gFSH9YPqzuuCbFy3b88HOp
txhGldvKgtUQ9lqAvODdmsjDVI7k+zAFFBoyOyK6zDzCBofo5/9WtE9+jgsgUpfOPUaKyWZy2Nrc
/tL6atiwRO11CcFOnMwOmTRC/b/CtAv3FS/9nJbOwsc6D/QLV1lRRoR9MUj67SlRVwaJt+aQgH0z
+cuR4/kKYgpH64ZhEptZn5pOKHr3euJvn6y/Sjgw18tXhI7db6+kJ5e4UpVFi/dyYyOfznfuAE+m
SHALng0YMlTCQcO99EDAH35sCkvGz9N5JDp6+cLQ5JOHzy7ibfCtZxnvjxJLEHK6PderJ+7a6e/K
9xjmkWaz5ldr0+ghOkgCB/cOoKDGAuPGjrGfIa+222WmqXj3M63dHIA4YQqKKd4CwnwKKMJH4Uxe
EvWjvT+E0zD33kAyD+XfgTLZ6/meZnJauMQhGitQVfQFEaTEQAl9Cnd6Pbx5CItuWfRAueqzPec3
t+IhU4xBGcqWPZjDYDTOdjU7o9m0c5Ee0BdVxKafOZJbPy93wd6s/ossv+EKyXHPDCojnMzFhjwm
NGBzuFujetQ6TEm4Ln2APAG6Cf3e4WvO7EFwNrB7AXvxdIFdYeLtddqIT6uNkftPryJE3Hcnp3EF
On57WGr8uqnH1aSkZeL4Ydc7oV6qzHdxFuyNLP5dJ0zdAX2KeAuKixl35agoX8LcCkKM0ADlP21n
tVl3ghQffQtMzP9py528oCo24uZB2MiXrx391mfTJ/eGoVnPfZL/hyXSXgfHpz/A/ZbTdumff+TH
oHXUBWRRGDWV/d4k2XZyzzbEXhfhfK1yhEdDgKjY+1eHJFRQKyKU57xK9q25OEo2JRcoHUm4gcBA
LSqzyQkshIxljOG90dDhGMqGL3dw360fQjFfZ2NstDaU3HZOHbfknkliuELO1pzoFOgwwYq/r9Qr
bGAQVUnMzkSPn0jdU3a5/cynB2bbk2VUu2fglmEyBia1JarsYw14MZjSwoZcy36tDNEb61WOedmj
qYWYfCMVoEgWIOrYZWoSTcz2PRdpV7JERqs81VUEyZoCkoJJgd09SWSv5OIZFRyF8T3uSja32Kfq
jc4D7mzeB/It950AKvyX4h0TfQsm9ib9pFnu32XZxpZhsjtKk4gsKkOyqKg64os4fcUpJp8DObRl
t9VUK1/oFOyOHLmuFB4gSz+Q67bjoZcBeml4sEvjgLSIXZUKasMOMLuQTfBYc7gxPlY3zblcQTzJ
/l6KxW86cr9khPo4LGELR/GIbtTG7//1iIZ3MhhCMrD2nrEpg4n7R6ERBwm5xNsLQgFfeEFb3K5m
54YX3UPCFitLOXbbjKSKImnPgJpa1rjz+1kxksH6iTKKh1l4+elb5McVuGnx9QTnNcGp9tA870U0
ThJxGxrmvSLDIONI7DIMjnOqt3fLKxstKz3CLXhtnthe40eAHXs2i5negOf7aq8cxhN19MuPDvTM
O0p69SuQ0hw7Ko+39s2T5+FXNtVI96i/tpk8jMNdrhRqZNpAOwpu5Igi8vs6FfotiWwNqHvOJCK1
liic8TBZJYpofHpuHJjhsyi4g3zIhT2LT5UXSYdjRvEU3V7ivJSH6OuiXoE1XWVRaj0ZtbIznuYH
Cj/2FPmuiWCd+8Ir82o0lW+rGoiDLLn8EBNSLeooCnD0jJkmsuDzdBpG2TowHKA/swYNW9DNb3a9
cT4cwKW73smNhXWlijehTHOhtKCWh+uqtf851KfHTBoUUi9pghuIDSxGgAxEf3ojUh2see0b0H2P
3fVHYl6HhUB2LRkziQYhxrdG8ScdNfxlwpvKX0jPj2ZDjxfFgWchd80tY6lDa1hFX26YpByYcYY8
cgfpr1Xz1GnaaLtwppkTxGHfqfFRaBM2pEnuvYm5uXF/A1w/iq2n8ING+jDVWzAgVzWGIf0F9Phy
KyP8jHFw+azTpb6alPBR29NEiW5uUoO6mNXLJXo4X5xH/HIpRc/kIiy2hug4AVZctzfVVsVjCHJo
IJmf7OjqS23bjVaWTN8hvUHv0ay5bcdFrCf/6abVHaL0b+sLaGuze799k8HcDZfh8Z+9Gr7KLXkg
ptTkKyqoiQ1NKsQMZj7NrM4ihRDhLHUKWjiYYXViUjQufpgYwRMAHjSL2aPCbwgjZ/z9W46YRKpv
rHkjpf8VtkJ9IEDJD4Ff/8Lgz/+d0QZTX3+N1Q1X+dW52hq21I5dOXC+A0oVOQqDgceQbs1NJK8M
F1X8fpGQv0iM/zQtgBrT3qPOTq12DNcjYWPDTHEuPl0yYEmEpGjEdRLbFLL16vlM0C00QPYsynAM
7ibYv0BOP+DyL8CRpSmbNd7SIeVK30N9XJoxyTVaH72dPSBvMAtFejlJT+lvBfQQ/pr19UABjYGW
ITK/9rS9/yomak3H1BhE4IPuCMlSdeQxpWlCle0fTvmvH4xHtKR/Elju80ayti597pYIOBzMNRmN
LIj9VLa4G5G6oyTN+KCL9t3oHXcXNlXAo+FWth6QQWj1MIndL9pR9yUuqygW5logSFQT+9Ffgsyt
PMLb75xdhgNSrY1FLrFQ8b0AvEcynHOUIc6/cBI06zkZRjc4owNaxCpH3CnusMkTAqKUdyfD1s0H
S3dxHQExz9YWLcCov98v+EZ6z3d6gg/HAECKmB4IEVyAuj9bdr+YDVz+wbSgVMDYyMaHsD+qYb25
nqiM4fj5h9AQX4kBTRgc5ftMdTT0SQMgZpYlBDZ/oP83WvVvg9bsNFdzrwMyeBawuSLC3UeOZNRP
GGpa5+8lS8i51kmxdfmN8UrSegLFMUoJObRTcHsO5BvZZS6+ABKhayQIB5kTqNgT6AW7yxXHihPE
CxEggWRRYyb3T1idbrdtJniQmDKSfDChhFQJNbYWfwRJbtzLwZtniNOFkrTcKk6Ex/xLKo9aSZkJ
c+6qSym+iAxLmkqX/RfRu48BAHsK4xOHCr9clQIuzjDQ2Wo3L6WHilkb3s1796a38kAZEud0cqhk
mYgY/UWqAnBd7UY1jDULS01WK65BvgvjeqeJbpawW/miNg5sgaKLTLpSlFdPklXWVtc2Z2leWNBV
RoguX4NfCLp5Z4/lXBrzT+QUU+mYa3qdkCuKsF3kcBcGX+eFDyMHy0Q5L3pcadwjzrRJrIkveHac
5G2cB3irH3mqEnNOzDZsPhvESOQXQ/tdgQc7iFPJvzBG8a42clGgy/22WrxAMiFwaGZBHIISULQj
nypRXz8XcXlBc41E6bMcrlQJg49EKWte2DR7fX89lpy2kBLNBMLMMjuDTJkuqx07cGwLm2Q/jmqu
6jsuxOYLAcleiqclA8Qo8Gjm4jcG9plsflcS4WlKkOD05dwt0R/s6d6t8dPgoctvbweyVL0IWECK
8uKy0IOplzAqj5M4NOVwxsA/QwDYF1tG3i1gOLOriQ8+jOJnVzBL/jxhkMpK872oGLbBgzVnxO0z
Q66OOlaaUf0RrpKQPhZNwRq1Rt6WAQTRiLoUzp1cTF41Qhpj2hgi6U5YzUPEo1833pq07l1Qu4l/
8ESenHyxKL/+g4ujicUXktrO/GUMeR2S5nXQNS7+pWfpd9id6mMmxj3Bt8lPtBfjscXO/JlzvOZq
K8f2bahBRYnoXq6kV+KvvTnCHy3tzvIrRItULGhcvq+cmFwxf1nLuEfmjom78RFOukU9WrcJdElg
+XpWX4oe72JI6ybo/ULqG1puEXcj2CtiOyj/8+yqlKML+8+qzqgedSU9w9PdbPnatxBKshbLXHGE
SWkg+APYoJJLPOG/mZUXQE6Qjg5B+mWLxvHRRizAANNWTJcmUpwHKl8C5y8JpYAVd2qtqMQYRUUA
NB+hAD5vJW09rbiouxjc3bGSdM4u9DGpeY5uE/H5eE2dqw4hNZFDZZKuI2h/ir93peL0rCMQJlGi
ebUPDYB1puQtj0dOzxRtrwgdEgxae8V8qB7A0vBUD8ia+rf4kJcCjBQuV4m8OyK56LylSpkiaVbz
/3pAH+VM2mP4mWv3V19PePv3nZs4osMNDf4Ckc8swcupXJPJHDZxYjSNxJb9XkQftMgAJB7Enjsa
fFleAAuCLpTEHCD1miw8klBZZ3RyR9GC/U4I3w45Wetlq35n4rQLhnJwOQRGhVYIacxcgBPdTHAN
c6Yw/0egaFMFK14fUsYhckfZ0OHTyrWgtl9FGomxbCbNOxJ8TVRzrvE7S1AQs1TfO4ZIyxfT3spO
A5jN7PC4VdYIW6/shFVvOLsiQwPxvFS5By+JMh7leF3qQ59bi91lSkRZVWDFDZdi+cNbIeo+2d2w
Ku9U0Tycs6mWUQ/3DySOm34/o7W/cikTYA/qwPub0H7odMSi4+tTE6XYR7GpJRCBOJT42l5YT7zI
AjTLwrVw4lO4ptwzQMQkwHvsvmkYKDtFm9RnFWLCoI35x1vEDEv1qtY/slq53y0QtM5vPDU65ISf
DgDeJFqo7z8r3e0rssqrNBwt1q1Webzu3aJbygFHFmmMtNGUwoIQ88aMHGDcnNSbhLWZZKA8UFmC
vTVtsn47IBfWTppWmzgtP3vsC97/nLiKKnqx5Q2S3O9dlpqzkYXrFuJIVOSh+1goauv4doKcDGQ7
vjZooFq5sAF18PkfJ/bYW0J/cX79ANaFLr5m4Q90xsa9HSVk1LrxQL5Cqwe94motnKJ0aDqfRv5I
ToazN5bJxbzhG5oHcipJkMGkA9bhpd/deJg9H5RYE78uxJo2Ymj2SOYANXLpmvnLb0k07133Tsx6
Q3XFFmU56Ac3i6+87EtAyRrP2nAQN5/rEsgQsMWFG+mslc8PejA9YXCAuLtapjVp+G3ZCaye3GSS
X+LDG3zkxtp4JyaT1upXL8XouSrPkOicwFGGcqxDBmD0Aib36wmGYxoqgGxQJbxCISvQgvdE/2Zf
S83Y4YHWPLf0dRsrAetDbICefxQjrwibeP0s7OSfqZMNwHGEvMnHjjIL1Ap26EeIej5pbRFFEIPd
+OBoJ2DC37q+DZNoOSGnuDINSLGG61y21aPXR/kHKN8BcoIivfoLfj6LcVwAxWkeNuR0y14dcqxc
TEFtwsCHCMR0iQbJ2lFQLlaj/Cquda2mrG6aYzI21ywxccG6236nmClCKVzt53SsCWoXGW3GUegq
vl46NooOtPICY09rgQc/BS92WbGP0Btk2wL3M1887vLpjfJ7/HOdYPLgbYfs1I4hU0SZYZxMudwD
emF/Mc3unzQjiwsi1/qlKjZznnBZ8tDsP+SjyautRBNw2wYjByv/TIUoX5MT1UsOh3ltdd9+vexB
YfhSUrDCsjrA9HUInKwZtJoeqfI2Un53fj4UevT+l7LCoEW1BfZC2GbbnIl3+mDTtSrp8luTkMAd
4aL4o7VPMvRKWCKerskdVQ4BNWw+KxhlBdFGX+LJ8SdLGhBavJ6tG0cpc55yYnoFeAe6i1f0x68E
80YBkZXsGthejesmPqg7IT51Hxg/+g8gXgdeY/9LsWB7oXc4Rc2WgLCNuB2/s9DhPWRurtVr3os9
yTl1dZuMdjsOagYV9fDLdNJtsgOmOw6KG+TY09wiXMFctYhzbdzWB2H4v6IQMnm5OSeUsYRNiMSr
43j2HNDmgem2QMZmaBESr7eyz7ytw0d0I1gvBmS5bCgjBhHjdDrxPbqbdANI5QUxkCZjZ+nvR0eU
NZ0UlUNcIkBbZbYJEDTL/AKZILtL55tAnPa7Rn8hp+/B7WFXs3MWiXdj/TIyvYiOgOYb+XMRhYh8
X7G11fwrxINjusfDYw93utgtt8z0pe6PSaEivWLC17oE1X2wYBM/NEQjZONBjOzxxWYX0i5mZSot
knbmdf/B7snmdEWN6DYFu6377BCTfRNJINk4txNKINNuMC67JDjYqQSBrxWikeQMkIqTvmSAB7qA
pyq3DzoC7pb2PZ50TYCCIz+EHusTBoz+6hQ/2qaLQlb3KPLcPYIN26j3pDsI4VrTI3Hp6kFPISeg
bNPAOsZYOIHzPyo5xfM6LUH/cvW75CffeMVTx69+Bjivy1QsdNhqM28zzf8VMBuF79ROe0bjFESP
DiRF1efFBeOUuYRZArblob5W3ud3KuLbEH8lDmO6xgNV/IqHLrHQxtsX7CRn6pvlDMuvMjEwHJOL
TDN+ZUeCAK4VQSwlWAbtmkOKVdpFxQsGB0UjvWAVXcQKPNMcSpYGsXV+axkfXxusffnuVN0eQySo
86vCOYTWXTo5/4oAQHFIFJbMGtoICwryqHLdwIfPNDLoHIBS+APN958bK0YMzTeJ5LiCrKeCI8yh
hmiMWJ3jy6+dTDsjv6GsM29X0GGE3WxCzB7eNk/t4O2kEL8z6t8ttQH6R9XUMnXjqn+FIJgSsiA1
jIX5F2avnGuas9dHsyZrurhWQsECTpo3A0J9Ntz1j3ZGbVXWdMg95jOIY1YznmCjmO3RiU1cyJyI
2X6VqpP88qQ1ucvfeeDqH/8AMajgtKhB1wumecJUF5ikxg4B3klOQ5S9XWc1yCjVwaQQ/nlsxBhX
s67OBDG10SQS4Tl6TEYnkaaNEqoKeMzVm/JvjY9Q9j/sbX0O3gBmMft43RdFsPqTrLs1fvbgOJ03
ttnPpP2V/RPsBy29BU4Q5/dTrXr+DSiHb6Ym0D21r+d5dntgZGSa6nc4C/s2CRxj6K+G8vyizJCo
XsfViQP7z4PmXTs/NfPFJi2lVTiOzagrsxsbOqXw1lwT2QBMVZPrfxqGoLM79IcUJ346U5jOPVDe
iVXc1JkkFEbJiY7N66ZG0hqM7QiYF+CyGY+SKwSezHUrWXZH1m1LSMY+AB+3c9oX1+DW/LIaFSrN
s5bVWoV4XDQuy7pK8XIo9QboKo+F0RcfvbYQCP7cHGbK+pmr6TMLaNakVokNnk783FCVYX70IbDc
6MKKyqZ/qUxsMbP2gWzPvM9nLu30n/Gt792CLHXMkPjiioKjUhbyof2bW8wPf0thUG5A2I5ncmS8
9c2//QE10Q0qiaPYc92uNz0trEaF25uAbLHNmWdseE77Y3wkGvoZ8gD9+O6ZLS4CrALZ1EQwJrqg
loh18s4fRZDEdKV9xPmIkljM5wi8otWz2rTU0k+9ri1LA+5qauLLzrOGr12hQ88z9UD+rZjjs+qY
thUQKILMG0ZjUWSWTlP8ZQde+q71uMcjnWwICy2E5aCuoPTdjXvvyMILmS5uxYfYaQqfLQqwX/S7
aXYNCc5kOPRgNvNnzixIrcvrGloyxnZsPe1GBSkUimvm2OA2OMx3JBRNLhulHOPwuzijKWFZMN/1
/lAAxI2cnmWNa+qEPhofCBFkqX+9CxGrqSKt8vnCQ4t5JCRzWvqn35i0ROUHAixchCIwcbRCAOqm
fBTYsQhLaXkYQI7auzjUjf8fEXo6qGONaPjvSfs0qOuERSywtFdUTyXE0kXV6QmhO771rP4Bhw/N
O47nOp91auNqF7wuSe7o93gZxj0SsJkfHuJJKRLWS0sSXXQ6hxHwX09W3wMEjQlxnqDabKJVy0OY
Xxi3/Y4sdag33LSFuDXMcfzI2guHfiQoz0uEMYlgrS6WjMWCa4NFAbMcPsadQA4o6WjfSieTtVPf
jJI3uo3JiEj6asjH3X6Zerr26yLvDUWjXBrH9ksEE9T8tzYXOVl6vmrFwmAMp7PEuLGkhhGfcqgg
V++MWQQep9HYuTrYnn7d4VbqxC+Zlt30vkMeb7mYuSi3L53O2mKJ9UEZUyEzFKHDlwdfFWarltNo
2P/U+NNo7lNAfg48yl11Afwdw633U+Ev1sVHynaYJClU99qcxx9z91br670uZxA44dh8JnnjJU/v
zKt1z9CDc7tMdeonIlJcvLEcseqi353JHMkyvz0HzmQcYK3sKNXSNgUJC69xiDV2yNBP/z/F16Qv
cQw5q4fQQzskmGoOxKekcqK/upPNpb62QEI4eYGhQf9DPfuDMchDrB+fWJONBcFDS1Q1VJ0JGkAl
oe6g4KOuwR90tVCS2As29azi87uyWJuFupQCvK+fTK7gZwodEGfT2J5n0C6b3HVRz0f700MzRO67
Lo/DPHHV9y76NY10lSQAmlmY89s/SL8Jh3CiLOS1RT28ossqkk7M68X8fFy+DBs21dQfbmjMZ5k+
cTtdbgw2sK2enoQkbM9j5gVcyWEiryFg+XlPrbSzrYd+OCdxPukPRW9VEZYM0RpAhhZV6uLTCTLV
UPnfCJec3bsDJ0s1PB8pbUc+OFnopM71kW3OXFUR70wC4tCimMcgyaTMC4ie+HmTe700CEdeVkYJ
CoHUroMe7u5VgYs4ZNoC2m2vRGp2yWl9Su2vRAr/zFb+VRX775aZnJrnf/WONeBF5x9PsnnvB9yy
2zySlfpG3suloitGAAw4Obu5/2cCpRzZpz10MTE9XNiXxxbphnNritj62jPcVIP85dQBvq5+2hUn
faqIQ2D2bIJu/4g3LmV9C4s/+CPzHwt7L5lEeKqjypyhHmO84o2RHJ4jMP/LUbV0zT53R0VZ6b0l
svgO5DjlWecDIzSHGIkAeeEMcRUuB8hu4FH/IBN+kyWn8Lb6lnuaY8BUlbnq5vGoMV6GOSvVnc2y
WNUQjDdd2oqu06HrjZ0MVGU7sVjXBGUdwmpzK/ItoMQT5iNHCJ4AjO/jeETJZBQ/OTrfbOJhxgVM
TaH/6VIqLcHV4wL3zMUftqOC0/BIT7XYX6JyKpAK2Qcv/wG30lVb6NnWbdyxN3giru/YLdVMXNkn
POYrRbEmLm9gvY059XWE8HKeODUl3rD3bc6CMXKIydtEFiTvqC/bgllRg6ieFF+km++gw+hSFBlz
NqLTOZzl4fdnoAhUMIiimoMTSf0sqrZF+ZGGEuoToIqz7zY4NgT3ZpAAMA/+ppCyFOtu4HFeJmI8
d5FHhSu7LkOVfFcE8t7ZODEvsbdzDDDHGSFL4w+IMZt76UNFmO0nAApkGvgEtoP0qj9E5JOoWgCM
0IAink02UqJlOaJIdfzi3ZrV2ObN8tE9uIbpQ7NL5bWSAdCet6Jbvss7H1hOWB/9y9FRH5c00Dis
+SK4gdpoM/C67Kw/4jylslWNYCmMrTRY+ihLr6FNHfVLKh3MpuZEHMyaoyjadNdX95Da6v03fHxv
4l0DT6UfPD1k4U0vm9Dv472pQLOz8B5Os/yxEThHhxo3zCq5ffx0X5exZcP5N+EUOYi5jG9dXcUJ
H+Xb5BFgb5eKtGSpnKaFvrDspQW74+WoaGV8BcXvqx3swmJ6MziOFCQRcOwRepRTMzAPemFRolDB
DhHvR87ZXS6umzhurppXEItbR7BuEKFpOAZS5Q8wxcuvmUkKD3ZfY8e3ETlxEpSixeqcs/dc6o/e
35GDHJn5cTwNCeLMOMART2v+KnC4yJfnVlClMWxvhToJut7OdXuy8ysdEoLIY3cLtCVNpXNeqAtg
yAheXZ9aLyceOVEW29Rl0AdVr3X2a+CeEKsiz9yCs6EyYDR+zod4ioJmUMDeOr095F+y80yg0BY1
Y11spFXnc9/kN8EfZtCZfYw4vT6aLgVKjdPQisV6Y/zKI1lAh1Vs9n891GaC6eSMpFJ/CfXOGEIb
pgmtrouIAtf7vANIK99nrabBYVoejgxejZvALKYatms11ROC3jt6jCehS1J7ZxUlDEd1fCBvGOXW
OKNkK9pJhXuMsMyaKvCkQ8r+PrDItlaG5rhYq5tnrS/gVCXMJDAZDyoi2A25TkY2yA6YpeilOWiY
W9kvPwoCuzU/f5NRHPLFBCu+g35G+rgcGd7ZXnzZrB31XVhgPGFRSCzlXloy1XReTlpr1wMRWt0z
nNeuA2m7UMurxsOZCExmxAAN5Caq/Qg1aF5RQetnNl7XVSzJ7tH/rxULJC1sZ5vo8xI9SL+6GOpM
/IJ/kGoNNYmW4us8EXXILoHhrQn3KFlGtG9idPSpwxdi/xhnMJ+0fReVw5R+PBZLvxaf+0ogk051
pa6Q+/IfQH7A3VCsBiSL8BIlUE/9qhnETFhjgjl60ylDctSVCWRVWI5LZ2H1L3Hylpyx/kyAQnNq
GH4p0tfTDR5atTdZE2hxFeWT8iMH2i1D0HpJBbp0I5iXjCoZAR01O6nQA0HulDm1ENKO5VBkCzB/
S0D1h+/oIS5QXkmfAr/Ew/rXFnu51xEW2zOWemZJT6sF/SJiLKvffdD6nFCIFykKCpwDlqzHUw6j
wygPDf4aTJ3ruFpM5iP4M56DogWaVTjFT7BFKuP0jbAN4Yp64PYbR+ldtjxqyzQrb2kX3mk6db5j
RScwValvy4JE4evGf7IkmEPonZzGDfBD8l8KC+Ye4GMB5hXyVTIjt1PkQUBihqRKg1Iui30xfWRU
sN0KtlMrGgFLT7E2YNZAwvGs9cLy8CfdExbr+//N/cTGem+WSw5aK229uQqhFnGl6Lc/KfWpcEP5
8Vzk2tQiTaLdswXnBQp0X+le8/OtecfSdK9Uy3X5afU6p+c0giY3bZsjw6yHOz8Se5x7Z/cXuJBO
aqC1n9+54y/601CS9HSGpLx9yvQ6p0v2SjcGMhokxXacY8V4vAnP5d5bMAWvjD9tmm0+KlTfzmxl
IdKvxLrIHJc4E4JaksrQhEztT92ZJFciWQD8x0NSlY0IVXd1WRYgUgdQf/tybFwV21t4AkRakReN
IfHKhcAuLLsALT4B+sPMcEwuWfgfneRmYZG6S2LSj0DE5bP+YNRjMpdpie72VaE3D2B56MTUFauU
PfoH2SSBGszHJhKNn0lhqJspyZi9U4in66jy4z1lOZHvW/y1EZvtrSpAnMviV13yVIR12FJ4Z0d9
oTYU1EjW3SnFSw+SqyniMqTbpuqbSTsFNIgyebJwBpZ+WFO6wpF/Olua7stB4dMtt68x+cQMGrJR
sUgjkTjnHLbIGZCiJThxm0asFCq7wqEG3vLD/AId54JZua4MWY/0oe6WpLZxq6kyW6iwewBP73zT
Rp+AjwW9RVlh45Z8K7PswMmakZ3FpzLYOwWADwtEaf0v/qvSKS5Ya4gjW7OGM98+oRf5OzFTmjnF
833u6QgGjG5BIR6AWblynu9UlQeOdrH3rQFAbLp/aBKME33ci6i8NbtOzyP+EiGLzPK+5PX4HFJr
GXlK3Dx5ie3U5DFQnLWk/8cw9hE1Jo+wStilRwX3aH/zVMbzyZ3t72uON95NP1YDqXs9g9T8AjuA
Mwe3JMw/8Gn4i5sq1rDfZzwoR1CLuU2/DPiJ0TohvYfSmWZ53iMGbW77R+uM6mV1RDaQkJ1m854L
Wv1+ksKyk2UZFKbQgJ7Lpkf0yhqg4N1l74r35ZQK6SfoqvRCo7hgrF1yDaiPg7OG/bt9YQ4K9C1Z
n+fqisEXJuHwJI1y7GiSzPk8wbfWwIslLnds621UmfXA+Bikc2+YwV1quOzNHtF82rHXEtRfXfuE
AwhqMykgTbzjFqVj1SPWqKumoB3/oRd/4v7BVqvaW92cGfIE5GMEUBImgy3z2mKO6TXCmxxDRMml
+V7JV2BQAHXb5qGY7gTe4bFU8LHNhqIrEqUCqNZLr9cMY51W7YZySr1aPK445zrXptN/ZNKGxtae
sNnUModV6fOvGnxFAFN33NxqPqjmAwmh8ug+YgIuPZp2yb/Z1gAR5qkmCcEF7xz8dj2bWN8MOD2y
KWrAPI4K12cPoSDUqseBP0jrLncShB1OtwuoMFRRKETzB0skSTVqpvj9dzqvZl8sVwmaQdnp5Ns8
Uzsn6l9JFjNsjTR6luUm+7tVUqLt7Rztbmx23a2zkJgkHreOPkW7JE8+NmCN3Cwqg9Z5L9Pou4y0
AHzgsAqPohgEXGw2fkOOGKI80rOjrQwNXOh2vnn4FL2hu8I9ZLEsamR9Aqhd/YQ8bVW97s5g9V0q
p6oBZWUNbKVUh8EUjv4vf5yK0ba5T9Vemzt7G/dO27fuStmE3obyGUzKJkke0c+JOz2T/2qH5Eph
p6ljQ40vqc3NfGKThzk1irRs+xkL46wPGf06USJNDm5RLvrnjKy4fG9rgt8nSReW3DYhIwzJiyM3
oKYy/GloSmsLKK5RY9nXsJlJOe4yajAJlijp0I936lZCNscwd/1T237XZsmhgqs9cgeGZOH4tlsz
qQc8x6nBhOzwNWjhV6LHdCd96jNgJvt5qYt6k9DP2sLqVIIW+zkzNGROjsyZWMvv5ISFRbfg+A8c
0y3Xo3MUFdZhbVWPZ3G1GUEiIz3yRR23NHITFRctsvIP628JEqOYJnzlepSne38ozAlnbF44LYTH
z7L2zkDw/yjDDNBi6UFB9p3rqlRd6HZvU+CEkbCPoqmG6vOCi5nDyq3Wqt6leHrsj5C9iaXCHjCT
ATvqTayhx+iGMp7tWyM7UeDPdOeA+dqwkvYGe0mmSvWzoOjoKk9rJEY20maE2zgKFfjr0XZOL70q
WMmSTEfgAQXGGkCApJc0S481UdkIRvHNL+rrT29fqC3YiKOX0jG99UNxcamfadELIK8u1YZPyz2P
MedYxIeBjjYIP3YXYfvUXs37id7rozRRQ8rO5BHXv0S9RQsIdciSa65z14nXksLpxrRYDD+UTtyS
+Ftixqe+NAaIU2WiUC6nZHFsCdjbKvLU8v+66KhX9qtNq8q5Wxf//nYt0XO1fk2Hc5PbOsh15wdk
hC7TDkmalTevnkL4zCBuV9qijQUDExzNgb1ozXb87H4iJUTWmoLxm33LVItq05L1q3vUjvXiCN+E
VoKVGCgzLy0eoeWoMcIhlNchfGDZbBPIPZvFrfq++IeU9J144V4SQQoVvkMPu0nllGxUlMHyYYV6
8NkIw4X1r2zu6ZFyM9nkEKPb9LmGlelW7Duw10Ai3U5aUxc+F+gRUQ4VNDiuSsveAt2cOuOsx1Ob
5cwcHZZs+hsOqdHgRx2cvMB/aXDv1f4x4Kjas/mkKJxVOop7low7s96tnONCvc4ffb39ag7TusDp
GCeJcxmz06HKALAWToG2WNtkTuaBRR6P0No+2/CMJOgPNX8+0Sop6EmLZFHNO2+c+pJXxEbeISkO
VJYv5RlwgcvG/xXHev4mTHY3/QoKXuiwyQUYW+iQ7+0zyatyY155upcL31Xoh+GvTT0l7SeyopTI
HUVkzOyzikaF8m8GrSu19nOGibIea5E0Y2gOp2PSBA6rDKNsyzsU+Af8gHy2g0AvavdI6eRq4XTR
qVrYbV7rNlQrvDsCCJMTd9P5UoGrl8OaGLo3KC/0m3G8Yd3bkHKP3kutzkz6x8SshN9jCwKwAY2f
d6v5SkKVpfFOJmxTt4Ft3xuwWa2zLRF7yc/JCtQqsQbD5hpGlzeFXVS/2bYkNAj2NypqCZnFad2L
IkMg20IPRVJhwBnojV9jEPRwibPiWr4779SCLkPPRdr4ok5OGEgHPky6lkMyyuRJ4eie/oOpFEhg
lqh4WA2hhIvb88lFZ5/kjruIWaAFP4R3DN0tgyAgUV0diKALw/qa3OrTfDC/CLjbhYbqtfMN8+2d
ord73bw80nrf1z7PNuYafxYWmgUgNdTbgOmLisd5pzJyBo8ikdqWTyZ9RNCCLt8k6pilsrdggJNO
xpYqoftgEeFIc0qbJyPRaT4Rk9D6eMbzD5GdXGsopjjlCFWr+80XCgXaRJpIkKmstKLjNXKW6Esx
D+SEv0ZsXespzcb7cQRoftRvYoJceHlpXKZKZcYhmfhdyX/enNZjn8OCLnFraV+AV2XI+dRdwroS
pZAG5ruLf2yvxIF7W87virNPxfwvnas1uinnQrKz2ZxMDvCNI51z7e3uuSsjxhYOgGgPVt3NJuwo
RGCi0OjZ4SgIIs1vQLifS2kVg4olHed7AfKwjhKT1vrGKYXzzyObu8qM1gKk4LziThZyT/720YMN
SuZrTGYHGqY2GEWVK6UZfRtwiwx5Fwa1Xsp90cTFQhwsWuNX9UaRVJB5zBOLfDWfIdc9Cw3cvKYB
Ec+ZswM0iH4m/9E96y0LdFknQahh+riz+P08i6oH3hQITvvXck96DR/Ch3H37cH9Ov6XICzePZtr
y+2qI9S0Hft9Ntqf2sywle3evZcQxuvmDzhKVzF99fPFvydnwVnWZi100F5lMRHunmrWvl1OUHrS
asHyyAJRaShfhIUq7U0ULciYDmqNl79V6vru7R6lmVjQ0ujyS3YABee7iDejpchw0gauE9Zd1Mc1
1deLVazF4nwmCeinqY8+vM3Ro52ofnsJSUbrGKZ2e14jqcgJAyIVY+/QKB8k3G+9X02bFn/DW634
Zu0tTRuvo2o5ZDx/jWS3G8M0pJFUFG8D1y0PSGcimuQH8IJusodvsSVzribZnFsKRuREb+Zk+YLR
19fXIj9sRmb3p8J9eS01fFmqcmK3LBHJO/5DlD0BpM5G42zlF7559HFXTn/HXswrDqhK9Ah8CTKQ
i5O4nP63dlEY7IFcxdAavHQzvdK3ITb10rigCs/z7o9HLgYirqnuZ73QV6zihB1wiECXDL6QoT1D
18mLrE04BZlGCmFKQqg7EbsYmB08mo1eM0RbGRuDYTRXN0hTuKXQw72z8GPg2fBtMP4llMCWWZpp
QmVSbkb8t3SY8thNuHen5GOS1ExCFAphdES3VowMKRQ7VzsByiaOdzMCe+F34cnj4mgPIH5F3T6w
LygZMQI9D9xq+PwvjKJJm0BKtstHgL9IHtmrvN7VPshL+8WHtnNL4rtM6wh+35Xn4NC1ZNL503xN
Iphq+WmDYrrTWJqfxY9f49NvzfTey10EhAdytkhkWwrHs3smefAwNcNGNqJOLgCtEZRukfg6xKOo
vaZOOBBxQhKWkAVqG7OLuuDHt/Ia+dITTGNVv3pjcZ+z8s/DDUjmQ+4KG0bwSyLgjBiUQnaT4nV/
lLmuS4cg0QKNuBTNq0M6XQakuH5mN2HgzK94MUFfUXAnCSKivRu14T5De90JvfGkU8C7IRiI0JlI
OyBklia4So99ozFesetEMf3+5dXRzKj8Ebsbjk4leftkbjqPMf9oUMu2I+4PnZaDUlsU1syIiRW6
Ml4ZKYei5s2TW3IaVq/pXnCUXcHJ6OmB4EhLJFLv3pYOiMmEzPtF11Yips1zXaOc52za2U1jiaxH
OiBTYQJ9uZKH1WLbcCKGllQHewS2iQrZTO3eKO3f+v0LDElK5s5FUMZ7BzQxoQX7kRYUWw0FKyXX
lWLzP8Kya1plPqAl/BeG8DyUbXxL5qb0f5D5hcOidRLXlLp0JTVZMKCyoQmihy+3PXvyaihTLmx8
EcIcZsTxXTD7w35zJ1ZXSn0RNrZp3haAGSwKalLaKTwvHjXtNo0hUad+QGIvfaNWupuLL20Keeyi
Ml+sk9l93LihKh5HaGDPjbf0XbrQ2/Ia9g/lEWj28xhNgPn88fmvh8cb1qtdS1z2vCBXkTMgf07r
AfORKOkC8OeTUxIpIRJpG8P1LMS8s516UOIov0wBOoXMTeDe1eG+u5VgEcFuB7NdMPT/9NyxPPor
Z2ExRY1nnpkPJ814YnOkrQx/wDd+H6gohaCWQZJ7oC/ceNYFbcEFPgEJ1i4Hc8Ui96Q2wC8Mxdu9
/3hD7kc3/T3fT519BnyGZBUEJDKnh7jBps+2MjFH5h0hH1DCskfizp7mKIpufilkpCkpkX7nvlRs
UH8LopHucmoMVC2elWupS1QcWncup9lYO0QooPABVLQ/Kvx5uftaOiZBJtdXcXRxQBryvy9Cqgzg
UT2Zv1PmzVYtjpgZyqgTdT6WaSo8iGklNpfVNHL8BIeORBiikHDVH4IbnckLyvXEpVBnXyQtZG4X
/6i+vWlTLrPhRJA2cfmnfhR0Wbw2Us7wqlRT6z+INZIEBFMu42aPw+mLVPB/WEI3IyDFdBngB/TR
pn9auxTVBqCYw/455jpnAVNBDE8ltjnN9Lf98TlndYx4JkTXJi1anKxiTM7L8rQT05r9RAc6m2FJ
IjspYNKMEyXXMf8aLRrtXSOj6uc7lHuqUcsYvrLZ8W+dPzoQWiQLz3pzjGZIF4Ne0TTDmgJKTLho
cDaOXdA05Af6IDpp3iHdF6NkwnT174hip++MGpKHwR2Eob/NdvBAuz9y1uRI+mqMlINJygcBepGw
5sr3zwmgr55mzJUNp1aGKybyAvUNQWgoi0nvF6aDNnr5pl7BqBD4+nV7Jo6SQaZfjKlnv94Cfy6e
BGRtqhik5Y72JOCwsfsqiFNXeflcsTxekH1ge1K8TK10JIK4cvGbGVmBmUW2kgz1sy14+yVWw/K8
Vp9k8UAGJ4ve88oTGiQncMN4eTJaMT0YFsE+CBxsabQXHhN0Gwm99zXD4Hxpd3khYFZyqcX5jkoY
K4gifr5clGj62VtvGFS4LZd5NrtIFMaiaLyH1506oV7G3s26xkaQ+gUKFtDbVJu1JP/jilzol2bC
PfN0fxyo7oF3XnONtR3qHi1RWHE7RBhmhkm00nBeONqiK1eQqdQb7Y8T3QEffM+TwOlGJRhKOpKi
V27wYQW6WHgdIxOSyA3XVd2igNwaHGy+r5FSBgCwd/8GoVcIE392zaMfy1a9TndHn5eOLtLCrIsU
R87DSsQqyEYUrKqmARSusLJ3LtAr1N0oOeIDuRryRHw+gs2Cg0TyS2GlE7w9HJi3C17sPFSVbbRx
H8lyda4m6vgeUYjlBUhRn80DAS/cfAy9jV1IzS2YhEaor26xcEVnzogl2qy7Us/FpCPhPMX3ZnH9
I8U2ES5o+TnQROwSeW8zaLaDHklhX9x/OCG14IMbdTHnNawwCr9zUDIvjIC4q1BaB5PrPMFoRzGo
YWXjIfx2ABxsXVoTiZfN+qKK2c5RPOEXwK2N4uaz5DofLhHtMn/bQBr2M/LVD3UB+42kDnXjeWAS
JZRNnc2pQCxxd+9di1ul3mwDZoEad7rpQhWFHomKrLhR4NZMfDMqJ5x4rx6pnH5TuC9ebmsh8BiE
4o/tIjB26gkLILv8q1wu3evMnR3iy/X5Qg7D0TZcDjjO2C/GoMlrhuAUjx2f9mjKZuF8t4Ha90/c
qhB2SswtJxI3gEZivwh7vMx0y0+6wtI2UrvROYI8mVTk1VtU2c0vyF19a3IHqhy+F3BL/WHulqEC
Vhcll5h6UKkulglNySzYsmTVXR/Gof8p4gvySknZh7UncfhGSISyUYHk9zXP67DnQOmjZZnVaO5Z
P8GQ7FLVKUY8KoKj7TcI5ZGN7o1P2xbxYu71HhxKnCFo9c3QAtcFUVP9lKAFkVgcKaNCvAqd2gKL
D5XL0bP5TTKQA5gIriHutldr0Rt2Ywxg2K0rMvfMuZNFisnY9cYnuyVH/XVII0AthohH+mkVQqyV
fFA3EQuEjkxJbz1QjCmzZNto/fXp6fXYuKKCgRgIdLoYuj2EfRQ+uWyumuS+lvilTcsSBQLEdczj
2Rtmev2jThr5vP5TYM4t+qxG8gwl295K1iZfogeVOcVZRp2neR0l7teO0Vr6y1sohf9KvwON65x7
ukNtxo+1hDxXPF/75RVsjusjtFaEo+jtu/k718p+XAOF1gIHT3OHlWNWpeH/UukkbOu+HYbrMlBR
i4uqOTI4WtsDcaLi9saF7f3wb9wKM9q/Z4tnp92KFICLEHHz0+3uWvuv3ae/Ag4sleMEfQ7WsrHz
Q2OtTEbmstbABxA7lBOGGZ+lK+UbQ2KBf+oprcJ9luDC335dwihM8yS0UnxSAD+3k6wH1k8ZYZbT
adrNapvs9bn3EIsq05y1uKo0M7N5aSI+9O6ROvFdlPsvQxWadA+9c0VX/gSRWju2D9kE0WsOc3OW
1NgCjUkhIDSbq9iyT7YxitKixJvDE+Pn9BOAunO/yxnV6nltOTIbADPPllGOF0Ow5Uff1AiFkuVl
DZoGRpgU+HTYnSBzZ4+7azvGYDzcos/U5ZUyX5/pywv+XWOF0s7rxaNp4FlVHsqDRhEVyuA9eVDP
CVLUMQylC824IcLmszbYQy0RWP2UWeKtfjcj9D5CzDWQxQ7PguSpSyEMQ48/GNIcXbqHyW7eAyNV
LkRVvyjFA0jteoUFHpuaYSDsCRnc7gvUvZVohIxU/RzwyikLc0hKOTvNt32X50eXefOOfNf+nHWo
V7Ml/dasTApHYyM0l5fvNGTVaUBOML4bCG4AkFTksCm5EFdKwANQQz3W8ykLeOUyoZrvmwDewEMV
Ifu3jPMG8cuPLXj+ChoqPqcigKUe1s0+Rxjf1Z6/tVxLfIzLnSjEY7CnY5UsTHToJnGY/biCd4NZ
R33lGO8mDzcwZV1cV9QPaBEdkl6uimzdHc3mGO86rI0QBZgiNegBF/+glZJ1M1i3whaQ6pEG3y8Q
WIqMgOEsCiaBJ4V0a0HBGe/lae1+JyECivoIntSa7TOtF1RM+ugPLXFfy/BW7ORHVzV/RJJwKkZi
pc4m2oAKwAzC2strMKebkuTuN72YOiuc0DS5wn23TtLyw2DGPdmfbdceAUAQwUN2+40evT5gZt1A
rIS82Zb0VUXVxa/Z7pVFS5WSuFilI2iGHLKUWRHcdPS8ypfUOPx4AYHLGcWzRSgAAc8BaOxKhYk5
inPpOs7Nku6VANH9cYQr+jXLgbXoIBQRB1dma+z3APvIgCQUo/xRjndgrghUOUWr7RvgWwYZJJIy
JVCXZ4QAPDK2NOx2Lclyz+UMZ+c3ecwQe0wvHAWUjJMBPiXJ/7vc/6aY7kGso9++CjybX3Dq/VLS
KFA7kop8JPDdzFeUaZlcI49RifbO20ZPWC0BzrrhnGST9pZ9H/GwA/j9OdjY7dAGTfrplRhrnA9x
7rlYm2oxbHEd+/Jc//uViJQ71AI9X6FAfB6IMNrKJ5bthkF1Jma3ymGYnrhoYXTiSzo3aj99ZsYV
HzPb7iCr6+m6qO3b7JyxLqSM11Qj1EejmPjDLrwL8t8SWMyYxGpRRCDmcUpFKjeG0KOPxCfMoUm0
YhwbMHq2qxjHqb+98JtkEAQUWxq/Tu7GPKWT61Apn9zhOq/oI1c6CsJGFnI0EVsMGCU3tJbcMAbM
wYmBoTS9M4sJQEujE09DZryYj3z4/7gPoinHRDpjnWQrhUVo10HRR/jGaZpf/K889eM9FVCNLSl1
seNwLXwhgV/WjElbB0lbmEpJkDJf47WTO4nXW/MRybo81//dvYT0KU40RyXNA3r62ppn2PKyN6xA
eLVSY4jDmeL8cmIp4V2gP6Oxki3OxbyM5B/EBApdOb/K9VnmIun/1d8iUjUBHVQjqQ0qiLTcb7fv
4y12rjystMPBO1OO0aWBJlKQqgzw4IFwudkrIamki7z5k63MjEPb3pD6+caLIKcIzrnNXH0xDK4N
pUQ3iPqA7oaCGv8zHCBxdNYU71eY7RbWM8C0Fm7+Y0N/77aOQLdx1QHM6chavmLCw0EZYkZ/0Sfl
1Yl4NCGTwH5BFGTX1o4F4dOmeKSPD/8d6/npofZyS8OEwaFNyT2uasZZOAaS9yJcmqQmPTzhYX/z
h65cvDgsxpfOWBilSRxZg4DQ5CVlZH4CorBTTXHTRCg6oDz1FQQzz7Pjz9hVTb/q9Zq57rAyvOWX
pO6MwwiyNPE/wJwkqzwObIF7sKoaboIcGbmeJju94athd0hNdQSvLlzt4Hd9i2V0PwXIRlU+c99B
glfvOvgST+yVeHSbvFO6b6XsZKaxrHdRTFCin5Ht1ugpC9jxd1bPNWsyPeG9ch82IL5+g6yyE8PU
VftgGBPrWQWJIuYNGRjxCxFlmzKrSLJIawfij/zRUeUfmDwlCrBLdVWm/LsaK8PcyVBiS0146a07
mroSx+0P9rBT15Qy+K5ueklewy/wlZyf7bgxTeFpz0aR6lX0OBR52dKDCWGBRDFqaNSp2JBli4HC
C2J3G0MTh44+mx+bi2rzc4jxl36swuuo+U0yA/6gjI9Rqko9TaqmoYPBq5ug0MVQ2t+vhYibp7Oi
pL410zH5fFE2EU/PDODb9fGSKbo8Wkp3hvnvc9rUZOsHRbQLGQnbeYzC9tMYz15aD6g92yCLAX5a
Ij7iruFtbzUBuMy9WX/9aVpo9zwWFXHwD6ltNJjqH3JVG9CL1Rut/tTiCUAlsONJf1hjn3c/1JZV
ggf+4KKkItRXyY3eSlxq1D1v+AZQB15pNd2DuIYwEr4EBDJw0+Jqs5hOJH+2BE+h0FXHWEOG/wqr
LGSDz17UDlTwiIWQ7BVGFzUppwF2m5XDpJMx36rVxyhvtZOcRTXUPexegWnn6ChOB9eMLrW3DSnd
0qmD5D/aLDGOK0Ysa2EWthEu3/MWVXV/S3NG8cNyBrOw0/DoE0UAOPPVKVka01Rmp0FyiXEs50r4
pYG4zQb/29IwCaIHXA/CVPvnVVqJZXoZ1utCfP7dMXd/B/NrZ4e7V/eVjFji5PxsEj8tNkaQye1A
9kkNoWmMCoZvcpE3YR7aBf1UdhapmT0TdvT9hDNOkdGjJ3PxzgdbF5zhi6JtauY83L7cypPYpUs7
S1rC8lN0QhY7XW8ZvaDFI39+2w0iscAgzYWU553sJVN+iCO/eGVCl6ZtEjx+krkSk2Xy0+k4aLhW
MA22/fJgn0/L8DGTRS1nsmCCaBSnpx69p2Yvvy/MhCDPkkXj8Y9rzMU/MLnAIaNgKGEXTPSMA6jE
N9KscyhUKHAqJ2rKr7+1HeSaUidiYfKkM7rHhG8qddxebp4DCVkE9v4cOtHV6T1Z6GBZMRRHuh4p
G2mt8baaKBzyH36Yb8ZdKv0GgTsMxAtnyxnzcSjP4gT+73rOox2S/IlydA7IkWqHiJ/2ogXroQPL
cDv97dLXdAqqOOcNp0HIp2MVdPS4tnuotBzBSjV6A5E7ezw62hELy6H/dAcacavaZ0RnetzG258h
sSIKz1+GPwGYfYbEGaybdnojybD3tMOTODHZFyZu9XaNoEc1O20a5mQULm0AKeBxwnCyXyOhmyFM
g6BKYqw0mWFvH6pwTvTe+Nj56YAIeV6pxPCd2YRldlucSYq6dd0mf98t7j/qxpNuoWyKInUTa6bc
vAtoDKxRYxHnuWXUDWXGyJTt8wc4OqcdNnsUfzSCP9/H41SqFfjBPg/DR7ai40tNGdxyHZUfAbuV
7G9vQHr/656XECJAwSMxL2MEsKerdQ1ndyqFaxvMwc2y3cxNGnwMLNKCFG572LR0hBx2PwEPl+dL
2tE+zcyhmP9AfwJgGW/erLv6T7Dw/B/wjefTVZ+Tq4f8OdHhhVb9n2gBdcoq1wdBcs+aJmZ8osYA
ljf6iX7rGgJzjpOLyJ/sd0r58xn1aeVvJZLt5krtlgL3wmo7y+ETEVAxethYbbUSWd3FV0yuiFHP
W+1mD4kBE+xCcsTHxiysnVNLtUdegy0nlEryuj48OEC0bGFoCxWn1eT0rT2ePS5AVMr5wpjYtUTj
P12ZjTUpiqysjTsAUIudacrxcxGQ6Kqh+ArQBSUF+IkdQbI7n97RA/77DfB5vzwt0N4dsh1KdujN
MSiUQLC0Uzq20t55boFJFtOlnO3xCajKzLes12FiE9ioRduDwef0QxxmqqsLAEgWTMGlqmYpmlkx
JRM8ap7/QtJvJzVgyfPuQzBeMIqpWsM1Ylu7rXejYJvXoauMnKMU4+0f5yynx6Bws48xQzi5TOer
YhTQ5TsrL20ygqgEH6qKGv1gNf98xWvT1sCa+LD46kE13rBnto39DSdFTknCnpxK9+h4IKfLKsPw
qsUCxh0xsutIeOBYcMQCjVuUuEh0j0ELFvvSquwsAbVNArEfKRCBxb/Ghk7KBwaRUQ+zDe7Vf5nK
bVJVrNFJMOmwvHc7sEAancSsHhtPCYlawPKCsmApY+KA8Xf7+RQ/QdUU/CkzvVsjWV435xtQjj3X
c4bKvWQY8UG5EOnzgv1YEe81XfsX6vHBqW6jXJvRmKWWSDu6Tfx0Z6gU1ugk360yA+5q50BDOGqv
ZQjotjNNgTSKlRM46BLypjzv1jXtq5CLaSBsNVZq1a8G1Wmi2sPiz4AIwR8L6H92fKCkvkbVGk2Z
5E7ILN6GFjzpA7wRYmOvT0MZgpZTJGMzkZ9NyDR/As9uaf/LV6jMJTAOlHvazKFTVWXrkKb/mHCq
i6YUCsGfPCEtQfYTp8yIDMbFwAOhLLK1hKGiTKnkuWPu5fsCsqNdBWpIsiaqbwWblV3qotdKmgVt
i/83p+d9EQTmPjxptfkCGpb8UwVQii/LFgLtqT2x70H0nSAc/E5aTMNrW1BittHwNCX5Wf75SKwT
mC11V7ySrYuEkudBbhLdnZO4TbvI+Ci/U/MtqwLz/dCH12T9LfMfN4AYL0LX228T1jzqVn9YMnIO
C2wmt2PgKoTCuWy5uiXobmVmhpLdU/LdVIC71z1oEHZRaXjLs6Q4Ytj0XDYNN/OvB9xvmnJmjMmf
XmeWF7JI2iXjeEaCRQuXd5oD8viG0AoN68y1dBHHyZkY5iMn/uQwTgriLjQtmyr/ccgkoAiSTun8
RQSvRBKQOFJgY1o5yuQTrnYMxDLR1s4nCHQwaA9/Mb4XxEbX8906mvbYBoikDm51pLqbre84hwFA
fz8XWh5ym+9YKWgGQvDdkjuuvrxkkqkzGYeDu6xeMuL5Fx1Tb11C+9Qs9EdlfdgYffpLhUx8mkc2
mVPJQMjiUyf0n58tEUF6+u1p6PdWBxaTGUvt/Yr0ftLdJ4IQ/bFN/jgios+yomWYXXk8k+MXoyXI
8vPUNw6ZoUNjXsci2+RBHJYCei0iv4MtPOQ4b+bTBza43d9rJbFa+0Gxddoo7eOG+7H3SECHb484
ew3HyxxojCkI1dnyLQ+9xXzFk/437bV2kYNg0gxibRSocP90B4tKmX0aZ2Ifmg8KIbMChY+KLUlI
sf/Hlib7cc47Fgln/7Hvkkh5Ceeft2euUStZet6LAkecXl/F20LukpqF5waN2SWOc5GmVypFPwdD
SZTjmtYJX2C+WWgEQSPuZXFy+YNarFBhRoX8/vxhiHF/EIqBUWfdWBX7xGJbyKu7D+8MWc9NHbUb
7zoYAdAPV6bvpdaMjzk2nKQvW22v4itDKvlvHdpXeO+jPqxhyCjlKUOdRWw57EF+9GWymc0LNkIk
mR7J1TmFQJoQs8C4HMduFFsf9/ilGqBchfKvz0/lxgL9VxkFvSz9rwjMOgYQOWvdpOyYuyeci86H
E6dYzV+uZfilPM7uLbGy/WTGdoOjCfW0tNXGDUjc6WNZ7Ilnstj1KHEb5HAZojZUGS/V48bupbTb
NIvOTiemGSW8l0H+itAl/lE9OGESTF76Fx8NKe3uBdg29y3/w7YH9Z7KQuUBZcgTyqDENsQpb1MS
g+6k2WTHrPR9VDBXveAL5VGFu13TVpZAe06n6EmQmOZzNsrKZbv/g0LOOAV/vwO1UswlVIVWk1g1
VrVdlUyL0vSjj1f2vi7AqVa6VP9j/gB5fOBCR2Kdn6wsnvP0z9hxHsAJhBUlWULRcMJKbAu5qxjV
36HXdNWunBAjDVPw18JPwHYzD4zan0XxhKeGc5mg9D02iCtvfBSQgDa7ITFTPUm+ysA1XtO86iTH
iHvJJ2djx/ri8q7gVEt/M91tD3Om2L5SJ4gmjKDHqXgMKTxYLgYoglhWbFV8bj2OPqyZfrNHu2pi
6Ti6veHmqHIRR7gouIoreHAg54fRIktKfpK4hEJouSqN/x9uxKpSQsvChVMaEG1kIZvrc24QucMO
l5e/RXkl4yJV2mRn5LXpJKbeuJcXQJMbGiYNjtyjX+g6BSk/LKcF1ubPQNsf1+TGqUvgBdeaik8z
3w47RlILX36r4wCArrpumVC33XZOFza45FizeN64ONbgE8+uwumyoQ5tehIOxfDNkZ3goHXpXmMF
cHgQ4XGHpQpI/OVeuu0naz+ufchjLjv1QZXGzFz2uMBqDPmogevNy3Hs0mXmptWTaDBI4aJGfLen
6lWfvCGPxu5JjlvwBY1V4RqLEkCQr1yilSYzkE1YvhvGJ1o+GYZgBmoYbckXB5BfjxWIhDNTEod4
yMC8NwgY4uLeoKmxs/DC5AYDIv7srDE1sy0SEQIE/DEPw4SmJ1ohXhKeRMcFQlddsf+V/7hUiJzU
MYqhCnW35A01sgBLCNDws6cVhA6V7araMr1a4YShWOYLChKvbC//bEEN7W/NpPH4ygLABCcuB5QP
UXgYdi/9vQD5P21KOMcQsHHLEHfhEDIz45cmmzdQFEFWewVTBud1uKAG87a/zpAwMuJ1/RY9/viy
0zv0gUUFWexB7sEOsNFbi7e4vl2abK/CZs8XjzDoFwBEm3E1N2W7H+oVDduJIgCbDr0fOUF7TgK/
RZCd1Rf+nQJQW+H1/ChhWmMnYeBI9NtFJ+TnT2Cf/B+hKtMUZT2RpGahOrYoYIsD+EP8OyQXLOgb
GT/jt0jHfDB7fh3vpL9485jOwGA4cY4QQx/EbvuKFAjH8snrN6kaw/np1IkIFBJ1UwBn13UMPA5Y
boK9nTeXJqyYMvDX41XaCNXoGqBS2b/VSQwh8xr0wHPfmTX5mZobK/MaizZsop6MsKzY8B9MnJyX
W0fY0KK8PS2Kb47sHSp1VVcF530Vq1ZLuf+ZRhTOwhxljVRqMNx9J29IfE3JLheGPebDCawRdGAt
VdnBv8ChzXHdqv7eWaYd34GnZtQNg3eT5OXrafhtmbJ9QTw9C0k/GbFidTnYyDz4/kHSFC2h8VDk
6Rv44fmMuolXCUqY4+IY28tcfOeDWWtVyTFP4wtRgUAxWmyaRCk9eszGAxQQCfLffEGnFm4YUo6D
/YHE5104wN2HxBeQTeCcAFFzs46ClZAvyfIl7NNfB3tBFliBDO3IJMiFTLTjmCFeb1MXN9taXUxM
fjConhymbPpOtSaIXlUZhNMbG8DJ6EKF6FTU/4T0rmcWZZS/hyY1eVaOBuDzGkPzEWnqQkBarDs3
L85nxeBxbwGb7GLzEcBdQJVeuiV3N736UldLL5iyyhanrITdveK1LMKF8OKMKnRJwdzXdP8rMbqo
l1NoVoTjQX9uFVFdp8UJtBJ0PbVqKa6R7liZXj5OkriIFREmMLEuUuUEELSx0oVPWwruEbXWmOuR
jtxWOGzNP+5rWRzfLquIMMK1nVhXYTTSMEQyXwx66cUrj7FgKp7aM4+it+/0RtDrlIURlhO3umKU
NYjWYYFe+0DxKa3p3c64hDXpAdmSmPHxovMPuCuC8QilDuyo+q+9uOjEWdQXtVggc9zmk88zL9x0
SzFOoxl6Gi5PlYXzmNsGxo6HzcDA87uOMwXXMIfOLD1iN+FaOm9VihS0KS0JrQsm84UqR52spEK5
chVKh7PTYhwqEOrwL14vdor8HmWqudK9gFweHdEoGcU3DNFUWufy6U7WG8I+Zizm221/w98muIBB
UQNO2jN6/1Du8W8p127KE4gfwQ8qQGaD7dsn2TuejwlZolNWwaEunb9Af/9zrgbB2R/2Uy94bdlS
hIQ/s4ZvTjAXv9i9ddUeDNSfa3QOxbRcZ7NAFV0g8HagCa7JGxDsjCsIE7SEzBdIDF4mIHKTmuqT
nrj3L6TWHB1Ej42cTcwfSMXOJEI8FEaroxV9XwDfg80hKM8w+7HGRdzj6J+HJe6XYWRB7HM2g77T
SuhFvPtF5m2bgp06W07INtYVYwqrPGjjMXpWl8OEfTlkaCBb0MB+DIvMXSqs5dOzvkO5N4kao6ug
Yw5zU5AH7tJzkrNmYXlPn0k6K1rPxMDvQzhP0vZA4cPfdLX9mf2fc6s6neLUdAsppUoSP0NR8m2M
F5JiUnzL8F2giCctFha9lpaBUzMypGEHAvzTFhyQFhy+xugKVsOywFuNaupn5ZA3SC6JSbvRq4Qw
eBMg3xxqbVSNaBbT4ukLNPGKM79TbIK1ev4GcijxFr/QXhSyeA7jruUQiREnhgSCa+ML8fytJ45y
+5hgWHBY7UWMU9PYd6vSxlxcvL4rjE04jtyMDYi/cFI+ARjw5/hQ0S335Xz4xV7e2/zLeGKA07e8
ikQLeEws6rrxEOw65jXKAki++ELlB+AoSNWQCXjZzWUzURnOnOE51WjDXne0fG1LtGqy+55KfWVl
QSxHfUnYcYX5uvP6Kd8Y9NHa3r51lMYEv/C66PrdqyxXehm64y42UVudZdXmCMC9RS4EslVz4uCZ
67fi0yqWmzwoTXA2Rm9QapPLDnvUqI2hyk6pZ8uITM5FKwo1bVH6IcazlOpeC3XaraKP5GJEJb45
ynTqBE8jRwoGGkJE+C/rxA7s6IVftYS55LFJGn2dD5HArVjFlitX2Rg0AyxhV6GolsN3yvVsTA2A
7lbsjP6e8PVu/EgAsUl4HBZhnWVbCGtLA6v+QXenfv/8SpTiTDKkmAr4oS2czAM7bTCBHEtTKvfJ
pYFXM9ovQe6NRQiRhJbkGqMF91nvuN9Ki7Np5aofF1RYPcjvs+bj9Nje61vM1JQQ6S/XHkxU+gm8
R/lv6xY/nwi1z0Heu1UPwZw06fwca/Rhd4R7Alb50RUc7tdsdOXraFMwKWJhtx87TPLnhOvUvaJj
BagGCgEt6Q5BAfVKqTmN7GwDvXQxU2O7DuBnbs/z0zJFM8Q/IJD1+lh0nIfL4EBn7bN1/+60Z1A+
WHwqsGfQcXB/Dx2G8i6ePUJ7y/W7B9OXiok0t7bh1rS4xCvsQt5/UOCgm2+E5GWOqaiObbXd9yfd
m0cvekLtGMIF6EXKSOjdnjrj3GXSkIn9zu9cPxGoaMDI5eJ1GgT+iXhraPgYivwMSf9HjFkpdKk4
MB8yZQaYcr1M/p/sdWYmsT+ubpd6+sE3Eiv1NgCr56YoHpFo3C91PigEDmFMC2MH4TIAK9XcPp2C
GClAcKqLqiqwRt4PE5oGh6AtWlf4AtPAN5GDFyMvmxDobeee1vb0ABLbLTyv4jFJ3slaR5YU9D4F
eJZzM7/zlJkRStbAT101VrGjZak5zFWo+CNZT8FLAMyt8sLJI6FE2xuFvj8onbnJ7jIv8XG5Ng2E
suaoIU1nt/RfyXcOkiIWv67XCcQ8ieqDguQpyaW2Xkb0YTDPER3Jnbm+iY58zZuJENEHFKgXrYoV
W2QTql3bSqjD2+IxhSkRounAb6UcQTcrEw7YqjQvbyvmXIw2PCphEhslUPaL0gzZLB90OGvUd0/a
5IWJfbNyouEo/THpvkOjIrqc/Qv7Rr6Z55s03i2NLJMb49b9eqxdcrdzGOJO5o/+DHuZKxflXCUG
R/D8Q9idcNfoymN+tee44LmgI27+i4yQYLYD7E99yOM7i0+zkrweVQyQFOHpLxoiB/XEa5skdjIs
/NuBT+wSyN2flV99lvksFB+luBSOYeIMVTn3qPgI2abNzabtUF4CNGcOmC/7S8YHXxPUnk5ru6kN
aqGIXiuLMcTVFryiGw/7AGnVv+lGo6GoZ9EDdKg3poSMP1aY3cqfRPrKuL0RvL554mOZFJPi7k9w
efg/ogc2EmH5WEeVDGe+Pbw4ISfhljikvA9HY1ZCW8ok2XoMbZwmFGL9HOxgooqcsPZjAl4npiqx
HLKiszaRAKotx8e4lNLjwXlH2WU71PJcf49zYm2gl37X115PNA2nKJcCV+ZFTUw1ouSUNF/zNL2D
RsWWhUVbWiQV41Bs7bkMjNBMbIclZL9NxyqOFCK77oPxsXO2epo9xCQ/7EEAJQHkIDEz8tShlPUX
rzdbB21JxbwQN9JSYYnYwPhJKSmWcvfSW3h7F6lWr+G2mulBeXBszox5AudnzW9rgFUJWicd7Nn1
fPR3IRmmL+lWQJfWutBO/8mKFZRrvAQ/LI44zEsfix5gzZL4VUFZP8DY+gpnT6TUKDKgCwFgcxzu
jawXNwD9dQviH01JcR9EbrFvXVWy9SJnJrmG1y0O7eGCptT75QF9iHkgVI3L8d/ZJFXbN+n1C7Lu
+tq89LdPVUaPqA0BD8Znv0uH7YvJm+HTS30vHHTTXDM0ZubVn0KKeWXPuabUYjQv4sd/QGeCvuyi
iwmMETcvF7fcQi3p0tWEjunvHbABXd6jThVegMju1se6PmHt6aEiFleDWzLP7MB8dqVxzaGUhaF1
dS+sgdpXIxy0IossG7a6Cda7mc4cM+tcSEtJhQcViaP541hDzOUSPOABIZmZumVUXg1HZmgStccA
Z/AIRZ+XEBQHavu6ziWnVEv112Sd8vSowohwcbgSzm2VZjJmjMLfPjXvE0iYLEKf42HMNgpxpak/
pY2psENUILVh9APyQHs0TMrvrbs7BugkAj8Y+K2bkmZ3ajQ/L3XEUhAtnTPMdsO/rVFRQpvjHKOH
ZHURC/0TJ8Xddq9DoZmYHLgG0ku6t1vsGrQ5IvwzFNrkY5HtDpnEMWDXPFY02Lqkty9I9DeGR6Ii
mvYBxvivuplwPViUZcHjv5mTePtSvHbm2eso0DUVhmw1ioAUU6irSdGl1eR1BLlXmzEIuahgW1mF
qQdnFkCwP3JT5ej7PUbRuUB15py2gMQ8N/DiSDBWuez5ImSBu4dEQEp1ci3Jms3Mjl5vjjua3Fwd
EMhXs4xEsbBMexde8eLCkZ09aO2rotyx/ufetHos699eaXsJprHCbbTbIxNCOwgdw3G96+rYhGtR
C/wSemI5oTJ1fevxn8kz//qjHkDomtxjfi4zpDru272fPvwULOB058+HvGhiX7baoSPVx5V4GjJo
MDvyysmn0iLfl6fq5k+Q5opzsHmSaAImfPTm4qZfX+8NzPgI9QS6GW+w0SunbfTLhbdW5mMz4vRl
YMi/09e6oLz2iHqsRoXpo1n9Qt2b0JGyaDfEh6/Rk/uF3mPB+29/WmysNhL9EwJUXEgAv3jY60Hl
sqnwUpzK2XM+syiUgqww/ufFlmvhEVr1vASLbuEAiv+0/A/tB7LfLFw20JfD4HpI7+zmOmLrAinK
dL6rdNnK4xJxckFVM65GnTib18MhlmFwPgLpfLoviZ63ezMreg06kr6Yn6BcnSi5UEMq19u3+/Dk
wvOoE7UDUqn9YNa7ZKueGAE6Bc2KXCc7ygizBDNmetuzVkUMCT4a6B7BFUAJ+HaJSE3ZjbkJS29I
DuwpyWb+rHACeofU5YJ1pVZ5AUu5whLn3kVI6JSdpZNsiOBmEMpjz38IH4NGlZ6d9C21UDoN+eXq
QK720IjYox+d5/EZ0w+fKs+EwY8ZVry93aMZCVNl6XonjYQ7+RdP7aN9VsgdBqGllDosQsAHz8GF
wfjUyIkmDeemFG2JIjzRwZ+VMpPewSAO8BW6CwqkATjUWnNK3T7s1XtFlepDLRjx6nKyQI1GWRe/
ZVz3t3rbH5qvtEplC7rwhqOuOMpQe08JViaMNnp1a2r2XGQ26b9sSmfkDt5uU6kMs9q1YPrknxgY
CuwQIS5zrE+AyNB279GH6YtSoBewyu8PyXnd1GTLlnRbdQTnyWZ+1qt+5MPbRgf1FbhCv/s2oltB
fCIXTNZq0Yoe+XaqoO27K1ZWuqZhxpNt5/TV6agmgK9vcBJiibiENFSWIHvgjdlrteCEriarljGp
iPxpFnE3dgN6yl5QNM45Jr1513Ao8Ne/g0l+G4fLyoFKP8BYO6lpCw/PU3FguvDsfRPME+k3L5m6
r7ElgxfoXDR3FULt9R3QZXgfRi9+bMsasLaKiFFlSJR9tXAm51LfNTLA3tdprj7n6KeIeZwqoB+N
HfC+PLhg7ezP/6ECe4k5NtWNpbQHSRn+zlr7F3pUIlS88ShbNpjDAiJ3AGTgtfmjtak1RY8g8g8S
P8GeGBf5beSpsrEVLvEzMLBYh4g+ec01VXt8yc08383tXypx4Sfy6hHsKnV2CNPSb1pWe7iClSV7
Excq5d1xDj7vJElH6+GNRbDm2KYWet7j/HkRt3ZGMvHORX0tR9GmFJyO7ix3pJDsAeqfON9N4pX9
FzLgm/GVdFKMkyCTOACFn0pgUe11mpxThkEgfBQDX4YG94paxbu+pXlYmH7VprRlPNv+V87eeciV
K6l838zozVQDT4rfGPhq04DXEw/OGRJn/Y5aeMjVIZ06mywFUWILxJLfRijN5vyE7s4aCk2fynOZ
/i3fleO2CrocKn650ZU5O3JAQYeCgTb1wh89/EqPENelHLYhzDqNa08UgLCj83VJXlmYEdhls5nl
N9RXTWFcErdiMAKmA53xWXxnfG5CigedmhkG0HKh1S8IzmYEEFZ0yz4ynF2mnXgLmFzbw0rD++vj
IC14h5pKJyo9Rsx+mu9KXp8HDcMSdYbKjb4FFF00wV1f3Aq4YVtZSFXXvrKo54med5cAK626Dcz0
GRC209VEiKSvkQjWxqmpsi5kGlkVczRq57WZ7Q2W3yc7ErOF3lYqw+dS+L0TvXCG/p5+ixAGAs1G
gFyTHAqmKjVRYi2SVSVNs7FEHBADqiyvfUG2SHJSETTGlWdHkduVs91m1S4Miacto/v49ieZv0BJ
Hp95kTZ2EuAd2pOpHprty8Y2uDM3dAuirdCDJCHd7NtUehcL+GfWK59ttKCzBO3mAm4vE0aYcryN
q5hWtK2pQX0DkFqmbe9fJMDNSVK5X5iwlRmNFNlU/Aohcw+juedJ0PPDLSEJUuNbmOBJ0dYjfxvV
8UFO2S5DCRRxHDHS6n61oJQHgJ4PHiYWCye0ghpH/TgEW5l8J7BBHYcSzwowjmEUeEhIPhIpCPMZ
ZwX9BtWaT15aTxQbbCKqcnmZbAlprha4Q6wCLeqRYgVI5MyzOwORXXnjEj5d0du4Id5iSvtgmm0E
XdyCXOdg28ICGGhxhz30oBjU9l7UnJpEdUgQxf5huvM7joinpueHZTISIFxTSu8wQ9L/CBESFJ29
rvm58YkjR3J7zNjQeRUHStOA3loeSV3ZDi5gy+u7f00pKCQUEbMwtsXJaBaixIRKmVaad6+lcaHp
at0/zmAhVfzTUNbtYlCGqz02xZK5sLMZjtcVcMTwBo7/jF6sqT3KoUPEFxNv9te9nR4n/I7TJ8zr
cbYSFXzGTKVrs3bfdJuojGOJWwJL7fjiOGYPOdK55VQ6+Z/yRNWDHyLfuZrEthM6sr8VaWzCtsSZ
tKK76HSQpRrLhToqLTkm9jwS/gPFRFHzW62oYYfVBJLYYA7v51TWCDdjWvGtUbZOw9IXocFGNUci
B93Vw74JOhw6/G86ZK0j4mC1pGkPTvkUcreeLQUxU/EgPeJVoOiN1yr0frye1LOU9nE2jooXcmP7
hW/Ba+0DGlYi6u6jm6SkozdryrupgCDKGCTEbb4BPCzmxK/oFtijVY4fNnYTwlW7WhasbIhe7cyh
CvoW8OGspf83lXITDPdgXilmTebHZ/oImOCmUK+iHWLeFcEMQzy5QEbf+oAqGgGIa7QrE69QolO4
7IMbH6sENpvcJuZc0PWzoKt0BqYCI0y9gvYwIIhsycULJEJ8nXSQr7O26AhsBSaqphzLXJd61zZ+
+M3CvB4Z92mV+vRAyud9YNbuiJCFkSPg16G3JQXPqVkW/NrCO7a0KRq3C91lMKKbHiJlzirRtZhJ
OIjSZtoqkslXAXw9qa4gJMTDyxICIdT9nlu3uVnCS+zWaaUzAnTO8dEq5tDvoAWfbhgy07iBvD2F
mGV56uiCIegqwsWRdKMW2XlcEAxxS2kqeJGURxCtJ2O//L5mLwEI/r2VeJ/mW85HtPZXjLam131i
Ej60133v4xy5OhXJkm1FBOaNhTSSjhqMiBh1bVHN8rTKWMfz1r4nfJ69sJXO+cI0+9jNFe3tN0PE
DafwSopFhK5L+IaHbUUkMHkBG16WP2gCltWS65dXAANDXTx53FyDT0hJ31mvc+8hTkbzZGO1DKC4
Msgws6BQ5Oz8YuJP59PsGypU+KO3Rj1ieZEWNWKr+ViXYhJIA/Shdrb7b21hHFnive6nimLB1F9r
qcHnez8sTFFqfl8vt8t7KbuzTWCytRZ9WpZlSvBuXdSM+izTAFyVRN5DS7wl52MN13nK9rEeysM4
g5+lebl/WeWa21MIFGyN4+DkmxIOkTZK9yBhFXpLU3xPwrwU+nfbVVvmFEnmbJDlBVkgOny6OJ/L
kD9fIiFTa3nrTAquZvvaYJCJ3gOXFFyRaSCcJ32ySjC6UXSzdF/G3NtnEUlUDwIUHiAfvvIClXYx
tjWyJA5WbuZH6XkkMaULHjwQ79JS6GKbVmCy274MXhvJgj++N7FXGeEJez/zNWiBQ0UCQzJFbkal
WpO/+CpwFqSsZ9f5AZ9lt1u7HvUV80P1L6FUKrM+fiL9b3M2c5mj2q5QGalyYADFlZ6l0u+Ka2Cn
9nDohCYLADlwRZQyg5xmJsKEy1DAChTPCU0OW/H4pbWl7SOLMiYmpA/oyQ3EElOZGn41wcd0bLO9
rqmFc3IlSxdlgdQ776CqGAFZm+pCw45sdvMCMQsYn71BROnmUSLfi2lU9cKH7OFINpTdE+7UjMvb
wh/shCXqV6GHj4szIL0RqVQkCL7TWOGIHduQst+ELANoNZ6xbHU4TUXOWLCi3Fn5WJ8efAug/0/X
P0v4ptmgU387IE32Ms9p1ZKVCw3WNPeU9rxLNFgoDPRk1wvgwsTJhFIby1e0CrkQS34vzMW4Ytlf
tO0vnKnhVjjD8mHE8OMAh91M8ErhgZLkz8Y9drAa4iR+Y7LTvQaPbmpUPsYXWOSn9/RQiSnYcfao
I0S5nstMqBRF16Qlqnc/k/IR1KpbAsBtREueQXSyrzm+SrZ15iFq59YgoSaUGD8KUpiCZClse5Ci
Yq0GW7O2br9XkOwE03M9tFMH2Itwt+1zIWxPMFjMEQ7SmKOSRDu9CZwmVeW3DqvuTtjgTy9DDmfN
gMrZDLQcPizlIKRBQju8pa2iaX53W++vCd0WYoWrK8HHaebuIbqWv2gfgWQD5mQfIbcnpOGjehYu
sDPz4xejB9X7ZTjkFSmM60iWap3K0b54E4m6+ocmlNXzGeko4v0TeJ2i5ZwaxXgR14IVPH1019/Z
h/CFFCq+MXrmWjc1mcoVeZpkxUFyeJCc9EJEiam6JwGQmbUGuFPVQujVpVAn+iW4AqYDulqEWoT1
1s1U+xKJo2xKo56bnEU04QUdiq3cHmjzbTCmnGOSxu+qmiLbSvGf0lWiJaIyvwdFCoyrCGZZRGol
PZu67A0dD04OfQUMvZJlF2/7igM8fAPgu2pA1UZ6rKXz601JMoxbWVTN+V8UV9rlTd0ba0E/2cho
kDY/Gwml8DkKZ/Vc5IGA0YCkeRc13aBmz9BKeC3hAOfmfMO1mN49aizbz+tz9oiK0MPgKRoM+HKD
T5latqORclKZEVXM0zWCh25jq4qJPD+JRSw3dPNOLLhc/COZ1Uh+bAEeIiT/M1DMLzexu0btXs4t
QamO5KWU9H7uQ+Hx419UgzvF7eheXJNpy48VXcdlNWEqOnh/9TW63NWFm+974QCUMQocVbz3CXRQ
IJcwcg/U9ZfC5h+SfFVQy+vEGorL2JvrlwnKDVt558xNo0zKp1lPNSKtt8vOLro2ZqwNPMZXz/7d
Vls/rmChnH36INqWcTGGO7mjtQYmOizLEZ1+udvZm2nAMtQoL5Xsfxk2Q/wIJ1GsBS7K7gv6legc
PnKaO18unHCq70R8cDJ26QlqNNbbtq8/FXjiSpedpWLML9t/2z6GLz/kayHhN15L1xfcLs5oso8M
LiK31v2fYDtB1+fHNl2jTzwtnrKX/9OXbTIAnjPUVoL00CRGYpumHMjoxWOCZ7+WzG6LWI6RGPAP
gXudWFyhT3vEMYlR2UoZuwLs2kKBGYO6eBwwVr4HNnyjkAyyUZAntkponr8KG9IViqE9imHg7s5z
vN7o5VYLXJCJnwUz3IBM8TJhvlQruWFI0ZIOcB8jJLmvYpqjoQMFH1hzUZ3KhiGw6Sug+BTBaVRd
38Dy2W2+KZwqmhcUvC5ioVSJREbBzNfFYlFYKskS2ZyzuKOljPdhHQO8Lo8OdoCoJt8EVL2zx+Yg
Fxo4UGyiRkHdWms/AKq45jDTuROS54fWrcg3uUfDv0T0cRqhBAhutK4n5AqD9dG9MKL2Va9YNToE
0Gm/6FPNeezDteEPfkl2dT+hjfqfgr9AaabrQp0V5YpnsiuGKoIygmEWU/Ia9/lMg2WZCgFKAjEe
yGh4wHC+F7j2R8ldGEXENRjiaG6n7dL7++yTGSJpF3wi6MkYJVxvVU19cecH/H7nlAaSCMHvZtGt
vdtPG7wklGvufvwLQVY9D9iZwW/mYBBloswzMbDpPtncrcEeQtx3D5Bl/xSnnWgo1XwocgxdtH0W
p45UAgkjk26vQgVJghvxAISIutttKc/hu+3wDHM5JYVz7fKKm3u6Lee41nPW7tiyEE5OitPKmjuH
tiRqBicpPQmjrxn/e2OKaZTE6O+eIfHK+4GjCXIJyg0JX7EI6Izb05qmKbJTS2uCHWAFR0UBHLxw
cYWCb0vVUD9X2rFumVD0VUmONeiJB0x8KqLHqvra1Lu02OsulycKJBCSAXapU7UEbsnRaoYgnLgY
bMDDcpa8Wy6uC+r0GKpJEBuMUDpfuAHs4ZWMT+iU1iI+JI0oydzOtce2e5G7c3Y1tg7DhuVLLKTu
ZMOwF1fzu0cDvaFGpiXawpO9VQR0uM/Gk9eSlXs++tju+oeSiwOh9gy9cy3lEoBapUfg+MrvW2IS
bX4Hv/M/ShqvRnwlJMGI39enrXlOyRndmJYGmz3cDgh1lLPooEkrnxKwBNDYvpzkgM/fv7M39rfP
xTDbTHOBg1S5cfkSbn3gARbxuAs2rkf7SAHP+RP5JNnPvhwt2yEJGBjW0FHxxDfQ9M0CDHWe8BJF
0e6av0teJhn3HJy7mdRUI1pabgwRtiBuvx2Kyba5wPLenBvO6fnLuC3bq7hzPLF4Nc5hyyCKc3FA
VP+PrbvvEKFOR5cNQ/ySRGNj82n9aVM39FX4T1kEe+8sJpm1K3PHahGMvIl1BvSd4L6QZ5Uu54cb
a/pCu+i+Ean0XcSK0/GPlITxhbbxwqEEWBYO75wiN+jXLEVlxCEDG97VcIebur/ipxN2nFXo+2Wt
dsAAFsiBpQm9dlV/1HIiHBgeqa3D3lteKbGOmQluuL3MvzPqhTamkTooxBRyewTVAhDOOHucPoeo
Y4fSHNv1Q9leFrKBuHWcwkRTewqx/SMzFNdSzq5t52aIPCs65YpTbOMQ2D3O/MvebdtsazSwjqCb
bEh8LmCFL2bwc51TGysSuou0UVzMFgZ+7Fo5XDZd3T6iD79FfNIrd0oePNiwrFjxEU5Y+0/1duGY
UFy40PAW8n1KqY7ls0bJ85+FLTNtX6jGvAZFjOrZXbQqYLZ+PCVW4K1XM8EF2Ll6SwoYZSaolcg/
2i7pLTWBOmbDCtxZUdAqzZHTBcn5cx4v29B3xL8p2g7KS/dxFJvF3aQ1fDH1gMUMAr70k14gTlUq
kN0+OTXEk1frgRPQfJHa3n+malmkF1tZIlOgho4itbRCUK/8BUu6lLBDuGI1Zp36BA73oz1nJ486
4mRN03mBYIj3FPD37C4a9x3Mor/QKrkvc6qQ7JZcjO9Moyxadv4cC0FrbnOsF0iKLhcVC76HgWww
OEBvZSE4VxnvJWnDGMVpjK7KkOEkRjVvXMsAgsTiaDS3rJDOTJPbpIo6gPBsZMKTBAhZky7f+6Ec
Iwunp6B8hTeQne+/EzU=
`protect end_protected

