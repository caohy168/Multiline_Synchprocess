

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SA5jjWkzeQomKPkCUNwPg5yR3xJF8sqCignVlCLm8CmaD6yCN+xgQnPz4cq10LpPVs+W5rmALvn0
vfEm/TySOw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jykHSjxjcJNykJVGhTxpdGlTrJwq4v3m4iZoyM5N4Fz039NFmJa/RKjhCRGLrnduUl5kmttA/Md/
PsuXf6/oAIKTmj+yR4+zjJ+UyIj2azCTxliCNkAZPfoP0OcJsBJwnYObLQD/pBx3Q0vl4pcVPAn2
XEz4egBdOXTnhm51bNs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ew0nQiLu4cw6hZkI/KX1nztr3s4cYyGFa34WSNqp8jgp9vwTLk2GBCZgEuyd16k2AfRRUF+2yLZo
APCYN3WVdwjEhq4VUz41h2saxnTVfigItM/zHMXaS283Sr0dmnydXUkPywQKOsqTC2pWGaca7gYO
NAV1HFhDqXzXYkBKYdQaQdxb3l/YAvXfPC+25VNOiexD/qezhyEtfkLm53X1sb8wHrXg/Hbnw85C
fnKVgEuZHLhw1BET2eyt9zzCpgLBUKVDQhUWdGXJfnQu5mCLAaQTHhdcaRCsFTiv1QENd8R8HWrD
qv6W/1E5H8ZQWtPtKQJnrHQmXdOJ+1TLJDg8eg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZFyEMQv9Nyj/D4Dp03zsfHcDeI/29E3JhK2MEp3hX1f60TinPfwRCuu1/vcrfcvEsea/eTDYMHCB
JmM94XAaNeJBN3AKdGT0puv4duFDxL9QOKgOjOYtSoPQvPNmL3Bg3efZAKLAvegbv5GCkjrGubYG
DhiqFFp8wRFzfGjk6H8gkuCVY3PsbJHgz2YhMLLMkp/r358IGVNuJ6jwUUJ4s2vLayUVGY2mIXU4
5qcy1pQ6JnT/qjxzqk6DpImmZr5/BB9gWWv49QuEnw+KuLCRchKsUAf+0hD4z7EfWPb2sWH/ghK1
lG2CrSttZM415vlh6j6q3XuocsZwNKQ0mu+z/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cB4UIgT2EOn0FB2NBI9VdJ+LzwNi8NmSjjL/kAceRE+VMTCBlYmd/+yQG6HuXdemQQKxKowqGuzq
BuV/FnMgQS2i+w/GQIKuINv20mjZVUwmlbp9O4wodbiNkBYSrz38i0Rj4ngZ3ARuguRewVA6m+dj
ej60sai4MI6lXLM8tYQ=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ql+EJLba6J3MSAHQ1wsJEGOL/eGh2gs9r2AASCE9alyXLRFVX99I3MR9PG2xlO+RXfHL/tgA7x1h
SmElqWDYEQ3V2xF1KiPEigvPfbls30D2uSXpJB1xlfVLNs/Phaz0mV4QUOrkfs2MePkaQbXQecak
yESTEWxegVAWDLSp4LAE77b2ddmeVCkzkk5AXf9zV0rL2JffumqzoF1CMbiluk47JxWczvg+0Es8
Ny0t89p4K2sAzASvu9iQPQaqGPplQ40LyzJhH5s6iISUK7QKCavdoPmwwGveF6WtahVY4WZiwXQ3
zSpPPWJIZpTn9UIYhd0G3RVVhduoDun3x1WBtg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cuqg6QfI5+mv5ahfGWpSepeuu6G1FGgaauc+hw1VIVvo4/yMdeMAQuzeK8jWoyzX9pdcibi+YzxP
Sqzr4X4KK019BLChmlrC1vJxAXKfzwoA7932l3uHfHeBBxDwhhtB1v0iZyULK0YKtH/kxgYVqz65
/DbifX3kT8GkQFPu5iYPXMhmT8Yg1nm9bAWSn44FsV8bxVLl8sAWL0qnwbmOKz9knkS2Byumzv/u
VENgkn0sj+/VuYmBAO7nxFpPbwmRQ3aOws2SUBBtcPW6m7Vi09ObnKgGbYe4agg7tSmSRkJvQ8h/
p6CbKKGsc1+8gp5viR9QaZVTuLbTX7L/OGeCzQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rb9Xrfzx1owXAfsqT6IWzypBN0cE5ufrV7ANaJ3LbT8ZLBLfcvp/Ibdc3IC6nae78pe6f4C67aNv
iS91WiwjunvCDdykSzyIIzpUu7MTys/WoyZ8tAlG/oGRgX5yo0dqTktYwo3fn1VsA5TMnWvUocT+
JfxEvx2crENoLnTguBLUVDyguMKVqdbNQIPJ/303JcOXOU9NC/Zp51VV/RQJuodh8RbXzpQiuocv
KEH43Uk0211XyyssOcQ/1qmXoCs8yuMrqunDR+II6qna7AjBgtWLbgSGVah038Y9oXi297VMF3iw
WAflTitB6wtd6X44nr5c8dhxiX3KXQnWM7Zrwg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ThzzPiLDNYIdxX+i6+puL26OlQDk0zjO4lvreJ3nf0uJlkSGIFn61SHBzRudo6KETOHAaXYD9JA7
0hGjseIy0T4JCo+xHtb1ebn0ZVe5aQfwKbIz5KHeCNU9ssYuL5gsk14+XvWt4iU9x5rbgAnwdxvJ
sVodnkvsP5KaI+UrTFyiBr4jn2zayFtdl+KyIqWBHih2ajuP2NaAcB8rle+rCLPE77P8GgYS3mOM
bnlkti1pAMRmAN4PGd+OS8CFq/7apPzhBHrztPevWlsnJlwL0SQW7S0V+YMAdILyz8vY1P4ksKis
ZZmK9A1loehu4zr3IQJ9KMa7AOXsg053pq8hag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135744)
`protect data_block
akzdfD5XIO2Ql4Gkd1Vdk63gy/E5fMYWl3D6DSIynjkedDOaOu4o2QW6KgZDjgkGW5yRkLoOVqkJ
/IcmirQ9v9p6Yz4D7nEZ0lkUVCTxJBWHiqHg1EgeQzUxqG0AXRLmOw2masRb/W9L/Y43HH90PdZG
iUjPOisgSMKDf9FEmdUMgNd2lxBtVjqG9lwqpHYw0+tSMe9vkxVBHEF4kHR1FnakhOQjfphAihkh
vdMERmuXHKjDBpWp98kYJa4R5Doh7BH7sVHK+oI34rHshxtwFhcNRSOjOJ5RluUluoMfbHk820xK
Vp3OpvE03ww7chTwcq3CuenmLq1c4flcqNept6896DuMpve+y8/YZDbBL0xoTDnh6limiQ33tBre
vfWsbI6Ss+mOa8UUy0ilRD+ER4Ve/DIUzTSw41b2iL/N2IbqVK2UZHh+SWxgmdPdcJekoEVyvX7V
AwRixi3ZPcj32JTSYVgV4tTs2eQqQp7XAmipGOVu3fzDk/C7/J8RtObJUkiapeK2RXkVF1EVGmcP
YzSmD01lbwRtGqncKrYWqnD8939kKU7PBln3JI0eCZZR1rVCAfWZD3LwMNRtzBeosQvtONLe8bOZ
sAeH/DBFvhik3AUXY2gm+ViRMQ3s/f+K5wpHymorA5P7Y/Zddd2uUeEvaP7lk0Am8hPanVnIF4B9
x08bYWKmfMJOhJOi3pJWvHXl0alTOqb/eK/iZNPvEP/x/5tQ8wokgfs7hRGHbphTi71T8rKZhCBq
/y/MefHW1wfD54FfBWunZCEKbcjR/rVuY36sHEC5t4IBhvdMnqkKASIc97q3ur0RAmlEOfpCV7EW
fibhovUxwIC2o9TfZG9HO0uEF2jdC+mukmoAiGQjN9MeBIXrkvSaodIVLxutq2J0otuhI1TOj4Pi
tM8JESCiBN4J6IgeNag+tUwIeg1yXiwOz+g5TOhsUH3Cu8Mict10YQPBGd0jqlvJ2MfjB4YJW1kW
TkK/owt8T4+srLnlCiJtJY/1x5T3Q8vBB62LaaO0tznGW6wn0+RjahbfiWhwm3r2DRZVX2jY7lL+
vHTqIK4I+PJ62bTukBs7hjEpcyG3NsSna4kTRdPbTBDg28ErFI+WXu8CAz2jeU2tia7hesXOUjAm
qayQe7H/ITZk3jkqLtUuaJpp2nmar+GConhWq88mqC1irvas9PyPVJAy5tumypRrUtEurJt5HYmR
Y3SjR5bF5acsh2QgF9ZYBvED13G5mkvQDFf4jhtSk9UE61G852/xIvBUBX8UsnmXWYW+SfIyt/fA
K4bR0jO0aQnuhSsE7vNG7AyFVUrwMPu2bi6T1zLd6E/phXfV4ysC3BbLn1SHyXL3N4seV+YGg0RN
YZAcJIpfCoGNIYvfOOPBUUXaBLcBy6ZrigBABaB56auyb5wI8MdBz92a4QZEUPwiMyuxQSqErY2H
FQwm39ehXe/1kdVm2LbmUzd6BM4RpkVjbEjHjmP1+3M6xgzR7v2H7z7xHSp7DUlQeGAtvC8Utbbz
NcciYSGnamEQhbbq2Cr6OkqHL7MuBePkLJJssT1vGCJz0ubuHiaPKJW7+98w8dffR/ajpDk0vmyv
WW5awe48C+IKik1DOfNaBK8teti8HvNZlLg51eQEOwLWIkN48FrRZuEkHM2F+06QoEq5OP7UtdyT
CpliMMESSQfvKrXxjWDypXkbPMbe7uvRh1lY3tnqfzqgTLAv+OItkHBV9Bv06d1jH+rmLA35Iiy6
v8xiNOHYDmEuJEHN4tNRtCcfaX48tjWHHDAuc4wYm5Hw1OGww/+geaC/+WL+5BItMcs2kVebk5JC
F/fHIiJkoL/5Ytn0aR+zAqvOA41exi+lhubxjYVNLORmspry3gqfi76VkaH6DBnJsV7zU0JSU6bz
1ERxFaAM5znlyiJ8CIDBZoRTrGGWd7Bw+NGX1gsha+AUPjFX0kyTU+qXZGYBXJDAsiIiZL57Kjlg
zVNlAUT6d9pTtbs4CyRUNmT4RDH9iIgW9/cMRo5JRtZtcDOX5uou1Y8WCjCk01/akwR22d1PG65Y
3la7Bm+BAo0i8CWawNKxVTkcmMK9qrPZLl61j13z6i/UoC/CWdIIknOp6n864ZppATyZg++52ElY
Z3hFrBDotV3KqyvEHjiX/pLgrExvachTbEe+TnmZpThJ4cPWAXz1H3VeSz/Wv/14oLdhlP0EHT5g
XwdC9luXlA0dZPJqell/o87kBDQKRQbviRI2G3X1k9AdWpwyQ0FNc/TgBYDvadNGSgR22AINN3f9
7ypFpWvGoDDQFcj8Co9JnagxYMAGOvI+X6RzGeAVLN3/xWjv7rKd4yr6fPQWB/vSxOQjR+IcGuji
wGgGDAtAkl/wXKlS7A54IDyQoWzfPlam2svNnRJgyiZEV5AGsbLBNU4fC5HLOcB6K+VQ5lUN0Edl
TawGEINMxp67cdd/q9KP7YRPh+Y05AJyYlX/twmfDI4B4E8mehXIpBOxaxK3mWMYGoFC2M+FK09p
+zOBxRTosDmDAo9YWKTn8+/iKzgYodPXhjgve/kOdrl9kggFOiJxMLr7Ndd5uo6sjKc6GgMvkTRe
3j2zcJRmVACIxJEOlJhrkC+GRp/ZNSCEtX+oM3Tht3eO96yujzo/UjSqoaHkomax7FVexWMKmnSv
oxrTQ0lc8d6Esx51g/U6gKWytm58+r3bXLKGtS4zvBD2o5PdPTjUbTo7dfdB7mTOWDsgBiahydJm
RnikHtpX+Z0wVVmMpXpGXwpc3LfoZ2k1Xe2TjAs8mPGcXVyo8WcPjJgHdzXtsb/BxfnAeemzSV/3
FEoBW5wv1q9pG4UNFzteRnZQYa0pHIkvTaDLY7GEEJWPRrxHE/L5kIAEC29HmcvaY2wQ1NAql3C3
qLc2qULLlMxIxroOqRb8FXHZRfZA9NGWpXbDNiNEOlwnRhIeqYOY9Eifo5YlNLvnmjpjFok3Uc6u
F2v0jSUsdCY1smmP8H24CExufO8uvMciuh9BKsBjbC6Ly+gV8OO4GJzkSDCwgHQSBL0a7JmwsiP+
ToQAXz7NBNfIUHF13Ej4sjBan5JPjdrIW8Kp6IamSrjFfUw9QwsGp8vqOIcmFhMYW7R6qKJtmGZu
60aCpb46+YzzjwH8/f/OizcZcMLQpByapHiATBbFaFfD+gOdtRT4vC4J/nxRQx8trGqgunTjW4XK
05q72OPx5xixxDWYDCmgFvIE4d9LYzkoZ/TW4OcnG6xHA2/vJofRLmSa8DqMHzzaBrqSjuDi32qo
joKQwtPs1RgTf4lgmklTtFkBoKkvJfx9BaGYK61+8Rt/9mNNpwyF+0H/O/biORa07ChyDU/oYU8K
0exGM+R1xMVKZ4Cvj7xfkp8fnuclNnoczpH7N+Maj4jBbGql6Ymxtqe9pwth9tEEJIWSF3fBVbK+
SuemyR0grSTVRcGnroKuP/kx0yRGv9m15q3Ldy12N+iN1lC0Z5oVrB2edoXzSf0STS6IYfaXF1Um
FlQJOilPo9koqTDyhEgXYVqiZUQCEgxg6KC/H87qps3yZdCxYm1X/g7/Qu0lV60sha16Eh4c5pRy
YnfceqbxveN7WRjbMGsXPY+HZf9B3CZwzglBk4aXI/mIPgSPWFaKm0roSHhMe6dW5d2lEibZmCfU
iKKwnSevFDp+vKgWb1+F6Uh7H7OCoi8cFIbS6RKOPK4M2hTZHycJvj+gFf5F3aiNe8xZqKYZUi2I
nvlsJi2mmIk5/3T1ovDX5g3dI07l4YGnqnBzVntKLDoRtLnRlDCjZpajh3/F+5nvRR9u4ugK2JSC
1N2D7j72vN8q2MdlBvcokNl5B1mc9+H1aIhlGcC1GBhG2/Cg9HwyEFaR/pCxbUOdAsc2WPhU/gFV
ZimHugqJDG3wpIDrCIkyekYX/p1HGrzf8Qs00U97l1136+rYRNZwCGm+lXpxEXgbCR4hDa3596f2
4rq8R8G3cOK0MlkGLqSx1z0QROgND0cmlNTZ6rr3lh/IKA/7woe2xTAqGTuyxvyvo5+MBhM1FC37
KVJ92O2YC34m0IIqRwhckZdRv3jW0YTWpw06PNMzy/0EfdxxwmMnsBFTXACL9fwZYuu8Eo5aPs/K
iPKj0a9iQXj8keKjB1YoKzSPQA+G/in73MDDnf/e9AYn0tqNabNJtHlSCa7tYjMbyyZjiIlBi+XA
uBCfeEEY1Xr/OVQNOcxqHsYFuf5V6chCxoU4NWvOYR0NkRNyjeMo6u5Li5xtOPIOC3THbiID82BI
JlyPohLPs2uD4nwH3JF3Db5uQiz3tNsRjz8o6gB4JHzybc3vTC3QAynC8pGLgB6vFnjblOCELYZA
vcVdsDX6hT8p0+dNvAfC8I9mEV4uYZpZXTY97Y2vzmDSxrIA/ySOVmKGBR22fDOcDgu/RYp+kXFN
5JCHFOo+R1Y8WVXV0aosK4Vadxn5PdL8RRxkavIqSgAs6fOISNWDvbhVcmy3qOnJN4+R4Y4ktQPO
abfovYPHWoAlZKFbfF/oPes2+Z2V0I9HaUCUj3Mv29aRx5BYBMk2Ok3f39am2d45zGjZg2kow5b0
/Cii3+3zUHSbQ/oT67t6T6H92eM1prUjgdhBICCpt0c9dBple/H/peTmCylOv1V9weR94dZBptt3
zbAbMNByQdLXtarg6+w8Vt6X3DDeNK9fNYR+dxGhcyDYPjwkxUOmb5ySlCNXIXJjg1LbV2JTDGAe
xGcPRFWFbtxvynT58P/XvetUQ0VuVKPNBSaHCHbaLnNgx4kp+jgXPrOWpFEpz6ggsG4IWw9MSuPg
0rhO6ybdTtnuurBhAHfrAm68q4vS+hTQcDUj6djIDn20x7IDj0LMvx8S88BHTMOv45uEKguTehQj
ZJvVPXefYAg9mUrTHmEQqYBW3FIBZzZAQjWdmgOtDcVXXXONYAfG2YveXveQ0QOXlaZBvL30WDFt
ClL+qNM6AxOwJdJRmF+7qGUQoKDEr4XQ9iYk2c4s5hmma4d0Vfx6AC/Xb2i8jMvo6G7Abrs/tfc8
214B3/yZyiFvCfymooa+y49iSgvOYxilyZnSB20IYbKb1sM3OOPChIPGCf89Y/PCbX22R41j87xw
sUK5jxPaiwvPcRmfxuMX2/ljNEpbZFEFdP4tisE01W7/Ww7hbCz1EWHyk5jSfHFs3f4WbjmZX4sO
uLa1k77kMGrMGTP9IZ5W5CLol0XR6y2zI7BUFmj8FL85rW43TAcJQspVPGyKJcsYaJW5BB1u//Q2
lGk3c9I/jRgk9zRuZicHMa+SPsxTLllTwarcdur6XxkOahnZCuCM3QujyRlGCps/dSOTZzj8rEad
fkzsVSVEtrGANxo1p8AGzj69H2h9ZIX6i2AOBlHfZahmQQl0VfqLVXVLmHc7PjQK7o0Gp15zsynS
IczX0ow1fC37rwJcdc3Lwewre9PZohtZJS+w+c1uBSGcMdRd+fCECa9YzZjxXKnknS/OsK+gTUyc
XWH1Nf1dVTZxVgpmrQIA9PKr5bb+lM458WN2YoCgCSHAPIb95CKn7ItMqChvPGriRt2bSfWiMhxu
63BhjAIBHJ50vgvSFCn/rh6700Xa+e84I3jwHh9AzhahF7hTc+UDHA3pLXPpB58au+Zg/RZeFg0c
iknHenPjsWPAhmr3BvdSxCKv4hbzfPsq83tPBxg6xwXXntEbymIgjNi7+AMjIZTA+/Bm4F4pK2+J
7lm/rGA9p4q9jJRuwmZKbvxmj2h0hEnAR1QHYDkSsDKnVwKGWgFnnUf0JmAqtFvE2TuQ5rul23zE
4qa+WhvwEi9a3HhHK8ZBiUSk9d5mrQkPDQ3JWCorQ2u5J0REa5EENwtDtZK/Q9Bajp4xHVU4Snr+
N6UyAT6GBtU2O/WeUAISCjM6CgpF6p/Umg2RLNxzxxz3c9Qy3jYEbx3oogBTumie2mL0aLl0jugg
vOlkTHJA7N5c/tCVfAwVsFNsxO3sYe87sVV5mI+wwUvsI34A6vaFhhkxonhQnxh8UxyPVcdbLBDz
8qSJKNvHktBKRxNf6wpn6RWGM4Emv1+TxWmCnwMYXkS9k0VAaL0Dj5nbW/fvFrzdB72jAYSRQJOo
gDTPwps2M27s4N9muHwfeNYL22Wr67c6vyzSErgZyvhsP1+7ocMfNMq0rwBeifvslbaORyaTJk1x
1hZfFTCRy/NQI792yB9ZYu00ucj1r7put3ChgPbbVTerDitRpUQ4r0tK8/NF1wEgq2d6rMRRYCZZ
zoMBlcYzQmVogX6Eq02yXA9CPZe9e36mwNCrtywKqRN9/reWtHGiaDAEYv+ayCJOgLCrEFcoHYbt
9I6Ipd50dRBUbPOQegKPl5JL+3mZJCXSr9X7Y2jU1kY61pEU2qmB426O0uMFcCaL/2LJhxQxHVea
E6BbnjbmuxgaxqIoydw3JNEmR331oE9jSrsCfQLBIyeGg5hf/8JNff+XKfRYczL4C0t39NyYRvWF
bYG1FKPQS298cIl5/NgxV2vR8oR4jjFA1oo5e1oVDsg8NoCRA4UU9el/rFp8DI7iFtjMPoF8JHcy
MfSsRmOJhlSO5j1ZYD9AaouaTlc/er7LarBaTj/7bCPmmv47mxtHOLfWHBuC3Zd+M6f7kJZD7cUU
KEnZcR8sMi2EJb00bqZThxGCUEQGpgWy6pRExuqgfLIUlibhrPwIRprUQ2/Sq2snwonsETY7Ouk5
ZKJJlRBFVQZOu3vQilHTNXlWBoR00dQ+lS8OQkUyCHcp35LL2WDE5SKo3X/oHYEs0rA6StDqd5iL
poflv28D0rEYeJ07ra0b0zf8f/EXol8LhSmHpLte+fZtKdz7KQnLVmeCn+tNug4PSJgS9rSoKjLZ
IMa+8T4q3KVa23Hrr7qUhpk2J1AWTBZjwLz0Qh9ZTAe4yzDw7Zd2I9OhZd9Zu26KtDc3IvxVsmdo
Web/QiAAe2C32YkJIr+W+sa765vPUwX5fxc8hMq5kujBFWUv0Xfnflo4oqBYeUrp97xxVFqm6Ccz
Bnd+eMXrzML6UpKMCpwQhtHmLBFKqW1/ZCcE8xknHff6mnwOM/yFZMI6FYp+1nUpYgu2mlZoifXJ
wetnf7ni3vJD89d9+MkO9ZprTaR+Lv/N0fMME4gWRmW8UbvKIPJxlWcDOhs2PLIG13dXL/32y5nM
1FNdGXyr4zZjjQfPgPwui3tbFgCxb5KoAAbYU5a4JsT1z+AynJ88WsaF2shTGkbWHW5b4J40ayJr
z99S3XIE8T9rWV3F60/2DPSl0jJw1psUVzlEPbFOD1w7eE3p0KHlWjUv1MajvimWAWHB48mMjSrg
5MG7RWLTwxcmxTUbNDviwhGtBbfRt3WbjCrGcrYR55iziZ6ucqdJlHAPs6ZWs8ErjKdZxI1kEZyM
BgHjqvx17JHIzqg0J0uoVeZ+gEWi6m86ntSL+xVrPYLCSZ4bG2EajdF3S5eJ72lJxtEsaEOOn4YS
odzkSW2BjAUOzx9/9i840UV7NJ+AgqprkfjDXUn4BPfQjZ+5AF0YFao3kF/4iTc6aMAjYMl2tDUH
i84cWKIFAYk4nA1/rDzVyNi17f9204P/uoJIz/zgKn0WkSH8SNJeFjLyhRJVpmdJ4bbspuHjL1HL
1QdNsLCCCzlG1w2QzlcfFhWeiGMnkNux8WJHM3Dz573O9S6zZC4xor1NRkIvNzikcYkclrQRsgwS
oALzM3QU8uy/xo2vvzZJglWfZeGORFNBjRn5dBdNbIzrO5lrFm/gHrb3U9/dBhX0xKCXh9rMf8g/
3Rvca/PoQC9vTxNxx/mL3AYVtWlKZA+O4Za2SRr7/NvOqRvLpkP438yNMB919XU/ilyGEsJVNUVW
QQbmTrvJ0HB2P7S+UFHmtWdv+tZLohHoGJaJkwzPLyjGoZTE3TpDIDsVUxCbwtnEw8OTuegUqRt5
F7GaA/gy2uF96Jpy05S4ndesB+fotDdPXrnnGwjdLrxICPvyOffkdw5jOMHThs5g66x5u1CQsGfr
DStADYNFOoOT71RHDSQ3h/glQvF7uHgy6LAt9uEu8BrTUInAvEdWJ3SuSCGUBVC063+u5FrkCUrQ
TH9zNbtZ79sR41Torkw9uSFJ0gMOoRl473qOZoCfNU1jheTzr7+rdHeE/Locn2Bx4VRYprU9tKEE
pdkx6PUIILbU6ooH0nHDlH+UaAbCnVTq7xP/OK4yGACKxw9vURFp84uZUZIBv6ElNSzVCCywDEVn
EaKxVTzgazl01Jhg6yAvXZwYxZW4y7P5yAXSFhG7JHJVOm5H1iXqJ2DhgO7lXEHxa76PRpkI94tb
6Yqw4/vBoo3TXLrjsg643j8ssYl+ILhg2VHIxrQgOFzL1wMEZE8Q84XUIweitLyVWIuNzU5VZuFg
Sd7MyQp7ME0vElP+9zM1egpHdQvQCT9FQmrUGQig412k6md/sRWbt+ONdu7JbmnhB0l0hOhzR9PL
WzKOGHPXs+IiFnrCHE2AZTRdga9LiswSKszYmFfy0Dc1WmRNlQmvja0v/sJXAYale10NdM+TJczY
1+0WaqlUVAYWDevHrV9Xhxyadz/61ajXzv6n0W/XEVToywimqwxoFkCmaM0DWu2Waae7tGEEND0D
wGWT8bfukj77F2QZOuwIanizavW4BTQwOzZv17y5FCB8KLTEXKxbkpLQDAUARRfXAgPxs+iPAd9s
gohua7MqZXdaEE9xb60Mi7o896VmVMYfQk8TyIC75r866FMOknsJS8bnnD4R8i9Pm+tDBUSuRMBq
cBPq+NociRnYvaTCMJrk+SgtedoRTpFkJRM8rXFkmR7M8tdbDyvyhRcutK5pksAZa5587wkUtvXp
xIl5SrgeN7u5tMgvjtIafGeZ96sn0zd0kHoIAXgi9BJSKETFsfMghemB9ItqZOtvv8LuNMylXsDO
nP6b+s18ciktSXdX/v+JQpFMHdkBf8U7HTxNioap8QXp2GibVsH86QtPr2p2HODbw6zoO7nBN4FF
YDu87FFB4j7zkwVXq8PG32uyJtv1qjhOFLtwqoXJgQ1deRwjbXYFGag16+AtdeBbpf8y0Uyk4AkR
tMTRhR3sB93gwawDWDgnRJF4VpKrauxIiUUW0VnmTWL6HLrRpXLqwUkkSo+zi/XT4gDorQAUhxev
+/yNLBPQe5knoZRqkpoeNRzpPTSGK7MxDM9ig4wzQ9K4yC1CgMnKByhBt++6W/hSf3rYniVlOtrf
afBzy7YGqNuRlmMrCrYurxyEScqcQ0m4mpyOx8KBHsfTvEdd7Koba1xhXQDEDstk9Osb3FUkniiH
3ThdUmXpUJ4NqaioVMM1Mz9le/b+grSjlp8OBoXAYHJwRhelkXp8QxC3bjn/TnHII/PmHt63Kial
u5+ckT9URWPdgYpEZqLpwZWJbLfJ5HBLUI1MJqz1AoaRvM7GN7F0r7rN6Wgurw9BrOUhzL4AkKf5
DRFvChPC/cmC+xAMiml2A3NvBsAPKTYKisN/TBKjVcd3gcm2bbHqjU6kNlaNYk2U+rc1pJf2EtYD
LWlFlwgboiZadKT1HuooS9MPSuMp7nHC8iNLmEgmAVGoWTUUrlyya24GWIJBh3IKXvwBAYu6LaSQ
3ol3MAIHuZJr6V5zmaX2Pl2o0+/kpJGF53AY7AA065ZEGZlKz5e4od1lWT9OJwSw6H0BacUjA1C4
BuqizL/xOM8hFD1n+JCzIV6qQUJggDnKs7y96FY8RVgbhr7kjzm/A0W4ThGdxCVfmN0VBqtxaMaP
f0q+nOq6PFyRppGohE8xYGV4J/INxQOa4yLkLLO2fC5KR9ArVXiDq4seJUah8bAMbXO51B3j8lS2
nFrZ0627cX6Hhd2sqkzH+rS0BrwpGq99+OvNz7Hy1KrplCWFidIF3BqKmQLqVtU3bALgT71QzZwH
9iY4RQSbNaxlBcsWPDa1T1W3FgLjzDBjCkdtOOEyLnIWAjkOOgiDS9fTy2xlAhSTfST6vK4zKCIM
ArnWmrSznvTOQnLU/wRrNlN85h75lHRNlGxEGfC0v9kztmARY1rCHMU8gzyGX0YqtVufdFibjFWA
M/7GgSyL67fmbTnDPtMF1ZVMlzkl1Cgf5lUgfwiZCZftu7jtEuKii02we61niZJz7qbpFfL0BSbz
oSo3FH5MqzBXHtyIMjj4APOxYMTNl9opTnTPye7zTbVLdOePIQvAqq75eYvgRHaZLcBjIuKZwT95
iXCKcYIMuX6cn72Nyueb6RhnDAvFcYeSw3Kf31h9Y4yveWkoW28RctxaYGNZgiUsiQKPIxpnm0Lw
5pq+Qi9JqAxLg4xTB7vQ8JBvMA48perobGPKOT32hF97lnpu/6/0kW0tHN2pxCqibvq0YsAOH6Td
D19GOqCeOEp3swOgp1G8++Kiw2Bb/axzynLMAbFNbceuRiUgmau/OCL6N8hM9jOQMk/+hQsVYYgT
+WCLJDq8zluGjXZIfUmum7K+II0H1FoWGUcnOJ1kjnk8z3nSP+qMysktmytCDbUlOyderciPTjQE
j9WZI9bBzBMyhryGW8DHbF8/s9iGCn14BHxYhOLXnvfYz0ZhJYfII7Sp+g9Sn5cErRxttL37Zy3b
Pea/Qb8SHoFvif/Skpt5P05YXJbPmQzsFmpNpO1N8JY7PV2Y/mDKp1Xd9SbqRb3SIinwYOxw2UUQ
05HuO3eIu4Sv9gF7o7wBxhLenBMElXlY31e/qbJunFd7Sdlth68CnHXY9qHx2x8oIO/BbCIrpxKs
xrL5QB2fSA+vw17lyMxzfCynidNG6h977yL+YWEy9MhxpEFTrBkbuVQy1a9xyYfc+rSEnaje0mJo
PGoVrg2Z2cGVcxZGBSnKeL4wUwgupDDPNI0VW9e6dzUroKikeLOpIcZVCaVfrPtWRsq93mTH9LSw
ZLRczd9JQ8HlmNJSpTIr86s9XXJuTruDJWtZMnIdtfdzR9mZEknRdHztnxKTTy4ZwN1mfmueKJup
NLAP39h/l3XWpPFYImBsFhPkxmY9kB2GEcFdI4DmOeK/SW/7dczENlNgQcQd7OcRSvhyRH87BHPY
tsXeOG7bmQVPJsK4/m/4KsX8ChLgtXyJfL00E38bA4/yJVjBSAVIOAbdadjjdeYY8FD2rszEQRWk
x2GddpFqCJzXM0ITSEJDKoH1uvIIO86vOX6SeUsQJhDrgSfmAOSmnTr6/ZFhqr8WPfY4VkBDK2Ni
T665k18NrEhcgMmTneyuHixcuRcwr0ziVUstALfX03OnACj8cuoj+o37Rt9ZKqJ87uCZLcq8K9/E
lamWeUlQJ1R9gnVkxfGK/vztHxlaq3upYJx+q1ASVt9JYjcEuJZjoS6KccF5lV3QZF+wO8QeEhPS
W0NgSjFLinxROE1zt2dTjbRamG8RQbjXKMiTjbe92pyFYx2Iz9mUMrfTVeXvuV6dZLud48PbzCF9
kJZsrNPPLUcFfgTD0w9QELlMt8gxkHoawmO5CPk91fGmQLaicfBF7eshwdH4a4ZE1S9vR8L7vPMh
vpK04EPjrTV3tYfJ7V0E8VkghkuOb6FUpF6rj04jRbTU0l9QYCNaaW/XbHb4vGhwEYc3j6dD70cP
IzHTNRsa6MpwrFaYLTGNuuJXSx1RAWs1Pgeld/dhl95N1f56Crg2XEDc2zfh+LZUqwpCPS9lQ+E3
77zIU/gxHt4wCX3neY/T+rporLB/duoGsek0+uyfTija8wJpMgbaUuc5ZTHubeqp7a2vAMvCrNB+
RpCD0LMTLwbYtrm4Hgkj0BEkxCQurYTmXSu5QTlmc4J5XS+mY30Zp8qb8OXtN49ax4f4hv1+g/h/
cbjX0+R+zY1S6NKWKsnZuP9NfBuPjrgFNalcIF46hCCArriOR5Fvm9ay5A127RGum4l2tA1fvQxq
eIjpUs3TISKQZB2JyNrgx+ITwxnIToIj/axa/AVcq8gtGoXwF+dtxJRIbPSDqOt0qnw7Zcbmi6vk
nprt3ktH9W08F4+vHbEZQmKvhB84ILYldXW5CvLVEepWkrR77dsli65FJZbf82axQIobiPIYbcof
ECuneJk4qamHSBDVgWsNo6WuALjvd/xLZQMSjbFBOflQFGIRFHFZjwYx3LJz0tNsfo3oqxNTCbhy
gOku2Dk5HNBflfSHJNXyP1Ru6AI5HsK7Ixc6pQ6tPv4wbBVtZ1I2pNsol5kdejPJfA2IWkFFv0K8
sloSnSZQ86xUfI13y02U0NxD/WsouHkdhnX6MzjVwP6EXoK2lUdmHrBfc9gBFInKl0F6mRWsFsXo
LU/sHZuzimmqIJ7kESasGg4nEXV+VJyFfo/jLFIbFXf4jfhnNsj+r0F4USYLFLcD9AKeBJPFtjYB
0kkX6INOVa2zfSl1pY9i0s81rsKL2XA0r/SjovKrsoFzgfAxde/FI4yBxiykdvIyNHdj6n7Z3BQP
Q4w2OU6Ce+jLTnLI9DzO8MtdSP6ZxXhF+njaYDcjNEPLYkZhuV10us0edz6nrXL0lQxXQEhkqBia
93+iYq2rruZimqwdYp+vCoaVSzQUTYSEt27gB1ACJ8UwE2laaJTVXu2NOA+xfLDmDnOykBnNi5q/
uimPDEc50+cO62EZGBSAH9ZkrzWKvBIH/vUe95EaE03h4Htb1s1a3iVs6k2G6ioy14p4pgUd0aj0
O8MJosWQM2zeT/ag+7YGHch3UokFePS2z84X/3DAf/uQBmDsvfeUe2PzdXX3ab3e3N8xljFwn6Mt
yMCA3Z8toiwxNXw62NDc8h96SNiCiMW6ivoEEncSl8R3/MTzr2keubdwfi1oPTED2nyUcK2LTsok
uO04cINu3i5gZGec8Z/h9k5nB0PRkRnhznUnRbOhi9F9ccrxap5p1cLT45lDHcXmwb5PVk/60hZT
oeslJPmnWqKN3cU1dMxIHcnQAB4Z6n3bdvgRqFw+HGuTuGqn0ufRo4qstxl26weVlG7qudcu1i4X
53JanBUIgG5vzTnVk3rquVQwjQyVbjn51RJn4m9ut9j8PE3Pz+v41BG3g0Gmi+Kj3cfs0EZabZST
m6xo3OJ1mGb+Mq7qXC3k/O9WfzgPD5S/RqtJlZ/YZrP10Oi8ns5+rV4DcVhCtW08eCIfoIqHrd47
QKaeiux96wqnJqm/IzzMjJIMgsaR3q4kTfgQrC5QaZmCUJQ3tzy3YOQEa/B4K0HE1Tvrz329P7Ea
cOFG88t5Mx8KiL0ptOK/z5RVgT7Jj5thtysCvIOsSyTS/v7bOzGvKrUP0KQgLavQoYIfHASLeE7y
jkAx1Mu7HlSdsOCTJNksHRxRcnkxTjfoG6USGhkovfsETb5g3XzUPZPt8yZk6V/65PfPSwDcil/S
g0i1JPCL9jqdDmpAvPbxD2KUj9ZlDgz19pVasMKEEquOhqYeFg1+/BmcFzqqD1NDcPM4bffjBygB
Yp1ggPOf9QC7KHxlJhLf1hZ3N4olTivgpXC9JFdI4KM35ZAbiWCPWgvWu7/SH1LZv5ZD1xATBgNU
mMPzIQpyJBq+RgpqxWTqcQdnwf/5fSAD3NB8oxcm95sF9zxyZytpJHD7xQ8fTCSb5wfX7sAu9EWo
ntc2tp46uyUINAen7vE+ozUswBTh+p3Hgmgza894xHXV1JTY9u1F1GLweKFEFAHpbuCkURMUu66Y
95zSy+s0EXXoLqBRj6I2xifBzYWLJhHht177Gd5aB0lJ/MktYmFLbr/XlY6Bh0KgQWxV6AgH5Ikc
DiG6TnTK2ArhmjYu2OdUJ0p63Kqj+JoS7M1IDtig2KgJ4SiMIdY7hBVwDFhl+DlUAUWYSxAUIgiK
3R8SNFEOXYQGuOo3FDAKCIB4Ft9quatNqZUEv6XmZpT8qzKeRrsC9lcN2Mv2ssyKeaVPHrimeWTx
pOK+o1AetqFBXJzbbynS1/8uJdGh3HTfuu6ujD9DB7qGrLsyVbzEGL4x4HiszeiH3/8ixxGd7C+G
qntOYv5dhaT11E8dyco5volJ5S/xJzy6mS3XeH+SAtvjVOTbg1gLCKuZOa/7+8lDjJjAQ+NjPjrI
pmgn8TpcMkf8Yj2Cg6uhDl4g14DWoAJ13FB6WumU1rzFU7oSKq+S/NOSmhQ41jdyvAHmgok7eYLG
3MIoyS0U1fFPvDy5KFh/OCjelNoKhWLKrNHNlnnJP3dke21tFhscundNISrRxV9dvjl+qx7nzdXv
ySaIhXv/BKUky1BIhQWhlyTqOwNkNHB8U0AVABTsQKFOjpX7DmHVMxDXoQAbYyGjw8XmLRWEkCM3
Znx2bJqYvOMcN3BM5pY56QiHKTvrHUHsaLUywxU1vTBsHAp+0EhHWQifaYlnIzuHXSEca//sFAWB
Ac0I21RiF5liAwYyMN/sMYoxYBrxEdsJErwx9JK01dcXXmHUcyosLV3isoqVZEiHiQ1xTmHegyDf
VeiJSYMWjPwGWrvNRGNcVp/4lmXbgK2F3jY83GRRv0XDqvWqKQNbh2D6cvFcniccaK8zPZ5xLDDc
VBXBBnfEUppcpBV9s6ogzTT6p15cjNWyCEEuBkeXMPO9Soyxy0Q9OzxTpfnsCk0j+1jDLmwVp8nr
ibBtGHURiMp7h4LS87u465TIi7x0/lLwtKWlQSvfuEGtCr/HMjeWzvSfyCVb2fHSNrcT6LxShK/h
eh8J88ezJy64xQtdNn7JwbiXm80TJ4+aYesGXP45znKEFQU77xW2M+rV+hAKfr5dfD5N5FSLOvvL
CKNdIcvLsIiZgzg/S9tsOEluKPAR1u34DOA8qhGZH9n+aWPLXjlzep2/OG9RUrBvFtS+sX961L9o
iic6CS5IpYxI280Wh3+d+p5uuqk4Xp1zv1S6ffCgD57hhLKjs4a0b5ImVHeWAsQkYK1M9PygipbF
j2ByLsNs31pErP34I+JAXSWn7juW1d42DU+HQYB56OSV+UvAH/eRmc18vXaG11IlHzRZVY9jylo2
HcPmLVlZTo1f4SD/r9WulLW+/JPVSoKGDQ5Ipkm6xoeRzFgJ8AS3izqqxFUjssF9QOOITPpXDk6K
/KQE2KaOQfEYLB8sqmGgghoLNuWASWfsDgLwtQmjKS4UhxclCmnAhsjBBK0qnM1FzqoidcVxRduj
Pzp/DfMElA/h09JWtuaOR2NIpfQPu0p79stpffzvZRi7EKJKERQpd1z3cTcdu68xnRGy1kIqiVa6
UEUmX88tAokRq12O8iQZpTrqrGO5SwhzjUPjZrneOzU407tAtcSMNTadPyW/J0ScEyxXy2r4xnQI
GRES30VT7pec+PTPukbzXH4jVwCnUpzJdY6G6HyNyYykGwVKL/6oFo0yr7BAm9m5OhlkTknNE4es
E2u0cmELpd6COsi7rDHB/E+SGO3UW0VlLL+Qmoitt9KGJAOKZFveVBYu4sgi8tbIRgpCjif2VYPL
xwvqeD+hYtnsYd4cl6hOjEVpU6dOwsTBCXKIwtfn3N5zjeOdxQ8VyHEtmeRoDWuYGX6u+mCdIQV2
2zPBipF95KmUSN+uZL2BHFKGveftF7LPGibXX8Pj0qjSE4oW5wTMhF8x4tMq6Gc1F7kW7qfgCYVG
gWCqPKAOumL6GZ7IIZjI/Sj3e8b+lG86Df6Wasxb8sGy1h1notamvu+U9/HnT+HIASVQq4I+i7TL
O9R/c6+ga2/kxJ1LyAvQ3PMaePGVtt2WDpp40RtRn1+XeIwoOjECNKpqneLT2a/XxPiTM2AY2k7r
NbaEUPUQMTwKj2VDOCI9RoKorc5jiY+/baTU3bW1ckPf9wAk3224TId/c+5jkO+76sY2ugpcwlDP
WSMZehRvik7cLtDxtVS2pMHav+IXW3/oG3fR3/H6EgHF6fuWDgZBpW2KB3qz0oJ/sCtCSzXFtk1x
XDsZ9GjjrWPewU++hOqnNCUK1XrkO3bSK4chO4hjBYazLePZPJVTrmw/RWTu4hSpQXL5xDJQ7LVL
ar/F3RZKsWuGXHgTaOymzsYA+k914RDA5HZpK5qbo1R4JmT4hgPNzuuR6PfILURWJkrAx2mnjBmi
KAFP1SoF8uhPcsgrFpMHD6vEoDo/PomxohkxBZMfynR7xBq6Wq8Sk4gJBa2y+iMSv79ApQ5m78kS
Ppcn+BDlOWIMRkYMDxgOyIcApZzqSM4I/uMyc7MHkFg4CFkaWT2I+42pc9yJVbn3Czgh8DtkQQl8
Ci0NG16/9NeC7ykuo4xOyBBQj6s6iQdnTamg0PTQwk7f3zcPkPCjATMWV3rHKb670FudVpSrHYvr
oyB9+PY8eX+cpS0haqgMF0txusKpkcTnb+iiIcWEh7vAlmBQnKZHErzQV1L62AHAyPQHWLs5s2vQ
m7zIHf6bbWentWSltCOwF04vhAMtQakTqdfg4ofqEV592bqeyBuPuwOt5zSALgI5CZOaGdomAu/r
Qbfwwb3lWUP+qQsL5RpUyBuE/nLSE24pz0p49ZT6DEJLTUWDuFrXVscHKEjt5gSE6P7RCtXoByHA
s4s1FZnBJ44vF5v9kSTqse8IWxX2Apx7XkFY7/Xx2Z1/4W/R47lCqteUQ36rSLsKs4PrX5QrAgGz
rsuahVVLSLNAbLXpPGsvyvcLJSZdwbj4qNmZ/84g8BRgtQKEfwLiWTHvP7w07S64HQTeNqxYRIMZ
FGQVOBCD+Ft85qHLA40J5+riP59f/lRqFrqYWoFsaSuwfqdbwFMQtRC/zmS3MNuYYYzd1o4BY7GV
c5mjX0HKlo9+tEvm+bjFPdjqFRPJSwB514CBOlJp/vooc+POGwKfWKMz88pLX+t1/jlcW3OyFn/N
Ocw26/n3bHj+PjqRcZQdUC1kFe0UPWfGzzBXV+SanT4TV4bavJD7Bzmo83+zl3D5EEBBonyhNQV4
7oRvM7D/3a7fs8wmf2DLFzq4UPIZ4EpIVwC1swS3IzERG5LWiuduDMJa8O3lKWacvsY1BEyXIWbt
2W/YTm00JQ1BBnJVLql/4dBoW7bHJxOWsJUyBSCCGfYA393F7QUIpnHCKeSmi/dTjgnBIHDoAU32
jAQ3zNoFx2uZ28FIyHJaU4gMCwzyr1cxR9GbW/PrLRD8aDRyeHJeW5ycLVrnYqm6tGlIko1xSpEv
3NEczoFFeXBYN1odg50caga4XAPdc15tj8Tgjqf2gbNEMTyVBbSg6GVaB/ALRc1vLP21iGvpHIOq
2YdAPBWvq578MVLBR1oiVJLlv6TjWa1DwKCAabIZda59zh2UsKmmnON2dsI8dN5PiOIdg8Z8ndZh
HrgQ/MYlEA5tWKzZgnxPoH5/NB7clXiXQ1cFxeS0yKbf1CBiQPnsgjIZ+/+Y48qnM0C8C/zRS7ZY
enPxNsPaXvgLjR3DQPE+W/Jpn6qxqtkWOJWUwCRIETrwpLEhiUqZQceHjvjy2MRBq3FNNdFZuqSn
1dJSxa/Rm09iuiFzjaBcjSaIds5BpCLgLweAQY8gBtIU3Hu7QsumSc6fFFR0pp/k85pKNGN1QkMR
bBGxZr1NszkhCLMHT+2/1FSZdtPgG+qnnwwicbqoXBRInPjDoh4aq8toLE1c4iXGfMUoM/Z/fTvq
Vw2ZgUq3xgcFFezF93mwMP0u0MqJYowqq9HcEvTqMs9FCbOThy0st3K5A5E3xM9XE6yx0f6ngP/m
DSSU2IzsKFV8bjdGyhKeYB5MHO9DtUoE9G7rr7WKtcC7oHGEmR+DVKirQjHLuBkqPRiUMNmkTdLF
Xpll0v36r6jb6Ck5EC73e8gxdW1OCjucfjbkj+6DIKhvKNZ6ha3qbvhQKuUT4FOJQNmjq93r2KIV
coBZ35MEiMn/lVMj3fhwmhue1gW+JR6894f02ip4WALmCG8YKK7yzCJVhQ4IMPAxEnk/JtnY2cef
iZN7hA6b5H0NRXdcb8Z9UhKRCv+3ZCSusKsCXmtXAqcBpMCAAaF6vk7elg3Qa13q2Z3AvZfccwBj
i3JBFOW9uyQNRSr9J9udl5QJwltxTeddCi3zVc20RIhyHQ734iarVMQHNSWwekR5NdF7uEPtmanM
92S3mbk87AMm3EiPX84wQC+qlUhtar9sd2zF4XbI6sMVEZ538apD3fn4EAoA1FJ7SGGbK1AD01/K
+5AkHvDC0TlCZQiqZ4rceNagN9TDBsEllJLjpEfKmVwLul0CBwHNK1zhFVc6wn6YrsgXKm9HJdix
I6+CVKiwdmyvcRuL71Wxei8a0P1F6JaYN4DJ94jZH8RnQ5HXz5tQ6fZmC7kqRWhanXrzpUFWRlU5
ohz06sYWwBB69MLdYPlyE1XgmAchKoP2UqwSwAekW3l9jfbVM+SV8MOkzMTUgCf4OabmhzNCXepD
3Yp9i/P2zuaKRb6c1s6xNqNSGZi4Go5C01XhzxGLWKjra2659jeNhHmQynrsceULUQaz4T5qz4OI
Erbzedx4HOH0C+jH2t7t8PUmyRDXZP2ltU2JVNmof11jBa/Iqz3lNsoYr8WNtXQxrr5mB25veZm8
3X9JqGhHrA95iHMB/3FmBunZOGhSs+oMqCpL0PLuc0MyZJ2vJGUeALaR5E6csFpNrKe59TiPDwgS
CJKFD7bpTi/ugw2XJYxRmgnwPcjnwMtSxR5TBbXHDxj/e9XyvSZFZ+7fgzc6JW7swU0vVl7LOFZy
Pbwd2+pD82eQNY3nuskSG4ot/g5TCbXPNvNaPk6ij6CcI0X27uRVzxIEAEj91nKA4nUXkc7ucpCL
9/wosEpzi3tZ2+zKsr/VMjMLTI2s9gwenK0sxFVrHDBc9e5XUqsljE4+Up3+3CSsPmT4+WJVlj+Q
m6S8gq6kOUa2wmqaijG9UdMMzdZI/2AgNmbGTZw3JUoAwRfEjmFxUTOYqtXnDjnD+29F6GiMQiu5
clhGmqPrIw3SJEWF10I2R9zxqq5hVB0lZ4FBRAk5rZ/Jw2BAK8mUF3k+FBHXL6Nb/GptxNIp4T6u
Oy/RYZHQTu+rIqj1RA8q6VAaNBmgGtyt9I9BEyEUmNgXmt15o52xildwG/lfKB4nekrLOh+rlRBC
eLDuSoJ0uKkHLuI3/yST74L/uujknfXOYc6c52lVwSS7Pg+hPeklZHxO9XkyLlyhghR2zmWBuS7V
MIySeSm/EIWC2rll3S9QdY62XibthC7R1WwmsA96Y507lGc7nwh0iofoRMrAQXgoOLPdNnBgZWqR
y4Z2/hEb6cPVt174Bi4Yg83Xpx6wASXSKVtqaQAiC1Q0Wws1JVBb2UYCTIstIaE6yKTap0t9GwXW
vHk+ANdS8JM3baNcNmJJc+LvEJllK10ec6U7So+zx24kZPSbAFJCgawW8pELnKoIE8KN3HEvRjne
TumPYDTtMLq1IUeq0xlSRozjS/weLs2rHW4gOiBMOWvMeeXzbQvayXsnB0JIbrl1jlBOmVB/npQ6
9uCC54yJER28AIbtNZPSMLaJdUOJPnR8a6PDxCNcj4zbWJ3ynNBjtBw7URkCIcYQXcNynLD5eVNU
rvd4uC+Xs8KMqdBBhT0tZqJ6zNK2c7T+TZM5OalW0eXum2Y8vLYkM0P8JqbQ5QtoUM/tnbMsLbvl
JmqMp0NbovI/At59cb8zQIoatFK7DRgZURbIGvCksYYQdXqVhVy2qhTRoNXVMYA5bezgMZ103e5G
AsvCIOYojsvnUztso6OzZEs7gEZ1rhE57HRA7UXRhD9WjHl08Li8V8XMp6qE6dSlPZrRNBxr2rDO
dPIXgqAORQOLzTnxsQyi67fj5EPovxjJPm1CB6zi++jsR3txzH9CWZUNZf6aev1Pplh1TXZShQKx
RKQBXPbq5IXMwEAI2KWAVu9Cw3Cd8EEpzHkQY+qXiRbFGICmLXaZjaGitYXgTdsq5LJgUfstT9VR
Jqm7G54grF8zdrzPFx6qDRck3WOFKCztWVWUAxajQ3DabKfq0KEbQN6OKT35gcb6d6wmVzNYLKWj
V0X6lYSB1aG08kQPwLmo3IlKVH9Yf3WS5xaypOJWY3U95wPMtcA1yeeHySaG+sm+rkwy2ZvLgqPD
1yfOwXvOvvE6JDsYWM4flnY5p2dimqzO39WZJACljTKXaui5g3UVqgiVVEdelMKD89A5AY8oVt3A
8uwr8V//HRk3XHEg8Tj5DQkVvldN+I9E424HNMu7VE1hzVzYeg4Fb8hxfpFIbqRF6YRjEFJlMGcU
M1s+SH9X0fGUhvrKMPc7Md4DrWbb+/2lT5OYlVc33KyZsJBAb6qbC0Qx7VXDYJUTT26l5boctkHd
IRt6jFtOPF01S+Ejm7YgZAe3Iba+IkOuQcsLu02pkS0bov5vU+Wei5TOt58GlZ6JrsaxKTO8i0Ix
TwC7Gfsdg6oi90M4dpY4BCGh5j/EJFJAcnRUT2LLI+yLKHnMfUmL7+Zo3+ONs+UYwwgt0BKcxCSv
I8g168fBkxir3CR7HpiQky9UoRktQIaXlSyX/0+9XH542H1c+M+srN/pPj4rQoT55YCTh2rChcqH
6EYznzbg4YgQDTE1QkhBp3/D9odgGtEeRZWGO2tRlh0cFB/LXszELj6m/R1tFD1o9PWq2btTKWMV
XY1dhLU+Uu1K5DMMYJa4xwnz8TqCswA3VMpdCcFbBfH8PjeH/lSiPxm5u5HlnUFx0kZ23Y/kPqR/
twyJsjwDM9j4mMpJhAR4TmKn5e99oF0DY//b/Vz3Kv7iRAc824Rg69tXUfVd9KGK3GUi3oDUMZFs
O0vJ6NGAnaPTeGgnc7B1K9eDgdmkuom4g+ICaVBZkMqOU43l0pV0Or9s0nRCC8ajbv+X2RP9AIZW
JvmdBxmY9EWQ80UixoP8Uui9Bzd/Jgd4jXaN8sUB50nNZ2bzLYHyfXmiu8yQEQxpE+RxZbF1RznY
C68kZXTBTsL+mh6T2gqlNj4pwhpGJo5vwa8rQkO8xElkOJYP1wDKW9FiCJLuGO0zlURmsXjyruNr
B07Hr9muCycvG8uGRm1KV2crp5zuZmYgYw/to0UVDcmqbLOkD5ylzuBIhLma/nvIdrT7tnG24Qub
zy7EVmbwCnxlNthKQ22MP1Kycu6jZAwBcKoizyQuoicnswiPrk0WHaSmQgyFNUa704IApHqUFpfm
rR5mQ4/6va18VIl0C/9LlANkBVuxMS/xpvK0njwFyT79cTSF2xft5u4eEFa/BRWmWgKjd6tJL9H3
LsqPiDto644Tfw+BSDE0oqWtTKsQMylOwWX3RihjkNeYDQ/N584h8ZiswWRDET7omThZ2YUtEka9
ZcURVNGaAvG9RrM76nmJazr4wdFxnO4fpn5PhDINp6gt9ez5434NjCQPHRUGKSTSWpWuZ+5XRGdu
IB/uOerXUCv6biAlnfEnf4U65uNwNsOHK+KBFolOpVgyMSFeq8d3rZS0g4dUW9bI7Knqx+VdhQT/
4ZadrBsrhAmriJqOPzLUPQ9nKkpucsIQj79ZE5yFyUuqh53l2UoAHECppxxUjVzxWhH7gjnL2ziy
REa0/jar0nh/PnwDYcP2hYJUQJ8Tzz4TDi7XETVs80QQ5BYNCalkc9auq1xZGY1NGUi8GEUEj21+
2URF89/RCmpYkshqS0p+bYpGMdySLw5K0URvESv1RqoTGPWUppw34IEgUYYd1SQqhwTunnnwCkWF
7DjPJj1u+6DDzc81uWNo3dmXob6nsAFciCj6wBORKtUvBDEUWbydxvq+OHKDfKpNWGhYPT9R/jPB
v3xM5iFdAgR8/oOst6Gr5M0UcreRTNdPYxZHAhKtfhGe++KSwT0/MJpMeDaTWL37w6+kNefGKJ8x
tVPY8rcRCgHyI0RVmpr7Rjwc2iC+kjnCUucKPfWzDO0Aozi2JfrT2HPpFG8QjgX2Y1PCalBrN0Ri
V9zh9y9tv0xRobLV8eL5A+rYtDtcFtfv3T1/ihzqaUTtfddzoHb2SDsxKZ8jgXq69iNIUYqr0IyI
dCYWswPeNeSOp5ZNg4qVjGkaYnPdKC1UdexBaAnjLBbG6aNRYv1cMoVFGlWsoDVcrIP7Cmy4Iqlo
G19c0IFrNJR5ZgTIV0aiby2Xrf6cV1x5AcG5fvX/gx3Yx5v5jHhgpTl/uw6JIL6SqCI1sbZ7WvVX
z70KAZBfCoc7K/1J9FxnX9Gy4Jn1er1qHlOXi7lvNBaryBORBIYnV7kHPntWwuJ2keHYslKjsMl8
IdB/JpxrUrCjWZslMt4kB8FrdRibvK8O4bNmLod3Gucj8jSoImrSuOxUQj8pCvT4i9/1vC2Fa6kK
48rmUqy2U+1V65AeB5Aw012QO8sHe280Uy82/NuK9r5VNf2Si2Qh3kHFXKGICmJxQEjsuLXrXTtZ
NYcH9ZwFMDaOsPfee7qZUK//lg5PVEFmHmPsqOC+fXzC+z60cJ9SXpLOPoLBojTNGIVAvrv1QmI9
QL6yB40avwNluUXByUwBsyFHBowXow97cG4SVpfiz/oQPWUrVKkxW7YapMIJJAB4c0FdrbiRvPv9
akRb6V3+j6XJuhuMVUugQhI9JK+ZZ76ePtwmvAivfSV3QdHKw6ZflJEPkUk8ODW6H1rUIFidSqoA
wuxI0n9V8dsBVYQYONwvKsLnWMpiHYqDjK0fIRjLM4+FgBdQB9gF2y+R9YOHzP1qVCL8JnFfhNAA
LHHJaznDf3ZZP/dHXzmEKGZFzyiSPtsUq2A+LDrNV4Fixt9aY6HvX+3+wKhV68AuqkdjlFntTFCY
t5MWI4ZOk4N73jFGZavJSszRiWXe+ai2eVOw2GVelK532yFQAEJcMjvE2AHLhIUkxcfFAhgbNdUa
NzT01EqRuSboxHqWzrvXqMehY8yQFpD0Rhf+kFdfcoI45JmJ9Uv8UxgHcenj7X7PeWVC0P+Mtjqc
IjaRKowH7VzEy+18k3QjtlnvQnuL0/DXgDuHSdXw22pHp0p/+kzuCIiaWZB/wI89UAWb8ekX/Grd
Il+/7i8JOA8vNsJo1bSYCU/8PRzzQFFAOWq74XCoTTyMiWVgbfmMKDhk9oeX1r3mz6lp19XaCEoh
R6x/avZivaj80vRH+5dmLMcM7bPnaV9IZPqlwE99g0MwYAUrGdlKivpBM555ytIDnKrW+BbSUp9d
7z7mnS53ZMqKBXvXfXjVNxo/JEJABbOsRQmE2OrYIDLZ+6vY8zm4exd5Sm0IRm3iZkzfuG0rtHfI
HMAMD9sRQlky+/L4kNpLAdS7x5k1BizXJYn5gTTM/Krgt8HKKmEe4myvIgNVmNJgUVhzThhjtVGY
wLT+K9eRddBaTCvQiC9we73Mdr0VPz7/eeEDx1klFOgJtQjz8Ci8UeCBOCDOho863IPHOhc6xa7e
4dL4SDzyvyFpSbkX2WbXKRp3DJd/+cJBTXiu9n/OS4BqZQRMzHV6EzL6tVcZGx2DHHnPoJ1Vq5fL
Qpv/MH3UYzvPhEPyXOmzyNwU2HoFO4xBXgjVTGiLh6R+3vbHplRdiVELVGu+YDkSEC1Yd2RayjzV
LR1ajX3jmOO6i2ZMc+CKeAYXYDvB1mScLWPq3iZbpx9a3isNZAi9sv9wUoUjN4JK9RiQrN9fVJD3
VvyqfLtFdPn10iZh84aUPNs8p6g4Js4kMCBmFor4bJJBinuDKSZf6rGFb/WxCbcBWRedYmAKFX/M
1DOVNDCmIoKCeQG3/DpXOLga7Irr1Gcn4zzC8H+WPMdQGcCqctWjWf3c+iXRBKAdta96SFTgx295
2DEguNTLMx87P4rlcm2rwhc1NtYXVNJeCI/bp8Nb/aq59zfGmNn7gLjI6JqB28v+wN29dz/q5BuU
Ea+/OzeOjq1y/h/hoiDBdSS1NkZoWUIV+VDcrTQ2f7130ZH4VQVf39z/eK5lddBdUWvb8Jk6iVwI
y04iSLpT75KVUOcXn+fa3GpycM46qaMeZ5MGfG0XnT4nmPX1CHL2iaT+BYLTAVcE69Toj0fwBO8i
GaQYpmteVHGF/ctTNdYJ/6tpUN8LhPKgsv+fsDxBJ6dGIALKr2zYsx86Rcve3fmQGj/dCEfoJrgH
D33XpAcODmBV+IPgY/iNW5O8Ye7BLtwTnFHT6MyYZ5jbhXVLjBIJm8veEZzEmpsPDQSO0NrAkitW
//BRqUh97PGxFMnd09yyd2PWNprZ/GZoHrJD+4xHWz8swlBcfZT5OUDCg1PJtu54FB1mftDOFHQX
LZTYbKxszR8cplNzXex0HxqWLmaSBQ2JUSXcpbRCS+M7EFM9JaiEC9PxIBak6GakQXURV0BPfap0
t0LXa9H//N/yhnehUNvHd5fYvpeUlB/uFElTmZpInfSkU/6CEUP7PcJLEe96vPiw6UE+8N1w9Icg
pIk7VCCmxE5qFYrcUCgy9XLQM7gvteIOF/xsUwCV5HyUqQXt+MZuzoJ2oYk7/q8GEMoDw9O4qtjU
s1qKgC2AT0ra+EOxSdNlCYsNI1ocmodyY8E3wq9uUlM1a6JbkFBPhvjDnwTBUQII0UGfvM9ctX8z
v36z/mI0Rzvl5s45Fxmj7+XH1ZHHjMT/uw0WyhkBMJdPzYfqoswUsUyur4MyUDPw7QdnmWMgMkPy
YSge/Gxy12d7cTD1ad3CmWQrHZYggz8WDXMjQyTy1GjaYiUKFbENcQdQLPuzvYfh0mMPYY3IJzat
B9/bAwB2bie6XVtm00n/4Ql6Ygy4rhvuNuuttAJbe/tl+10jE1g2pQBpWXzc9AguNJn7L25IX4O4
vECzh2doADtNBXOj4JGsSbamtcCA0rv9MRwZoTYIrjP1mHAe5KuDi54KNHPnvfsQHFKi0fPomIhN
/iMDDOYI52DN2Slj3j625HV9rdMeMgY51fxblQFyDbAHXvPtj1ifk4rYbBJ4L0F5E/jaRQsb9wSo
n8/eClQBVQEHcEpO0trrj+onUb0Vh+2uyRkTCWbVVvv8lu1vUMMud8vrNmzy0VqQHo2OvkyNFFYz
HUOoVA0Miab1Xl0rPGG8fqv/UMrG5RRpc4uDKGufHAjD6A/I5f7jBgby8M9H4dbdLMa8l4VniLk5
SiwCKN6vQ724MQVn7MLpGzfGb+6m+nAbXoU6/Z/3whw8wZ4wTwC1TLSu5S2UjR28DPJsyhS17ZbI
bnTzaron4xG4xZnlbMQIJ/T5Q0Jsm/kcY/NButD0y0yPTy5vXqjyvyvbFueCh0K+gU7QJIj27YvM
4oKeP994KsXhm0BJRFd1gIvPHRMctjuCFGzG/UExNApc3Wz/qDr4e089R1kE8QbD4lRqbj6YURBG
5C3o+pnbNJnWwdT/GshBayegKVq7RfQnrdg07rVY1RxSiiPwjUe/urkgPdCHTL5/prs63TMB5s4O
PR8vMNLZ+4n5gAiKxrp3gdlqg74j1cgMIwIHISO+JbDBIXOPDhB4Sj5AK4jj3c4RsCPHXUpeWWCF
jMVsGg+8s4k+lTxAEdSOm8YvVTXSvmX+KI/Tzi8E1nL3Gx1J7h5nduj15MqF6nlr6zHbGbQcFEaE
zsirGaNvf+h2LdbaZpN2d50ffOH3neV0A7JnvHqDNWmPtDHzoa17CiydpE4gef+DfmJWr+w9Stfl
f9+dgwCfjIZ9fDsah87QqklNX2fyuuVPmBazIzPIY/GvqUwQjSxgY9oJxcPB8kj2sxprj4L6LHpz
ey7zQgluS0EXhYSTyZie1F+y/91Z7s1msA+uI/lg75cPtV/wcGrwkuvbIfsJ/JJC0MpxPHbmsi8B
g/a+NaEkBkwh1oUQJwij8wW+lldiZiJ34N96qmA5SKGxdbxs36LHwDio6IHYrWibjtKQEAGhcIzu
rEfiEL2rQiCqCEzIWstwOz6dRIJONBSfIWCT18YbAIvobKRzb0F1b8nNfpduRxpA4GMRfJrmXc7Q
2gdzOpfpIwrD3kITUOke87vFTbimfIvoYV4w06DKuH+BECr2LVMRQy1PHmAaBXiRumm0hfCzmeDy
Eog3yoRB10mVyd9Fu6zPQBbBDGLTxsSeYRYPA/oO9DeHPUMhPsOQSAtxht+evVRKl48RBrgibKpj
3Zs0JXKIL8jQXzal7kv/ypClCqrTPWfICbYqzAtRAi1UJEN6AXzEx+7wXzP8Ay3hK8ifwyJ2iaRv
qk5UZb6TgxyFsAW2ADY6SaHHEEFLh56/aDaVt/tGEewQsPnAPLNwAJnEZ9h6YPP6CwUEPXdf15L3
NnJ9/jHpC9QDNnVFau2JWApG92NShoFSfKdtMY6Z1djIg0ZzyOgMHWy0hqrbstlPXAsJJJBbDoCm
apC9N4YaBLUcXhXEbgEU++a+8mT4aHpvpjYt0J7rYwar6VBvVKq5DbxekjrnElXUd1EjybIXxq20
S4zmerzKTGahQMTDu+58urHD+ZplAwfhR4r14QvSVrrQ+ZBwUykGDNElHvSdX8hXz1FDf8QYcFYp
6cGL118hz2FQrPSC+0nbK/BQaOH3w9RSrQAQh+iJvUeiTyWV7GPb3mu6lKqTyLNGNDCAzgwOBbf2
cvDQLG8b+6PA6TGi63p3n37o2xUxdYqM9iuuSuBKA9x97l54acKfWbLYfGMCmcCwIyXkTTbF7gKI
/sJKWaWYLFoa2bKR4oO3P6FAHG6hk8NpEwPWsVRVWfirgi5UwP6IY7xU7RZLmuNH6cVBTbUhg+Oq
3tdvIrDiKujckIlMvu8ki4cMPYVLvLiA88lr6+VYe2ga8MFPB06uG4EN7Z8/e4ydIVLN+QKY5NDP
sj9JNFC+2W0b6Yij3WAl5o9gKMMdaMUkvMQraO0TyPDFtcRKS6Mvner7cf1ScFfUeeDevf02xDo1
ZPM5wuMEE45+cL/zCISgmuutwG9p/H7fJxGkpXOfbcGp35UnM34iwDbPxtDaKnXJcDkZNRqa9lhI
2fNMRP44lcE81f6R1Ct7J3QoWAWoC+mKLvYykskhEzRcnB+EUQycx5DoqVwZYnnfVEScZ9+hJREX
tUXlmMylH4ZTFGgg7D9U89H5VLDpcY7eEYFuzxtHSk/2yiyOPpeE86yuUyZdnVy0fUq3kS2r1f1V
lvCwn1jkCXx+PQqLw6L+7LotG9mhmtGNZluiWWbwr6JDPwZt6DHnZQfqXSgpVPCUhaTtwehfJOZH
qtCf739jVSk00ovrfJA1mAbXOOETpDGC8KQLtYg4ppORMNFQdlH5GoL1v6G5T7aez2Qj95Gm4a+x
nxVKD7JkDKlo0LSP9990l9JK2/RaY0qQDRURFjjJ7YhQaKgsXChexLVdCyVsjfbHT+TSwECp7HW+
nW8Q3Ub5WdDqrqz/yb0dVmnnfVmG1c8QjzqxXwBY3Ul8QqjudMtNzUg/ErJxxjZaQE4SVYliY0+p
eJsXtfN9KP5GRIJHGluuir4oUAzMhY3ceNfbzK0ZALEJAJJkA4NTxE6gxEtVqE54ALA9pktvpQ7D
8y4RBMCROTR1Ebf26boYplRTdaj0bMunld5Y2RXB6Tc07mgRiZdr73ltU5o/tsl3W7lXWVa+SNWj
UzYWrKxSQ9oIY8FHd1d9aKCTq6ZUB9yjNGNNJRMC59oeCKXA52Ier2HVNx1ETEQg/lbNrs3mUeIF
k1Cp87urC4I3Fwd7ihFvZc+T1FdA6BS5kvdv3GvN1b2xIRNlLF1F079YjrKqg37TxB99N7qXjLo2
CQE/1MTTLN3FuAvo8v1UHKu3bCXudWt4bQ8mxRNZ7Ob1Jv4EOsBp34fHkv52W02V8ApRWhJxhA+4
KlYm3+rh7AK8vm/dQXazcDS1Gk7QYzf/02rHV+CMLMURa1MgWaceX0SaygQeSIiMsp9+wl7rBUg6
6gVGbsz/zTiZU3Dr4ulUXGk5jrUQzlW7NdKWyuAVxYzYe48GMBj4lAf7pESZk6yxb/xmlEx8egEN
FOEHopl2zKZIEdaquTmwLK7+3DfAKINsl0C/qgq/6s394MvUf9bm3bNqIwcmPKqTPyZorHT0RQ23
WCTHl+zj5GXbhhuq4S8FMXsNsXpgxAQ7S7LsbNPaJbGUWuEAL/2aFYIkL1Z3uabt/7RfqVHd4WtF
9a+z2vEGU5H174/kkv8QcB5am+MV+JWmBUDyAGd8/WWJK5CDyso8UAECNouuGzQCVy8mcUbF7Gtr
E/X+Ok88Jg50rcRZjmzvMveXUuErEg7BALeIjJQtm7f0kBwK9eIMaHcjNSfg5ohv7w98ksF9WSzj
LMiI5HlKcCzur30fCh5kPtFdyLYSjRtXsvc1S1beOr2vbiQQej0wSF7W9QtqEBcpp2vjJOfZvogi
W8BNijSY4yvnKIGje4Ld2TmOVvh5B21tZWip0eY2d51K5n8+c2svJ+FuUc7N7srOmEQRTs199Ike
OK62h+Djt5/TR2KGjpq3IstdkRJcGJbYM8BlNO+yqsJSy8wKD9xIXQUxNhqLpH1C6ctyvz3P7wZy
fSz/aFdEStRooEoRccKNTpSN9sZSXCJj9/bOc4OozQirYOywuZHbNmpDBrJAzS6o395OUdZ6QYsB
a0tCtnjmezfOaUW9/xCfOd4HrU/L7A4yDNO8qADJrEctmPp4TnTdMYlPBfMsBEggwxSMmnW++Jia
o2Y2XLY6PiQc0Bc9pmfqoNqs9pS/BtrUYhLZOiKW7/y92UREofVbyznJNypRsWNjdx2CuM2m/xfV
3E9BLZrHqzQClbnzHdEqJ4sgGXRGosIL6Sy2FL4Mt4CMp5i5mPjE5GXZVZyJDMzX4ubvZkPXkqkV
JZnDXgjKee1kFqBPsVKDhKAchIQ7WIVHNXsWlgkhRhUaeYuQt1BoPW4kmNY9vJUQS8jyHIC9ITld
3V2+I6/UtC6Th6rpuA2AhEm5Fo6mkLBIyG9ttXG7h6vLcpW0fT0fIYCvEhZMMvc0FiGkQrIRYMwn
yjEIqqWMTWj7GJRCwZgL2qbbtu14KEE1nRqvPiBsZb9ml57zotbQm25H0Qye+7H0XwDrCJdZ8sYH
k1CNXrr1Flecb1UKEA0pHfJVGLnMygxmV9kqMkRFRODCpvT5NdNdinJABWsjHkvcD0ytBWKHfwrD
3SsotWyzVHGCtKGpmFktFY7jIJ/tOIDbMExwhb349QS9MhDErblujurp76+4PVZDNVNUbyrWpXFU
34HjFw0qRjQk7Y1s9/cPeMo8bFFY3ShUypecLtXUg5B/mefyOLCriRw299NENiLwNLMA7DMwa2pV
8l2U4Y6rMnt4zaaKHgRHq+ncrcvh9Ui0efLFqG8J3h0rpJP/FQWOjCF+Yb/evlmcYa1fJA/jzzkX
icF2wsDrPQdxi7ShJf7acLLh0E8dXFjtQ0nJDgUC8mbUp1Elnw/XZC1Ze6OK7/eHYk+0/HtUDdi3
DCRbhUTiPNbqwNCL983rtsUBbhLfp3sfNSkUB8gB1phOuCIt3k5jj+FM/rLQ75UJKDZdfTHtcxjc
ctj2OWGjMrooeDyKX7pmZKimH4OHoDGj+0e1FkzHK/lCqNIzn/N8nnbwY6cTip8bJ3SfR9Tv1jrm
FiuyoNblAMDvxhQKHqypjKpqlcXQjXTEfiIBleh5TkaQ2A/VYpVsA2+gzeGZgeSaK15W8WwbDGAp
TymZQWiRNiLFDUKTQv1wonIFCDoT1ZAQQ5waSht8V4stXAr0lezkYHxvIKgOF+BCEBb4ins4RgVt
ysPnEpUcijgajgEUbMfC5bG+Rik169U8NEDMjEmgzD1ZFVxHNQxBJj0XW1V3s1Cs+e2FGPslgahT
qyI+TLLEbniS5/3pbDM5cyeFR1HyWi8c/la1+Cw8aPEml3wafU1LTtmGJeMrDF/ny4PKc1ISZ2L6
NiYbriwEkEg3XOxRFDIehJsi6a/+4h290NdNvc3kF/r4ptGA+WHmaORMzMZdepaG7UKe1x3ifevL
CFoxDAiFYfSoD15YyAyQYaEKopyK8lUbuT0ys/aJt0zs2ZCHOFmkrpiTprlWSvzovX7eeJ1cI2oq
TpiizXSo/zzJQ1Hx2Y/FXUUmN11gQu9zysVXIeDkcUXydOQ8iq8WvpBO/rsXknXE82GTfAmY2Urv
fWa/g9xe3/oNLEpEGZ5rOL9mVF8Zys4azWfpaLUU5ZK6DUkJQrNHGgNmYLUw4hwSyjFa2QMIPfP0
R7CeZNIAMt5q9GnnT2iGTXfLSmnIj6lljjhtMBJGnvYVFdFi6cI9bA4vuKIbh/Cwc9w5n0hm0Fpy
WguSuPnLxwwDkAgSexE+Fo+HPLCF7q4frvDxb6poMNaJdryuy2OqVJd+rdse8m9hR7ox3S3T5m+S
ardnSRX93kNWd3ygpDIkeRLFLPxpHSa6TCCKzDJ7h5AOsclnDNRaphALLZFMLq2ONFenXGDpK51j
VhVcX44tL0wjlJxftc0R78S+dUTNyjOffM4Le/OOwTkqfYbvs4arzWwte+tsc5qyYYeq/pEkRXKC
xjJfO7H3lMFKds1moKN66oQPgjo244fAnzjldUBSChM+p7/qQ9HjlxMWjHnBIjdmBjmJwDZNecLx
r90f1+ZUrRerIoI3It53hGUTmKFUCUWZK6Vkhs+pE3f4jt98fbl82FWj3ScYOCGB6c74I4xHjhcF
k7E6ld+WXQsyzJ7nownFoHTcEfbaQpBdtDaAEKgVI8AHiYlSnGPD3It/5lmEApERnQWlQghix1bT
SpsRiv+x1p1sDx7LChrCWrWaYL5BkMlk780dHPfkBXNfV7uzR+xaFXDuHpm/EBPnb7zvxJXC8Mmu
BIjgFoqL1Vy/axTcsBa4kyZoFQ050YCUSvWqA9PjJSKtF4A4PVr5thgU6uMd4sTsv1n6bDhNlaB8
hiCodzvkuA8MLuqKtBWYtaWTMNuuSeDK/TTo0P6pGu27rQowPVhLHMOKRGedfgwsXdLdxPbPSGGm
8/FREWmTLNdkeitHBOAdxRxALdaRVBMVePpDELbsGsQxLaMP0G8w2JTqRc/hfPcoArRRjWSwTTYr
kTwTynvmLMhtcFngWn7G9/RLCKLgi5t6J/8r/7clkIzKx2xs/LuTEjdVN+6CFSU3QTRmo7w/m4PZ
4VvcSuHGbBBvAjTqjYMkGYsFQtEJEkAUR3QQfwj9p/G39xalkip7BIQZkhViRgnvLL6/OPm9o+fr
gcaiK/TshTj0vXJTteUK8dwXht9STDyTu262vEijF86dSpbf5/UBYbouIM2O5zf2h8hSFJH3vliv
pNX+wz4GzjqD6r10d8mPRY7Yj4fLA/o8Ykf/N4d2l+gl6YldyPKefOqhZQkI56yGh1pxbdcmdOiW
4dsLo2U51452yMboOuKm8wJGORmtxfyAq1aStQf0GKyXOkvWhLDnpHQkXG8v/iKPSoedJdzAYkzK
kzWjRbUpCZgRc5/IpVU7KLq2Cieg/FzsLVgEqOljRjAhVVZtx99truhaGwcpySe1BuIgK3pJXTU+
QyxI2zSoGBB5AfLDJO1vM6vHa93SagGSeyrT9yETBbdcBo61EfadwahMpke0xeFyZop8YdPXRj5k
3I8COPP4VC1bMu15kjdeNz7GhYSpO4CtPUU+nCSnugZrwjsQtKZxnqmEaTE4lmmP/9L3/yMlh1cS
l5UxFIXjyJ44TV663nmcXYQaTT9HOPWPzZx9BlwNUKr2XQGN/jqzlXIvnsgXQprcXFAACfRSPRC/
Sz/pm1Y9HZgazyxVeTLPqMEJdRT+IQIEvuL16V2NOLAGHhVqcRlPymsJscRBdPXXOb9JG88A2Px7
1Mpt/MFC8VunSdl0rqO2TGGr3pSQvJ/YJSJW83FPjEOgRqumIIXfbnKXAJfatiPkNQyQuI5Ael3E
pA+JnyF/Kp+STHcm4DQJNgahVk6iuJco6jROKwSfk2G3p3Lh37Lk1W3VxoVFKvPtWDYrRqmCZu9H
5LWVlWubtzkC6i/RgcuHRrcjsmWQgKLQOzS4EV2oiKOf1aTzaDy5S3pKKvca0U2wmrO036jCWQ+X
73cDAvD37fjmB2FxOUyBoIuRyAlPZVD8C+iuJvGnRT2o4f3RLDSCrkNTx6PGWdqDeMPbs69SfyiW
XpPazNoQq3Og6wSQxEoq5bShZ6pIAQbvQb1bO3jj2JvTeEHY3+l0ooW9RqIrkZZJd0TyIsMAJnFv
MZPOq+IsYB72UPyVgqfWZmJbKdgC7hSt9sz+xb9f2FRkbB5iP/0TqROA/bszejgPRsX4EXGzUraT
tcX2IP0jRl6JvQX6ZmmT2f8r0OBmhppmjbVdLIQ6FHZI9pdwzcFM5bCqfSa6bQI4Ed7pf5PZIusi
5ByLkG5QtL/9LdS1lNj1MXsKGihXH8DmH2XoIh3Xr51/AzP5C1rxnnEYEbY54mPPFEqpvrRJINCR
fe7bM2a1QdKRgjL1WVXjnduXuVPs2DzU7Kcq4Bdbxws4cv6eTXxMk07gED6SJxRZ8TKg0tjwmc4f
yYLW1y5faOhPvNsuhiuHeB6nzdIfwE8WwY+5WedCsCKKmqzEPzxkyNdTzWpQ7asrrT46m/H3AMtw
O/m0HcTG3b4PbhjhMSOE/kzxmJiBMjNVcNzanGyHoZ/tTm2uyZuVuKzGUD5pY3hB3PpeuRrzNE8o
iRgflcW61EPo49hTclq2+PAupBL2rotKaW3mTzfiemV6rsSx89wZOzjjRwFvf6EB/m1ujlJB7dXx
Uyplesb8hw54F80RFL4qlH+8SveUNl9/yItZZAbA1E/9BTXOljPP2BkSuk71fgDWBAAFakLa/LB9
CILkrCnN1i1DgEqfN6ef8ckUj110q9mOFEJjotXModdIeChGg0cJiNf5437dYGX2E1ThRuiMkyQK
xr4JE0c5GqG95JUiokQ92j5jOAcZ+4tC/9LKTejrJlpzdBa6W2le0xFxRnrWYygzKGIpUhyDSakl
6syHkNMtwtflFAVbrX5hhnTgdXxAcoZJyI+f4gDQpNqlAnKYGjgMiMv4k+xJCL2vi+5fVthhbWI2
YKRcJdYRfk0qwlqVDNXu5ZDg1UCWgdeyEx//BlL6Pl9bnd2/7NoTyFTL88dWnDnQcrShUOCxYZLY
yc3mMotqZCtF+0xSqFZmiF9h+ohakiAqFHeRjEZB9VQmIWCwAuntt62E2XbQXZQV9+FMwHrEWssB
PzO43ZbGnlreXikxBuTzdpbRQvJxRjSwXLIzbz/Crwh/gmZpLxLGvbfIlVzSlwDgeqtdQ1KgPFWq
G35CO3u6VCu7Sw0Z4JeYC+VVXz72mQEo+cyRz7aFHAhY9O3q6S8lFnyzA6eRe9egEwl77o32mlT/
mr//2j6QHdGqzpT6quLnr1khfD8epOLsbg/qgQ3V0GK+FUO6g2tR30NrRz2d7y2+Mdq0f20m2Qli
q5oFQJySITvxi9zJAywMmW2E650XxgQxxyvHSTNyqeJS1Zult01yF8G6+iDOqqyKxOfJPUb501Il
HRNX0NXFmb8vOi3L4UVCWZY9YFNqXf3LJefE+YMVesuikiNUGOg0ZA8uLp0KxYbkFzzQTMkvhvVe
junK0RddXZ3MGv+xYNPtMq20UTxoShbvlF7GdoKoF4XK4OiR+oGNF1FPIP8P6db4XDk5OdFxKGwR
dv8n4Lc2940zFgQJyLSp+OgRJvUcj8j8vJAR7e877byPFSX6L+DGmi+3UpWkZXLD2IfzuEvdJJGS
63VTFmcU++BFmJWSd/3smC0OSEWkjqfkd4fzrFfyKDh37Y0zGfgsv8YDm/FJP2RrL2v5BZLfpq92
e3CO+FDiU0Q6AKsdq1x7yd9Xr9ebYyUAiz0CQ2nTGaZDhZFcS9MQr1ZTaLwiTzoCt4UwRizg4JrQ
oa5TSmrWml+ysmx/xgyGw+fdLWe3xMNe3Iec1Zh4JDs1XgrKW5eU5kf1rlS3562iPAbIvO1UwQbP
al47MA9YQAZaIBognBgEc+7L1zCYL2AQmCjckXj6UUdqBml7av8079Lk1WQ9wAObkqA6C0iPAgn6
UUKbVbAHM9dBvMVIpLxL1KQnbXDjxCtckvHlyMMNPUiBTdq+UOFPGC1b8k5oN2dRDgOycX6Bu/kY
CndJyMgPh78EnxJvliZUWa432H2sd+nH/yUuGp+yvsbv3P6o3w01HumAFYp+3yvVGTomj7djIOTh
3HH7A2/+iqu2ukLyJVHH2hxf94WJEdc4rDWYf1ZB1aJQD4mQAOKeokQv/dMcJikGwZuXnpWm+eMB
C5qZ1Ue3QlO6lLZbukIT+LAR5t0B4/cMlvOlnZvDOkaoJsRQLOxv1W2macO62xMngIktlxMH0tIv
FbBAJUuf53uy5JPt0TQF0TxE/Y1KQr+F3ySyHIx+/3672jm1VEDwRGtYyBqwNJK72E3PMwqWXR1U
OuRGs4pTVGme8PkeWjnj74R8UEAIlvz62AAGlnoceaYguIkfPiwuoBiB2J2zWlHx5/B3o2N4SLDh
pOmUu9GRCLR1D6ivu/cTJ0MSEjq4Wa8F9aLW4HgALQ8CGP5ea6Jo/2sk2KhDPY/4hcutb6XGB409
dzp7dEmQQbcplmiY/sgdMCkg793mmrbGoizRS1CU9/bitqnuJmaJIHfb/xlbePQZmR5SaAmxPd4+
O2EqVzofG54A2GZb1w1IcXTtjRoEhNbGk+i8QowymTAD/Ha9HLD760qXsovndJCvAkzJ9eAnlyZl
Y+suO/j9F3H65rEKVNBWH3EaWx+zbtVMsjrlkcDAD9jkjdwKpgBvrQjTkujGHFGP1jiSt+x5o+lN
gctJwvSQcbttIaHNLhBZ+TGzm7USJkRLXTGnnebb4obhgIyfdd4ojdyjKq07CVAsfRRP7AMOnxYH
VfQJF1qCJC42nSF5bvrniA+DQSeGq7ajOEK+v0yvX/jepDy3kQAbyphCeh3Dywa6tBg6ADDMNN9F
oBbWlB2rTgY8rS6+H9bAivjlkJYnbGpPlCyYH9yZgc7nqeSy7dLV8xRkABrZreu7zIYS7vvO5x0b
1Dqhn2ksiJvw6CcKOD5QSAfHaujlB3jA8PlWRNNlobbQIjDaEyj91sSuXhHw2wpA9tJAVxJ6jUZF
iLi+4PYYduWolKj3idKgdsTMwz86USzVeVgjT1udozVB6mmDqJKhA5RR0wk2H0Tbor99YEEmVLQx
H4O0bntxX88qBHp8c+6Zysf6pfGv+qGYoEppbTOBGVGDzTCsH/eu1iyvcwaXP1oMzUJihPz6C1cc
ym0VyOZWIyfvuUxji6Wov4JI0xJ3RGF89L5AynSuKkMYcma6y73uBgMPd4Ty9GBc3XT1iP6nTzUx
5qeuXXcZoFWE8hytj9USyMlok0BcJ7yepA8S4Q1iB7FzWxqu11UROzHOPIdpTfBKscyRaTXXBLi8
2+3vT2ENgTWDKq/czp0JVdPWZocSPAydALrJOidLs0no82pDRRUU1SuySrVraQ1gD7+XDESAOK8b
OrC946ochEm/Y134rBXqg1ET/ExKLjr/i6xsREuzC5SYqfUi6Fq6bqekSfyINzdYsH2sKZZkZX+y
W7PG/ohM6rXmOH+uESdfK30cHCdqZTT4JcpiBkzs8syIc57uq6DRvcxGhYq2qWyJ7gDu/+qeWXlo
GWDBc3iWf6SwmXG/v9+Uub2lPbNPzXXr3CC2zy4tBUjzUQOkY9Wbzjl4gVMbWYNAzcbuV0JcRUAx
noW73yZ4bAeOaeWeyAsvL9gS/JB8w0CCQkpytZgaFrKHLQYMU99QF+hGp+AyO/2TcQ4dQlVh0Ra4
dtJCS11NdZ5jIKJ2a5F4IwBgO/E1OUYAocfUGhvsSCbuaO/aPDxEfhYNtJuEfRvLRCfI38EGqukM
fhSYsClZxqNqzvKk3U1GFcmazwgxfW0JhCeggMarUAywBkuG7g/ZkCE7C3x/FNeIUW2pjB4smJyS
+3dCunh/hO3bzyMeq60iCXXLICHYLX8C9NHvT3IoOZQUZ12t3zYidqTy8uOjfUoLczuqzxbmLJry
bii6BGyas3u3PAbY+Mj9+rtyR6k7cfYnWBQL00AGlzQhm1rZ7+Wg1s9KIB6OCzMrtSrVKUizQ7CW
jeMP8OmVpXgd/oa3HCVj32XuyjRai3xoHpBYc7CT5YzFkaP2SgyocCN5coOEm7XbikVZHUD+SoLC
3504J0sGzrUfcfK50Bda7C6GT/p11G4Kcic1PQGHJRf3skjAuBicmKZIEnzofIaBOdh0JmsjW/Vj
vVP8JK0asVJKrT2OoVtneOI96S+RRMNvC79BnpzwnDAdwXF9Q+fVXK5VMfBBxbyHxVdL60p7DuUH
KVld3rTFLrRFEKXQ8vu4stEbjJzjnGKYEAmiDk5pviQOTbPFk2IJmAK2n3xy6AdKYKJOK7INoFxv
X+uolyLfFAtdpgdPHMwrCWdhwmgVSdHyODk0OtK4CjwfV6yJaLbgLFzxDghPA/SSWR7lbvpo/88v
39BsH4+l7v/aJjaO4uPl24zHpheaRMcJemHN06ddzYnXIOy4otjJEEuG8d24zR52sNVNP51aXndj
Q01kMzo79xel5Kao5iK0la+XAlVZ8MqbIxIqz3pjTRGqBfhr5nDkeziRgjYJFx88QbmR8oZlEBFP
3nVhz2SxK8B+2NxZm7i5Nj6/VS7TtX+R8quWMczVcfb9Nki3Q3vYO9RpH/efzD/Y2pxaEj1q8Dw9
vBzq8t9eWtwwogZrN+H2WiKQUv8B7CrnBTR6YDDM6815VvxS7r6K/Dtnt175XVe1MmKEKMShMtDb
PPNf/faHXKXGTHXV7udboo9w7YmCuB5lNG051A99TUhcoG8InrCH0PT5jLbGfSpW3D4SLfltgTsJ
Uoq7eG+alwR9SxpB9rUOu1gOshjztVYqiYAQIs1UMolgivAPYUcIeut5PWfyxpQda/3rzuDCMPKt
Paj6Dk9ujerDzPBmbQHa+XspI2hjgG8Pe9j/f3zazeeB5CwK2od+Uf7meqs72VzQes5Odgayfd/u
TxZUW3tcKwu8O79osThQLlHK09DiMkgcdnAepYjCXHtIf3c1fh0esGzEAGaNw/yMtXd5RufPQHko
IpZ5Y7JkCSyqfeplvffQ5yjK6QV82KWreIICQTPYQYXwJ5L+MCi2ZWX1sprTcgc+pTLtWTSO1cXv
4CNuqPp+xue6v/CsEQGBUPm4+zn+tG3URNNBWMh7IanuoKB+R7f8KPzz0oey/tcrFWyScbA/1+JO
/5w+g0miA00SeA6loA5W5U1MYCwzMn7mOLfvnhiRT/uajliFjnPiZ551aoUl9cbKbZAutGM/BbzA
S9UaJ6Qjh3RejhOJ4KXmZAbc5btGsvaq6yvFTZ6CAlZcO6uGRGntWwHhAu7mSbsMl3Wt8jd1Vwic
kDN0bsfBoAKN5iKz556i2cqNQcnzRr/q32jfkS91A+WTRXQ8vkJh2qXHK9eV9qjByKYdDJQjS8fs
I3MQGD9OpWayrrcDj+gq4JRIMJPWMtYUInkmTbEtjEpb8rmIR75FdUNb6QGAAN9HJD1z1C4B2lyf
rWFrc/wGRtHOs5/hwsbfSTeidHN0qPkNFuA0jnlaMLkBh90KEM+uJ6+LdFO6m5fXrJ2hpL71EPnD
fWdf9ss+DmsNcRVjAfl3hoXBgFJX8OUfJRGFriFW5pTWn4NasmmzQagWXFzVyW5Du5hdUTEdR1vu
Wes0+uYsoHmOwqUUCWTbLEvSwSq5etEfBYAREV22FmvEGA8T7qKmuiZlqXvVSYP7C3YflFiSBc0u
zhgqAzMlfXiAOl+vmlseE1kz+BEVPU2MupqUAwTVIHp2ygb8TOle3OxPYwxrqimrNJtC4zT/cKzE
NIhRbhz3+0ygXps+atCY79B+c8+sbH+OvowmbUcwi+3AfjTexIBSbeLygGdGRDy51YPzyYwbmmp9
/AbfENCm0iLZvV3bZmnmUwiLp7FexgEoasLqloKxdCUhNKTLs2rDbTqIzOuBQdgOhTyPxkmqfik8
JdSnuOFfuE7JXHesARLbWuMgLOFz8DQcRJXVIOjxV8pR2EKVJ8SXBRdcWr2uDze4oHGZnbgYpDNv
r9jaYjhh1JiE8fqKbCiFGAG051dMutyUmbfwCGa9eEhzoM6UH4nsD5dbUIt/2zCX5JXRcnLBBtvp
tASX/Yd6UubDp0vNBCtJb+vaqC+AtHSdjZIjlepbaAoM9ZaRE2VM53otAu2nZ5QGl5bAbkZLd0F/
AkvIXVb++C/gUAFOQTjE0gKulf+jecwEefw1TbMHvG31+vgbFUDu7lqKauVeDplssAq/pMB5Lnoc
bi9COdZOGRLHqvBxLq0FWh38uO3/Ji/lqKTTX3K0H15fkxnla+EklF24m2Hlz2MsmBsbluVbWn/f
jfcQ557FkdwVTuaBqZeXcv+FJrITuQXuHRDgqHaQh5YMH/CYAxCk1BsxX2lmuAdHhkI9i5SoqgQu
RY18kN8EdQVUtsp8hO2HcuuSGYBsXrS35U06n4FKuFlp2Me9sJM1Pb6iC/CBY5D0l3oTgCl/F5AZ
5zhDtaJlL9n2GAko/boPyWJDqSkbV7eBtRHI+QVzLzPNn8AKBl35bv9j+SUWyhpsgjTZO7xBroh7
MTlqYjxfi9Avv3nDBe5rfCV88h1ue7HbUCLlzNzgwNxJfdzHJSpxRnjNHuueWoZ1vggfZANkp0gO
6CAjzGBVEJ4QfR25QzVeEnsPAOQWs/DNMOi99Li1+xfAgdxcn1nha1apaidkg0RzRbRg6ErYqY5P
Qt2YralnAC2j2nQTggjKHnWAweMSncfK4E4u+TLKs0Ce8Yt01D2fbfz5tJGFWNbBS5m88ONxw2pL
OOr5FUTaiL00IU0fvKBLQLbH9+4onCLdkHgpMhQCb71AaryXah4LRisAtkaroHAiYgPNMwId5B+u
0mNKlBrLAaRA/yiho3k93T5ywIFIKRv3ir4jfJPcs4RnrMtjshsTDNf0+S+x/UtbPVTvgtGggky0
r5nVNdOCAbOzz5mXcaE6dDRCqO5+QqIXlj0cs0MsKYKVjVhwMgGFmp8h6tPjGpmftu1Wv5Kgck2D
REiRYPMP7KBscAvaubN57neXc+D/v1pu+8I8f2GCFGaOf/qcG2L3FW8uQEevBUfd/FrrKllLEcP1
Wu1d2kuFAkQsZfB9/yRUEu5O91nlw03RD+A4yxizXJkJSrqwspXKc365PBpVeBwk0vO56W/IUZlI
nbV4JfJeeSbxdR3F1c0/SMHzS/zzO2Ld2B9gWeP61qiu38E6mKKTtKZGgZDBnnWlM0XOLvq95aKG
GIQWlNmjgXVle5b1qNNbiH0USKI6/hQbVDT0LUL+8MNowFTpSpNC57cFW4dHAWnBN8xTEwtrFjBd
+UlVBXBg2SeayVQ+vI22FUUijUgJA/aaQ09uFc5vWfVrzrnP7TFu3ESzQARhluOL4LnyRSm2zwNn
VR5C5HQamG6VtikRthxPgcDNw5zhOGGwA+oeLMGY2Yt9fFyPcQDSJ8dRxSt1k+Y8tI557FszEd1z
rVfwQilzHTgJok2VkDvV0GBBr4m3TE8Xd38N9ymIaQoULhembHayRZFGEC+KIPJiuhtCyon+yiEh
/Ki1p881bt2jRq5HCRJeV1CeEu5y+1tw1IZ34dfQthMAuxMyF76IEV6quBrx4d+Is214F8rzf7Bp
vq1YRYmusskcEEUa9VQGzZdaLeJwu9LtM6RFjiWrU21hHKwBcU8aZ3lvPo9jQi8MAr7xrD9hWpmT
ANNyuvO4p+Ap1mqs1FZ5tK2BbVEx81kjNtldFq/QKd9P5NFxhlaMVeK4dTRZdIVir22nuzYrgpE/
hb9F4KutsdgxW1yfjAtFKlootlgxP6b6aDwZfK4KOW8jK++Lw/awZLddgq9Hc3LzDU/OdAnLxwAH
qV3FOVLlJdvCUfWxxyhoXZf7f7TqIn1uBghvkIePo/mMAyaXTr7whJsLTuOxgB31UAmU0Tdt2aO3
OB7XGoj7CpYVdHo8VLY3vbUg//OJ6ibg43rZYvnW0+CGJKDlaZKUfuprT1OaYIYd4wCpjUCsGhRY
z+I3QLkqgVgLUOuNKez9Lg1Zbr3oS/15uHgLDxhmI2jK7ivgya352s54idXr32LXEuGAQDUXpHeQ
K+vklE2o/6cyMWjpmC7K8pFOmZ9EW9K0/NxPjAYNIKnGZVVmlt9GCPpCuQ3H2Ev6aBr+KJpUcEkJ
e5O5EgRB0o3f0Nq+67JvZD3Hy7pwFxZlLwixA4kCT6bGzpXUZ78omMfQAklaiL7mL7gAj2LzSaBH
N1MuW8JgBadJPXTsOZGLZemgI96zkSNukUgNqbECN/JG6m+9P5S6HmNEib+0JULx1VnGbDC4hGHi
2CAvhY+9IKWMcawh6HcWmhWXWsT7nd1/6hgXss77PyjCSYfCSfswaIJRtXEkvIarL71UENhFAX3d
6Ly2gfOs8P5crw+MCT7a/gPXHdZvm9XPlw/rW1LYXdQJGRskergOS/JMKYsAWUkSoXBGb/4JP1BD
ABQuIewTcIun2TFW2w/qTBpYcz5Wk14+LArrdUORPMshsU194IuobmE84ayJ4DP/LVVqmsVj3OgT
NY1nm2LXPyHrMjSbEg5YYlBy7J7VRvgyxt/No70xlah18oSAv1mk3Eiwe0dUuEAfhkz37AbcLX+B
QiUcmwRvIfa3AceHB+5P82t5S65c1iZ2zYD8Xt851P/ZomM1/DVTEJhvkQzv7HJsUP0y78wOb9OH
ZfajfhabVqiwlJ0qxQXinWI2HzzbPmCh6XuSk8HR3Ih4oiJmqfmllmCkoOarSxfVkRTu9PFqoPkf
fnLEzZ56rYSXEKf9cQ1CCCmSuNLKXkfzN3Npf/U4zqQSXs5jDX6ZbLGDPzreQMi3110ukul8Icur
a51i5SeQacUPISMXxFWVOzVMy+TKNvb0xrNTbionlsLDi+6qUfKZAWPlS93vGUG/jLgR1kdg7+AZ
SKbjZ4ZLB3fUNrNS+1USIUg94oKiDPUTNGraOAnKTxfu3zUG3O+S7eJjduyTjRQX3/fZKPYzL36r
LEKfNygaBlSHEhuAf7hUJLyvtPNU4DtTdh5dDkJmmZjYUDSX73dm2AzI9snaWeitkoOaDlQ2cYXh
HySBkl0I9/wbBPX5vhV4Eq8M06HVIWtQ0zb+JYx7qnxFnnUiit6zpZJn90HHbqdhyA9n0JGko1Sc
LVww9nCTOaD+f23LAXFHEebg2/26Xx0akCqXvhCRl9Do4FEZnzp2KRZvR7b9Sm5pZv18EkJyB4jp
YQDr5OkA/5pSHjRMJjFxGCRIugqpmooP7T27fwPH19At71yI9DTr+iGDDzQ6Qm/AumAZYfjzC7ji
Fn6gxAVu4izD9Giva4gbmP635CYoMVeFFLoSyPMpYuF0Uhrl50esSr886ao8KbO+fvdCfaE8/7uP
WO6hElCdCtuMMF4VAvg/1reu0MGWuFvBWDG9gNThpfFaN6D3drujbXdpiiHzr/D3r1gIytb3VhQW
8Mn/C1LixeVFzLbaIok4RaA/eG20o7kR8SaaX79DPRV3ycMGJybffrx5Est8MYi852Bbhv4g6vlj
bq8biQSwi8skAJx/f0LFmmDIdmP/sNqc0s/Y1YLNPBvoX5DVgJP4KeJ6X3zQsnGRB2xl4XvVaZ+F
L5zhafZNnuEsJVXbnafRHI7ZOAnytaR+dJsehqyBz0vBeohJUncFeuL7OSK6HfU7arZTY83rBbfg
MvE/O8yNQQ7c24QIrpy3onA91esl9bsLJUDYrOIzC9iUsYuuRiC8zdIIOffaN6L9AMem+nbVKq+F
nEuLmXUpvLbVE+TWyVYuwv/uuBiilL+Sqxur1dICUiezEwKIctLhp1fCMmteW3RbaNfzT41qILOL
+VajLw0o15Q5yF9rqQI3dqJq5pTwyusOqF47XfrF4BJZV69OAF9pBFCKuY03N+rYBQD4vddhlQPq
WssV4rh3bZQG4s5e+KZwtw4a0dVQUL68iui/KvT3rpSA0n2h9LgLGi3pvpGSkrEB+cx5vinyGln5
WkUnpac0HTQvJfC3ixPDI5EFBJzrz5yIKRNAyZDshytCr3Tq/hPKiPgVYyL/19vtzrttEOSIO3re
bzoeby3i0mjgGhWuO0yCEmeCv6FKlpPC/xwASN3JNb4WOZdjMCaIXa/hSRbWoyFWz2o3kWdhotvS
ldOnVHlNjTkuE2ChYT0mSXe2p4ReD3cFASgZyg4nmKGRuMVqvNQupUuXwSZuw+z0ztuZv/7qWRkf
/b8InmA7TA31bThOwXsiRfLgMClR7uOMuvBzY0CDRImVYtsPLXaYBO+r0YBmEsM7FEOpTJj5J7Nq
KVZXF9yEIIr2ZpbYyaLAp8ux49Ta8lBHi1HFsxCbAuTZ7HpyKy2SvaMvnsRiW9RcWhr5KmboCRWi
qfCF/TeoXO3EyrPa9ZeRLVbXNbE52ZPn8zMzBjIzalpXX5cTGsXcO4ROiqIc4nd6X/9Ms24uqVrD
RG7R/7TJJlND2EPZhHQRkv+j7UJMTXLND+RZjBXThY8kdeq5u1YFEbBBVkmdkmBVv8T/XxqWhmT8
uyie8YnB5/HoVyQCfm22BBEe3mmiOxcV+Fe8pPDMhKEj8eBeoq8swIqDz6+6WOZn9FKydQneyxp8
QAvwwciwvQVBqgsKlLGaLWRb31n7EN2DQr6qv3s/L3skC7XBSyU2FW3uJJnFMa7EawCsgca+mrz4
TkMtfqOZkhA/wzlUEg7KqGHzKz7l5G5xuOxrhqwhFOizQy6kYVoLpNYJFJOct+ec58xRoMeHDvnA
wEuem+IjmwuJWeO6QLWNN5NKch74PZftibx66/i7PLhN82TEY9MxIM1SCX660C4Bl5ZP/+++xIV5
eySrGgLryOmpNrMnwjESaygDPQOo4ZgyG+c++e0FY8Do1f+q6vBn3AgaISQAX+US4YR6Ym+lF2s5
qXtioWRvwDX91mz5QiUvHb06o6zX9apN1UxAWY8vCAsoeaYYT0lC+40tthdE5vQz8Equ07bGbhow
l8V63W0kjkjyu0y38Eqa3V8CmsnEVimTjCYuB9Fy988GKhVGynftapl7t49RBirjg21l+iyJ8U7/
Yd5vkN4NSWoLhbwwbmXZbdir3K4R3RFJYuNBs7C/V3cJ0hBDKqCdiCc/uxBRpjarchGWYBZqAZtR
gbtbUn6DOq594O49+xLlYZPLcihAEhpRgUvJ1hgme+KxcVdC0E4DdKQ9qy9aQlFwW3tbyk7zKyCT
AeViHmMZqDQU0WKXPmplyuiubFAYMyy5wPKrhCh7lSmJBO5dHJS+F21hWhgcW8ZxgF9Nhtuzrg3/
tZOHwfsUWSDhOUmi3lCB0e1y8Tupvmlj9FLwX0zw3gEM18omux7Cl0ji2hquwDOkWZ2K1rzdHQ83
sJSOlx9sSozUeNsqJ3qz+svE/uHjT2ImS81S+zcAuEFtidVNND10FOy+ugUxNyy8NMW+f5IjUL0J
4IlTWLhTFucwva/BqZj2lvHfbzs+X95D+pFaxvD9xn+VIg/buWd5lPfpoxQul7Vu/uGDNdpeI/6X
Yb0mXP+W8BE+fLItbWZeVeZmLJ0hA/UvzAVCoBikzaGrE6noYJ5+KMlJCci5cZDYjc5ImIwYC37I
EykXSe6KOXXCszEye8wQI2oB0f+ekDFz9FF3zU8FnxdT+Ut9c5OR5tBkoNNwPAJ2H/gnGnPeMLUo
KWYJQERS2ZBRzrzo2r+eeJmVHIcjsxUdvd5Lv4u5ILdzZLNyRHsYalCbJaK6XL9F/wAx0Kk28UWb
Vg/e/jE0F9ghC8Udn969ARVQ0uWFdGiL/TGzB7OMSR3binfuAvUnJl7TheyXV4ARmBQtIwjgPEH9
bAYErTUfeS8foxNsXucbxFdhycCGJKLg9xEX8bixxrlQuyAL7ewIdUmS+ncxYQ4OzyInJmXaGpzI
zfRewOp6g7d1ncG/JDI+pWqlf4PJRvtoPv2f7vmaoANQySZr1hD8a/Vq8gthClT9hOs4Z7VIGpSY
tnLQ494jKEPccrvYXtMkpCOTHsx3Htrw/vHGvWiAAg1c5uYz8nmjs4jcd8SzmQ755JSelA+RlYut
+rZLIO6SYOVaNf+FAIndh+rlCA7X7seznVtsWKavBx41njjQsRWyAU6yhuqOsYvV9TKTIOwWc1IR
+dbjaD6Pc1a0cjoz5XK+aXOIKV6xJziAcXiupi/o+oOSjOQUX5XSt7SegRGDf1gcLu4/j78KC8Jj
dqIzOR+RnJjMBdZNAG3wG03zNeX2vhSgLeKBgh9v0POB8H8Vokun+piHzdaO2U8x+3bZ7K7grBFI
Q9xzg9cP9GGRHlvkWB7V3Q/lBFrgBni1pnyhQuzuPn9snI3qiT+9O5y9re3n7PP9MD9PEJKqNRhh
j+7T1r92N9i82vvPLKM6tPNvwonN3EjDBJ1h3g5z13lGhYmmOD494zyBgbS++GVNDFyKhD4lYpdA
QumhwZcMavos8P7iWZQTAAeUnlZfixK2Qygz0eBk+ct0/Y1G3LogIweiAu22A2gb+QhkOevCW3fH
1sXn41iO1jFkXGj3WGqNozC8Ss57Vnn3H3cJ+b9WtXvRNDVP8Z4p+emzy7epDWZFJZbxSC0fse8v
emkISN+sfARwSwYOEVc9wnm6S0VUem4NY9I82l6laTSLd492SAwOKVT6YmgkT2S8BU44ILtWpkU5
R08rdYkVK2NgrBRbuI+upTpJL+dU1aCevUJrPn9Byf4U12hkSghCbHialTcgL5oz6vEjbFLRDfLo
PjZ0dEV5/3qKb+5hyxQD0doaTp/ZuRm5IRSbM/3kTJbIN/6ZtwJuyV8uQ1AmUx8TTBjjVPxnuXNP
Gjpv3Awl6LBAMm66ixKh05k7ttqKzuf/LDiRkIEMg4c9VrY6k/Tyf6LCcHwl+0KtTDp9LR+41v8B
fHhoNxfmB8re5a9s5R/YYE1Q+2HyJejeZVH6BGBB2C3omXCH0DekrSJ5eUxsfP2lL3KYUgjflbY3
wyxiK6jlWrp71AJ07ukxAs5jeFhNRpJQLc0Xcngz4G4Z/Eb4aqrLuDeJWvj+tOYlT3BQKtLYIfln
0MjblMfDYPvoBqbzF1+VjvfbYG4wmfUUIDARkw6vAsS2poljL034K/Do06q2MnTZbL3dg9CAiTKq
Waa48rGrrzswbvpy5KkbfC+9tIHl59TjRWvLR8BtAdRb3wV40X1JH46NEryN7uYyVsa/7vARJOMt
+0oOhanGu/TJcxndTKBYTYo6DkaPPNNKEGs1khfTsMbWabrn5b2vbAl4gbLxgMiKNLMrz2UuMtBv
lbJTT+Ew4IUQ3Gml6yM+XwHc0qz80sYeTh68+WfDwKxvMd7JUurBW4k4NNbyrDG2E3mnNhFKRZD0
OoCUMninwv5W7FT9UHAfwRFBJVtdQo5j0L+TKDJTWAlG1j38i4T0MEM5d5p+VW43qzT3SwMxR6YF
W1ht1VOHJmxrXHOYrzcq51De4HrPwjxhSXW4jPvSNxhfv1MMLjg93G0ltNpT69xQ4qeEKSmHIufc
ZECd6VWNeZVZy+wVA1Pemdsg0C1C+bkSXBUIDS4B4Xpp7Eeu6hUEm1kMZZ17bPEfahS35hKtNxws
YkMX2yQ59K5LGPO7CLzTg8M3rvngby+IQysYyWESZVvx7hJ9wt5LB3HDRSXjZEdM62wc5WydD0AE
CbJ/cX5DS3J3d5iLRE4+e+QfWgZhlIdREi84J6AAxsubrgUWef1Jx/lwrwVRzs1BiMke4UsYLDVa
MwHkry7vHx6/TkrqbN6q2iiVo7i5Eze40xGXOOHcjow1mkHMF5hnsQKmNAGNxTXZsbuI6iXJ0AU6
2Cbu6AMW34p5J1+cepTOIeIgcJQIrz+AQw/DmW/qfH0LIDbaPEKbjYjlHwUyrZPEAZKBSSLSxG3D
XrPCppMrIqXkOo1joYFbpLDVtARbDQKN5dgPFkRNXf5HvdezdkvK2HNCyt3OsjEAd0QM4ZAW9ybx
NRx3hMzJ4VuDfa50roWYGK22fkXNFvaf3GlcgXXY4z845UFjs8Bb7xvCEFjtKwy/bU0DytfLS5dH
095OVuzWYPWVYmF9BFUWSNomSZY4SV37pOSqyoKd8ZtnNKG5JAR8Q852pijX0gM2iwMn3WL8jjqo
UXw3GvGrZ5LTn/4zxW4aDqHWIiUXHVzHeKiaMSGq0e/sqXLHSD5Gd983Zdi+Xv5eQHKss7FivVL4
/LyydAjFuKCkR3mGuFYIAarWGMY9//t5DxLlIW8r+wCQNmhSjETkInikjsdm+Ihfy7FbQstEb88W
1OxigrcGM+bPSE7a0PFdgjj3kuvHoINwI7yhFpWStjaLyKtNbwfuCOG5+9uvhbMQ5apQKHUW07f+
ozM2VnhPBUuJkFCi/brvOSQyNrV42v5Z8AmpShAHgYeX4Jul/jXDr0mkaQfLWlGzQ07La44ciMU0
e6nZ0ZCInQzTIhOHaG6bxOn8cUBqKjlKa5UUg7Yx+czAQk3TtKKOhT4R1XtskFqrwXz/tqQWua0A
div2jlET7wezfKFXH5muODMuiD1purgFtk5h47fRlpvEcFoP20CMbw+JKGVWQVBFxahifY5tlZg3
3HMzG7TOGy4sE5a3rncQ8hxhoVXR7XX2vkCOavTBCUw7irRgOrgTCo/x0y8Ix+FGJmWsg9qwyFpv
hmDHm5L5K6s504Z3ygwrKR2yKR/IWuJ/AivP7g1Zx7D/7sg9XHJb5bRTUeZzRPCJpdS89exuOQ3G
/uq1jjA56HHQP1y55CT3q5MjFX5kftGhNqHjrdXIS5ui+ZOhOhHCnJPlEhNki3aMwMq/4JYEqGls
h2PLxZd/8xkDGTtAXqQlER/T5U+MSBofEMpdHovLv+4TkZaIjTSmb916wjbUv1mBQaIea/VEA8f+
gMGX80nDZnbzzaXwHWdNrpwW0/kMmlWROOaEFohRylQU6CwZicVHkh4+az40ZaUZeaikVGVlceQ7
d5nEgQwMOtLlI3qCLSVzCJPiMhR1csus7+z/CyQWW2YggMNVgq9Gdz63ExyOIDsZ3cCw17kl8C3K
APb1CG/PtUCQwOP0w+QM71kqwmWo0/vJnFFfggZzCOt4XOLnSpP5cBtgxNkt59fBdlj8SHecF+qm
HzvRAjJz9lie2tPehbBxVbN885Hrd2oP6BlEaROXIOxoc/ZEeEtPer19+RP6fV8iCsgkWuOjqiUU
5RfoYrIJarqJ5YmdJS2nDOhPU+54FvlvNeTGd21sGsoNbT7N6DGz0zuydglAOMgI0i6Ie5gjWj7H
t4TRn8YMFgoFcPseHV/t+YY1leo46RMFC9J03cG78I4jVIYvyKfuj/9V92gQCmXeOdJO+plU069F
IZeDuMpdpfsHywQ0Hesc+F7pOE4oPBJQ4nYqCe7LeO+vX79TEiD/R34TKKrL7qLGfqmzi+6x8jg7
ircVj8W4rorU9jodWARrrROgbbMKhxRReQ11S3p1SQge9X2ExEMquWcMkgboghdJc2sTjv3LAy/q
rgDNPlQezHF2kwoSrYeeGCxYEwhZCuaqYYKSdU2cR2KAUvqjO+Qgg0jGNyrtwDUSH77CbjAy5F2w
DEHxuoX2fpm5dbQ+kisQOmTL9q8g0k6d5cgZKYwWjikuNdY8AxwAY+BPzUnqTftjLUxn5JDgQnTO
y/udvnQE/TL+R24VpAEejLv4WazYRp6d9CBNif64RDdCULzgXXfS8opfV+7fFj2bO2kILE6mYahy
BUSbdyJ831oIhslZfDGqWmQQMpzWB8OxQm9GgMfc6rQJ21mGFCGSTxTYK4VF7hjZ/Vln5D+VYD3m
IgOKVIQiyEKzDIseL8RvMrlQW9egYfz2iIZrK2AhCbW+jof1TyOKmyYlY/ylJTf5pGQLzW3sSIt8
AwiyczekmXrP2EyzHEuc8WquM+uoJueAhKGsjaX2aUBX1gdGxRsnzD/pDauf080KXrSfgDM3cRec
pVAS/PRSpua6mNxQJv5NsWHXpBY1aOwlPVCzKuq5/zbxqKEiAjq+jCSUNI9HElMIQ8Q1DJWxMqBE
TnsJW/RsEeUy3r0+ESAIZei305GCWNWLlb/5ZJl9PJmpSmRxATA1D4e8NekqBIiqOqqQGqsNQ0kl
1cDSaBst/Gj9nzqg3wsmOZZk+hD8YiyO7Ph6o4kO+aGucLkMCj79UX3rwXOwQuMdkhXwM3ZaHQ0K
+267Po1iD7nxSsBSuFBQPku/HBPhqM8omMyxiw0/i2pU1/cW//AFWmspsM9Cssbs2wFiHO5aT8ia
mGxUUi6/5G+QzYmn7qHJU3L6B6GRKd0DEs6HxHvo4VWFUSkiUOpYJQfi5ydVfFH0gBMELvaNyBnP
XLk5/45A2kz37kimBJnOy4cTXvSSKr/unLcb86Qbm8KRO4nlEA42X/ATAS4aVfONgXrib+q9muIC
xXR0wrsPGhtwZDUcIJZMY0espz84eVDSbnG9xM+Db3tieh9C5Gpq4bnLwnnZvQ4ZhWH/mImJzuKZ
P2aFVKmxKt0hjbVpGpGu/JZD/LXcgym/bBgaiYToSIzOGa4MwErjCXeTv0K5dRPevy0yWHScBEIy
bYYpGKfTPaN3qKgXoDpU0zVhiverU94OLMOFowOIFc829Z3MlgbxDfaLhidQiqX5IVgXjfGcbz6n
xbWXwzDej6ga94+9VErVqp6BWEcBEUCNvllTiRnnjw9EMxUbVNMDeC3CAPMMVOCHtzFzxg5SmWNE
+/Cbi6C7MkqGUwvoWPtVJ9zxidc6ZwOSHEZP1rPOaTcvN2vA9ItQK7BmCmL3iU3F3zjrWAP9q0+a
GUsGKCVAmDaTGpOPNnFump0Ysp71+VAtsLHe8QOdw6rcwFREx4f8a+3Yr/2np5xKvr7MFm6cR0lB
gcqZFF4iBYbvDAPGjIY7x3C/tAnOMpEzP4a8nu6bm2tYCvrMdR0XQLtk8NHXllWxntrbw+9KFWjP
G3I8tnnajSgm/wytY7OCCI742/e3RvfYivfjCjE2z7vOYCmKnShLID9G9Y3la6sVXvfsMT+1iaXW
JpYH4LRhIDoqgNmcorI/es1RZ48Jvz+6NNRHv12gHM53ftHZqVkhdeI2J8ElUPghCTjlEvSL2fEt
qzxaLmelIOeFSxN4xWE11ScsQPd1k0tM3alzE8TIbtGs4J2CeW1UotBBCSN8KOMJekwlba20f2GT
MfX/RT5ada+ZEDvX4zNXC9lan2+b2J9xiGcTHp4OzA3mAl829cGxszB9VoHjI1P0/YC6JUiKxd5n
xfisub+tB+kiAu1ikjXjfCczWxOjRHv0dM+8SnyHOoSL0Th1ZZNCgCUNCMJ/G68qs7ZcnM66XzFD
3ARNkOmgfQEmUepdrFXG6HB6TydQ/GRnS+MJ9lOFWF0AsZSvGQHlh3xEkDUzOaxHxHpCv6PKBKbk
5OHjhogdSydMd1ca34ausjVbPZJbvErHCpBf7FzZ/4vs4zPl+fRwP4WRP/HMvDLOIQvIItUg0jXy
cftym9vJ2B6RhKrPqkK+FUWQOAls0KjhH64Hpv7Os8r5sXZCvW6jY5KZ9jEkVWbC8CHZac3PDB4D
7CTnik35UHvuVeJ+pV+H/1/Pre1V7SUE8wVO+HPWgKZtzYEJXKalDxk6Z3O1R4gEhrysNlFJpk3W
5Tl3dti926yfW9A0o6Og+txuYrsxjvGhOlxFNHGhvEtPsxCuHY0VuKdKf/Ze7syKC6klOdcN/mKH
AsBeGHhiy/cARwSf71gy8ut4ov2QMExmsLjSRCsICSRJNXTZ0F8DzI1k7UxubB6xo2eAxoXqTD/F
w77QrMs79dTrDLT2w5vlRrAH6sTk1t5WawsZO/so/pEi2ZrWjjasaurcEzXhjp+0mEKAaKS5HWXu
Uc2L5M6Q/sGLl6XS6DL/3IFxlvDwnPc08hqXNIudZWihWdz2bqcxu1vM6ay6AggFTiY7aXvPie5G
T9y3UAS1NRddBlzjd16hxyHsuq2Ff+XwD4942q0hSA0LXW5+52aiENBs4sEHPwUEOki6mHBO0gl6
dIWJb7/ffsaG/yRCLWe7b8U41q3MgfbjnMBaZnbYpAlh5RET4YlLUxKEQE9OThhm+ELjd+664rxm
4JGJL2AuK78FJlfL9kKEip7jXSsJLlR8f9oAS+wMLRc6dYfqm7rlaQXevST/DezvTeKm/LQ+reIc
n8l1pb7nwX4WX3+NZeXS0j4p74/41qcWL2RhhZXzOqyIww52fTQPRMzi+YkgL1eblZ8TbvwS8Hnb
H8lygIZq1E9cx1k8rsDdPuI9o5HZ6xX2Vl+FUW0tw9eggtth3s0fst2oHVbaUWr1dm8Hy64s7p17
vZpbP8CyHPMg7dvXG4MQWNT6+D+kAu4/aviKTM08NOXmhYowm+ScxRhQpMJTr9Lka9j9hxIp+nQs
bcYOZEn0KKQb/h+KtGKER3I2mCuLI8jTmNNY48Tk4zYJUYTa8x/NZBlpmSTPKAtQ49aRC0PFm4iW
kh9SxFeSOlmmYfnwSV6mAAVZvtMDvdAy8MD4qL3hEbBEOjxOdy8fzoZD6Q730/UuGvBCGrVG8iTU
ze+JL2YpXx+6F7Me88aEHo3Ftn2LNnf27pTmecptaEJmG6AV4Ttb+2PFRMuVz96ndA/z6eu02dLi
URhkJ2u5bdaqd0pfiEHh6qDCf3y3a6IogfHqmE4ZWA9IKz1/+h6JcwSHkt98xS6W2vHHdy4bsW4e
sSocVvT/dC6rFuu6vb5dUYBztj+W4pIEAFT+licRK2aNzyv66hlP+6flonT2VLY/QVj8HRj2Cu1f
poEanIu7EusTbViSUttARKwMFj+f/z6jzBm43hVU5xes/wWK44AU4D5FqLmUdqZw7amlM69t0WoV
k5NCkyN6+KRZhYUi1oJ/sEi5X8xnevLBF0nGGMbyHrmT8fvkiaveZyCMFHJXDKG1L4vO9DxaOOSc
hGyRBKxAOwEI8PYLqaVdGU6ShIwFvEMiOUKoVihHrovV0BHy4A2aJ4EmDWzDQHmrb65XzTaiAlNr
eZDJe8Yq4w2txp7DmAcwqs8+XkLfJ3gDFW1mauWTLpgoiN/hsNam0L4HQsRGFCowQlxaXiVrc80y
Sfdw0iwHYochQ4aXpGREVL1vPujLaSX7e7ahabkbMMDN48zWXx+BGj1tx4jfvNw7WdYSADQebXP8
bXhMBE6huPVvu3OU+T6iLQI2jjDM92oJrFf5956DgcgKHLa5pk2HOLHRHVXkHLh+KM3QbofJrEeG
bIiGJSXLYmIZTPv84ui3bBOAhxV39elqMOe9iWrcEwfkEWZi98ietkhlr01k2XxMTpt4UF/YnhNb
0RkZbQvCVubxYjeyFUi3E4kpPDJnKIujQhkzxJz3SboN/RD5E6kaEwMBaW0ZAmMj81OxUclsMdZa
P2Petv9IDnwtTfpJWmN5py0Sj/B03wFATHPdmGA3d91lnHFHvb3Hoyi38L1/WydWFJxGn4b7yhAM
wCrOQIa1kugd9VZriehEYFjgxKXffJ0TNLcpQzIBlt0nujwEpX61GfqHxZN8ly6Thdva/uPBUoyL
2Mk6bKtNg6zjoWA2dUH1e3BiWJyCFNUqTZizhXMelOrZ0Iq6uH0k4IuAbUaYREIcoGK/FMZ2k3rO
W4g3rAIKEkEzbrr4pqdYPZxccYC1Wd+kaKCQ4QtyQRYkXyHMXS57T3l+hlTtqTdgPhzanC48WPVz
nr91aj50jn0HJkIYaSAoeyipr7iNyTxxI6v9ZOrUm8vIr6LX4sBi/QmnTCteN1X5+UlshZKSdRRU
NtxMYQqt+myNSPmI+UnXNrQwjf+96dCWXhhJWrcEeca3OiL4pgSJSYrNeD+SzF9sEtQdg4pgjev4
4hgxNbGRZkvPLQj2tWyIo+ABQu+TfttGqUrwkzWNVBotvX5x9QxTFa1vgiiMSaHQn3B4L3+cAXX5
2gNifGro6r/Bslc/EfEH5/V7qrJhdJCP/sW+v/m5JaHWcYs1REMeLvwebd9x6nGnwaYNfmQGrJZL
jU7w6sCqTl3XJQIhEeN8JT/E85LAgDH1Gksy9lRlr2tu/+whmUWaFVeunQWg9oavd1OqlVB0pS1h
XHmEy6phAJWEG8OUvlu00m+sIsa7IhtPCuJ+VuFL5z1CtGrmosV82uqBkeus89Crw6UmR5OiaVCs
HHE6iY8AHG6rGjy6ksDNgneuzY9mGhx4O80ZLS387pK+3GLjvEZNr3+CbrlfbrcDy616fTVv9uv1
Op03u7EgSo+u+gJqwyUCl8ozqD8n0S8PUTZyVW218jrNuL+yOI00hePCO0piIsFh4kPB94GBYe9m
qwx0j8T+De1qtstDCPQMuWN62XbOkkDuI6DZ1awrFcP6gZMMSmrsVI2hmWMSgNWjGKtDGE5KbUSA
BpsPfkP4XZLVEecz/Q6d11GpgaD4POy8R1ROM7K/d33S0Qt5H/8mfnFrQi9hrW0LWzZhOUx1w5Zf
eX74fDaX3THKKUSC6Jhc88p/tqaEr44ErgzjU+4xCEGrZetSxoBtQ0DsEcIXkG4G3VC/JfSolWmL
Uv+o9retDCGf1dL0osurXQEPuO+0NKTFGCEllbKsJmkpHLfhUfu+UtX4g/WhTKBntlLo8T4+cS0t
rmrXHRFldsTmSptXNTnTQfM3qalHiiNnuHBNMJwVqNaTNxCFHcUzgS0aTIqyjMJ20DUxw1vewPRJ
XjpN35m5Y8DX737FPeVbak/hR04soQBh3jVoovhOpO6O1OhPQUqcrVmCfIN0YWnGFeULBRlDQQ4v
eFqdYPSyo525uJBWrH8kDUt3KSrwi4KTvlDEOC4q+DGt85/GzeWO7X75EMOlh1IMxwxLYqcEvVa/
6T+chNXei5rMS2yIorAvzLK6D05bUh6BaTAhM5DUPdIMFdiVE/9BTi5N8GixoWbmNDxSSWEnDHsW
sb4W3XijRWmLnlh9iktwfscqtVJnl+UCRKt7CBY0D46KxXQ6GNxWKnL2RYB/SdXULuslpJHwVJBu
uV/BpIs1dL/PpoGhSnwU9VcvkTnwERQkTSIqHuBgCRsvRemdr78ozwrJ+SkEX82RzD3zn7oMNvb8
d7ipgjKKaB7/8aO4qXEhAb+kCRLy6yAueDre+/ti/FWAiv6u6NuIJgG6pHKZLqCbLmhp19hUVkwI
3OsD2eo/iYDZl2kkOmmJ1notbFivng/cYATKynWFPYaSod2M0g3H0K5SHk07ZRaafoc67nsCl30V
IhSsXlz4WZNRXIfJTyJ2qDbMQEC1VW8nvjrVpQepodjxGhJEoY8PHspyMlyx43Lvowud/36xBfW4
+kUnQV+liliuU9nRCEmxq/fVIjIczZRNEYbJxKYH/+XTZjP7VJaPik+cgDnZOA8hak+KSrFwv9R/
4GFKLA3K3nuBoZnG1tYbrOC8GvdA5rF6PEdC3YHzqkKOh6MI6tQTpOu9dDFNKwHk26v98E69iuI/
tVrqe2P06P32GlqIIFMVJ1bHOgo6dLEUN9Ggy2P8WYWfkJO1+R/28a0J9/xUs3zPxgD4Py2r01e+
CCwJzFxTzks0P9ZFz6i9qabLU4wXGn6SUnoM45ZtBpBgDiGqDlYTlNGBfx/fDYKz9mBn2BfaNt3u
8L9/1hQVgDPgJHyuqC/1Bo8ntLB90TxZOSnbS7zmUlAAuVpUihtD+zMJ1jMPN0JCiKHSCs8s1OJc
vL6dQtH8ql9pd/dGHc3edyIa2sMzbvN0JSgrCDPY4VQOcCYcbhANPTBUeqD1gd4MRGSf8NhzjusY
pTNW0bCecER43p5/ltXyy6tXKJUloWBJFX0MYiCTjb99Uy4fCmyqpDV0OEtKDx5chIQU1hmpXzG1
fAyzmHd4HWI/NqfvI7yPVpp2an+v913lkXIKcy8X8QCsfRlv4r3fPBPKYxb/vhg1z25CKnRyk8Rz
RuHSp5i+6RNQvnk/nyhpjUtcaG89MFTE62Bmr9Ph6bEdFPqCwpe5EnRVKAxEhCvxl+2NRfyWKMBW
bCJxHTnOJkv0yhQHKqC8ODGUm1hUoqmxn/jqhof0V6cHWI0PZM++24iklY6eSG3tT4+DzdA3wNQE
MRuyTmz6bt/8ZRu99xFdooa5rwVvqNPEzViOIQ2VEe7X3nfM+gdxQetWuLH51WPA3KExbGG9SfGm
CTPZlfi4uMC4sOpxpB32dmZA2Owlr/z1Yz2O4cBh4NjYRQW6R7YLBNZKXu5PqPiDc3ebGY3i15jg
Mo5s/Oze+7n4dcbWdJRQ1h+v1fPsGxaS58Jgh6KoQ5wtsw30LwZI6iVb68TZE8W2xPNwcILFf793
ztYGZyHLfugol+5Pc91jK0yH9m8lCfPJ0j727GuZidgWqthxqBiC83Pw8mEoi78Er29fjiG6t5pi
d1i54EKbqgWTTo16VoNq5R8+h81fVXk/7La17xZOQrlinXl77Z0J8Dp5eWh3xMq2CBY6YC0OBTkL
IiOj3P43IoAz7YgxyK60NmneKtiFFIq48oaFeno8uR12rySJK8PCHDWDG908NNaANyLJRfE4iKoR
bqoqNb38cAMJpeRkW2yTBJPGi2+GRuQFUPE3QBhxHZZ9fdMCRpk/l3+IKbM3cedwww/DmPO+NLgf
oZNcPVRjOl2mjKCZ5eBz3wya9WCp7Y7OrYxMLaDbvvuF4STts+OXw/L66x+ZrgS0bBgt/iffFo9O
QjgxsQuK0S92Ul3eAFvuyHEvp6G8Af7F/YHW++33uk8+0Edh6bTMz6kkbptInHkNsf0Ja84aX9TB
H25MDAP8sTGA+uQYXmtxAY9bUcNccy+AFFmgWet0tnjpzhFNKklwqeyekmtcGWt5NpBTW4DLa0d+
fR5bNPqJSFDwBQPEL7BllCaN3ysWqIg7g/tArNbhGQgwOgizrUyTJDpPEzqXlwf1SQ7p0SVc4VnV
vZvT4FmCnjOhuRNGT1bRd5VgW8w+rECM6iDj1vukTdHGgkOPWegQBMT2Q3KWdbh9cWUPL8vzzeKm
H4UPah5AWVN2H5d18pGf4Oh1trFfmoW2VCy6KrfEq/eMAuadJx8KR3HE7bqBTDSWBeu6hF3u7pF6
FOkxQ83yU3jrmSvNuRrohDjgeqeemrAAgWdg1Zf6+vbNSprPisGZjdcWbEzA96iRmLal364Uwpr6
zZs4JGNNpawCJs0Pcbhq9+C1kk4+DPKivpiSll8PQwWKLv8QR566S0mz5LTwtwKsQmc7wWXqMI+b
EulgDXyaIHxVDjd8NZf0Vl6madHRtivIWlF49MdmnB2VhIknvu6vJB9vUJVsJct3b7psjTQJuCiL
ZcYTe5UOPMfwaj0upeHby0LBkRng6vHjjWj3w0rnWVk2NDKiCL59Gy+iUDyGTcl4pufQhsk+98q/
QJIN4DyMLjTNWRo5+0teOvtE7PpHS/by13Cvcev8ZRIRYJy3sn+mcOBqi7+zm1W1mTje2WMtjJJF
sPNrvgv35s18jFNJ9wY1mV6zXN2unxDVcaN7ZucomqdQGbSxDDHfGR0cnVVaeA2zUcVXZDvdg+Hy
X3hb4YezaI7agyQzZ1jPUaAXI0slnCPZazW0yDL74IKZMYEycau+ydVD0zNh/gI0W3hrq2jwZWg6
hg3OAnVEkU9Z5ezn3JiY8F9FwQ198ODGCfhi8eHCVfNPQQ+KZkeKaJCAMxZt02W5UUZYW89CRvNT
InUx10Gzjj6k1QED9petQkrLYk3Erife/CHAbWgaj7vHNLCSkyMf7MIbmqeLHoNSzEBQkuLXt38j
miD6VkjWApL7tew9949wAk90pYc0SnOUvpkrn6HxT1H+urHC3+WmSx5PfuU1egcBKCdVdYVJF9jw
G+9IUo2+RhkQIcCe5/Mtqnb+rgrcyaUS++w16FH/tHufXGNch/SJcCIr6nxrODkVakq1SAAhfdyb
TLkEp0PeuIbWMlqivU/QRpCu7b9Jod4kQmwusM2/2JeQfrex+7eSHjuNM0tUCwqx5ZDjud5t03sy
jaoZcOrA3EYzLMYGc3hlwNr6qtnQqeWLM/5BSy37VRQDLd9cHT3qzrOmEDZOtM6qp2ge4//wqUZB
zbfTkjY2HnJe5uqHJ1AwaqXg/CAq8wtTycOEQF2MbfkGTNWPkjwjpCulnzNdqHgGgQ33z3+qg+DM
TL/VydPn92N18ML6hBgY9hDbidWf8lIHHWMVv6LfPdUDOFPP34Xx/LxmKR/XoTvYK7vf8beMMPGI
gSsGBMwTl7hnHEtssW4ayTwqbCmcpjlkxaZh/OAcyPwk9DNP1X5wy6NUW5NUJxVix94Gny6+W6DQ
pPsLHgiJ4q67j+eay7Yl991gKh7+q710RmgkY4D0mPk6JCrm72C2b2xBt9UpSwf3GmENfet+o0Lz
OlwXz7NzVVbWpFBO8/JOqbO1H3yF2yYqahymrTDqKTcwOgytCHg0fWvSfvcR+QuXQTLh349jSINK
SGa914PlDKVGPDWOWH3GT+g8PdC0mZt1Ri2zLcNK0QCl+9LKeuROxiKtQKAsg1TE7pemSiYiTV4x
DkbsvaiFbpjZHB0EQRHVPhlCHzQjrQszvXbtJgjRFqNobNcGm6EsmnDMBHgtvyJ7Uyqv8cES4tTl
9uBCGf0pL6TIxykd+63QLLAaiE9K4NbcwKgfcnppw0n+X+k4fhjGjoNJm3ISfQeg3T0jYS2N4xJc
icQfqLNts6Fhu5qcBSlPTVqq1STGPs5hzQEj9S5TIWDPntC7BR0qnf7xP0TDuN6NB1mt4uKFPMep
RcJJKn63UVU8XLKp+smh5AJ9XnBdd58O8MYAdpOcq+h0XyR6mW1cTf0S9sIvetu2ulcmU36oB3Vl
F5TW3kHJmRZtH6gP7/Ub23d6eHG7VCAd7Ad9GfFWPhICpzV0O3m2HgbS918tGQ6BoJZMG1Bv/xoF
qRr4yFJSfu70fYeBHN02zEjwEIBpzt4wfYBtUAyFE/ukaAd15f2/rpaFI0YLeJVwn7uMlguH1jTl
9EkEC4WBqaTsIc0/G8T7mMMxBaBtd2OvT9w1HZ00tty7QHdHBwEEzl7xAgvblQbjL/cgPo/zvdKm
40OOtnadqwQeMr1lW2Z+ArKKMmCTjF5zLBc1HAFxKMAMNFFAjGZlEAL5U/uRr+QS1od3etb8nLPv
9eukpQRe92HXawAwhQBA79/OrLGjJv7Z7FX44cgoBpARvdBnod4ICx2GEkeXgGT18dnpci4uma6t
tI+iHYHUv/IRAMtVu9HKI/JwEOivHZ7NhjBp4XChv3IZGw1XXbdZtbXIBeSJcGOn8urAkuT0esw0
3Pe4yPShXb8ZL+iaz9PaNFbnCKz1RZro81VZe1EvQeVM1cq5FX9NrRmsl5Pk5px5L0jppXtn6d6h
RMBD8OwmBIxsDkdarhknzELHN/WPWOaSNuSNcyxP2gkCcwy5svmqpZ/3+kh8MSIvivriHSxuKABL
bMFqPG4/S08VVvFTHwVmjk/75Pr3nbR96bd7onQgxidWUBHZJP2xQnvvHUT5zXnfTQyHR92oaXy7
y+EpK7SRMTZB1vrtcW01ACDG2uoUc4SjxCRE9RZGp2M9TYv+Jgz7x+OHrjuhevkscRdO+dndsAYp
NHJ1ypaEXzp683ptZ3ZO6jfnj/YFuBlQyW7vNbJJRV1SmrgkIcZXlTkge3fz3BzdUHFUGngrTsuJ
0HJoOcTrqkKO5ARnF2nJuLQ3mLCHtfud4DCmSV2hcugjHrtZeFzdcs6+kp9Rm5dnoCdfak7uL6KG
caFrtQIckRVaRdSjVl2W8875oHFtCvXhOtTe9VXQr3vyDaE0QoT796jgjP6veO0QIpfDcTWGsTCt
zlzn/bdLuhaT9pwu4JDGnpxPanwpA3RFNYAM1TdCgXFUcmLoBS0ak7hEAqQqnsNdrZBo10OpdEtO
zZroC+ANwHptqg+3NGNl/xCUY+RYXIbZtyZYMTwXemjZGQ8htSAPtGrQaK6Z2yaebZQYHA4S2RSW
iWArv0gCquE45ZTfMEJUVnMyy4uK+CtXgR01UMy19zUYi0XLnZPFG/3YaRXiZ53UDnht8BoEgES+
PvBeH9xz8kKFGswRlJe9TmhPiP8eHPbnYZSkuaVqotm0dTYZBHziJ1TA8vAOslam6lbphf+Si49v
7wTgCTTjE36Opjpy3s8mS6vIc4YEhGvxzePeJLFl2Hpo4nUEBdo3+mPMtXwRjaDO4ybjJQ071gcH
ifjy68+mAPK+ipFwvCOYCNZmTLenDrqBNgQyY93fHx70MqiohT/vtQ1SbfWVJE4yjhAT85btOw2N
bjOMWzpPzkkV0YRykcAmZaBn6iTxnWXtOm0fBH2WKWZ7pDxfMjeHoKMne1j5CaGUnqBnhUICQXQQ
VldoZQMjjPdKnfcAMVbJSdfzm9H0NS3Y+DDot8qk82UcNQbKHqDeUSAjn7lPyIs14AFqLwkJ6EAr
kikF/T93HDdHJ1BzC0nIwJHMm0ButYKNoJdTXWezwbfX+qqUnUI2rs7nmtuIrNBRb74mUN/QoQt6
SlnSjg/RHTuSNjWh/YS6BxLmN71Gwf0QvydrwLwHXhao8luztOVi6b84ZHdI38a473qrNnRhCoer
rO69odVBJvZm6lkVMrUXLxKItgRMxycROPIrp5JpzcPUtdsoOQxb6NnGgp6jRFVXcB37zB9CzO+P
h2vkmD/+IyFU5bGZbmZTJR9fT9EjruPo+TggXwcG6Xlhuc5ROC21Wrk6lma0JLRLPoz5Xxy5ieDh
P3lpYN6PBrF/ZODZoTi2SOiQIRBGAJMAf3+Z+e9TNfTTVCXl1et1qw+zaUQita5WkxdXmelx1NVZ
Xr6YIp/7OjH8oCfgRrc8vKTWd0LK0X5AhDggyDy9JqIqQeWm5VM1j2oZTH9yzDaIgLGhyZMyM7ap
Q4e5obR3V7yhUt1WiNrs5SysDQtxJuZllqBLR24S5mhfnQtOnl9Jlp2xopnI3y7JbKVzi5u+dK96
yu4IvjigLzYncNEdLCoKc/FRQpG3y/yTRiqOCG3saosKHlMjNK2FG5bz946yr4DGdvA3Y+on1REo
/ombrHIYJ4bANrdG7mqSwQotAJ0eQCkbSlqow28sQZB7TfgnSAVHOBRSsGFt3ro318jRT39AyZzY
Zzu0Dj8pYBHj7Fpe3Gbw/fOFuzQaU56uP0cVrKv1NUkTi80NhzG4CwMZluyZ8OXn4vu+vF4QyGh1
l0iToTyan3H1JtVqwoWM7hfIMlIZjp5f29njTMKBrWx/PYfhefn7Z6L/nr2hXm5m5IHDYyy2RZhp
roMg9IRBUNtJGzm8F2DSk3733I7obNuXCxDV9gnU378U+iqeLPh7+ScWyKuLImyAhXG7HBkYdSfu
Ctf/JJWFSNeFv96nUKJfgJAMbdOIDAvpWUi9AzSrj5NyN8309VVM/FXw2LBh2u6HRgLQs4gZGZkb
MRjSlyzF1O4gsMZjaEoXLw35YiNsKStiiePC4m9cutdkVRzuHvwDy2zFm9+EdjVybbtdW4z/J7BV
Oxja8/hPASzw67vHfxdBg/wEnZXVitHxcG9YGcmg+d4F9KVriDxgYgVJ3fK/4jRVCXv8RSWgkzp7
T1vgeSLemVjUI43Dqw/cB4Qk+gMBZLBjWWQhgO8IhJL5VxUJ/+r4GLiealOUSYLA8IZ+hg1KtHb/
X7UX9Hi0jdWAp81JTVuS0KCCZg7DxDgwAYQOPrUUvhOKYq7l+mvKmyHAbFdWvUFZZ+OzopnZ2tWM
ce0S9SrPKZYGnVNepnzbjLlRAkTf9YHrkJoSZOOJeGhexlYJh4boiy1hhmHB7FjtJss3+4v2XPjB
009pERIbE5rPGfiPZX3gBdPxE9pZdVbtiOxJs2om1yy7bnMdWY4ZImcMh4cfHZ62piSdnkNsWzzN
TvHCclnQWzqtxZLHb726g440/yZxgGFSTwHmw0bWRYySz1AX0TkUPSD5yw3O8sXoKsUZnhk+hLS/
RJ6BWqbNVYu71yiiCoCDjaju01VfUI2WVkIFJOaOXPEhbkoJCQHs0Ucz/oNz+KpiNz/HS6j37vGI
xnLmq3H/xyH6qqzbRshCKzBHntcov9SyHxe6ZAWnCtWY3P7qjisKfob9/S7sQIoj3cbjYl6aZsfP
QM9DKqG8I+bKzT6qyAyskcWpGalID7hC/cFot1a/eM7b5DWEwCHWKh7mNLHm9W1TOl9Fbb7HwYUT
vNA40Qff+Tz8EFdT6ONT8LOkCvoR5xy+0xbEUepJVz4FAeCojo/rkmgUcI4Zn+OOy9GUYDUeqqVn
d63KsKudkuFklgcsIOLYuNu444mseUFbMyoR1t4ZmAVhPYsHCX5DufSGLU1OkNBdgKTt9KZViHS3
X89OLabWiS1phTkeNeSft2Zx+YDCot21SvGTO6RTXalxmR/k7yrHH0xsCHUGnZsmVlE92SV9BVCi
wlKbm3QH8Alc8uRsPnKTJTl8xCZ6SEnG8i7njJnSKkB2dWu1CCcmNfUVNs5wM1PcBFI81KyXucG0
dQZbWSUXj95KctmBkgP1fdIygufPo6VhJDiU+dz0490hx40hLv6GD+B4vEPL+Y54JKADabL3810C
H+ZRGWFrNCgMMrNRulzeJa9N6HL2DtT/PvSWxu2Kjyj5CBjRvU/GucA4gNamB/3ydMXGYXycXBOm
ga7lWKTULbeGXDCb/9dyWwxCrxpX1B18LUyOq+ryLggfApPfcUVMhNJd8g6S2VJXX9W6fpmqQvgQ
1Kj5u9RyaLxJBMH7vEAzWazGkjnkV+CTsbR4Mo/0TYuF2UyoRzpGECbXCAOaN/z2FX7Gc+CxgyvW
0xaeLgWLzX6WO7Pib7f0q15xIAGnkysYJDHi7Km+G1WIm70lRjza1AvRv3QqHWISvR96lXqXppWi
xpeuJwDVJ3qLi9z2KS3F6KucppV9hDHd/sDtF2HT5nwoQyPk0zhgzoAs28jXOKSMjse92FYL2v8Y
2lLNtcnR3kgXDW8POb6uU8Ri3L8AOdiNamqKi+fOAYZjZpS7MAIk0KzCb/8bbsYsbEpxlUse9wER
1oNs3VQVSn7r0OsqwKKZeM5kXDW/Eg4Jthztmq9enduujgqBo/70l41/m6atU5RNbofZN1PdLWOV
Vrw4wzIWGE6n8FQB2mU/Lec/WiYk7pFU/wM54xpiiaVheBwY/5LbA/IrJG77Y4xD08j56waxU4kE
5u2EnlZ88QaL0C7P3kAJtPtYK0SI/msFNQOyg/vyQU/hJcq2083lBaW0s0iDAf1i+jWIcqMant8L
Xs74thMMDzxaM06a6fBrWb5aoNTHIeaSIZReFV7POKpH+b9GdagxZ63J+T1l4DlMkYbLYtLySx4J
YmY8999PzrprAQ6i6fMXvjHaEO99LfqgCcEplNbu3TdW2vy0aVszGptnxcPb2hx6fvv6O7DsPMNE
Dypog9QAm0fJVZFgN/DYuzjAVTSHumLM8gmBNACY06S3Ut0AnxT3tQO3p785L3Efr3lItHX6Y9E4
PdQF0JI4PCTX2Lq746Gbs8WlBU4wMSl8dmjdsuhME5S5R0iD+3SfpoxaqD89P6RtMv1QHDXo6fRx
06Jz2FMbUcRiZGS3vilVv//8MYGMH8aOsmDqejr1kesveSvCN8a2lczaIOOdFvAW+w3YzVRp23DL
S6ki+I7FCfOlMEKDJQl2yFqGIaIPf279J5W/b+QFNgw04FSrBSmeTpxieRuTxfaxfW9qCDXGU3Lm
H5radazL4d0USf90oCSw+vx7ZU6AzcYoM5hHktH/UyhnzbPSyYNEtEkRXt7FmY6cwmbVA4Rtt4/S
tx3STtZ5qBHITQDx729Lyv+fuVU1t5d872i/I7ImTfMoUp7MXUb12dGJcIifR7bfpnjkSZvMAoWX
CC0jh4ry2pr8GvCRDLMFZIn9tpkQUqT/rcKwesWJUC3FN/rIWUUGWyJdyMHk8PAg/XlgRR5efYJ0
rwM7KgEox3/dPlMW1nLMHckIQhjfpJlXoau5ENGbscVYeSrDALsoRqwDCpZh4xJs1jtEJvAu8RXJ
anUkjeFRpN/FClaT/v0xC3MXz163Pz+Uj8w32nItMajDpUZnExQeUuON1+kky8t7+f5n4vs1bnpH
mlHXgyM3k/WXPJFT3dxiIihc+zCdDfGQuPSNQ4wn3uuwgVF4+v0vbstyEBsKuYLxsgp/MRAGMS9O
ISxAPHNes/0fyTdnpyAt8lEEawqywKHCYaF99inAoqZjA2pUjtXmuJ9CCoPRhE4TJAr2niZ0JwgZ
Vf/s5yZZ29YOjb//Wm+a9/JjOhoR7lmfuzHL8e7wqa7NeuF6K3Bzca9eDj7qTM1UCU6ibCbAd22e
JVDvAc1UBtTifgjUmDELbTr9vhlwPqQu1KFBzPdbmqn52zdRlY9MWBjPeAT9E0Aea/R2WKAV07cB
Bbx6sNY0w9OHgiNzdxGVbTCUQD0N8LGb56gHV8UbCOueGY8pnjHXyomxSOFbFA3o3EFCchCQ2/2J
Ys4cmryRnboI8IRDsRMlppI469KGWgVZdeeHMsDhncsqy558D0HH+cM2faKITrpdCylLJHrZpFMk
CxFh5Q62SiEzn527EMu8uWVP4CNcqVREWuFYKNYfnpKE9gCS2BUZFBOs1v3C3abFbvAzwMPButrL
/xUTC053Es0NVROAVvHWNeLFQ6nTZYCI957OaP5XAtoPSxuo2E0BuAjprxVmIy4VfytAJTRcN14m
SxlfUxFrJ+byzTHMH/z+WyyXF+8IfUNmrVaej9dTi5lZyl/2zWcDGV8vJ9uAyVlNKr3PKMA4dTn8
VIsFZn66xPH0YIAntMdknVsJVampItSY5eZ4vWOhLdv9Hbv0cNjHdtO1wfB18ljTl2HPl6kacQH/
CInBmvX7xDxht9ksp22/HJ4FVzUVdZ86VFERl1iuH09XrWpDq1lkNgGrJyVRsY5gKqvxlSD3zSv0
xSuk898GTzTvhG/UPMP9JPqaxhyLQdqnU8Og6Q84HGPr05D5N/300nXQeqf7uV2OvjpsvQdqbUAG
2D+IBQt7R285XtftT+wlND7z60gKVNn6mZd1v6HFFdA3wu5l59xQS3i1csE/y7SVNfolmuXT6Wky
dgnh8VZXjt8PEwZjvtw96YS5lrAaHhGJSkdl0V9i7RvCvP3UP0cVWZazIBqyUdf2F7GQbhLHHPor
S4c63P7ZH2mWZPotGD7etRPbuAiPg8xg0hcWYcLSFOpiBnMqh6Z98VvCzr9dF/JLov9O4FH4mW+v
KQRuQQGAMLVMbzT69a1/O8q0jjL123Xt9VKQdvBS07TQJyniJY5tGfrTpEScSSZYqcsc01+78Ult
MZYeg8xUbYArhO5xbKWR/KKu9Wkcyktai79JX2IMgLIFJ+ycOt7DS4dlWhu2AA83NqDC+OQ+VKlV
EtI3UtmkNtKQiUppUgVYm1Duu3KBOhgRqkFqMFsRU4YmpC256Q/HRx1TFWymkqtLK0MBuj8YCiqu
LG4QuFYUKV2hi2bfUy5muFcPDKz9401cLtzkXXSTSFXtPopLPBrVkY3xeqgMrf3U5XVq9IA2FevR
4wFhQPFueJrwoKy6zG54o3AVFUJRwUoVmu2TW/jBzi7lh3yXiQcAdVu5rCuLXOxf1wbp+03UB+Kv
Gs9T5FGBKs8yKqLsM6vjnrCtcv9GzqxkvCFepaPHLupxLr1UKpYb8HWifOUpkeyhwVfQXsyf+w1w
rVhFzhUa0eS/q7bwqLGwLFRCydBAP1KX8MwvHG0Ynrfm1eUAkFmHRqDffY5EFs1JoZ+X7fXXmWMu
z9v9ZUhVU8LSFr4po56eDTyU1NTfK8CpSH0NY4ed0Up2xZKgm0mju5qPCbzMHmMeO5YC19cQlGPy
DKy/PHWxvGq6Vr23GUsHBJB0AyANpNE6rFr6WxBRYsU5XepKprWqONITuy7mUv2vOfTVGsg6Qyws
c15qi63sTO9s7MO8beo1SnNMCNU93Al+X41GOvyLC8CCNavOgM2iFhSllokuvsNRy403kQuWMg5v
YamG42Talp1r4IjFc3X2rmOWQ/WnulwLPtpC3hrAcHEof0pClOKEbjxMxI36Rfr+gE0AnbV8GY8y
LMYRuXYrZYPsuWvK85AQwd7P/vp+YLSMsPL6ie9BIjV1glIExkFwWB2vSJq1J8XIh1r4i+COhHnk
bUojLcTdazH/cg8CJVlBuzFHHRt8QV3pooyuUyghK9pFDO8Ualibb+0jSJ5T0JMaYqw4wjKmfLrl
pMhKhdSjAKR3fKPmE9IyguSs6HD+Kv1vqAsX2s7m85Jg+bQtoHWRA3tyeqFvSTNK0zRLFZoeJlpp
YeezoNnIbah7HuTnkSENH3TCiX0Y3j93A21qHjEA7qdok8k1XClB7E7nCo0Dj1uLxIo7vndjF+8F
N9Zj7/dATgU+P71vlDmQcUqTBTeopei1/ZIqm//UN2VGIIlzo3xWHs74eQprYvi2rPzO4wQY0oh1
KX3FifXaeemolCUlimbaeqrNmkk1Gofy/yAHFpyTERO1yEpXyx4D/9sabI3fiyMYQ8zOMKVweNyB
zPbBClNjDRcfpiu/ciQHLFbQoj/T4ONja9fKM4xmLVKLHlJX+IEDNZDLSuUsiVlofkNz5IjAax1g
S7oUwRXFcAzJntlbXom/i0si4WAp+NjpkEzytfZfRA9RdqBb3owDQkIk/TE0h+ehA6jOz9hQViEz
ByLXFdA9FCeWjGcTAsWP/pQInAM45Td0CcsHnh0lHBOBJPSfyqMnKuaZYFplMBlkMw+xDUyUuUXm
x6BanFlrdWdZizIT0j9b+bYaK+3lUmamCAKm3KPgrUZ7wtw5NNq9L/1LMUFR+VH6MOOIYA5vMCP+
WmYzSb5Q+ztmcXI5Dt2U3M2klTXmQrXHalVCn3bFAeupI6Bw3Mn6EZRbsKQjOzyTo2NBJ+LXbwm+
hcUAqC3xjf/+TZEbWFwEbbTGINfJoq6uzNW6R9HdHqkvPYGsC/vWUKL8jaAruyezDosTSg8xqRWM
oeMQrdMOjmOY4X2HHoEkXDoBLzial33LklUAlUe+Vqffco+9JlZ7rW9R0mxvM0Oo5cIY95LR+xQR
jU0or01wzELgOdxNDkxfzLkQRWb1k6u7b78Iih2iktpiwknKgvQ66gjuvwskA7/FM+326puSV8X6
RrO98KhvCi7VaezD8V4dxmHOS+TiIWJlgR1fwYZEkClbXjLfPcbOlxNz1ivyA2SwBcZtBAhfNQ4e
DhEfaPApLd4xq5lCMcpDnqzb4PQghYcgYF46eHGkbU/233FO9x/74dj6xIRMnDJTDO4kkDL/b1c6
ECqtwUjO9L20YfSbxKXYoG4xSDvIzvdxy20gqShzfuETnnZYTBekZOdarWOwv0MAaQg7ug1FommK
PGHIAJsYn3oZ4bKZJ0bluOi2oY5zUhoUmMlC8ZHodpAbmrCrxPXnbwZWxtH1dtTgkflBVnkw6ROi
6OA7qhpncJG6ZD4HePDQ87tmu8ZGgVYrIkimkxe/ADJHVP9hnGSrx7ofUMQvwi4jwdYpXm5fq41N
3lWSFKgRmQ+XPm3waNCNpTALwnT7Mml/BBL8dfJ1VgoW/9m6eYmR6S1sR4uA1lS7gfaubinJ01hX
w82GUpXAfJEn+ATTl0Nz71a1GeXR4OUgq/ioeYUrm0mBSww+QGiLDqkLtVN03Oni27Zb6D2sItLl
PHxOEDVlLFiniJmV2ncTlhXmvhrkFy/rVf80FxSdnkT2B4h41QhqxGMO9AfaSgsmYAvKzLmGGyiG
fjGK1Qz0e6aHrbpfgP9bAy2iWbWwKrC3euhQSqxjVKXzto9Zapwn/eRyfYUeHTgNrX3UVXcFwZYb
OaJvNfjFwH+76WH2s7kE4uQ+pBfQo0Ne30jNz+GRC97hx+c7ahgCPAdiyGKO1qQyBXYgdFWJLs9u
t6raJpio3YTp82o+uILz1kY9SoOWnv6DYluCioZhW6XTVoUfceO07UX3J9/TlWXRCFf3MtVJ2nGd
whRJ/v/emLp0OhWDtLJkCLKilrrvb6V4+1Id6mTGq3r5tAbec7ZAumBTGG6/UulNnRRL651ekGjs
GzOPU2h0Pj4Bpul7Q+ujJguHlBGDu3mPC6bJx4BHC6bXh2WViRkD824ZWMFmJKaaLr6pl4f6fXYG
buosEjAY92RmKaGV8+gech8k0yPzxAl1RStem0TdcCTBUsJac/GoPzNRGBr/Okx791JXY/Ge630W
aaoO1c32wOXtaiOL0uiaj1t/W3t/gmByMoVr0rAfSJv18gCDDEGQrrRfw6A5ntONy8E9RY6oPk+h
5cLpY03FpBfcvg85PcQRXCOnLifXWgFxTiTtAnocTxSKSeEuluSEi4BIrL8uny1kcVAnRQxH+qy+
IBeTwLR5cMcMlf2Wvtii6Y1P0vAg1ebgFwrM0x27kSaDWlrmXTxaT2tqv/RXLi0E4wbsYcEWZ6AM
5lN7XjRbqfM/FyHvgaktZtbBpFAD9NXUhP6NOyOJZyh5R71mgcvyV5WCUWz824rbi9cfpmLiJsOy
A9ddzKzP0pbFeCGirzToEmgn0JrIueBjvaK6iFQjPsJUYyVG3uzNJTpg+ELXYLWQHc2H5ZxWD75/
VAU/OANqCrMqTEe7ZPJjrqOavjKb3FyxiY2lpNDN5hk2wZdGn7CjqrUKd/nQN8aQmefF7pK0mt/j
vaw2e+kk/l5qDFyovHww32oxHz1a2p4RIWKQNnNzrlSXN7iV10mXzjzyB5+zidBggPZKWCF01rDn
thBpYkq9HPUX5yJT0u+5IMUUNsHTv2ZU48gkP7TiQaM/xtCkirBB7w9xErN4dL9WKvpeV6SW/cGM
+eCsvWybJZoujqZZeB7Qsx5bbj1FGFG+0qqYP10/lb96R2+6sF2h/LEpE6k2RK3tL5+RjgrqArZ3
fSiSzp4h/L6y166NyJi/BfII4uncYNTgcgjuO69w42NDIEOvwIuXXvmzEw8cXZePaIxPY+9Rap/K
uiy2Exoc8Z6QicPdKnIGPGh92lJsyI3+4kgCNhL15YfnOWFPvZypaEOc1vTnrG1aE32JagCr3qFw
ESML95eVOclKjFaEzY6PUCNUAy/gpsu4pKdmIQX9xWtJJCVmKJeNYIRY74Rf0kRG+49M6QWNgKsj
sxJiHMYZ5eXzrCw8N9FJGsfmjolceCJbQ04S8dMuAxX36W38FB45mMS7EA8x5Prir6dKG8joNosL
1pK+lw+GBkjdBuwDBM/W5qFulKi6Czi+yWgy+9n6qPLj/rGzxMfjwXiiFOO+833SCApaVCVaVGsy
bqctdo3XUedwphZKua+SlgXQJgexTZ1YvKSvmhlIPiP29CpI9OV/XfSZheC9LRG94aPwQ5g3Mxqn
V5Vyvfr8pL0w5nDhz9rRoMnlC/R6ef/n+iovqHZfGBvPVBDFwh4XCi8fjfsYpmx/MRCJCuSYPFtr
Xl343qOT+znkgX8VuioErqRvsPmeMrdTbvThSOpEJ1TEzbibqee9paX0UfKP6UkZvjGlHblP3UXt
e8lg+rUFUOsArCFfCyVP9NIoOXSkTLN3UPrZrWC2wxQnEwIW4HF7Rp7kctOzIHoGdQYIjlMB3wMC
ReVbKlA4B8q0JFQM9KjD/EMtOsPSafl8Ax7KyYKA5t7SJGuTTMkDD+oZFVVpRV0HUqIChNAk3HaA
Bw3hW5DjcuS+Zj9POrtna41HIuWEPfCnFN10yt1/60GqWFSDv7noYWyEART0E39SV07YXHhsAksn
E5pyNSTnG1bAMvLIwNHDqA+pUWRjaX5dl9dH9s/SxqMnsWksJu7O9MdK6+oZdyHApK/qoqK7V4kH
VyceoRUNYzI5ooPRnCK0CDQl+HcshEuJ955MnJiBxshEMjd1x9zgnUK6vEncj/xx+/D57Q2G+OR+
Y2ZU2Jgi9MLYoYuAwBu1uu575N5dP8oxrHC5CmuJVvbjiB9h+zE4xgGdD5A4C7WFbycRT8tqaFNr
r7AhXHX1kRV45NjATBeb7//woqPks0FniDnzOl3+wOs5h81U2bLKBtqsGq0kYpZcV8TYKyuxpBJe
lpdxtHyPJ8Gh3MEUFOQWboO35dLEOYBvwCLJAV+k3ugmCNmdG+6Sj9qolJhf/qGFUeWxrarFTQj0
4/fXumuEfCI3d53wv5i2LUNdG5fMBmXNp/3QW59GkC7nN6q0WzKfJz4Yh/nhXUuNyPxwvNPh40aS
W3ljWwOy1tFg+xFpyHMhjj2XPgB2xk4LYb3xIqcFX4KwKQ15G2iG8BG9Mpd5Kui+T9EaUjkg5nz7
ORqNYnAf/hdKWubb6SsEFH4+lAN0EPjcLlFiXYgkBXamitdQEc9PzRjhN+ZZYfpbfB2Ev8U+uJ/Y
GB9uwDEM1i4OdhxOJm+uz2BfngWpDT1cWSxd+7x9jRuCj+0VWzGRO6uT3A2JWX2vYiibFRdKVKiu
yAkGZBp9JzWiikDrGX5Ns2p00ytuA5MskDuCUJmqDm/R3fe5jtGoNxZJWAWaCfQQsDN+4DWnsivQ
NgYD9L/yKArJzzvdrL28QUsbtMqL2vyDFWwWrMklzP/9K/y/tQM+CQviGHac0tH4vJYQzp2ZTies
adaER85kbPeFWYQ04P1yVXFtZT6VnUkIMEH6eItYKXBA0vn6C5xCqLRjLbxUjSdoPgguHCqccBaW
PqCTqf1VO/GsicNtRCYjTX+5lkeA7z/ZhbRy45AVhQH/1RgCpL9XsT+cmbyeAzsYb/nrr7Ld93k7
nIQdBJu8lVTAzroDVe/VN2RJiXOL4+LCklHvneVmO3qQ8Lhr+MQLa1HpWL+244vdrGHcEfh0TTP4
NFJT+XMgGT2eSJIIFea4BlMfLGtI75JiW2enXhNmBTB0gXPvqpwkzzHm6EviR7fX5GWDGwWCUHYy
LEJuhKNkbYrDr67WlWnXtCFhhC5D2yA9jw3j4HqcoQfSqEgLYRXdDU2w0ZQIOS28D6L61f1GqXVF
VG2k61k3HUd64J0kPtUU9NU6cXV1ADwVdW4hFCMS7Hogx6PY5HuWMUUnXmnrPtY7lBPnekbnahvV
ta1T60IVGquvB6eVJ56UP7u/3Btr3yEeechE0mjJego2lL+SFfIvZLM+i5SmF4NNDilBStwodDHY
BqTHdLXn+Oifxt3jX28xkZwqPWE5GL3+ls8PldFXwGakm+4fJo3hP3hlgMniTvZM/wjDT8fTlTvm
HQBan4rJ5QdFYFDaoy/uXOw7PCcleqpylzoVRboZMOjWcTX0vvElxga/msxgz+9sh5sBphuNgVT6
N69yuIBCq/1RJtinTmO6rcUf3KuWbf/GzapVPe1lpL0QzJWsSUERq0s4Qz+GiMs50fabgqnroL1+
brIe+R+9F59bEtq7w0wYms7cprnKOv5TXmny8aMw8wNjwCZxKvVCycMbVFR5wMd6uQWUFUCCnomN
HOv1lLqYa855VMXBN2M7mu+E9lXVfI/nQxTWXa87jlCzBkZ2Y1n57nMpuVcDkthTZ9z+zViAMaxg
KfHaO0r5TAbz2wFndSGoe2oJn0SzbJFm2KN55EBtncPcH5A2s+WTvXioQX8OYNqTCeAe4m6pM4z3
QpN29OHeMqUbvjahiKZZvEdpPi0pwQAwnCmsty+IXzTtYRbC4FQ1eJJoPiqSJ6s158dkGT1COdws
a1+p9dejedsY4Xd7mk2zxgCPASjiuux5G96l8IuU4KWfgJ4Ss2eX1onoMy02SuHCKd57uTb2k+Kg
9BrF3hkrEJAPGUGXuOhadK2OdqPuubPqweUan0HnEQIAmr6OWie5mCJp8o4ZlBHBqkoM1WqE9pcz
7+q73rmAQBEsfIA/ub5ilE4NiUvoCkDEPIyCNlyEGkfqfnJfam3qIS71enBJMj56iWBk3LELGcc/
Sxx+rgu1iWS6CahDhT4TWf2x7Ijx9to9jzUFKBy1d2HD/7/6v+3W7iKqzlAsey0NKYymdrzxvFDP
nTIMt+buve+b8b40N9qqHu2sMiOAZERpgh4ajOyb/iIpqkyG9GkdXTMH7XgA+k+czqfE5QG80OAT
qXsPdg0HrWS51xmkPXnWe/vfsxZv65Cd16fhb1Te2OF/baN15OSzf/Imr2mx1Ebx2B4Hhz3JMfCJ
7zF6hISceivRNqJSehvz73Bto2xGBVFFz0e2nGxXQeHqKEofZbuM1jYu0/5ErDUkORwliszEVG4l
7wrVfm6jJjZ5M8gCXGiOENc83QTjV89hmCpXipHWoBqvzyjhl61RiyAY90qkaWs0TiBG1PPu2PUU
37toIdOIecKarOItq2UPK6O37SLeUwXux06lZSzLMLRgKB63hW5neEzg1REKaTNgZRcFmOPPO2oA
haGSNS5lRa1dhx0JjdjZJAljWZVvJJUrvPWmnIu9xxCYPYrQ+fuWsIVdIYoJdQ+1fQ9vtmacFwr9
p/5bzXJm74aCTClUWvKnRbibYn5RNP9VtcasMFte3w5nmt1X9gt2yRj6vng9f/ipROh8yK4Fr3df
ZDhoYnc/epV9fdjVyMcCgbEAdQYLbY80Dlx2k5LL+L2HJB9G7leaNascHIVIRk9TvCvcOBM5fVQ9
Vjs53HXKlnirjduORYDg1Wq5kDAA4y8Eo4YpL/r2GvUgglUBkZG8Tv+EEEKYizmRwy41vBX1lJT4
kxWpYGBvnCa3s+ye1xAmBTaaztHOD32acFBGfRe91MGYu4vJ+oohC9PwSrrNN9dr+f7oE9YpDBX8
GcQipdCjY4u9KwmWFLlybpKae24bmgbrCtWhAcqGWSHyIyMAcpPP5QWhoELyaIUJV/RzpPb/qm7Y
Ju3RoWbpp5LMX/XkB0AyA4Uu1MwkVeKI4B9sjLjMHEH+PPoObzQxtNQtn27Ca+kEv7X09aXkgMQN
8wPcSb9JQ+LSdy+MP37kLyXvRL0d5tLfjhaSvt6KDgGqhu+Dc2+HrGsZj6gFS9dqDKlYPkMtt8Ps
bMK1rR6sEpKernlf5jlrYfbeqOPaTylImzv4umS8oOjghNVVkO6tWPK8QFxaUsXMeJZ0lO1vMMHX
D2gOPFRksPZ9Mz6dc7JLGMewjbTuRmLxSfrpk7b/+v3UXcRmFS+CFJJ/bEsD/q1ltNX0kBUY2iJu
bxt6+XOpqrchNsVOUf9Oi1I6h0c6HT2i8XvJalSJCZTQD6JIDMLc9rA41HgqWz+8ClMbrgShgIRc
E9cRehMmWeXkqZKYoK9ho8c6o5pQCY7PlnM9GPbrLl/BqXNfohM71PDn0JUBOCaFxtRdzRyf6Kv5
MVkxDDdgQ7XvRjzs5ed1Rdv57rZXZAPkDCeNIQaD/q4Crbi3r/XcEWfO/Y9BAklNMlQphkDQqlJT
xUoCx7OZcDEj60Kj2mVfeN8fmy3hyJhE6D0BpgFchZKkKRjgOU3IawCmbID5sZ37+hMANE8KKSLZ
LW6jRic/1pYH4qUR9DxRPx6leF8wV7Nty4R3g+aVePaflTZfM1B1tzOfxewEIaa0xqZmUbTpHy0H
HbQ8OXiKzH3wW4HnKj9GmLjpKydOAWX+xAQRqwVHYNYeyP+EUJcXm2DKnqVZXQ/pXMWrJhEIm9Y3
8z99shsyXk3gJnuqWexzXNdmnZCsScREWOe4XmHox1wp5adBRjBBh5on6s8aCgaT37YnV1Ma8Hgz
yp2LX3u2Um1OFiaKSokb2UtRYySp0uoCM4MC+OyOvtI0C0JHwxzTzPgRtb4ujqagBh6mt5op2lUp
kOo0DvrcaJllTjGX5RPTxBkWuU5IiT+G8IXGbuo4ih3epVS7VY2zpW964KKECTKZPrXQvF+fyKfZ
fwh6HqkyFXsKQrlMnFHrxcMHgmJENKdwRzT20Py63L4XrBvpfo6XM0MmuHJoY0ZPo7lIPebnWpPk
AJzVD2lp1V7I4GPn2AnsCayoe5WOfsDyWQgjhQ3jjLQzt+ReffzXBFMiJqTLaxOxG9twSN3ajxL+
wHK3958KbZkGlIxwzeZSdQfdz0NVMyBwguu3RnV9oKvaXYQbQcIayTTHqJZIShuFDpMyn572Wcbw
y96uGzD5haGYgOT6ZOhF5G1QcX4vJGpMh4Vm6gmZLQuB28GTV1v9k8IFZyYXgjNyX30wbKCOkKy7
ragL5KS5Gy1RQu+2ippWtFD0zYtZ9O0vmRmNtLr/w2Q9+aYhyvq4dhdRWq+Hczb0lZeQQATxdiba
HsNTuyH6yDZsCclWsYESiK4uAIx+Lv7ifWZZmGLxc6Jwuh+0MlQ/TSfS2z8Ughnc2rS1aYsVwarg
qtDS/fKfQCrYLgOpa/VmOkhOQIV13M+V4KZhxMRGwdQvgXRMeUue6o6jHw0uxdaZkPMvu8I4VQZh
1L7DJ7v8oZ+3IB94htjAMMelUfDVcmdk+XGZqGP+l2h6iwWa+09Vac8GMY1aazc7rWEcC17wX2Uo
3aEkdcU56Ty5JNpctgi91qBC+Qg76m0cKZAeW89e8P2WOrrNE3gr5pQkg9xVy1ikcm2nrZS74eX8
SH0UX8qjkJh2k12Fg49KTBqbUcueI9laNpGH/G2xc5nvuw4a1QaIWPNjNubaiY6rlXL69wEoG6Ka
SpEpXWtEaaz39Q8oo0/bdDkfTLw/jvArYzn+L0WNBIHNpj0zAVYrF/SHwlS85FhCSYiSMyGd44Zm
naJ3KQX6DmPQCeEwuFKmCdUBN6/sf/cukxDcAPAmCC43Ldq4NR74f6bIey10KNBfOWtNz5KphWYG
z9sceDyoAkdODNfark8Mnr+mGJH1KImIUycT/zEFWhr+menU6FIael0EvjIEaMpwh8Mq4uIgOJr2
cEcES7iAb3dsFrkdPH3j7LDpEL8L6rOl3g1GteOkJ+WejpMdUnuKIModxM1gm5z+LkP4eqhu97LX
pakzcsXPNL2nN98nhaZo+mhxZOnWYnoEa1IXoZ01fZrBZw0IUdSZZ1/3GqcMO6vK8GsZ3v/hV9/Z
j1xM76oHBlT2p1vi2Z6nbz+eH7KVn8Q2rNOE9wKUFztXWm5Bi991paJJ2kbiabr3cRmE+fmricf3
0txXd7Q8WDhuipny+BN3A8vLOOsY9v4LhveV/ng9AWRxg4XCrgmJGaIsDDrra1W3wUrWPizEj3EA
BQge+qatc+uj/zUCT2J4CzHH52IAXV47F+utvo+pQvcPJPC2NMFqkxDUaP1EONNpORy088YSaaeX
9NFcQBq2Aejjn6AcPQBN9YGrdMsbWuBhmnzxaeXgifcJ1Sv0ur16rEWyLsrRek7ZNFz+jxgAhB14
1KKtv1+8Xhsg2QtPcr9AJQbO1n3aR4HXA9s0VyNkdnhhqFbtgpe7y052WTQw8K/4EArWKtf9AIIb
/T/Ydv4J6KJwjejgsp7ACF+dcNkRmzNpF4juxGxGRMc6VsryYZkXzQpHXKQ0iVHgPjwr9owaIVji
6c5SKe4Y1PhIAXTew51UbvwRcj8yxtZBMoFPh9vSYLkA2SdY3MCzpeIrXQDEx+0uiV8/pXzYFlQn
niU2HrSupaUhQ+9U6bODnGv7jZLRh1GnB/6CfzYcSuMWNSt2v2p7T4cbppP+jFJ/cBxm+kB2i5UO
HLTvjmSGh4F7c9smCQWELU6QBoeciL2fcAU08sYn8iFmMMjoFaqw0as4wfEvh4PN0acdEZYNymcu
u1V0yKjbpAnZFx+1OG2VjClZvbxK3Q2anJ+ek6S4igRQ328/Z1H9dRWFh8mhaEVnmTchlj84d6F+
sVu7ZmB0iqHGywVwvhfRBrDwv7fhh55KzZzwGNgmiqTj7OCGWJmIl/sEF09gYj1qrfJ9oFZMXwP8
mEToUYwyrxjb3O3EeuxH7ExCsz9YarFBR2mrPWTPMrDbSX0vwWuM68mFGm/6r21YGpRmgo6M2RKg
DUN4ERWonyNywh5M/S3nZsbng5p+550XaMwWQBFopH1tNChoq4J3L08xZwTacYZpPztCdOBsVPqQ
e2WS7seUeAmAzmGsvny9jR+6jaeBnUhbjN9HDL769Yb30e80kLx6OkILXI/57a7sigofF5XdW9AQ
fIpEl+LVhlgj92mXD4fxBDxtJbUpEyqZnXydtCp15eBUl2hw5D5WOA3vYCUBYDL1ExoWghmyAFJu
W2oOhQT+19JRvkrLhRJRwPN/3JqdyXGnIacMD1QatAaxR6UlJcVrHD8mjHJB3xUKU26Ahq0aOp/c
CQlXQrHT2D10UFjueGoYu9cFtezkp25ou2KuqAvWKNEPIat4aKL3ASMUEw2U12tWZIAGnXtoLtZI
sDS+0s4ZSWMnlN8baTTzeG6zMaC8qXPPGrgD4QinraLCkIDjdEYLic9SoPLZbBqkevGUVrlFhu/4
4MYhV3RRC2cIJ1/IKNnPH7BRBuLa0Ef55HaOFSJkEuJghIJgNJWT48A1Ab3nYj7wDaQrdR6KGRSc
rrPTm9sTYu0R5R5sLsz291DJ4S+0UmW1sHSPO9r/SM8wgyQ2TeD4vYoIVFbq6tEUMozWJfcThw+5
6SIFKrqLeo1VdAmS9NfhbWwVfWMIB9fEAAmKsmal6kaIO0eiVJmeQ8T4EH5QgwFxFYJd+LWnsMNJ
h0bH1rTE/bjU0qbia7u345bChQ9ebIANq6YK7btqafThBoZH6npaT/wUhtSERrvrQEtkARd7q6vo
K5y7dgUcNm2kNcKKQ7w0l5mA6IXw9Zb3GQqSw6HVZVYUnRKurKJwr9zGY/HqiWNNBhDeNoLebrcO
iNkHXmGLOiz2QiAxQnzSR5uvlOKCDVWuH35J9EON9TB98Yr7qgTyxa/OycpEbIMJvGs/hc86NjFF
omHS+/Zin77Ik6VBL7G1W6ThO+gZIvCCdF3drnJmwFedo4qRunXKje9Q5mZki0ht6ytucOfZ78sw
i5Dw0HF95z5sEzNPg6iBJW/w/8F3+Z1akHztGlBqawM6WRF39I+E/88nle3fLhkti7y3eUAHeiQ5
13lrqfQAUhYyyxGW3fAp2ZgYJ7p2ALQtDdoT6kiA5iUbrkQwpMKb25WWHkcfuRkEErrlxG9W7NOS
mMwjcIC69c5UWr/xvIWVf9r3NzATDIwZtUgXKMGXkBi8ERxr/q+sYjqLE1XH2aXmYJsFb4dZywkN
HmW2OAIlxQ7SQTbZf2oyH4XbDAYHwS6TD8FOuemqcBsIagM9Z3fSw+zcFPHXGVtE1NuQyBRwZgx0
/TRdA/0sTLuM2RLI9QLVgcT646TFe3Z1xpuDnHwHKqv9/NJOuj6RMqWemoUrmHzoMTYc96+3tC50
yB1PsT24WVAzGKgNPY+DUdcdt84WoJ7XeDooYMzYpx0JUzwFChDpMRrIJROKpnE2WdSFryS+qCfW
rBpbpSTDI4vRzQi+z0BIvAIyyZ0oo5S1blkOAWLZ/oix/ShmjwsJJqMfFb6n1HSBSjNLBxpK/CpL
cMW2RpCleyePsYTk1HRib2gQxTTiHHJ685i2YAD9GYuhEMHsOhWg/1yTE1+SoCiYPS3fSDVHsBhv
WQYjPvjxGcQ3v8xkXqXuQFjag06DTzHIhf315YI3QkifVk5bP9Qc37Q+bFcB1KNqFy2nU8FBXelT
uUXZ8SKsAcP+mPdN6qR6xiUROshernZphmlvwru/enige4zTHYM+NwdIAU08fECHSKxDVqD1Wo+V
zpleao7h2XELEamxXUNqWNO7yTSeLHgE99NWscqFJxdyG5X/QxjWDNXKaMRF8uUa/ESWabVqTB5v
j+N6EQKL7nqLjfhI6+2XaTNJyGo+rnhoACZdRcYMvLUqFauAjcLmQ1n3jx8F62iyLyqlPSUPiRPf
dHg9Xj0y8l99IQff86YmVwUB7+RIhM4Yq+Uthopf6AD3VAa+9wzMOATJ2bg2Klmii6zJJ0CJN6q9
f8p8YCbgyF5eldqBQsKBO8JPeidku3ebY7i/lrz0PSBn5V5uMG2pJ/RiNZEy1BiNIHwYe3Kwe4qE
tp4jsdeKr0hPbMXNqx4yy0sipG9zN6uyxLTEIkuJ+aLuGYFs2taEo64taXvY4T10fpcRq5XMoiDy
hSeQfp3ruIpUEFlf/NhIoepUieQQGrv021MXeuH7yUVgBEZ4V8W4MhNb7YrjON0qjtNMZglF1zkC
C8UmAv1SPfFzEiRPzaDqphtN/s0Uj07IXFbKx2lDJ37mtlGjxlwWljw9PcSEcGgGg0mfI4LsK6cw
cfjxIJDr/Uy4+dRS7R/qni9wW+/bFLAbg+ROI/dgeidBnzuvhv/l7v1lTzVU6kax0WRCmVL0z6cT
Vny2j6XHhJ6UNxhDK8iy7Bl4XDb2lkEw8K3//ZKukb3t/EqAtasRDpH+p3YldaqC5EJFQgTcBJBu
mD63gogvnDplTnuduDRCHBND9w9SjqHnyR6ZAubAqKlH9VDiR3XCn1/aOC1hPDLblEYXwinXQNil
/1EXFTpN/kUIbsUKprdO3dDIC+eeUuphRXdDz/ruUK3vOyTDyFjkZQyZnuGhpZRmxRNh1ZqfhyDf
nB+bb0TnVslSvAzhONN97IMzKQhGaDDf+f3zxSWrL6RmOL+wnZUMS3WQL7i8qBdCPuGfiXtx73Sl
T3F/1cVfoSF3EDf0MvWjVYmVSLSGqG6c8JO3lrZ9IlldU3KGBeASEg0w8hLb/fRBF7CoEkDAu8Q3
+IDAD+rto9m6nieyy8lx42SVizOSOwb+9r2bxKdQey+hKgbXAYqwMZ30Efae3C9I8qdTG8bhUTzn
r7Qf9ZYBWIJdDJ7gi+6iNpXFhDawVrK478wdutyg6zxspLM0Ih6plsfdLSpBmX853I63IgqlugFI
xSPPiSEgjnYBu+hwkw47RS/qQAiTqLH585XTaEHXfR1VJCIDfr0O0QEN7IKwQgYW/73YRRP3Ztug
lI4ylxuWJrXCzSZlsJqnnWiX78gaiP7wIu1lDgN64mrfzFdfEiFAn9GdwcBOCh9YgUfQYuPU/vC3
zhZeEXI9dRYaB481/Om2988wIr/FcHpIdnwqsWZMeTb6oY+60BkZGXMNTHBJNXfuFbZgeP8x1d76
PZh7Gpp1apoYX1oPEtRuymzWKp29bKBpKJW/mKlfJQKC4i9i6w4Tun+9ZN0V0BMRdLuBgtzkyo84
faZqBnKyjx7FtPba6oFqJHVIGIC7xkQeceWbt1vyEIOPTlkKs6t9L7jvGGrT8z1cOm7wzg9bojqZ
fzrh/DbV49DngMv6zZEjSxdU0EE9h9oxawr+fUdvmQgJi9oToWROfcdZs4/p5cg8ZDAiUsuJWWhU
bmA+++vWS3ezn0WeGJPTiI5/gA0bukVZZDySLPngLZbX32F5N1sI47iwQefQy0wrL0SSW+kPbf3Y
6085vi2aNPQCaMksyH3V6FEctnF56X9TRxTDoZzyPCYFd2U1FIBoqGhdDes/JU25MpX0TKWuUdFy
VuFAhd/GMxv4vGNjUrwpPtaLc4HbVAErg20I0GdL3vFmEyz6+DmJOkl/fbWKNlaQBPfZfy69jiB4
ZfPq5PMKEh9rekaGn4KFcXyasFJPiP6jWDvEoRDAxDzkKw/gnX43D8iRo0Q6kwuJpeleCJLY4Uw3
Ew7iLGLZLa2QK2bQx16kmDIxeUhfUj54SYTU58OHc1gfDHI3fqBbXa4mzgCmR8Bg05PpVRcZOsiA
HDUckhMCx929wHb8tBMFrhtNuzC8vPkCwFB3zLuLxcwNWe13gvGfUVklndsxArpX3PPmpmxYUdE6
RbOaQPfPoGSIShI5L9dU10s5bTstvqxAHnTwfcRyhdMNQsXnC/zW21SuDCs0g2Dxh0zmRUIacM1O
MhY//Ms/ILNvbVp2UgPm2JS5d1oS2Rv+GC+RRv32qKfu0okFtNAVuXeZxlh+USrTWarppebFjNKB
iVtcbZXfz4nQTuFv+Y8fpu/CZMw4K9+tbf564Fcp5i8eJPHlxZLF8NsFMW63JSHwgMp+OLMd+VQM
3+iYUB522pGmVFjFLU+w8pnoI9mwhzvIz0P2kHiL/BgKClsCJ01e8HC9hazwIgbL1Mc0rfQD1cJt
9iwVqt01ihynlCrjtxbgSGQCW47+6VGHngQKQb6k9ONWpu+aR1/xdx0vp3d7jm26Oj1bMHJ89tiJ
wc7Pxpxx+pKeXP43atmEYygZGcC2VizEpRmB2qSEVCtwKQ2MLz51I2cHacSBCplr3y4P0mYNEabl
/XCdL5PMJPRqKYiwItQHCjEDPQAOSvY5/LhRCGjVMZu0s0JMQ/bIhhw2aiOUW+UY6FK3UOTPmLF8
b9O49L4qthR29hTcJBwIl24TTz+WX9/mHct6XT/VF/OFyGDwdZSy2ub3AUljQJVdFW2aptGZ5kkA
egzLwFvNdGEIvZiZBXVpaJYOo7tY1P5YO5XaHREn89Owb7lwkKx2noYDRg6s8FqZlGKakpgzrWUj
y/wNRax0MIW61yUzGEpzqouAYyIMcDNsntxXd7ncUrQI6JxIGvNHHXRxaNkqB0YzfcBtR5vTTwS8
YCjmo3n0JxA/YaWLdiww3yxPa1b8QwZEWPwUvmRMLpSwglcLjMXiJyz+N8N0LwlkO80qtIcSBvKC
yfmr2LtMPht0hMgV5S/z7d42MU9lnVCxjLcnLns8irR4j0qCK/tlvRQQHjLK6wZeqAaenmG3sP0N
qkyJ1tm2sGFxmD81BBTeDY4bF+3WqHLll3JRGsuVPAfIlj35psPQcVTQ9cOIkN9LG9zvbrW0q7Vk
fL5R6oFT26vt5P3Xro76sAJvgAOZ98eSPXFMWC2CpAdtT8VL7hHIMPhcpV2IjspN7ZElQopk/C91
Emuxpr2mHI/SWtSlbWlYWjwf35csGdMMgCH4t9TLJsEq6T+vLpiabScc/LcTEzFGU257O1wGnWPd
840SNIYx/zaJI9cjYHJIdvurGY1ICRWeYD3KkBb7rKXDXz2H5KJedNd4R65Dd6mUm0bSibS51kH7
aImBiRnaacZ+emaSvJmymyTHe2gxrCwFl2tL7n6/DQq08Q0+NixaN6iLcuCLxsWI5Zj4rtljwkFC
Ow4ioQKizCUw0Szg3pjgErGLl9EPLTA9fOD9rRSqN9KL1vjUhiuSXxAmAtfey9qreHXx+okWLpHe
FN4ygFYcQea2LWC8OBzCRk8P6vtEbg1y4JVAceP+g9KQQAtTwNIGdD84RmLfHM65JqRdbZZ051Gc
+dr4+AtjNzAsVApzESqeHPH73ApqAEJzsQQeW8tdDZl68QEuB6i5t94S5zE7RgMOQrH4KsTfzElK
eB9vIfwmJlnawVndIfG/KKAHtqwOs0XmJ9xdzoZzlaVcdexWrq3kiZxQZqfOKRxyMZFEAh4caJ0s
nzMteH9Q0jD3PtsxFAQvS7hqgj7qbmlGJw9nN0zhvmzojQBy8kEXKgZemU/k1NzWwyVavLp2U2an
eRIb16kUy/bZoqbhQwOTRkGpsfulGCpGyuVPMuSRXpjm0v/fHfEj3H+XRzaV0dcGEkduUdHv6Vvi
bHJpkQ7OikHVDTU6d3RcynEuRgSIovoFq39mzk4cUbjNZ/RcKojiEYKR7IU0XR4UmJOCUDheW5Of
KRoxGPNS1n0n90mH4+mKiZlGh6HuS9DnAkUQRybJr4c5hUQdWBL1BztsE4hfTbLZcMvCjCFhPm/g
o6CMsf7PkI1C6utpOYznCK3ViZPiv3ERKXZWHFiNb/CyHbotDrXMRHCYdDK5gdszMLasv+e4ieKQ
BCrlAoLfjjb/ujKu24RDEGBMHlNi3ZHMZm4A/cSvan/ZhU7VCohbB/G4uceG5DEkHCqWrEbNVbWV
CLfqCAml8btquDVXLgk6Qzfl5EaFW0t8UIUR9EPn/gJFsUKNJqljA+n4FuMnFDmfZ7R3o1u19gqN
9DFyp769cLhGkoqULi/V5sdgwHrBkIETSbjO4vvKp6Up3EwXyZNN0q35dEKTaIqcFV/u+fqGyITo
bJ0/iAYNp2Yr5G/lSBsmX84H7Q/Gxl6AtCwM29z0ai749WPwG62Pj95oqbkw4o+uoonOjw5GZWF2
kOmHCIvkO22XkKTf3uJDILmLdrgPDnBwE/lqMueIkAI8DwSNpqY08bFCdCl+RPZmv54kcNKWWFyx
skwgITqeoJrZ8y/P9phbsPFBeHT+Plex+2JIwrAvTudlT8kGSSI7NQO6v53FFsCrDehEBECj+Qp+
nkudQYaJOmWKTvAQOomIYFNXW5jwVzAcHELkbr2afdcqy8k2vd+aK3locFN4BA6+GyI2SqqYWGhx
QjJhlVsz6HQUVOZub/jEf3/wmcoI3JIhQ2PfITiZVmo/TMZi97iFOyfAJxy2LlqJQ8LONvl7kg7M
UIHbBCX0+14Pb/iyM2HgHC0B1farkDfz3p3eOU9mgFU+xYLh36CdZHybKw44hPOr0rd7byUmY1lm
EaQj+tCrrN8AG83JsRs7Kd/aP6HmNkRRvwjawpbRyvH+hxX9xdY8Iv2VMG7U0HYl44b1Zx9F4Ocr
csSQx1IvO9s0jjqF9XtKWl7e51rFUO6oYbTt0cnDiVEjeL7zcwlcjhg5GVSAWTLZHOAfioazijyb
21HE9bchFgyb/LifduNS+0USuZfxs7SPM7jg0m8ObfFycFhVTEu9X88L5sA8K9S6pLrkQ03xDmzA
9A/FEz7J0xEYGkQECpglYddeqzAt3oztdAlCyqyRX5EtKtCropXp7C9104oESfVc0dGfAVBO03tt
25zJzHGyPmlPMJEYjkx313Gg2DC3NDUj6RHWCigNtDS6+av9i7UwrozoZICwVIPgWEWYE+9/Xtc/
6Ax5J46E/Pgv3JsNaGyx3Sh3OsRiq+/1O9vA8zw7Re6qWc937J9QZK9f9gJrTCc1MAZCeV146J4G
HGQmigCZQqUEnN/uLSLYILZ63wVf2931vgvoti+yvwxGwtWdQn4CX/c56BBLQfWETVG7iODP7c2a
kLNopT/zhPT1bBTVvzZ+3DbitWcvYB9KO3zdMMicQHb4QC+DueMLodQkuA7qE8jBknzNx+AsW6Cq
g/ODNI2LNDeqmDdnlm7GDk2YL8Waea1sv30H2hKHruQpJtoiwr5/ATVhGJsrYtAQU7699Zn/T80J
zNjcmUq15ZF4HtrXpG5lNpeJLSxQJiL3tMAKWr+umcR4KaLDex7bP9LeL0KEQXCxZ6oY8koHR/C7
67QlEFn45B7NVCt0rSsMCNSjXQnP6p6qpywfinFrwXJXN/O28pOSTIu4G9Ky663df4UwzysxWCRB
BepAVJ8vm94ybtxVJ3kTv0fHIfHn+yj+zlJhj7pDNBIz/1fGFIBcQAEIaitYUaeaRmdTzhMX5/WR
RiTR+F86R4O/Cq5Iki6gufUyYhpC5JGFutXQea69rKjpLUpjXDxRZ0TZMil3AhUhuGABfENZMkwp
/Gx8LSHDqo/rNo+UeCuZrlZqIU26T9m7yAMcBkT3Ne6Vyl4MSNNDHfGHffoP4NTvdhosxjgA8vg2
D21q8xYv0BzKCjz6kjrwduUsYaFEtWLjOsrcR3gmAnMW3Yvq9Mz3/9+5ZB5nYGcyVfUBfSZ2VEQ9
GfLwBCFGg++p45qY2M3TVhR0pGx9PLNv5XYk8A68qr5Dhor2mN/NIcWPhzVpffBWcm1yaFtMKLpj
jxtfvAL+huospqIalqaWjY8CvDEZzO6WDn0A1lvMCX6Ift3ITtFbClwyImHFdCkbzsUZIAyHnOJk
MALeI3bWXcTBaG2SuB69JF57qWwtiv1uUnlYXmDjj68m0QyCvrrUB4jYg4gDiMqOTL3G7EIeK66Z
EA+9QShQA1M5vksrs8OZsCj7KhPXA9fPpfZq0Lv7Sdi5tFc4frcv/NZj4POUXaqafEBaw7TIQejG
NQHE1sAycjEAQwLB9bjrR4QwdjJgK065d1ezuNTYp2cStVuW1UormWbmMdy0WeZTkblF21R4kb/M
dPpdPYKq03EHqkWcF4POaT8VjA6ztF48W/oIBqhH0iBRNwQlZXxCIWpa+qr8T+aulO/UDtgdNVn8
ufRSqwCpDhkdMkSviYLykUWvA/DK6PVfP3acCayaVgSrm1kJbyHlNx/dSQ7BCPfFMQiSTlxot9dP
1pJUGEEAgSZOkHnZ4Y7FLHeq6a9UGXMr+VRIWChgN4YJMwpYohDwRADEFb3uQeqCFOucKoPzW1KK
Dujc3R+9Kkq55AH0OR3yOsjvHMK2HIlGnxN+izfr7nPbOx4ilILrNvlRhqDv7L37nXIX/238yDPO
YECerT2QeagFPZnQtqfOge+YYeTiOq1Uw8EsBrsvEY39FLrC308t/F8Q+Y5f3Gp0Odr+aH87AsE/
tGnzadwiEzH4Rn5BO8fib2WkUScsno39Sq3err0tcSU8tivYQHv6xKXYxlcQ8qyZpJS93Xv1sj0L
i+6Ow5CWBxuzVJqQSSlCn7WPhEMk5kM53AmEqMDloGu/QolPqvwOOMxeDS6EWt3ivjcVb/NocalG
WIoFWlj/BxYFgxvKQJj1HNICcRLpAY7HwplzIxN9puacZ5PE560nmSnt5ccblsbgBEdp5IZwrgJn
/ATKXCZ/sUczmHdPgoqtsDK9eZ2+oxYK8Vf/Xl+Qd2gi5202Aa5xTQR7Zw/JTyu8XdUQA8ariAIZ
iIivsd4Fh6oYPHa90aJoBKPJyik863FQcJcMWZjgfUoMfcw3m++OeecLeaAXr19xmQYs7yh0T911
RVI/hOwW38REQimFfJEJy/DI+kNBjyoE5ygE2mU1ZX0Gs9/+G9XuAJPTgUlFGkCCe4vOMTJeLSgG
cKTLYM8tq/UJxuu8QMCvPmCXvPGJ/kKsTiOy7hZQ8A8+OxAJhi8LnQ8+OEksZdz1r665NEq5Mtd0
s6A1NUBcvqe5QRbsC//66JHNjaui5KxfxVMnjeUWt7uAegkB2OC+2JSpmqEChdOj9m2KAVby0mr/
C/+7TbQkbatgXLGVYRvelUubN5lSvIjeS+XfhYhY5pENmx/R9kIJZq5sXJScnr2rJaYNlqZ8EsB1
iFEV0duTVA+wOhLLUCl51JpgGowg1ZZvyd5zJTb3EqFvmNymL2cSU4RvYVelsURUjJx/Yzk1Z1DY
XTPu/zXH2R6HELpuiHJq3XwZbz+4LGWA2Xa3v2OlfzlEEeXmFNZx6CaY8mdITjPKnoT1GtZYwXyd
hckOHQ5MKAq54k1sHXMsI6e1JFa1EkliWeKZdvAAlQxdx0iUFtuCoKdJWSWz8TyM9swf68ERdrJn
gzyShF7Q2coZj2yY/qw9J5q1fh71TYVZ4wuirwmVz9KacGJbCK9xI9yY8ZFbRb8TeRwRrlXuzHVW
+5Zoqc6MOIrbQNz14WUldqeF7yqgSP8paUl38JqC+HdMG98pSjlZG39RQCavpYpBgCbORkC+Eu3I
bblJEF2KR+/L67dq5rvO/SFDuC7KHb4sKGtaCzFlEqmyXGIruXhxM0RFqcwYVua37+8ZZ+33C40P
2Nxw/Kw/8pqlZWnX5xFPX+0c8EC/Pd7wKoHGfNQBFPo+WNToOZo5LyIo+Wcw2UEqqQvaOrUB51tX
R2t28ecOON/zutUANEzQRdyH7w5MYxYjcK5gYBe7kmKfw83lsZN44OSVnBManIz02TkvE934NvOD
ERkKOJavf2FOZEOhxKaKobfj5SCoTxWMlPj7Kxwy1jkgM+XbK6x34mB3Cf1J6tHwDWIXqK0JAA2b
y1h0ZxZFkJfulIgbzAdF0+xjH7DWNODnij3NNVT0qQDPEhlOfcieqI1tQZ0entLHn7QNr4hFqpx+
aRwlGI946WAezdoSPhim+xsCLEYaEP3R6EVE1MXRBT1IVXix/V6cz3oo10M7za2wqnzx0G/U51JP
U1UAMmM97lb93UuG1r5vCZwMBHr9JXJ+he3ohFELV34BmRejDA77ujFYZCcY2RAVxJuUYWNfwsZn
DHz3YvHzEju4QkRSUVTMOaH40Kj3sP4vOjBwn28cHZslh5Sp8EFt0l+cnX47XVi4thH9vwqc1H4c
JGREpEFBCrdbOmrsq+DlZs06pjXPQ3alrRqy8msWqdiwgva40iCLSrNE32DLfyLsZkbM8q76lcKj
hRAK2pVvlHsUJCShFQSLZnvvIlKaEVbMwpFBYL5ehivN6BAEq8Li4mIyrCCV22OF49u/skiMpIhy
E3lVocv1ET5oieYW7A4XSHtiqoM7ZFsxMUkM+oIEeFw5NH1wVYIJrFSJLNA2gnJRUcCykujlSq5Y
ko4TpRoTPOnjb3L/Bv0FVFNzT8QBnYzUAsJOaUCoSXXoeOr3khizWAhpHAWevZNI4YwGR9JIGuqU
uHT9HN90Knhc/m234uNFg6eoCk91Cb+1zkFuElcZF9gvNGGMgjxUyX3O9yQ8uWKC5kyWSsiDXond
eD7yq3RqokEJ9Piv//hIS31cw9iCOACzrxuLaATyhvrrVuQCdJ0YWzpJgsOraMqQidh1vNwviuLV
rh7YtcmKjvlMOtDh96wkKbMfs7tkrz2uCMcpcnnJznv9dVmcfkL/k64saBXUP2hHFg+ZcoY0Pzut
4s6j2VgblXLUOwh1c/2uZVLYhkD1lNH+XhzPKRY8G5T6d8K9nDOBeMnswtIEBfIN+07XplhKmR7I
U0gb6qq1eTN1tMY7eQFB0SVQShuKOL3Z3nbUd3DZD2uJKOrBMyH7uegpxLrP5GSBuvJxAluqV2jW
ticB5np8ASBEKSbpUOSwShnXfNyYCfZn4OGvJWJiHTEUk61vdiKC2CCaMF7wd4i7ZuuOYoy0sqeL
iJdXQO8u/JJ0fUekHvYwdKuUDwhaEDfnYxeDlG7b2NjEnI/RsCVdowe5XWUFfraObkXikazVAw67
Z2t1d1eijDVlgL9/yYG9ytjmOdP50ujnEj/J84IWjJoQ0EQUdmPMJydhxF5uuPMs5iaJbWaq0G6e
lkEdJSx8lUT7OH4YD8q69UyWx1qbNpGLR1pt9jrGHuiSzl1Uz3zk+LbQMUTH6X7YGM8A0aMwlDe6
rLIklEBAFxrC2VXTPcojJkAv6B0+PhSrNuLOrQF7hefrSMGOQQNVe4FDStCErtcj6NvEl0O4c/XU
sSkJDrwTwunLu/O4P+4akTHfEnSKTH2W2AyqVeh1PefQTO1EX4CY6XN1lJqnrBrnZy4p69ePs4Kq
Wfe6gIrupOEKkj2yaqtmegz4zi729dczksX/5FP1qdLezZYeQe3ncYaxkKtnpJBKfW8QG+TDV2EA
ucRkH36Q9bmklyRKj+vMvJqjBEGfAEOtbgVsX5EMjZijmKBWGGdZ+gjPfW+vGspq/PVbquP+TnO6
hDb5GUaCARxNoPyvpXDGXFb4wOAB1ATSfTedXJffqSLoe7F1K+rDWaUMgqZEf1AIIEqVVcISwRDd
svR7lAGVOfkpQQypr7DTdVuG0nxMcxtVviu/y4wWkW5f3PqeiKVvl1Tj4uBheIJCwcwEy+OrsEmq
N6V4F5rNhWPgG9INxAExIILubJ9nlbSg5e+VSNrfTYlj/64v9TaddLz406SZfs7eK3S8cfAp4CCI
+x7T4gUaDWF1hjEL8HkUdRhnRqhaJRYS5HHjX3s6jk+gsHy934xsp+Bj0MBx21lh9AKYWhINdfjn
rKmDchFwW5j1WiIjp5DEL5QVAnxdqIA2QEBeAcILA+GQsr3xKyVPpnGMFJ8eGWUJ1P4RlmGiYI56
CfJ9G1rK1l56puZavzZHF5T/1jNwRmmOrQnhNPIKXjNL3oVQC7Mv+tE3QnlhYizKb02n4YXgBfGj
qculyY8CvYgtTJlId6Utwb7sXdKn5LcTSrgU6BKxMqLPgxg9ZCYJ1Alr1F1jGw+uHPzvEv9V3xay
IlBCJ1xQrNVUsJkTGZCdUJ0nqWfgamhdJy0EHMBm495JEpZWrfesIBYa/5jTWykMGBatlxo8FxH0
qpbUQmJ+ar+gBeki6WC1A0KCWjVD4qr1k1VNHuYi+RMVqSyBdR3qndbjHlypqAERjdFZXFsBGGMa
ALmAJ+xa0rqaMgeQ5x35d2gDBLbzaldHjzP9Bbg7iTtkF/V1c/qxo611EY5tl9uyJ5zHAHBTf0pH
Q5dmWa9j7N64MQOYT1578sd7k+gsVyoe/FNAc/uudSUSto+CF3bRVJROpxAvuGigvs9JtQtwpoAp
TuDBgfXi5AUyjnFy2+VTbDQvnahSaLU9amP++W8oBV5vIhmUusw9NL5jqOCqG1wHs8le9H6l6B2a
4BsxkBeOyd57XoUYIfW0ki0cHt5NB+M6eNZGxSvUzPMaQz/rTZ4RsoNHG35JkNX3BUSx3GhzUV72
78mwzeb3t4mSr5igleAnADaY8ppCOxgkf+/quY1ye19m3PmKeldGep7roLcn5jMmTQkmbPT5y3b9
mbsO5F9EFQZXxsBygY4ftPN2A7hHs+5Qu+p7+R7DOkMk17aLQeGZfyKH57743k9uWy3PukTK5CMV
Q+465Y9y+FUkSEoDCugw+lgFPaXaFtDa5qcIjYwGTrKIRTcUTAKdMURVK4sAx+LiyN19lltHoxJY
LNkDJ/LD72x2gR+ufCJ7f76+Y1XSeQNXwzo10h+eHreaL6KQ2KbT6Z/GzhPsPlHe55/zqqplc5KZ
6ezFSc1U18KUvhXwYdCzqKHH3WFmK5HNW5lz77IXWuGcOrCruQsDXRnAJE+cT/WYxJy6dAwAerlU
OKDf/CjtTgSO5hzrekSaQqbhtOsqe14NaR8+62l2SqN0gzsdN6UdiJbCpizCvGy/JdUkpxR9bNiD
BsRLiC9PQjbVwT2kqc3/QiofTeIJFXKUsWH4o574Q9XSPnWAP2PM3sflTx6E5oYaZ5dtVjcKRJ9X
A+VQKyHF9Y5LEG5L0tFY+eXWBqW3cIQqkEn8rGGNv9hw4FLeNdC5fQxF75vCtnmX73tNgyRzNCof
jaYRtcGcUAto+crf3sb6A2Z85xPEvCUuvzAmCcR21NnWv1sX7o1hEg9mvQLMLhLYUjVm6o94z1V/
PvUbDqFiwIeFcb2t0FyHM1OOAYcyqUKKoSNOfhZ4jzJP93MKG9JM6pF5KBBOq6X9Vi1J987I8/FO
nMsV+wDVITjIB17H6q64wjSjHPHZlMOF3B6ourTp5Nuqu6AwmpXWGkkEK7Tpyjbdd3e46SihvZyd
HfXIrmlxuBznBOhlTaFfPNAXXmqJybAZ8NPJJthSFajpXI24CFGYyqeAGsHSCIO74YoRntO4QzCj
dfvJ1rUIWmq2mGajuRG+gzlOjKNtPfYTTVg4yJ4wUmYiXqWoa/VGdqL3+FkAKGlBHwj3M8J83SiM
P2Po5iOBKkATlEu9db4Eg9UNgHk2AHVKOhSgcLZuERnCVsVvsutIaU8ijJ/WiIdke1CvQT+FUh+k
PsglBC2lThyVyAo8E6BXu5G8QUHBXo19UZu4IcYiYRysgXHenHMGQvVoZ2Oe10GtmZN6jOlu7c7r
3qpUTCkx26C0z2S7LPG+5lL/koIp1cY9MekFxO9FhcA6c9VaL9IbnN8+e9IBo8/QIl7jlcy0YQ6P
azmVISUWOzfq8uMviIjp+86Lr+5dGGWH+JAgioHP1Owd/RvSCVdYtzgooS6zi+yeYcofbrwMXLuX
jPdt66RsuyFIp+teAEDrvw7inGv5ZReGWpQF3tDAHOmS6pLi/oVK1t+A1yrOI6jwMK6rSnbU6ixL
E1Wv8VxGWFHacxOvBO1ecVtXIOKjuULK1+vt6FulcaYqj0PJZNblXJ6Rf82QbKKpvH28J3f9tFJt
zfDvFPfpeGN8Ui9A6w0w6B1IFZ+8Z/DJO8ZvIcYzY+n/DukUo0anZecb120i6TttOKpey8GJP7sJ
bD7akrF6czQRdhOsyT+NPLq4vyljEJh4AWffd8maOqOoaXCSYhqOR0yoVS2yQTC4/Xg/jNdLK2Uo
dQupPmryGmyUYwDLls/qhRd7R5/VAuw/OnXMSj7NZJ5UNw3uqLvmBf20kEajY9RxVlkCAwvHwcV1
fD9RK2bXi7uoY3rXV0ek5iticlf11tjx1aIpRkclGVkp8J7ixwMsU2ZiqhHaRx8trczezgC55Hzf
xGC4OUtLxu4ECWcLa5CHqELhxfsolAc374wQrxKiAx2sy0yOYH93Q94REsDyQ7WC4Zpauy4CRSmL
NloLlU18Xtiker9qgCjIxLGX6z/5s5xmaFhjKt+S5df9/JN2p70QcD2/iXfLhOkbH9jCK3pVmxCV
xxTez2KgFhOSks/iEhnyMn7AjAbefm9sCfLwK5B5nrJxrwtduU+OukTv1gFmjePVqhdHxxgceMny
zbiV34xZMNhUnbFGpokfosydjZDJRLpKqHpsd/TgbH9fsv2SYdWYXwE6JtEEY/jSKiHqC5FQwL3I
m4Y/ojNIhX93LFu8Ip5PaPIB5Sn2m47rluUGxqWwsw1I/hs/LOiM4yOApi0BcQLZUzhkedOjTFBy
RTmg9sH+kS5KqA4m3nmTZPR/H1hjuXNy7TNROL/RHq4vbbvYONiHNgpIi3Fptr5dB+InxiqBjfBG
EoTCZIwL4cSh04PH9ZqEUNhlr4FSOvlut5CL0TiX1pot5U8e1ELN9CO5bsEF+1oI3Bo3gxDgyLfK
Le+2T++sxDG2nRGmEpTRhsvUstQhupXOoxAC+mMuEffjOD4HPoY603CO5VrOapB7GNcGDK96JjUl
nRX06dKQ+Pc37bbBhyLYw/7/hrrTD8Ba7YNS6LbUo7D+TFlgMESOTp3+zNFCZIKvJef67W+uT2Yh
ygsuTK474YIqFbgDuGmsd5E1Nv5NyXp8mNBHAQhebGMFpHSN8ZNB6XGIZxnM1KdCIZ5n1Aw8Y+nZ
CejR2kJrcXPoHSScFOplxrrIo1T90TTazkM+cORmo44d+ysvge2kCvJM4ZSIzgD2a/0WIfrBm5Xk
2SWvZC4z77u87tiq1egWG9jEbjqzqsiYiXiRJ6vUTzEfnK1Wh8F0AUiUEM7Gy+Pr0JlYEEy9VIH9
vxKaKFbksg5Qs3BctG1zPQE4Isqk0uxsXDwWirorQjwWHp2EGghY2qoOX/X2NlryTyY1b0uO/yLZ
VO8gIbJ2rjj35s1iBYYS0923NpqJK/nBxVHqvKyxaliFBS7kPSsq8dtCRD30FoMBpe001MHLk+fD
8jY3n1DycSmweAO3Qi7I/m89tfgmOdMs6otrfNub/joeFLgn5PqdEc+wyzM7m2+V/sVAhDLdwASP
pXWtwOf8HpwHEZ2V/TjzpxS4/t4vLwQ6vWqgBH3ACSa81Z6PgKtQMpQ6K9xOAquYrR2oXNFd8F8/
s94jOUgtmm0E1ZCRiTJzuUwG21tNWP7m97qWMe/OkCNM/TuJlvUT89jIpwnJ9nJvOvl6KN+TTrLa
1M9Axt4wqumSq/ONkBEn4UWxVrDAI2x+UpjbrFlJMUHmHZf+urrKSHtVjB2uRO25yrWNwTAJM1QF
TtqBsft76bHbrqzz/7pAAuU2oEoGiekVqkRzTBVbdXYbiw0MtX9GzShLoJ6+ftfDu6j3FJKWu/yV
5kpKCbYMxaPvvNnumf9YqC/rrHVcGgL8WcG/xWZojSVjfhh5Rbo7gdYT1IVb0w2kjbfBPX/TpRMs
ooDSJUjUOw4RVQHNo1NZBYDpWd9+2NWjet9EBzn8tZTU5UBjZakeXn3bWETo4W7jyE0D7lL8Ww3B
s8ZQaHjcNUorERxXmlkrFOkofLqnE0+R7fTjz1O/JmAshB6A6bkES3KKmcEONwdv3//rucxJ8Qyx
F8frgphccfknLhyvUww7bYKn91ENECFJ5M2TF7xl3yZ1I6CIc287PBoQA8Sc4KTd19MfdElWIQr6
d6Vf+D7PV7fLRv3NTTwL9LfjvG24EhW8qDCHtpROlV7IQNb/EsnM28MBf+Dl2WLu/rGxpIyVw4gi
aSckNbqZoJzmpZZ2mnfq7zA3TqbcoFxttiva42Mk1qrTMJ1EGrUuGje4m0LNGrVqjDmLViuwOhtZ
m1+TeYi3XNmhnlr5h1zcWzrUdOZSlahkvMyyVq1IBRR08vJT2uHbqzOQAcmNxtlXFKrG++QDDVAX
arZzlhMRsRJDBu2397iQ/JimCfEppO32oB8iwAmAZXPqlFuPPC+MIGWTuUgEM5RxU9zEk/CKhbLo
8Ozzp5mZPAYQiMmZn2/SsGiMSqJqUcQ82pb3g/LNKj60S7ya3sVvxQA03dPMR9SzOryAQfAKPwEa
/xQZjjmvDAyB86CjEVCKi4LSJrFRvamD5SGZ4k7kjKNyGk1wMzGKl94s7lojdpi2XjhaQJ6eNYlB
JQwyseEPzIxz+fs5QJUVxapWlf8rABJQXDfdBMlRBY6NxX1y7f0frZqvGa9yoAM06hrlFEYHHZGE
a4Qa8O8PpGHAg5ciKMJL7ICxmyE1eGlyDQBQXxhDdQiybqCQwgkb80RpRQH1tqkMwEb+d+FvQlpW
+p8FDDPR/gExjpOKRC5czL9w53MqucaCXX06jIOepCG1TyEzZ2NVD5voUseAeILZnjBBp+FmXlSW
nv7ZkwYMqw6xjs/8B2BxTdtXBoFem12N98uRNK44nUy9dQyZnb1aVLrJhtq7LNcPJPDvbyMOUc0d
VqLuCUvOOQsBdkxVho+k8tdGz4rbmLpKLJ3A6PmZuXV9+OC1CKvh2KUykg68aPoWJg8IsZX3PC3j
F+u2TK1ynKLJY7c8TTk+qMEnPB6SvtBc75zB6c4EizM/FJUHf5cFnYo8TsbYUuPf9QkY1rzWAKh/
gW2N6aFMBsP7/6CFENzrVh26uJ8I2LEj7E+XBPsXIzCmlbPMyXlSzaPt5kin4+ib9o195oAoBS2q
Uttf022dO087J0G0y+m9+OVJZX9jmrUOs3i/571W4vfW6GbQGGZj6J+MsfwY2u0Wl3IoarqTs1H2
cWpgYrF3xiivhgchDqpNvxudjplXat3b39nx0HbDcc+glM2TCFxPOkDqld617JpP4hk5Srxr7VEJ
8BhP2oJZJGJjwWXaX/3NPRIo6oQRcH6RIHhp0qRygyZ9wpqRu5Ll1DnZgqh6B8b2HBsXune3zAjJ
6FPS59eKREx6A5LNnacs15YgQ4huFeNq8+oGJRX2Z0G6sM0IOtYLO2B1HglR0O/LA6YkP/FWLzib
HiyGz48bPA0TY2vmY+qLROYJXlqVvEGkWh2jPvH1T0QsHvJdwpTKCLnj0MrJMxF9r23pQRL9mTvV
8o5SuhNWYQdiRtl9okFbdYUfiqtOaJ9LT6YLjQB7GLnwlqOzTmnXO4zs23JG1MM7FbaZRgOtm7lW
8kEWktSoomoxpwrWUwaomLIPdm6ky6PxGiFTQKQ93IbKF995hUoU1tL6fSJ+4m6cktieCDud8cp8
CgDLgmyqJVZvReO4fE51CDZ78PPJbRgEGbSN8eio/b8ATli8h33fYXuCL1jMl39Hl+DTWEq197lW
4MN5RPSPzU2Tz3mhKoyqbiyCeQaDp/7P9mVaDSLkQR4BhIiSUUL9SpO7HfkjU7KF1sTmpMMM413m
1R9SLBmKmKvEvEr9sCeei0PQyC/ie7Po3ZQ4HaSBj73vpQit/2SSCELwcj+FpIPxHCv1tH42vhp4
FfhL8R7NqR5COXK0WS6pr5ytcWwfLU+I6QaqHZKTENG5h5M12gZoBBMEtTMImzwY/6hgZkJTjucm
zCTd4vLpGYZe1ykMyi2qs9v3ZYBThia/W8ki9740c+TqxCFWONy0PaWqAFjDCIAZYmyImvcpl2z4
qT20iC24cDzJhFYfvJOlFXOObCba7ltC/o0OEp6ELwBAHC9SCj5ymut/g24GTvXp+NBbcZxCShpv
bx+STgzdTCZcZWWYfRtCXwi5oHxX9FMMZVmetuQyNuKBfHOdkhi1oubDvgeOK2aK/XI8sTGcpLpD
MbMq7qyzuLqUfQJqy3bILGZZ5HL4E9nvjKjcZUzQbsIE7EZN42zhvRUO1aQRwOS2ZXEf/x827zkl
h8k44EMnJxG2b3wO3FDrPb/tpinG/kKBSXniMW+87FPfcCfm0cSuLdB7bLzKy3q3VGEqN+0iBDpz
RDbFpD+BHRs4M6cod6fXBYdIPcD3mx7aPSQC56fYqQAt9yEnUSzRTuDFX89O2jc05nap6phg8boK
rpsW8vds5J4Y+xCAEyovuHoHGC0gJa0xrKKl1IRgJalptFBK7UivkZRyrc5rhSPPi3TV2VJrmRvA
QnYdMfQQetlnlsOZsT7xTMOmJl2jSjtlMZEgiq1Al0OY4TWTXNsnPD3tSek/poycRdipJbipv7SE
i4J8ozeRlaA7F/qNlGJOy9c6OEVtGk2EGArRMsDdubH3tGvpt94rGHeBs4qhNT03qlzxjBATqL/p
RrmDGMANvLvb/lS3AZFOJJm7vAR3ahH4Vsla05tobmUF31AfSIUAXfMaxVxs+hQYYBa2aZHGhZEE
EWyXJLLTkuRaysyehLczFBwAZDHXxnxuYE/eOBPSvi8yKdpGP9Yq4BBBhnUtsfc1lL6XSQihDRjD
B0pZoAI+3PwICKlbi5bLKZX5RuFcUeQXLFTGN0AbGAFcTvqEFVbgfW5PR7K44L7JPnc9OugT6Bim
hhi0eR9uh1/zaz+7YfLBRoGK7+xcTrgk65L+5nwCyiov8cE45Su3WKFO0OgNYPxdUKMo8ya0oABb
VdOwqxZjC0tOIAcEJjC2li1YkPpMofzj+l1S7KyEunmXh3RRwBYfoUOnW7lbEOmVhWl9tIvJ5Ojs
MbKmFhwlEsX/6/XxC7QhPKhi3t20EjXxTY4m6FHErslziC4ykeAj/JYBfe9nIGuCHdkA1JExTUX3
7wEFsgrv24GAgcHhOVhEO12ynDz0RradSKtKhSRpSDdD2u2wNGGLBl470T5FWuAF60BMANV9TxFK
OJbgz36YK1qN3xPKcUKGz/ZoQgIfWR/95gu2lm/XczyLqsqyX/c3kMWGSW3sZ7QWD+knQpytplzd
M7LI8fozuBhcgYRWwYZpXe4PZZSY+UOhaa9T7K4/RCf/Wb3Dvy5idGVYxxR3NNR5XWTeVbGYBAmf
cAM/eVbdPL+DQrg4cDBgEyGHXrvEZBk+MH1xtFVDuxWYhqugs1RNywmwLZSo/3u/sRFb1/E6qsdk
OQ0TtweQMQ0TIZCXRl6R8iysHP34oeigMBbAiuHLt+25AF0cRF3vg/apJXFQdpqKYzqhojnHmdJO
j9rNDofKW1Z9vzYe6sxckHq9VE+JOJ+0FrIihyucOvCzwjwKNY4TUvi8p5uHEuHDhmAnoTCrSuc0
zV8kNIVXOTojRe7/7O2ht8FK+7H7KCoDcNNpj0woNe4vpXdLCMNdLm6P8/2JOSIKNFPcutxn8VWc
p+A+l2usJOiBGhE6l2RQ9OLFBuI3AXGP/+1WpNfGbWUb3fK5vpPW6ts4py/01ckfsDTl7seRy4Ux
dyd7A1/duSqm3QEydOP46SYGbB+koYX5Sld9USLEZZubBDPF8wPZffVj8zMHZPNIC/tUuH0e3MHX
WZsYd8HKl/1Biym2foLySKdGJI6hzVvGJ9QGWf1SxLznL6Pdr4T9vuejiaHyiaTBfiaFYXg0ExYf
msWDK2WDGuoLObmJIcyVzh07WHp/QnTCp76UxnFu8wehDoIxTYdKLVUl3ga++wHIl5HoS6u5DMy5
38hd/d7mU4bQTnWLdsTbs1jxAKb9w+7f6uNcbsYCvsU7YE+JOJhPne4QfgfUB+bzeSpwGPqAvnm+
PObtHCVfIhar3wY0LBHxvvTgUdHHoeAkU9E2xk8ZvyJlYiS512NZJ+JxggLpy95L2XvwBu1iB/jV
Q8HGqFE9A9fZHRl2/DWfhAy6W1FsvWj6lWMxnYr5NZqEeyt6rrVGUZavOl89LlU342LIybHFJu8b
SUhKghz3kxoDDwo+0lCBdByzahzS6LZrMVbS3w4L5jWvFwe7CAEj5CZRDnIYYBbrLacY/9QAxiWv
bRxZ8uOf+gXn+k80VHJvfQPSacx9vWrSUh2VNTlhX7XzVT2393Yx27rxhR9VMiOzyKrvcX8h9FGR
MHO78BImt4zZPpoPqcB3DlcNisa018tk11PScFS0l1c8vDaWxrNhsj+rRvDbMBxps7Oa0qX/QARH
q3iZz4A+WERRRknGS0te3DwWVQ22xm5B47+u/0h5oyoW+YLlrvbfzg7J6+LZ0FiJce4pdJ2WE+wk
zN3Wy6yegIAmfT8KR2MJp5AZpgGYy9yGP3fuyw5lJWGw4Ag+JYxhUHnugw3MWVa9X3v/Xzy0if9/
OvzR2Ga0Rqh6cFQg9+eegaheDIxCiW+y9+G1/mGEuH++Lq0kF6q8mkUcld5/KRpAMye5pEFWDT/f
ksI3ACj3E1uJ4OMMrTiuFUPHVbS/xku7sljId2bH3ZIxFLALw2b69invnPGaZWbbuBu8MK0jZZJo
W9KBLYlgpr9G8RwVBWipC6p1/1++lA4ksmJnxkAdnQ+oKvD+V49qkL2wqyYq3W/HOPvK/D1tCCAi
he3fE1hwCVexdn42IRpoLXgCqRJ1VLUxBT/65dnivsgDqCp/VpNxmCzgo2lmT3fvwptKSvpqo/qX
2UVZNypw5InUSB0D7zM5TVI/lF+A7CHhCQMqBc5CirQciKHjkkv5EsrFajc8tXw446ECDuqb/FW9
KYfILayBeHrG64ay/Ku26idRDszPebERJAoxQ7E7H0Jl8KU1ZCu9+Yj01bjcORucO9F1n8utf95w
O88/BZ2PiR1JlfwLiSUV7tvW8Lh2uV59CmgCIsjDp4K+UuRQ0ttjpsnrEdqZl+J3IRSEaPA7qyUY
Oz1gDGn0UX30kLxCR+KOyVxzdUo4M2Sa2xqUonSj/QZqMezZjECHbP8F7dTojfWiLHfnqyUnZ1nz
HKybJ+OI0mhgAevcjhvJuHAx3/hxrREVKQqNgnhQ9XlhoDOvFP/lDtzdOrY1esTh8/WEqzvwz/vd
HeM/qwGXob6WmBMNtaFogMJyDvz++brax1IHl74kWLAWOH8il7Gv2jy725dlc1zo0u3k7sdXcUUK
ZqRl/6UgSwzgoM0YNDnMUQwwgnbVKdvKekmAMFfOn64ZV/yL5dz/x7orbu8rdHs4K5q8/W0YVYoV
j5l6HaGiR3p+y9KWkJjZF7k6ePeTXDO9FcI4ekO3018guPEd5t+9FAheZn+tugfNoCEmO0rlHyzz
C1hGjnomXywTmL/+YBVRuLlDhTVLiqAHsQE95hCG5Q5Bge87YUiVh0T45zPTekXCwZUfV6bNIfia
ZnlR8kURzS9jXWWyiA5KnO9DSQnVSiDYrCL7FleHGP50cv3wfobswVCZZqWh1cG8huKt74gCwon5
UQMUaJySyee/Ry0keUVCURItvJ0sfYGtJ41TBwGjgiePDbeYawA4s2o3z6/1yoW27QN25cJOz19J
qDajSezkvjsnRZOijiHzrFDQinehNUN8n7fQKcmAjtXrAQKlBYwRB+drscskoIeFrGaQvlpSr7Fx
go3wwr+cqa11oRGcJGUzorVyZZaQbiFAgo9DHX2VduDf0EFser7OS4Qv3EHKLt2IwPgdg3UETZXr
4vOSVmHDdcFjTFNJZL95YrgV6QZyDBUSemTiDPO4aOW/mIlaNiHDsfnlilHK6MGS0/BTTam1/m2h
+1Gl/EJuoCn2lTtx6SGogF70Ngs8oy+igPUZt3wCdBzwcj4vEcyHryv1v5LCSWdNBGQO0nf9k14G
TIiEY0aHAD+UkLwKN7KdamgnlpEwjTA2/XpFDuk8z8L+BQA+wLdM7ePcyVl7An8RkzpleXcbYP0v
BLtEx7Ev5DdqabrW1g+rgSzoDgcbkDME+rOoH4scNMY8LRw5EFgnxDgAbAm11xBAl4IxZlprgk10
YmdYUpr/dVLb/zlDOePwOD2Nu6f7GnbZUoSNc/f5kbhQANZcjTIcK+Zb0HaNVQPhjTmpYmwKxmRZ
ZMqMHo1iaE07pyrPDOodEdbFaKaW53Xzqqu+pVijXAtA69g+mZAp0qfk0WowX4Z9BhK4H22dIn70
JlXLIy6wRLz/HbYjSY9s6aOahi7i27SYUoHAqSjALiCOHJpZos5xicP4foy4DuV7GBl4zOv77UMw
ZyHeAaqdr90sewXm56f+AxOL4hMyINWjs/CXVp2qYVCUPqA5cmfIbFBL6LP7wPXqw8kb9uxJabeA
A9kNoEIM7PB0Vd2zdHUsQlUql4sfFXq5ExrZdh5Yj6Je3FqHR0EeZTdAfm4q8yQoOf9faULdI1Ej
LSJuZT6r+LEy8uHG3vmr4QQ9KLcYyKkHA/3Da0vR490l44ISpBF22u6K1RjM0TaSMLEQVjm397BB
Wy3GOqb93EvAP9gkfokNfR0/ibrtCqE2NFxs9dWEhPl7K9naSxEUhR2HMHCMrz/6thJgf610qp5z
GXLMC0UPYnrQTjL2iMI+mWN5LZFKQ02kgFdGEYIZdnmWcPq1V/P0sZp6ScR5QOXP3qXa77a1UMT1
vpa6TIZ38ATetqekfvHUQQRwJyIa9lyXZhvWkrv7EiKiP8dr6NpXUcKzq0qle/sz2F5oYUcCRTGX
3lar9mIahm/li2aIwZhxz1n8BqQ8qDXWK7moCuobghoZOJ8Cs/KOkILHkS9Cz29lUE2TieXzoBGb
MRKPiu+iPeoSEGLkDyd/V+jyA7nKjTcrhCplIPMulJ5lEgJXoRwfk8aAgU4DLa8SwXTZ8gS61ItK
W3jVNWKtBMb1uNnX0o4WQCDz1jjazXfIGYdZmQDv5TePRl1ddfL+arV2o2qTHD5TMPPwemCzUcd4
x1Y0OlxBzZvev82CQEQvmxnRrQ8dJlzeOUViiVbSn4R2LhrtAVI68OtcGCJdtfZgp4n9UnpFoA1Z
qMnj5+EN5+Q1pvL+PXQZ6hRs+WJKMurHdUyXaJtRts0HVhOV6oleZeJtcq9MTRW5kTwIXG7hq3Q4
6d/0JNf4bpa5Y622H+mgZzc3cZ/IWeQl3Gh7kWrCpL4Yr8J4Xg4hMUN4xAifWp1/qkvM252eZH5e
glFH+Bi/wRw81Q1XGLCE/Xg2i+joKwJi1BXrBfrGIGB7uaJzH41E3nIrQQfnaOnSKeJ3X06JOG8w
PclVQiVUD2B6VCqpoWpfiWFnX763WZVObT3jIIcBAuO6vRAaLXCSyGR0w2PiM6S49gqr+pKRtPxj
+H+1QtdGsLCBzmdqJKCKH8Er7f58LIz5YrbbfIXVG/BaNM0CX+vl9CNM30SH6ffVbrNq31EUT8iB
8EL1RBNY3cJNlu7haAI6sywmORH3lnIm57Rl+o6YwKzerWVWEYFg/td2poXycCYuKltcYNp+sMiM
R+2X/7RBSMyEAATjc69D1gDIuG7vH9QCYG3OYQ2HY1xaqnG1TBSleEKTIQy4uZTU3PHNrwtLpmSF
PtSCpNrwvmWR7wCBmGz8CSmBbr/Q3USzySmGcNmRkOzPGxxM80b2oDVvjwKhB/cfda9zv/AtaH3P
R+D2RHtnRUcsULTtjFCmWzsxUzbzmlKTw7EljlRURX/F6unTgn8nde9VKQvRao9vSShQiN2vL4gO
iGPiY43ZcwGHPCT1jRUByEhwcSm/ev7Z3mKNwiVAjdZnN0oqiFnQbLMnvftPZoGR8r8rJ4OxjBMr
ZJ4Z+3DGnRXQf3B3DDNFcDdbu0becfRP+d4cxAzthQ65uiAM5hKsvb2LIRiZfzwP4FrSDzEfoq4K
YPHih0IE2Z5gOdTbDg2AWFVPBcSBiFS0T07lLKWIQcFVW99ZYorX15dieJwsZ3tzK0TBm8FzMmsJ
a62jjMlxoDe1VjpvhQvDo3AuUYpsjOp4rgokxclv4aAfo5DPKkptAtaLgEpzdtqO/vlI3qeNDY1U
kd8QgNpTaNSCQOKebjQSOdfa8pxKicl3Rya95+MFLV8AaRj8kFdQFMueVCyVUSr9EdXKli90iZvW
A9SbIvJu4X1YXMbjDM8rNuCf5mCHlPZ3Kudcwn14R1tFNH8gNY4qDPixJPmPLA77jA/ubEtLHhw9
maDFJmu2F2QMyrnnFWbvpBLyJ89uRqR9lB1+bcug+7A354gFR4t+s6L3RXp086sO3d53YVGlWqTp
bEZ+0tFHub4AIgBPqzGC0HqBsyjRLrU5Kep8ZNv9lhtjV3TCBtmDhsIq4ssMhJmhFMT9NcIGoxc/
9smn2ScdPCObAdfIY8kQitPWEsaa+pPNo/laXCbW4BaKdWyH+/dXViuQN7dhj36SLzIjDG+hpZvF
NNmqp9evHUh9nOQd9KRNNzshlgMJrgW9Uu1zHUCn7SUBN5fJ/7pzKLEoegSSy3u3nBTLjvwKjjnz
/taWo++zQQx6Et8JHRh9n1zzLgxopJ9F6a+xoTygzzLhfUxwO3JJ+9NVKTcGFLAk6wKfr2mK+ryt
0LrsGOKQCjtqY+a/qG5+9MxnTkwRlW390lXZjCWbDzBbQI+PadaWZi3Q4mkVR8b3KSOQVYA8RyJQ
WJAno2qzodB8svu/de6JZ3n/bgubrhewrF8Mz/Tv/vB2Xcr28c3TfRTbvjMrcAN+bPlCoIE9BcUd
X7eUbHEcwNCJaKBXQCajqjdkGMyLju8Xxc/knXjLVKh/EYyLwKmulBdHhxNjK+EYbbBwkRGqpuvb
pxjThypDvy0P6NTK8xqZSDmYMk2Ku1AWKY8nPkTF3cf7926PJQ3UV64wsFpCIavJxuIEpJSmxRDK
WKQSMkI0GfwxwyyA/stBRoP84HJGICVqkfV8eB6FeOx1vXzX+f1uhn2Tt6xAwe76RnljpD4UFnYn
Gd0NEQAf5uCMOHE1E1ZkCuqUAWWkidh45lEke0CQPM3WOPTayXOoksweLVqeip+G8FLJ1ZhIIYPS
ROFmBBUYPJASVTvoHB6n/nqMx9mFtZzdbR8HhAwQiZj9r3mw23iZc0mOckmEkZkXfAhcUVgBTGvO
b2YQC2wgi2QSQAsyA9DSmcyKqzNxwwlq9gbwIRDVFTPeN8Fb63SovhOEB6X0csV+ZC00jyI218Es
yG8cy++pOwrGD7IRle0mK2dkk7hYqh97eOLCnviP4UXjISrYPfF1vPjxfRgWaGO9RdGb6XHtrGzp
5tlqSDxMWq6kkqTZUe7lJdKlXjyOVVhHTpauTv7ljBZV20984O1m2xQLxqnmHJIlFOoDWpbnIf6p
/hFFOEAdl6JPyJF153B7tjnBuOKniWdx1Xo57Udz1WiwHW8aVh+wN52ukbLnTFK626O80E2J3m2P
cDJTwYc1XgV4EjCfE3wpjTvuizFoAoMNfv4T82exmEiDMApjiLQivktebWrzCxpVcJC6qhGhJJTI
qLPedHa5sfEP/mf+OTKAn2K9F3o81AUfAD+tRTmTgEYPibZ96ufnsmHqkHvEJJQjAbs7mTDM//dY
eR7EfN94wvIGhoPWZdoWQp9bX1SlESsurP7eOjm17qya7uV8v9xMCnNpdgIBfM1VfXBiJf7Q6O4T
/cjcFkY2QVelE0nQ3M3jYp0H0s6wNCNUzs/0ewJ5CAyHetGuPgb4kxqgJpr30tE2loM5DQ+uaQjB
xbnO0XV8g0t73Lp589Ot6GjzmUleEqvXtQ5BMxVbQN1k90cjr6H2bL/0RxsU11QvfsEC+cpIzeBu
uYc/M7KApXnJWx/9l14F6lkUX1AfT7v1/GRl7NUbziSrhNmaHeP/aNe0tRIZxc9sxh0SCTzfpXzs
NrG/FmY/cpM4EM4ZLvAqzRVrbvdElp+Vrim8xMwDgiZQR2jB0MICO02kmOkgZNyjf5Oeo9/f9JKY
lKef8rwe8XaRoKQZYU4iuWpZskAH73Sqchsvv1sa8BWYPwiKJ+fCEjwpFW7rWUFMC+oMYIAI4y7d
a355WXZvKdWhBxbxiU51694yr+YtYU3zPKno83UsbdStjzh1Ncoky9EwROo+nmBPJz87pNwHPs88
2Pkzy6X38YH6QBj5RtvCv8sGh3FCSueuHnLbJeXooxuYKFXtej5bvZkQQtRxwveVmMQpsbW/4+ex
Puc2V8sG64HeILsFyvXS0/WzOxqqyyGCSNRAr3pk/93p9rk0kkTJZaP1f+TCpRBf+tGMmTvtZlMe
o74CKPla4YRWaHQ2GNQC+ArhW+d01/X5pZAAI58maVV0Qz1GJPOzjOeWz4ZUbgpSAlL48+bRXkDV
JUKt9fWieBOfajMZUqqrvlM43vHR7+pP21qhOZQYvVTZiMtZP1oN6nvpP+98/k8O2ceFgFOviB5+
L4m/M4s6wxA3Mb0COrRaAr086H9jPPe+L3ACymoYMVfHR4asKcMI2IGYUDxNR+aamw6M9MhpYp5c
a0jYUg7nPlmJpTI5LSEEJQpkJDghzfjID8MmZ/xolIiNQSsKJiKoYMjLngBzdmJ9owjoBlaoKc9N
KS5qZIS2G9lABoIMwWDRT3FwWDuuVwpzAh2ScMTJ0M3dX7/UsbU6xD1WA6ZwPZFCqqamh/+jnr0S
N/r4EXIbs4XA9dKf0VAC9zjLb6z2sUgHd44lY554E/7l1AEI4GDiWRNMeYsrCZldunJUMPVQq2YN
AClxgEnMj1G4ye313Lgn6sAcHN9xVSMa6HEqZv3NsMqhGJwkRb/eHJqtNOd7S9psZdaSMLu0JnYp
vYQwctAIlW3lL0Bm7Yv6KPK+Noewup8VLZOfdwQvmA4jUcU2UmEcG6W9vjMc9xr8IPI7xfziOK1z
9UI8j1REiVPSnQcYfNBa7z+xxUIzFWkPlOi1Osxz4iFlZpJUXfDkQuTZnjcK6FyAQsbKnNMHVqUT
SLisKqes4vFKMeE0UbtuztHCqakgShis5y8Ew1SyEDAU1jQKIEECvjvXNyjfgxaixPjdVGvTzZsC
ER5GoNQlwdHEdGytqiNTNjxOUXpVrzQMADdtvs/8YqJ68DhIvFcCPRkI0I9Q7+jwvCb25YDno9fG
UXhMcfGdKQWn3G9ioHIrDYXO44alz30hz3KmxhD5jdxBFIWcbLUW3YDV7FZNDmdJqA/pciRMcysN
iuJ2cWgzeloUFPYvdR6lXjbZ6Td6Q5cLIAhYRt5Y7Hlc5KHtH9xquFziuJxFg0JnDrJdQ7QMrG8S
xnbZ3xBc6znAMCv63LIwZumAc9KtQ41HDUmM/z4BdXloI92wY+0k7pr4Hb5JHO9bKgcEh9mapzt/
9uJRPKkPTfKLCwgO8CWw9+Bznl66mX1IWNklafaWYyr2CcCsDAk5m0nsqfs/SoUDjODHyqdo277u
ZtfPLDE1Qv3FBWwLuBXC28ETx8EOKvSN5Guvt10DQD5TqJyTII1rwoQZh+8bDEZLyx1M1IVEtXfy
+EPv9bQRlPOjE9EmVVghXFan9N6Rx67agghTmK1WEKMPosZo2EkA2/4oWHlbZG2N4y/UWz+2iRg9
tPTJM2GzNSbnlyPS8Rv0vpuZnB3dqTzapBmIrOriClxzxKoIMtzzIP5JcHD1R+IyEOVTxcM/VN9J
n3Rmnh8Y8rBJ/mG6yehYgR/WlMNWy/oZBRGy0CaW/Gcpkdx8cJF4yqsq9rYsY35UwqaDv6m07HrD
hyIYjK0OqiSS9xrN7fEWQKKVRb7woCc+iVtsfhsjhf4qJ2DKEVO0Uk5DJPXABkO2mkEUFKdajF8H
/hvEGaXTRLcdoRRu5p5clgL52wFq4OxBlhzCpw6u9QJAGM3w9xmayAX3ykV6lBBAdQdjnG4syBNa
lUKXYYkRH8cn2AJvxyevijg34UNP/3UdS9BITqfBMpRvCjrCH8eGKfvn1iaPMA1ylBElzFav4iUt
WS+Wf87kqEd2EeUeIlMwpWi/74QZi6LYaIZWbD1DHLl6chN87f6GVYORI+mJcLJ4PJaXBo7gifIu
h1Y0ei9DxFjt7rIgwaE0qYaxbv20qUU/WvPTRF08vpSel5jcThZ388gcd8fCumooHtrk3jPg101T
jd8xH27/VDiz+AI9UgA37kBKapiI8VUz39kPWDWlDNw+9AqabEpKfxfnO1D7BXpMnlTUFyRJ7l7m
Xz0mbJRWNEHm5HFjWpYkPku+oyaUw1yaRNZpy6IJGF2K612/M9SYjHSGBFayPSh26cnqUxS/kLJZ
vY3THMrzxPAWuBU+BcKtUsiO0lYkv1Fzj2ZDcMh27tWDXqQYlpZzmW12qiLcxjWKnuXQlCAU6+mo
FImXgCXf3pGbySGlRSzKec07OFTfeisPlIi4WaDywDCbAbnN2+d2uGu89bKqgwP7OIFZH18ZnZ9c
g91sWkOT5DaO3ikY0a2pzzfADXJYx3D4w4OY1Ilfa7baqpQi9JqnkGr3Tp8sxrbvGgVIDWCbGqgQ
CLfT4bkG0OaGzQGiAlrCw298Reu4Jv/Xzljm+5m7sobAFi04U2PWD0b8zn3kvppWFZAoaxHkb0F6
GMQn50RCml1r51NFjtOFl+XbHP4fB3WE7YXmykI5BzP1j0XTdgAgDj6ljsfRsjcEljl35yhi5Lhx
XKmo3AVpezYL3henWFDciq2VYt/5tsvCTsA3SXMcxGZkMPN+MPybltGAONEANpOk9RXcDVQuNfQR
gu0cE40o2hkZ76+j6FveooK7n2ed1b5xgZxgb9nr67nfU3MRCORXrgOBZxtS63DBqeJqq+3fY+yl
/UFpoDM7Wtm4zUtksad///dDtrDkEFmFvciVY7e7qhX7qFsPxfKBkToLz0IeUZe+1hD+sBsLOUzV
ZLpxYqP+Niwum1lYxTLdw7sRxjd3Dulk9vXBqpwlcpcSie0DHrLYSqmaHgEe4nvgQccTKu6Hfbee
e4djf0JnX/y0/HkoQMz41j/peaKs1PKB99Ut4kwfUQ/1cobYDrsFxGnomy3HMha3/xpR5RS70K9R
lrVjkuS6gzySX8TNLnkls0NoxLJRXtvE3k5dAUEqngSbNWeDBAzvaAl5JQFlMw8QS0lUooQwJeS/
VpXXTRrDij+uZDbB1xiC5t7M6GB7lU/zeY5lbog6E7yA/xf9QGxxIXvtz/IvFpCpsRlj5TabRLdw
07GgipDhRC/q52PrQlNt2NY5+YMU538J7t9VxGw1MQfzD84sa0Oc2imPzkqLgQITPmDapWQvT6/q
2ZYjoqw/9hVpOai0tm6iT2H9ynXYsvkxTjpU37v9kuhuQ4il42tRMKhPF5f1xme+gNyXCEmklzVm
aYJd2Pi5R4JJyOYfvOdOurvqWc8tBelqhUiZu1Hv4G1RKAgWWi/dtirrXYnZqIDLA6UZttoI+nvY
fU4Ohz4j7/xLm9WVskqtPzJoed5WDfanqbMMelEOjTnsYvHnaMC6veFgkdztP7EUdtmr++mEXNzG
4WXcO9e83xXDP0bNQmZjk9Y4ZXNGzPwo7do+tk0LBijH+lm2IzZ6i94sWY0fQ+IyfBaXjx7Oa7mf
Dhbv0veq8Ngp8JSV2Ksr78nESslm7x4Je7TL1xefaox01Q57wLdt+u5BsCTqf6wZkJYO7/IYl7pc
os8qUvGMTsuOjUEoVjLCc/9CBTdQshK8j432VEWwc5qygxo8ePOJfT1IDbRVOtaNWKuV5br6Ujo2
6rCW4TFCrdcK5V79C9da/vw2u0yN9sqh/vY4DVcrQ8afiyjE2KRUFJlAJ3sATcOLDMuMwaIAezBz
NBU6JTc0ghzM/xxiHpTiRFQOn4t/nVn7IYXvYNd89/o2CY+f8vTMylEgPqNG2eTKz/us8dPsVkHY
oTk8xHTOFjOY7Rs7gEu1VS07gd8yHONga43DZ4F7FOsi+y2nGaPM9fsRpn/XSrpiBD2U0GiFQgw6
pLdMOGxrxGfV1Ou4AfU2JBvU0fNFfWXTB74ZuLAZXwT3EAyP0NpTECBMgMsUxEzjicpqKutzTGkX
T8SlCwP4CEyVFxE78kLPwqJvdTQbx06y8jU71q67FEvR6fFhzqpfZOt/Je5kCosAxE5pBByD1pAw
d+gNrW69Vps1+D109f+yntHWWdUUu0m87BpCOKV+ziincUmIm/65+EBW874EwjzwE+MaSy05PUNU
acTsfdkABSLCB7WYsX7xXpHTgHtJfUBWTAmNb7AoDMomSvV/U7DeKpKeBHhZAGmn9ydmHFsTC5uo
eBG85agGWsicyQhESSBw3zXhaPts44ASnAt6rWn5WlzeOVr0f2Kz1tQwERfk5MXJfQ0/g8QSNlip
iHAw1n7gIzQAu+aGK+PvaOo0BdKo756bph61U1enDUcThIzamQzLxlUSGQOIQwegCrqCXNHfIc4J
619Q7Bf+C7JQyyrn4PPQoTNaGVu2UaB/pI2efZ5yTI51D24ZpvvtDkCyxqsUCzSVZzuioedTDLFZ
gufiNklD9hvc0BYIv1YgVMDFgccSrN1i+v3i5auS4pFLD2uSGhr3KiJMKq+GAEcfW/01OFGEffna
hrg2lVZNVQCn23m7YqD+3oemdV67Rnm077xlnm+d4P5EwfgtIzRRGRNvk3YZ+ZrWaE9bDvwdfiMP
8shqDOD5oH7udcS4a7QVvt1FN/QGOXYWqJVzIIT9r3R6sD1L4C0sWtFGC/wR1p27ggVF4obZCEO2
0rI03yE1WBh9sfm2sTHX8Z/xCCTMQaNqjke8cuFPjQjTzFjXrqclD0MTQnndQ53sTAkBTL9UMS2z
DN9hiKzDGwAhxaQX2Ah5iETJNb5/7zZD4dvVqle7r/P+3uH/+5bAt/gYp8sSE4tYfM2GUg7Otrr4
0pPBSWqC+U+1T8lpzXffcEnv0ud6/mk0B7MPlCe9rd0wIlX543pu7R/MbC5Sq7w1XL8maAs2ccQS
hdHAfXPZuaOL+xx9Urnvwxk+eP77wYhdPxqfw0yCMQu3T92DeOaW+GxxN8gPm9BsJIqcdAI3irDB
T/0GuFPok5Qh0SBSEgHabIzwUUhfbku+Rxdo9wjTRDGGZBszdcr5Cu3QKq8/HClhmHO9gZJ9I0Ey
7V15f5S5d0W+WL1Q3X8tmVKFubme/xmFRo6afzHI4BSIKfqreZF0oIsS6eTKMHyQfHSvBrfn2FK7
Tmwudk2XV4GLIFd48i9kKUK67i00UmT7RBub8ZeVtVOSKyjsFbfhbIzQZxMxEq3pelHn4MvR3VCJ
l4pzPbiSRJJCsmS/DlwXiRG0RpHax95ekCUyeRE9S6drTWQ7YotaxuoTms6XSY9G31lAwc2YL+7O
9Txq7EIb3bzoJR5geGMVcVkcbJMyJfFvycjvc3uD1/zHUw3+xVO4IdC9bkk6od7KFMJIJBSZYB7U
jpm4yCxJmK0Ru0VVYrfkuAHacJet78P4ogYst0JyN/tUNV4CyCbITd1qNRXXyE+XK7oYeiMobnjR
aqGueGSNpEsCuH0yaHyV+0yNoqhCo+JIiYc4s3YReAjY8qtAgvxxlSGAvJ21dQr/wxPEVy4HoJjE
yYzkdSkDvbB0HzwKANbLn0zd/rHubDvUlKqxzfV1zZu9DG2ORPF6qCMRWs/wNCKziS1SwjM0Ehqp
sXwtrXqziBK+a1/69gPvB/+Cp9cJ9wEaGWxHDseqbmcVoIoew3T/s59sCC1xJLKnhqy1Q6muJjEU
bnypta6GbKpQE6IObVRvyYny/8nYBpCU0kcjiqiCl8VolquaAQEjPKHbGSsDb0oibSSvyXE8pi/4
1XFcdmxNicm4nEbtHYuBG/W+RTlL2AMwGUxlHhy71MeqdyMGjfxJTucmIsrZfHnjnNtxDSAKqV8S
W/970u2Rm5QSkRkK9LOEGxtgdefThUDWUy+JNtvqqr2a+6PZ9J0YRZp6AMnXBFvxFLidZHR9giLB
uyyB6TWuQGRiAHDQWKNbR/FlHN/K6/30UU2wqvw0h3FJKVVPd5f+w1fUAIaWvoJX2cpkMt8z2G1i
r0ieAL//K+kssXTU27whvI6Cxde5GuFGUOqhky0bAQNxfTZM7yyk50WlgNK9RkYwg0nENpi2ptgf
xdwHCh8vffVJSMB/m8Ec6NzfibcfyJbAQ1tlZvFPfAEprIprOZhzJp+qEIesXCbCmjaOkR+Ok+vx
wgHbiVMwqWHfkqSidtcf7klw5mQ/wlZx3H/ANI0VseRnvP95IjMxqwTXZB73Kabx/UXOx843gFUo
hQfZzpiGPye3G5KRidOoCUr24l7KWYBVsJAL7YlaFoi9lWJo8CklA7BVY6c6huTUWhBlMd61Ez0h
p6Iq4tVhM+rOb38nrjnIwRM94Oq+Cpnh3DG4lxciyN6E+ZWKGVDcIN+WT+MO8NZUis5dNRVGpS6R
PJ1lFty95NEGNtlIsBnWUrbu3szvqJFwhY5i3vy57BUsSGvzeYBRuVknZp3x2ros/jOFc94fmFKv
QvaI7w+jdUqAF8Q5tHNNavSje+dD8YQV6+hwts6BFi58MW9/S1iEQlCNKeQdlo7vgGdSDB9bQytm
eIIl5OvYcY1Xgg9vXcOLN3tRsRCFCRSfM6Vtj+8EOWTw/8OgySlQz7W7ybKtqifdergi4HvPsqD3
NjyUsUEOLb+WWWpQcsDuEIKOa84PYCmYIlh9g6e06GBE/A5SqwrVFs8qIlZTOgVvhwmngManOms2
MMLWhoEJ3hUbxv4EiZe17dpUFlmRsgYM5Iz6CcqHOmSobd2y3PlAKAlSOmuJZLKkqkvUBAGXZU7P
uEcNSPfJQMAsHgoxTihLTmF9WOURLHUpeDBema8gIuBrE4oXDxjr7wyVlvnJqn7o7hrdpv8aZmW9
un8h/LRRd2z7roJggP5A20+90+rc3PvJ2nPSCXiSQKtIrVy78E5ZftLZDANcGFOK4yDmru1ywmnU
9kehKL7pqZmu8M7JzqxEj3/EEhnjoKZk69qdL1VLfpqBRM3GZVYfXJPp8pVJw6sBKPNg5Afle2Fb
fvmHPr1b2C48Nbid0SAOyL3l3CcKJcunUB0elohwnxcsnpAJVjidsCj1Fj7t25nwElrdhHoX9pE0
+gy8WDMsdQ4WJ2Y/M9h4F7uBr5TLA1yUE1HQzrA09pvrb7LQpyyGn8DdBkRkQf1d0EhjBePIb6r7
QF3oAtoG/DSfi+sQJdiohENyttThs4mrnwi1weIlgzv3rGsTCyHTA0DYhkfqmzUZWg2inNGlIkEJ
6vfyg6Dt2gOHH81I1XekwTd8tsQqnWrZ8K0mnDjLIRmKeNO83hiN9Eak/Vz9sQELoceEAL53ql38
HYsoZef0qZjG/EFSe3FWiq2xc10iemJ8UcyvqmIaPUA8r78ybKmnFoi/tNRh5CwttYOsGeqPegYU
GvorAVGqgCFzV1tiLlcKZt88t9N0FHWrK9KZyAZ1+vn80PClr8Y+qtcqwQDGKTKrdgwJKVJl4fw5
+0nvTQx9eHVU03O+quRs9i/7nNFtCcQEly79atVRHPE0PdNVaCrcWccxGAK21PFvte50PMSX57/k
8HNNFwZsA/UHMbXKF5htr+7C1hrsWh4Ua9oNRhpT3M4fa/L/4ZKMqnOmZHPkgZdNfWXk5++G8Y30
oWv7WzY07SOkQQ36Fg4D5sIVndKNSDNiODk48HcGf7Tx0kQJdvlciQdPAhirleWyAjCfIl6Kr0V/
pyWpSP/CCVFl5B2B0udPGtYgxcv2hCKNhAL6frw+OGd7gFkfFBLiJyb3xhYn00z4z4/7u2LILQxX
suupEZN1JbzkCltm0jFUfxdQmgQpblAEO2a0lwIp1BpkqjiFzo6GD+fuKt61G2N6uFa/Qj9mLdF0
1oXYflekm3UXdikKydTDkI49p4Y16zc7GUV31ukW/8Pwnn7sXs2AMaksX13TEsN0ZC4/qH8d9R4U
d8rATdiiBR6F8Ma8LpAQtOKbCx3i/BkXJCmI0uhWErI+7cg2lc23E4jh9KxR4K/IXUob/WPplCVK
IO06kW2oWU7gSeBROPRbarQ9GukvpUKAa4VDKm3Uez8pZZlFv14VYzlY4y4Ax944fzHo1vuQGZFN
ehRKAZhqrumBIzGTY/73ZcAjegCnqJ4K0TGpEKz230m6RKIGKdJHyFwew17A+5Ti3cLQXVdxYUI5
hW0NhhVLcu1fN8fY8S7t2tWxOyYM/JQL6EnU2uhP7tMazK/IgF9shI5hT0NceGb0hiIAK54diar+
dAs/WS/BP36Ev2tb9xUSmWaR7ey+nXKdASCbEfVGeaKYrkbcET5/ZvWmaJMZpjkvrCIfEfGVpu6H
E+t9JLUdCJXgv1iezr4cw/6ICT02ZsZ+61ntZInrcDmMaOnM2MZ5yGQaXnDmlRY7aFTWIVGiLcAy
KugxzSLWDWjQoIAaRRaDA2pmqMk/IceL3SqZdBtBipTRASRYzBj9m2cNeJymI6v56yuzOLWztVHE
8AobtWt8e2is+9U8dLWI3V2uSQE1zlqJWnVa59XOhPdhTSRa4nE3TuwJMFyozzN0GEX396wV1c5H
RhZDR6bXKELpqLwC4DxxWohvl9xVCffkWwWyA5om9koX/2W8hFaGeuGmXnKyczS+IR2C1ujnyiHh
XliqW9JmRNQkNm2/EBrmLTC49mf2QBNtP5thlxQpnktlMxGiwmVq7IPwZqySUzLLm0m5WE1LXeIV
J1/gE+NoNHjqqv8WuJR+lZLSiMuUSSkEpKiDpsjvR5R/JVDHu97sGabF14H1HwxAieW+z/yYpdgM
rPJ08rJjf2g7MsnI2dn/25w2gyFBURZkceYL9YvfGFUV5aI2k+dPd/SLu3dQWlLK/KgfPKvnaYu/
GTAsF463xlLRJDvcC1mYdaTNUtZLFKrAuHNAnn32RJBGkAJQ+9qbVMVJn5b8rZeRvmR+zTzKUGgY
BOpNX72Wmledjz8EbyrMFgwEW70aFVMujg+xOp4/yzVx23CxS/x3Deo+AWujAD3EwWGYsr8U8XHC
ALOga/7M/PIBVcuA4JyqUSC/150IyGHVkKQJ7SQCRIbYtzWfGA6rOnWUuTerOaUceX5XdxO2fV0N
LgRNRzjDr2PMoyE4FewR+xMZmea7VAb7IaHHpuBbICJRrceTMKqqfKZAh/5EJrAPnQ2Tsw3LQ6x0
fnA9antylC6ihAlS4VIUqIqToqNbH77XXeS4kOo8G140CtDQ6qLEnFfm9m61DdQ9G056PxlpDpKj
sYHFkcRpmqEn8UzlrLFNCpFREOY6o5mVWhWaHi5z8eOqO6iWmMeUFRrmT45ojtFe2rUrbOp6l+t6
+rc58+ptr/FO2jja60EmlpW6R2DzTOFCVO8osLvj4Z5dVuSAMG3U49YANGpl8Mdz3SckOJw6nInT
i1uLr0J0wNpAUPfQk3NzTxNU5wwvJ3dg34/CQPItv3RohXnWJcWYVSKIPjWda+j4EBVYAvzx+rV+
8UNylCaOKWtHWZD+oEzfno7vgf8Y6mFWuLMT4koxqvBXs8kNlJZXWDwMtSqFzwg3z+bKcHIlgvSu
jBy2vnsrWdTuwihP+j01D8pCAatRXSw5r8L0l8GD5M3ilEiuosuhwSAvP9NqgE+BO+JYDdnI8n4E
hkj5lTWFprml7tR5Njke27fZNwHOm6IFd4QG6MGriiS5ehHtyq+o06AOa88wsCG15pctaVdnhySU
vpYYb4euHgOUXA5gVld/17dTj9ScAFqp9JuRRR9p6TjWi5U2HalQmU4ynZ/4TzG8lvO0csIPjTgu
dETPmpzzM+4fd+U0fZVMX1ZLX1P6YgXbRb4pB+qBZPEEz3R8qcLsaCV/XAoSb0lfX8CmqXfuASpK
r6SuNkR5HRrbTrfjp2WDThNh+VbKeuemUPeZEeqi1lzJiNn5KwiqWB5OpenUWsfsqPgyMkLTJfAy
lIJnLT27VNMrwuM66Nj+hP24SDTk2QVcnTbPx4mJCiaOq6oHrXL16XP/NPLfjG3G0lYptVBDMm+6
e+IvmLkRjqzFD7GplVBZ/fO7+omzitusjwXSemBIHZDPSFVOEo62G0q31ekqDPHpdchGDgmGMKvK
/nz8ekMSqUofPAdqeQl+JWofsI2aZ1N21+OiZWuZv5Ae2i3Hb03Qo0FDtiQ/SLK2+AjMHgOj94AN
9++KQcCA9nxL4nz6TgYotLFHsZ0TBXu6rkAYlMj/xzhPzm6o6bqDvd1AcdPHhGQBJBhquHv168gH
L/IJTz9Pefs3+WF8Yqe7Af2m0YoNOdaOi9Rj1ZCgjsm3od74ZLeFfT/gyC7uVCmvIvNGQ/ThSAOx
QGBeOeyjo2/iO7nwwB1ASPqEsDK9z+QqQwGZXBWCtuBXzsZse0QHyGs0ZOCSelZsorLqbiLSxKRo
/wKoAGwzb+6dGPA8WZ1DpM6qp7kt9Hl6XwKEiML0P5d/5lfziUVyWuQUqn4hnRHjRj0ibA2wD+6H
Nu5TWj+c/yhZcYmPuKTDL3Yw8zd6yPyj1m6XkMekpAfI00jtSAofkFtJ/i8CTB/+Urh9akLIVA1Q
jtFvbPq9HtSO3wK8XOlyW/tPECGyR11a8OPy1cfCv6Uq4L59YhJ6ZZMntazsH7gq7Um2RiaVVERw
t1+jinNTkGYsaZQG6g3V0neN1lf0Dx82oYecWYqikfLwR5lO7Q15QY7P7bRRrgfUFDN5yhzeonQJ
iKnU7JA9fa+LgC8s9H6WKwDyapq7IHlsZHbnu5eWXv5AAKhWJv0T/WYeXqjptufmEMcS00dEePOC
3H9DxbGtnY78LMHAk0FuE4ZYxe1ccZxYunuzTejRzhTdZ4f9J05L3JqhaWZLzHOxx6DAXZZ1+KMj
Yhjfpl0zinUPFC6s5AbcS9IbsIHT8YgPr7F3KbuQo/gfDYFk+NSvsSKCTG5LdIDfRo2I8DdiDOF+
hT/VIcH9lDhP8a21gbt/R+LPjb+eajxtjlJXT89YIt03WhgIJKSgjnQn4OxJMFHTVMf73FPmOWLR
XLpz6YDjqDUZ5609F1tS3D5wNi1ESV/P780Ycgu9qcsNMMrV7Aef0r5oQ760ceox8ZicJ5acA+xR
97TmJrm6O1Em4hiUXkhzuWFcJpKYt05gx8vDH0K7Iil5on45h5oaFGEt7EWr38ZztKWl+/8+TLik
m+H9kcYF12mU1K6kdClh8qNjJs11F0RigO2OZcAoc1roihIUFVyAM+5SDuOFzoQS8S/vwpD/gbMQ
OsLdDTM3V3woz9kKkVr9GA/NZOrcIkgBxdjRrWSN/XQW6j0AgC1stjx1nZBU3gHFFbhk0IBzcrfD
cOQMqrRt0pL+VJ3uO5ay7I65pzKJmab50nMYNgghoNt95JUcF7aYLA5wFXKsdGt6tOgkDM7kb7dg
GLpK8BR6As6E+g4s0F8ixdRzxH7K2mvETr3jvQ1a7d4AHgcXLDGqOd3iynjvldYnT+JyX/pCCzAX
OGZZ6jDrzUVI7kXjclQYnE4haUIbiBhlk+LaW6chaagamq9jt5c9jrhoyvvI0RqZYelH9ab/UxaO
eqdjH23e2BX4eXunyfh2+S6fDBlxqBhSbs4x5RqZ16FFmRgJY+yfPRqkNhDGbL5nHUhjgxruxjrg
PWI1yfUj1kym33TdwT+XUuUpgUWxIsPHKFp44s4c6cAgHifUTxVLFHXr6HzWGBHIJyBGfW0uCnQn
cbjpMjNQBFxgt5IjuAytJUU4ontrqEXK+GXjvLwM2gnHQOhC0Ba6Q1BBycLwBMItdj90plbqyEZ+
HQFlCqNQSgyoOaUpsZ+lI/u8o3fSLIpFr/2SALHfi6fiiO37ZbXvLwcmui3qtiDokAxnu0wUIWEO
jK1golCI59DvsNDd0GSB2flegZN0vLm9tGeHBfAxbMgWm+/73ti5PBkiXuDRI6NLYomGH1+q9ZK1
OypPgosDY966Zjy6zVyvQWDVfD5nFMp7/q+Af7UH1Jz8CBaZB3Sn3jgXNqR4IzQmAjXl1h0XmJlE
dymfxSboKb4/XcABKDASdNl4xVjDNjq+Rq63LP9xg/CFiw0dg9dzKSQ2OHD4AOaEbIcfndxEr9uX
fi+36BqEkpHJgH8tE5Yyy1KAWZl4X7+k+r5T1MjZfcXIx1w2cDXa86WHAvnGWT3VCRvpCoaVjcXP
bdZ/FYHZkUx0uaZh3vEyhVUAQJcrAK/aIK8/NV48hbjq6grs2dnS3M2h5YDOXcoKcovBEj2RWq7l
zR1WsvMo6l41PTPr4na3OM203445gzrYX4v72MgBc9jJb1XNTvT48A2mPelcFe5cL27T/tx4ptAf
+D1lZnayXRVukNbGyk4b40QWCYwSN4EHRbENMBEZlpmJAb8n/KxrUxZOcFIVOBhF3P4bWcxoqbFv
zT9b6CHDUwY5nVhM6CZ3MmT1bK/PMiK6EzNoTYszt5LdWS+MwEk39I8mBa4p0oiYvFU009IpQV3l
ohR83jUsqx87soJ+U6LyKsZn4u3jIwRVplOLtWwNeZQqvykNdWnxExxgXhOe+8LmYRuQaOR07LSe
ef1XrvK0A6q2fhYbl7uVDxEBXFitd4brQRfinfx3hQ/9PgIeBLrueye83MfMAi81MaP5Yik2ydlC
TUZdQafuUeRMMDAfhM3GtRIz4olf3ozIutwd28QPeNel+5mSdWWlrMfKkjSJC/c281bQyPmfZsQ8
gqOp8b3E43WKC11xEyrujXbJzex1lBkL99gx6eWNvGttfqmmQFH3EOJQZ5BGYrnHRkx6hYyqgfsx
yMPnz3g/athZLR6KuC8LTkqZQthndObz5QE0lkTD2BnyGaxwZQhl8SpIFi5Vacswkqxh5WGpjgT4
pVuy4dS/Pz6mkqqQO7lwa+AcHuGKJyPD5b/SU8TQqAhScKFguZowHR8ltTMGoqnqL8vOyI/CCKov
y5EBeeQ+TIat/kPv7ykKc6WPKbW+6syjyg1Ek7f3xyNKGTLsdtozRrK14Ku2Q9iLbch1LV+RI/Uj
StD0ny9m3XJ45UrCcPe0lki+sA07Q5+6NLToeA+bYF2jhQ5F1B+nmSv0dHA10Ov7SEfiPhmigsHk
L7Tf7BP4lRcWX0BIBREXxv0826s/N5Yk6l+etPPD+urdJpVXc1UrCBZ0C7rIVGbyGB0COM9rYi58
dNPztRW9+5JwEm9kcEcHqBYyqSEFK3HjYIwnL7GErI0H7l6Hi7kbUQAFZ8c8KvOJfS3YMibyfq4S
BAkgOqC16G5HmWvPqK3yKlZCN4iFfRk2JpqGzezaf5QQom7VO1VzWhu6THAytu6zHGdIsPIzS3Xl
O7/zGVkYxBcruPiNxVrrKVNYu+miqlu9yMrSFojFYsmKnInm+4UeME1ZR1hr0jNCwlpiG2xHySAt
wcdEIExm4LrLtXttbucEoH8U9SXnpcExMn9E7wV73FEBgZ9FLu3Fz/htzD8dMJOeTktbbmJIp3xy
pRGPBL1AWaS2qgipQUrf0I2q3cBa9zUHXA9EdU0VcHBNWYsVpdYgsVCHBP2xJwcQsNDdm0kXHDt+
40Pv5sBhwL5CFnLx1e443evqoddalnDplQQV9QkNI42N7dsi5GaA5FcCYIyaTxV59N89jDmO0M0C
3evKpJ21gOr9/1mP64XoGFBsJLFE4x3i3uD+O4iAW2xsdH1SoFF8VWfbrBEMCzRvsQdNGsKBKS2q
A8eFwtLhOUZF59HN1JQKaAXpCV1/wN0UnzpUQTEjrN4JxMFjQbpR/rkWGzzi0OoLW5ti4j/A/BJZ
lU4UlPcFznYrvVGKwHgDCAOHsFiAsOdgvhWzVawCiNVr77BK0WUCjnPKYPsC5+MiJE7FP4VimbEB
uoT142XatW5jz8LyKd3cR77E5/vKQW+6C/XW8inOxe6JFuwtajOjBqts2KzGAdtmkePgmISTIqR3
NmV62OUhq4LUUdBdRt3x855AixBSG25bW60E1urDHxZ9NwpemoT+pw8C3vA1Hh7+L3aKy2RSy2pg
tHFb6D3nZa2rmy+7AOcmQK8Ty+pa6t5SDMdyp/MjPWqQ3+9Qg36nmA5nz+yL0IojDurPIgKdolq7
ik2UUSmyLyOziotAVMRDefAVlWfnWzFCPWP2o9qs2KGiQZfJ+3KBtlkdw83oMio6+2ZXtTok3QMp
9Sq61sIMEDsezwz4d4ik93xgTmao2v+xRofqKycIdhImeioLyD/h2pfS+bWFWTTmzVACcGXtxlKN
ieyy1V66OaJRGLlXwak/pl8m5yFPsFo3zpLgxc0enKnwAWsYyTbelUhGgHoAIthSqp1gFulUiu3Z
v5QCHEkSUxAe2AEyxAtMjEN/ZIx9YwUnPL2F/n2h84b/w4M728wBmc1Ls3nAVtjeYE94NBWjx5/N
UdyKd1DXHG8l82mz/C5eL0P3l+RJsOT0oIqPPmIkjIUSIDAjmZJepxKRi/CLxSQCeIOFbZkyUY9M
orHong7z7PoYGQnG/KK4yrjPak8YnX1gno8GYrIh4jb1Zs8nErATWT3S4NMR5NSlwYC8s3z4HJO9
1galqcIoOKaUk8bCXEbZyS156bsoMmpuFJ7O/vrHbrW+lenMMg9Xk3cQ3+lubwrO41w7p3DtVHH2
CbMm70yLNdVMCmjNV9PbaeMfKumOjTPYv7m3XgnjvGpZwGSUInkaMa4PXAgPJps4XlbuK08nPBY+
hY+R+LQ7x4uwZaMuw02iQvQCBm5fUw6pf/Frgp5Yi+eJEk2n9OEeeSZIl6iIHAxi/5bkkKIENovF
NZt6KAdoEG0fy5PAPZh4m9vcfb4vRjzoLvstjIrwCzXAPVOXZ9NwSrMFtPR0lFqOPKZXF1WROHQb
ckApxaSIA77/aBspzAv69L9nr6QHEPF0EknWeVBga2S6oj7tYw4/q1tZi6yMJeGdJFhXsRDf3mze
h+A0mWwVNDJNal/QR0T/6WPwFUokpIaJYjvKOLvSWRfcjB75mhwLNA930Dh8Od1Z9gtOQlfdCni5
s9cMTxAlPYxOkbtr2s3VDT7MnN6c1ayYndBgZUg8A59VpitsqhZ6YOz990t5sV70nT9JoWxRpIcV
eGB9mkOHHo7xv3ALtKviJBtREuAU5eRmXHHP//0IbT3HPRwtd3BqbIoGNZuh21cPjLO0vsobG5Z5
zTMOgZTeJYODH/ZyLnUwOzdfIyzf7IPVs627w7zjze0rgEzy8Ijl7be67TK9mpA927YOo72J+3VQ
NtgeYidQQY2VJy6RTqYxom1XU2rJJYxjFUTeVQ43R227A9AjBuylOnMgMmjA+JDWV95cUFkUzucU
ivgnhrJajSm7ixeHSRBrEbolC77LXJwIXTyK0gDqYMcgKCimrODmt8+sL9ebawSaUdMEbUR1Ttof
XAThclJg9lWYD9GJ24d6T/Zk5vtwFo4QAP/wEmP3KS9TayCpMc9vkT50AOJBYnf5wtIRtHbfhzBh
bOiwg0sLjPCNXOETw8n/zgW9v+YWnCoqKIldtw9X9kHGDbBz4bHO/PCgs9QRRAGvdFATP8w0wKYT
ZPfMNL5ZK56VNpmRoa9kXXA37X0ERfccZmMNdXAvd4IeJXUeAjT6gLChjyLbRQ1s+bp8Urs61/8m
nBvs4GUZ/DDtr3J7aBmf0jJ0EE1aKYf/APMKOTlVXrGtrw/OgSn4hgJzkIORRXDmRfswR2u71NQb
jbFUvdkrb+w+5hjXtkhyKPYlLHN3XErEQTRpIPwbPA6crOdf+PUb9t/b4Hy1qVZuuzn+aCGqm2CF
6J4pkjWhs5t2y6gsykI1MQ1b5M01wcmByTGyCjmWlOLkSoBjkUDLrZA0W+RvsU3b8V/aU8eUj/G8
q3irYgE3EVd6QCDno0/MOlZEtOjKwRTSkDUN+ONRzW8Gr9yKOJUxUplYpe0d2X7rzEkigTNUxR9c
glz+zPlhV0v+GmcQfe7Xk/Mxjfjdqt1NhO68lrPLh1gMcRgZcSvWxWAp2pK8hri3TLnhkJk1INyc
yyTR6Y3vuTaUsTT4+675n99N6+OvXp+MF/hWu/0B0ZzT3BdYM0XUPGO01KgAEGLt6e+prdHOeKUO
dY0XmNrzrIUFbrJLXiy2b2bpqWdWvYWFV1DHJBhGJGT/CYEmeXs6bSATPUKCiEBnc3qgybmx6UED
Bgap+bHVzNgrBSEAyVfcTUErxTRfOrbuKpBHUAm29qffdBwZJAHIl27DbKhLpDqpwIlhhbMW3xVA
iLMidtfZNkm7HpkhvyTb+c7X5tnVHm8udGH2p2vEb67EIsa2ckWX2g0/NKsB7MBy9hJdvOYAT0H4
1LYOsujHLtntqRk2sghbvgIDNZKGidysVPtGyC5npSqlbWdvbc8Q6qoKlBE84OULcyOsM0FGkuuc
zyTd4suzBiQF2ZjKUC1uSj4YaPhvzWiIAZp+4GOP8DAwtxrcIjGb6xxVPJ6UiBbHCspQh78ZD3ll
L0a5v6yRPnasPqcq66dY/o3JrnOIEljHMWCOxd6bXV4jwziSLJFc9PRqoiA+ez5n2rHB9SbQOnNu
LoyaazYAjXaRAQprnT0esRQUs6cowazL8GEJ6dFRxk1Zl65RHwcWi+O3FsAJLkDrsYTKCaQvqcUv
cuwdhBtmcqUYMmiLBgqWn1BwVzfEgBAssKCBjToBET38/ku07JcMgqwBiR3V3LiX0RrHpuWn7rfs
WYLrSdI8G74UFr888CBH51ptsNlhVQq62x/IBEekpdsS3DBeIM5/bbD5xILh7x+cmhXVyy3lmgfP
wJKVrAs3ntpNA0PuzzAxK+xSuJ50cehjgmuK6JWFwW3e1CtRtJWH9fttCkWN2ID4Zh/TtluVJJ0W
cRiHqvxxrR+5zIOEYFwLdTboPsHrdVkbSdwGy4ZFz5QO58pIDIbVzV6Sbn863STWn3Ht7098DzrB
HXa+BZHd1Lyht6oMc3K4JQ+StRlj5De7MySLQ0gvLWc3xoq8WsFYX7XAMUTGmRpjfoIJvG5gqL+k
7VaC+GuYF8DY4mUnxvUzuMHNcmfQRdT26sDJXiCqyGFR34aqCGrRkqz2t0cVCuhAfmJ+Z43ZzXxH
8nYnLJ+psy9WCRUZ/gw0cucKKLM9yjbxcVDsOXiERBwLCvkZTMEbDQoabsmObA0kpxvAeNrQUje+
kHRgMXL5Z8/iMMOKR64/iCcuwqLU5hm5MvKvA7WegAHp7zKffcmOnRwDtLx05XR8uV5u+mhyvdK0
bPRbQfUFE00ga27FSMM1s1HAm8uxjt1GauB+VOlURBmUnHV7oZwzrbYAHFCX9z/z3SIqfUg1ibRO
crKGhUzSEykSrxN4RI/brfW80piEWSzf0CjWgxGUXtqP6OmoSbhaVH+g3AJpv7BhxgXpkwDCl8mG
oq2rCMb/bct0RV/HJwt1MadgFWADhnKZNzIA5y9bORX0nkbUKVuNOoSNgnZqJkO1sufaCH9zDm3E
cW2saOADNRD5ooChxvGIYFKboFK5F83QeU3MLBR5j6+arHmsJ3rYt3wea434rfuqxkN2EpGeCdZ7
Enn/TaJ3r8c6zw54CSQHBtJ5BjrIWmDUeFXoaZTpybLaByOdIzYv6HOegWtFFTUCcGMNooA9ayuh
E+oQZAwnT3THgG0x6Pbrir7MGPgioYMe3QNvFWMHg5moq7WUonot8t3Wv/M+e3GdI/YoAvl04W9z
yWOzh4e/Rnaje9cE5drxTMkQDQbVpJzZ0FIuTqpz2/jzGBCYTPCmQVR3UMtnZDmL2+P+sWuhBACx
LkpPhyOgBnOaHb528A5gdTjrGSgoPN+xFZhdBcbNJKAdbPafDpzgpmxOGmHvcl2Plq3bLua1011N
3V6NOKrzDdQ34JhER6zhIrb22O32pthSs3NK3QS/qV4Vq4HCaloDEdPo56mYhQoNn8Nwh/LRv71b
z1QlN3EXKJ4HUutQXrf9pcPm9TupNGkvRwMU7EzO5kRxWzcShg1ol8qjcW9zu6KwTG1NjkY9P1lG
uzDq9hXekuUtduWY1hoPmZRyPTzlkakOE59fi1IehGyc2wvf8/JQWG7LRbMgG6EWlx+cMHizYt/l
LKA4m9zX+t2JrTeWUX2FyoeTq7ui7bMjMllyyKBjVcss2crSwHvKr2ZkyMC8qAvINvn1AsTBo/1j
FEs9rkog26gCQkz189SFNncWQmlhEXxiBR/FRvY6/iLHnIYJgQCUnt4s671Emc+xb/AbvwO3CPYw
4626UJlkPCaJ6Ih88e5pwFKl7HiPGxt36T+zqnzNDTjoB/LBRp42iCH7toXDoqRYizj1l5uCb0W6
8TAUYiIJXu/8AmQ1astgQZMK6r7r0l/8yuXJi3j9V/CQaJwzk4TK7GydfidF/oZ7PJ/YlAw430kX
iHB+BBS1ZvobTJmAQNuDRmWOnsRGhEuel4i+K5dldjSwQQ4deGYoQR6owEEAFeYsft51gRKv7ERN
0IQgp66Bd28w9Lk0IL/7WdfmEpVHBm+WYSq5n0ktn3IxH3AmzneXdN8BNOefdXQm4cQO3SNQjVA/
YxR7U/tSjt8cYnhVQCg0KfI3DIlNSe8wbQeN15uZemrC/pQY6uJ7yu6KgJHBFCHIgJqj6sLm4DQY
IMzWQ2R0/V4bUK2A9mPJBb9RvonmqZtrzWkdRu5kcvXDZTClqE3KfW+PacrMJXOh5cP9S7Vi4d0T
bJzXEFKC3Rs7isaV6PwZOL7nNwZcVzT3DiAb0mEC7nF0sTy9AP1aB3wbA6BE8KmDgqNPvpsjyJJw
jwtnOB0OUrBSGBkSjilPK5PLiLdg8g4TgCg8PDBySVLM5Cfl3eqefPjziq262O5r7Kqh01BNuW1n
+pwlupwaMZD3Nir9itTuAfKcWkekcGg492HoE4zzBNmGKjUbWqusJoscifeocZ9jh5P46aedI0b5
PFACX0kLzKGBcE0Nk6/99DmVqgxI13eA4brm4PKvOVBpOg2F/fB/u0tIy9deEpsigDBaxJ1cip+7
B00f7k3qcLWJQxkhMEwp4xNXeR7fkgpKKH+4a/6TExep9EVAtOZqm4qbjxq71ODXzsEglVdL9W/G
pYrWfZ7LNLuqDGXc3YenVsG+TYDTxeEE1OIPRvjgDJOIE2ghBPtTtlzEUHTFKdFGMxUKGy9tiN6P
GGYbZRFkdMyGB6HzhCzyaUmeyAMBxSKsJG+HzdkLtZYNWFUzmR0we3Lk5dQkEsZSG1ox4Zao4MBy
KFq7fMzA8XreMNU9azLBAxMNxXj5yGP/D2BxeLVpHVwsoagdJ6X+VWVWd5pVV4wtrtsmlxhNIwaA
pOTC+0OtYsgWCLSd056pRwJtmkhK7+j6etQHb+QGE5PJowvR2L9v91CrdgFJ8oY1t77yCjH2/h7S
bE6jbV0mpiqZO+HmdkFvtirjMrot7RgZrZuxZYGbOON4AzRks/5qiNJGvrMMGHxn7xJnAdusGOx/
53r2HpqLZz6GECAPo8CpD7ZyWFpCy9spr9zdDPQMxaneHLBtW8TxPA7GKVc5EMbhWFtvRu/38n59
td4YVy/m0RsVf/rMWPu6XNebkblEGRKOb0YPCR9QeGGRWmc6lQ9thGFluFciyUwpeuu0J8PtS0+f
w/AsgaQABacqYtdr7ITdiZPQokpdTRI2xdL8RRS0eqoYvwNaroKfo9kRAt3wOl8Upy9+5IH4VFgb
bDWogwNYoxc7UK4AZOhxHHsKjXGTyXevnKow11EZ+idUcRRm3ea1ujNTMrNC2L0kGfPCKHdCJ12G
pqKbzL8mW/3n4UJbiH+jBJhFQUgRAg7ASv9eF+6T4+KaTXoJAmAK9L6DCTT7Tm/wSRDUih/ngvGN
ip+xipdBgrh9H/VVId18nLP6cnIWrb4A9J6fuaTfp9shq/Tm+br0+ngrwu7FK+N1jqf3zs0y4Bkb
XIqtKQ63LNSGWh+eGzy2JIwcUvZujAE9d9SwZteJFgLmrdWXXy+Q+0Hkhs0/C+/tE3vrS2mfhm/o
csy9KqKS4V9m22xDsXv9dDtzxmTr0G38h/UoRjm5rFpWs1ppp/dO4OmKXbSGIAJopztJpNIfv80C
S9LVPIXcTB+zsLDp5n/aHb4kpY8yGyARDBFzHm8KIEnmf1MEtojVC69yBDHZA6G8rnrj+XkA+X9C
jE2jPuQyjJ+3o5th//nBZV3+2MVgImt2s48gkH6kz5h8UVy/iFvShcDzSQtgY6s4DJcP47wNh+Oj
TqSFkXy4mkEojL4WAr4+paYo/SE5kKDhlGODOsnVc9BaGjDGhLGHNMwHr8Rd8HL3AtvTK/aEJ2fc
qNypbBKY2iU7M1NxaljOv5M9BrRihmxteEnTfXNYFXbGVJI4Zf0+Ib77LbNMXAzPSOSZxjvYGhZU
D0L5uB8koYTFXjLfAXRpRdido38WHmWQ/R16Yod5Jcy1a1mfNRbr6g19nR15aOLGZ9q2ydO0X5fy
bay57U3e69oFgD92IxpvdSoRUUeNrqgzO0sw/RHaIahAbk3LwtSj4J0XwWeo2YzrzRY8kDAOsmxt
9Ym48wHn4dALUiOdJgzOAjyS2QBdOzGVzh2xR7XxCtdbgICJys4oJEWUabU7hWuu32O4Mc/rlvyb
uFzkMEUkWDZZlxkOE74WIkgiMEHoYj+XR9QgD+S0PlvKzBKmOxdkOu8O8uSixD3Atj4CY+J3Y7Hq
JuT5k4KcA53afrKQ4w+NwmpNQe72rnJMUR2Q9nhLfir0/2ax5+La6w5RqVRwozUvoEEC6QnT6aiK
1S30ee52erV+foKF9ppizgwKBZueFqDO/bJ709dAInVg8kBGInZoAUzj4ZHTaskIkTBSXT/VD5tu
6EO4j4Ow/qhrarm9eulx6SiVbNM/RRy/VHJ7rwNvq5/dLLcj3gnH+PciT+AOM8+f20XZwhwfCoEB
293YhOsh/elb4o2SCcgn4Crlfr/QPkGurpbumGpfQ9EGsoINFHC8bzkEA76Iyej0R9jA/nGXboqs
As3y+AXRJcUlD3NqxMp/dlx04XD77p2cs34g+x6HtdwOydyiNipDTRId87AE/Nwr+flrdy9crvwC
Zs/w8dkKZLcGyFhKbqmWiVJ3lbx7ym9maxNBAdFxnzWiSkw+mQgNSzSwVGVqIf5XKVlGGdqy1uQh
CfwU8umOT7dxoYo82EiVyPsazkhBGgYxiytJBPkg//Cr2O73ECWJNxBhLFt41FwpGJqn444NJmMJ
1kB4Pls3gOFyBKVGw0xKdBFwvbmhA4twpYpWSEwA/R/HbJjic91asks8RYaslD2zVhm8p4MrZvtk
PW9fg9gJTxJE2fgF4VXhgqnFRu4zM84ahgehDcRY3imRbf8LAmdx96KaVwk5MnjDW2ZgCAFVdQ5l
zbzCC3/+QeatteCtrNuwSxGRyQji1ImDHci4lzqqDkvRlJ1iRdCeAxgtd9srGhaal6mIigYikSPj
SeJw1Ts9rapC7EwbGwDZRy4qDp9E7fLg0Os7B1BK1sg832k/wda+14O9Td2H2YdsXZLUyTfVOosN
J7JgjUzxhbLEBBcGueI4Fa0Fl3BCR2hDHZh9hIJWUY1frJb1AgXjP2HLimDVEKulzDHWVvjk74Ao
UCsdTvg0fOso58ogJlZJH8ofRaOWCaPny16myZwNtAftReY3KMGWBDj1C3Sr7uYuBw2hv8T+k3uv
9PAuJ2RODp+myA/zJ6kfwSov97UX/f+S1uGIWFo/ZmT05qLH9K3r1DZgKhvLmuTugHN8qs4+hMS0
SdmZn+Cq5G4118lbkcqGoyBEcrWce1ijp3dItHyoHhxXY4uqGPWazl7QASqTuG3aumoXbPlwPpwd
EQn3lhodbgNmOamVbPmcvwgy+1FRXbc4jVJPfvML+NKJkGxyKktgZXm6FSipaNA/XgCqg8E2Lix3
WQsC33wXW0rOTLQO0zB4OvGth1fByM9xVWBqpE6tWfAk3eXp5g8KsbSOACDbO6XNE5QDkfO8cJvN
1lcOWS20x3rwp4bGAQcqrd1+lQvrzOnSBKUFR81lCbXg0iuD4jv/opkV4270MnnuoqkK+8EAyse8
LXPjFmS2ieNKgSZy14GcQ/PAG12DEompGWmCVDn5dZ93Va8LI9b5heaSMCFCz0JE7mQfntn4xTkJ
bAwksO5wkhaSXv74ZIRi8/BBm/bWkDjzeP/NVWDmTRlvo6VSTi3nEkBEtWea95mGMqb/phUvXEN/
1X1YLIuyBxBI4iD/4rdBhFgk/yAsml1VgJDJoLxun/qSUbk/LoWqmRPh3y9Y2TshaY5wcDg/6xN7
DhMrpD2p7bW5+AT/uo6OkchlwAyfcjC5Kg9nLE+WCxjxobIG8blXBqM16/hRwvhmUAutwjRlM922
C81fRJ2TqR/yP8Dz1CDa8u5ObyGiUCS33d6uBNOJJPEJMurauiLx0/JuXYO6kNy9gOTSbCqYmjJy
dvw88bhB9Vodlai/La1ZqtUa+2Bs3YndAHq96CHEEnS8GE2hBGVlYfhxoAPv4n+0mE/phCqVEa6a
U3yd3yq1ZzgZ9rz2HUrNqhQz4tOhG6s8VmtI6BvDOPSMkJ2o8HyDIBziCfDOJ28Ne9abryZZOe6W
TbAdSv7D41L/sNTO6ELMFV7AOfh5ONz2J1dsPxUn+4c4xGGrufd+rsh8iHHVEIxPbNAWtd+n5rdE
cWNB4DDqox+bIFr3pfhopPSxOCihPz9KPx3dA1tA2lWvYQ/3h6L6cuUKHrYbpfyT2y5TBIEwKZI6
RIvBIKQ9IOgGmnOleP7+MS/kNxkBNUVz3whvbQJrw+T/3K9M/ncSYaTiWT7sw6m9TVwUwq0VVDeP
wo+lQfwDLXfh/nFP+yeUAiS8ZjIiM85Qcix0XWRAwBUAoU8QL7+DTOOKir2FmvtVLSUWbiA4OhBu
YZmnpsRadr98cBvaeNks4noXtmcgCwHz0LyRv85cGsk5M4bN842Q2eisWFJ7ZiGv+ZF/LnSYnuRH
RXdhprg5XS1dQ53Jg02l3KKwwMpbQNqDeO2auAKcePjG6Fb4FqrTVbyq5YF6uujamtY0WIQmlwmo
dJzEWc2ZnQxbae6CxyDJRfwPBtbm1IfeAoqWSFSJ23HA57JGC3hrO0eSdR8aY4gpPkv256ew97l3
iBaU35G4tfchH62vYsNY2wkOIDACOzhXeRN37O/3xufyc4lSjQxB0JxJyM/ZygAHxhN9E0W811so
3Z5o5tAO1zXlamBszOb2pUOaI16SbdyCqJ4jIdgCFYCIMBiaP29ws8ODt4T6a8tqR4Nl1VjFoofK
+LO00R9LkpVl3U/AcCN1usxc8j+QdeCxg3+wjkSzLzKCo8wzSLZpN3cpHly5JdeBUqbzCauufqfn
uF+OPnG7NcKv6FUfGo+X4LdJcRVA6vYv88Zesnb4oWzkJmMBqwlCY9xNsmkTaDuU26pP6t4KB0jQ
LvSyk6vqd3O1uCUjC1wvRf2OOSB6A/9ryCT05duQ5z2jw48bhL3O7SwNxUjTHPdqJz2iAQARzym7
3u+Cl/5GGFY3C+Ssg2CjkozoFDpI7WEOJI6qaFYtx0hZNXF4K6ja2oWvNkEcP6ZbZ9fxQ17zG9hr
WcomfVGUfDxsZaKuabkIJQY1Zd5m60q4DJjupdNaTHapmyzvit5EyzBWWhA0aiY8sK1X0VeSKInC
QN5tqD+GSqjwJaOmKJae0sJOJWrv//jhzUft1X3Ps/F64ZlVCK0kryeRUBMHsDLw/9SMgKuReyDr
CcoCPO+XWxAWjzn5pDvEs16lc2lWAaSepJUI0O+7UN0OuZmcyMAdinKU1EB6sC+S1g23AtCscq49
FdmWjX0AXrA/ZNDC4UP3ONnznosqzO6Cy9tMdzZvKnoQFxkkMwCN1SGYFqdWpM+XKWTwoHhsY/PG
U7IauHGIYQNI/fkntdnDB7YE59TgMA6ZYEO2YgoR+IYDvW1eXLuq62FOg92eKHBo8cAF3455PHvc
N8vBgZA7KTPIwcaujxA7NCNZMl4v6mtqcLuu95a43L24EqAo9Q1rNtmT/Mo2ws7Lp2XXua52J3xc
Oo+VAq5cVdtAQjtybcLsh8sf3sX7QM/OzJmJnpGNM8jhE8et2LgnEXv1/dTJheK8YRvnDNa0pXbY
U6SR9J6G6zVOtqWMMwASVIX4sDLc4bR0/aLxDQAuzf9z9AWc1kTFrubGRYAopambKD1CLxpZD/Wk
cmvR5g/O4HSjBwLLVsNXgXjOF87x6qI1XYnXM0w5JCSuDKepAPanBNz/IKfON/DwsGJZLl8ZPU+a
JMzV4Vp3sc4+dHK8VUs7aCi14JLsluqRnPOuEDPOSo5rgcP84MSckVz2MjI7lCFyCwYCd2hrxzUK
geHKFYnun5EXKqZOeZn/3nUqUSBKWeT3dw6C7W9Gg8p85uCgA1pJVNPFrpGJumfmV4Yu5IWDc8qH
cpPTQgDTph1LIW+cL2BqUnjevFb7KQz/yYhtHC9HSqVK9tMZlnhYeeybG2n71rK4Ete3qFklFfh1
inD7AHATE0y124AyC/nNjzBNxqtQWMXG1aK7Me9q2ILP55+u7pSRBfPtLBIJKz9Sal6tgMUFssXD
puTH0ctnD98k0iiJXkJwxP2W3ThwwrPhc9/yw9UFnluiIZony3DGRsbsgMuUc8gzZI1hSHjJX3r9
d22bI2ot3xwQ26tBeHM1X1c1vXoPLXYBCNl3yljCUg4mgi2wMxHt38IosN/pHQTne5G6sT9dDPN0
3YcXIidYTtZ7jEnWIg2AyyMEvOz/Luy4bfGmSsM8eSK4PVbu+Cs4lKI2/VeF5zccHpM5ghJKvDOg
e5C1gsskpd8NHzHLqe7hqzM/M+OZ6YCtrPhfXvCEc2Yeg7+keIyV+L9rCIRdn/qTVFv87v0JysZr
S0vCRlzBxyx/r9Xliiwjh3q8ZBBkzdhkLWCRfH+2lGFA75fiqxr++f6SuwBb2OnlvOSoKfqM2Ibb
bH/mcK5VT//7ii6skWNybLJ+SH680LLSBmc/Qkj44s9JoP+u/GWNWjXhtcJCFbL8fx5ORWXw3zR9
7kQDK2S24LXpXKC+0NvRJ6wjrGj1/ojNt5hWdG+MBRSAIaY8RhpEltqZNQPRgCfgRoy2fQFWHJOm
Pz8MxUb0ihlUlUxepnlsQ5H5qkWCuYuPqCWGdbhHRw/RyFCWcnOsEkQE4uMZ3OfGf9mu4yqOiPsT
3BOYj4RaDJOkLcQjgMkZLna9a9AtJw5JCla+vKnuxzA8JXIC964nq6spFK2HuoZauJIkt6IrTUjT
xNkeoOYQDYHyGgS2YDX5pMKjY/D7vc380/PZ6UIOJ7+cZSAVZ4dlilZ9dAsh/4KUnvcKwEb1KCjI
JldGIL47HEFaGXcKGA9e0oRHsoCDS2TdeWj1jkUJaDQtAgBWHcBHxuRS7Pi1j3y3wIPtYvKDt4wd
RT7SS7A0KoVP64mROrHxl+8qkDhwnQMlJk8vOxfkX19oP45Q25OzBixGlKrYeXWAggCM9tnxeiZ9
zEEokWrnw0S3wXugBDo/iiNcxMTvN0WSTBmsO8jLmuJRsbtV70GWmclaN2QquBGSjeMAoKwYGqp2
9FA33JsTX8dXNdIiNq1LRmZB3MWPoTdnrTuOoWPzjfLzhStzXAkR3rvfxJd0ShSpmrmYR9LbEUAS
vrTDeQekp289l9xzVt/tHVZfSQ20A1oJ9BXknk6MRR8MVbAUNRxupu9irmm/oSq1B9PYeilyKz1p
AGHDSkS+ehT4NI1ZtNS6RhkFZh+oqmwfH/9/EZb4DDrrL7dOJm3fMDUW98eIeFwjbvt9Z7ed45Nr
4xRZb9sNqwSPWRBy43wBq70vE0IelIyZj42efolQxMSt0hDODZCxh2LvRZj7wJ4sRrfGpjd9fZ/j
YSzVU933FzjX6YCLM/L2WHin+H0RPOGDyIlwpMMBI9dab4od2KfCQm82WJ5wuXPaXdTvSSD/3YVK
5l6MBW++hGZQu8EHSsn6I9n6h903MGc5nv3ev1GvuIKlYwbEU75NsV+UFDNUlc6PZ3gIpqcNj8cZ
QO8TM1sJ6ezrEgJt1BdH8dHxi8ELlYOMh3JkKJQk/8TT3s+ejDLtzKzB23SDArv0KEEe4ag5ASdl
7rIgxjlfKTTVvcShoIerPpEYgTxStHiWxz2TyNX2nDPzIAuHDLHh5zb8u96hzTVXFvXKd0O8CZxf
+aZOu0tMWOGV87A4ddNvY2ddZYtI1D0W6Ur4hDq4HDKkUluNyEHyR7Y2UxPL98QXpK3A1nH3kbdw
SkupmuWrQvnp8reH5nGeR33K+wwKzMvl6DjIsyTktSmfHp8CymKWrL7qJeNJYSCHYrnqBojCYEvp
WqhsMuHFJagRGseS75UfUaS9qN0FL2vOlHmm6X1OAjI6d7KExgNL2BSANpvb169zEI/7MzuS5gbG
3v5AqBYUioqMtjtLE/ReaEV1IVq5eNMhOBhXVD3B+Wzuigop+gBZR4N+2YhJzI7iCcL3Lxsu4sZh
d3UV4g64yguWyN529ywYF5gsTy2IHH/FnG1IoOuzQ5ywLsIB4FVfqvqxLpQ/M7y/hHmVSRR7/fYG
tQ2vOLIBUoqsFYmTCJFDzqcEJqVvuMYW/6w0ML7rr4eGnmiqI2DQF9UXhpcxuiWF8+BQh86UEevV
WfhPwG0x/p0yIfhZNG23cVshtvFytAlcOaBUUPz01BYq7MnC9fDMbJ7pND/0zp3FSCpO7ua7bVe7
76vy2UGTmP41GTDygF+E5Q39wXtJ1laQkQQxtctH09wcZAaVX0XGGjs4WMtw+a7s3QXNIiclz10g
sZGBMj1FjlMIVszrJj/eXP+yA44g9n5y1H7ymONBTpblEO13uXbAvytiqE7vTP9f4txa/MVOQd43
yoJJqv1wDkwl5qD5iAlhHAsJNaKExuKFJS2xuTbOAawXWHZzVlldOtb5Oz37Jn0c/G1mMpGVcBaf
fNFgMoIUaZBqCWmVtRGuF3CeLur1RlETEcIV5MF67eVkVb63a0ez2IvPxuOpGBRU/qgg6Y2hoJr3
wneNBZXMwyMXQFnCG8iynTa2SA7U3QUXgAPqO6g2MWsPBw++Ds6USXsEO2shSrGCbZ6ls7k+Vl2+
3/Wj5P4mwVvzjNGAe0al0X/0ZX4dqtIEY4XmGjYbXyAEKvsiccSosvvWN0Lk/Dq68uiyjH6JeR9S
Uz4nTbP0fIC0o7Yqay0poN4M8fITl7YOQGOZHT15/Rbgl0gSgnYYxzKAX7puo/U8FV55PV4gpXSX
EdhCUAxCW191fp1Vo07bo7Plr5FZdRo8sHWvYG44pohmGhHkPwU9VKbLI+zMLxPkq+GOyR4Fe7EI
h2PFuHTvDiIa4lvsnHQMMVFA77LoNtD9ne17IORtOnRw9bTJevv9Tw69v/8T149V2KHjSkVerP90
oIB4GgmFy7xGgRPDa55xflazSkNalE6+TLSLy0pAckNf0ToVOQBD6HhdfoDvKLCq5w6YogPwZFqR
fCPDkIYoP0idUbzOsZB+PdNR9N+iCa/IwBaTlxy74pAkIlNhEmdF/Yke9u0Bf32ORJvhIbVTEPoa
sEh9yMeoXNVRRGrDdkkpa52aD5k25YpFNMINlE1i56mYYSNb4YRBpDqgqFY698qgnI90CJQB3g5j
Gqrx5Vb0UPCVZeDsxD+y0VFvYmEZ+W+qd6r5fCCZJCCt1G0EASwHJLHVW4pUvjrH9iEqDTUkwnIz
LWZ9lILCRloKdEpGnOVHVDoin5EiXnLk8T3JmtQNFn1e+2COg74I9iQ5bsGyQtzbthDgP3L8knZS
W1LO8yzLyxxVehTJqvmIjftFaxeDftbKVVscSbsHQZvjkhlEnHE9Toy/Gu1tqCCDkXGybya9EDK2
jfy1jTbkPqdLs0nBBww9p5XcispNcD/3aOrmJRGK6vP4ekvI5ULjZ1lBpyynOIjiEiDLxGA8OXGO
ywXR8GK1QPUEC9oWiU+arA9XYC0jlAcehypOZfzX+fjAN/GVi/x3rZx5PJVW1dxRzzxB470JodE5
12pX6/tv9tEcbmyv3U1oE9RpDKEJKZuCk6OLVtWG/duE5+hb0zNuGvYwymjOYs/LKJ3Da4vplkQM
RUj/fucb7fZNoialkbZYC1yLD/IYr2TkSh+4n2/Tl3SUmyvIUpK4twnMnTLM4FMg65VZ3bdEdHyK
yZydXEpdG58X5UwtF+gV5jLLv02WRxurZF/AuCtk+JwZKbJpMPfXBpKCN3Zd80E1e3IlQCqQRAiz
i3nbQqFJBPtqYtKUViP9t+i24VfsRi/iiJ6xUi8ltzCwBbZS4jfVqP1S42euzwiRcS/GPCosa46r
Tr9/uklWv2jRto94uv5bWmEoKX+MDme1zv08HaDgGdI1pvl2W9Y7aMV/kdEk5SE4AbvB/qsjIUB1
LSPBsodPnd8fRlpV0r9ovMTkBdMJaPjGc1lLMtlt/C1Q4GV/gXUXIhbyygDAFiILZBFgeQ2hm6IL
/stX1Xh0f1abjMG4r9erSXOomK2r9XZ0b2MnnBdPiQmI7ldgmVipsmHmlasOWkvysmN3sSzUhmfN
rNK2KBfLkA+ZYLyKCwROJcGvM/sggY1z5iMmBED8JjMt6dSXVGyQOSTrE0auIGHSo+YDSvp9dhYz
LVlCvROM9O0oDP555UUpy/BLWDhvNWLUXjAwlo1g9O/L+V2BKpJnRJauEvZEnIcHPFEA+ju0iXtX
jcUb5U9vLTvZBbRMEcuA9snissQvIaASfuP/0nu2oJpwO9SS23MQnnYt04shHouqTL4IHeCdcvHG
32KcTBneyrHOkOaJySfjXP8OlcgzxL1gCMlwOFQa2rT1MNX0fPACwwLsNKTww0T+JVWRS6PiVrvj
b2H3CkMw0BxqHCCDqGUWFJUVB5ogSeYJaUVwNG/O2CRGWjndWGxmdYTK7Yi4KTmaW450XsmOGJD+
PwyQhyj/X++ehuypb8WP3loUkJpqj7wIvB/qyapsLRLjTdCztS/D7yijTH7Bw02sBpVcZz/oKSkq
JR3eLxzj7vSJTCQ5eIxWbbpD16hz9rMHmd3/yJ5E6tLwTN3aMIXX9gjgL8t6+N7nQxjtAUClI5OB
6e9qUhgwN5B2u6EbTpRM6VkTJSDRw6cD4xLZvmhItiu0sf1YG1netFp7i3pjf6etiQAIrwlBHTg7
/PiU7xn4kItWn/Y2JDnNVHgV1LA4hS8ILgzy6yTGwIKWdedDZhoIIMeik9twZ3DTcLMQN4IqDt48
7mEKQ8k9ZlsWLY+KFYD6XgcQWH5W+NdWdowwTmhLcvpw5UnP5tP7AF2zSWZ511+Uq6T7T5eBLKq0
3FHtdaebNn0ajemvuXEGQbBysVzIkYbjS8n6dB9/UrqLynwRUynDRUMKO6G4MSZ4xVuKncg8aRZ4
6BvVSCBaBO5cSVhtShxNosxbSKIQ1xNRul4hsE1+dfTt5ELlhLQfUOm2TfjmAetPeKmNotz7W2qq
FyFfOc4r5mMDT5LvsBXdSdQWaoUFzUMXlp1kG0+BlqyABZjcvfueKB9Gtqg5cou2QzzdMzDCHOG3
69YoZi4yI6OAxve3LODbbLl2+3EXREpufHp1mnj6mUFBjhocDWHbNLmV4jax4M2uLtLcOjWTLxcF
dModztkmS00SXldUWSPej6itog2UbhinT7jwC9qAhle9PXutkvguGHyU+st0dh0Gw9f+Czuynf4G
9H8nugWc3ZxBe/yUd7pwtKC3vIQgDiOgsLCNfyppjwi9+a3s4zm8geVy+K8NKb21xOAHDbdz/pB2
M22NTjfD0yvAK9QYwJK0LLR9OdsqGw50nnsPyhBdLKK+xyNQQC/nmy24K/Lj0hEjgPJAyIIhKmQ4
mF6YxlmSN8Ys3A3oVePxGuzZaYEY1SOqhO3CXCrqXkg0xNTBrV89YfOR+1zLfh/AhjQjBrp/BT+k
vQuiHmKHWDhEs/xFWsFZhdasZyOoNLUK3pclc3arjXy0MS/6MK1oYSbE1foPAYfCI6D5qMVupStN
umXhqNZt+LlcnVyARXCgfvOpuhX8w0wAhaevhtiAJmytmoHKx1UlSimJAFXj1FKIczEC6ONXijwq
egFl9MSMcff3xSr1wjTslT8cNzglqp/uOrwIz+qCTXOvAVMjsdC1mig8YBO1SSY7XVVHwFyhGykD
T2taqSXB2aLI/ULTpy1d9uzlmJJ6L4nBw86rDbwR43H062RXPDosN74hyRICdMaUTNilp66mdVky
TF/rBfyFq3900Pfyg7Lde9wY8N0KdHtHR5AP58CWJcRZk2y3Bb3jIrKGnEcIb37Y7zT/LBeYvgka
NCsmSU9lYZAfJYSvUQGR8vxk7Z+1RPxQZV/KFfvKkVMHZi8tYouxBIzxM2deL6++PcJfUI/Boa8P
8WjtxABvgb5fpWORz+zOHZE1b8p2IlR3nHyyW+UNJkjv6cvD+20puvQ9tluGMizxDSVvdJBwMllI
ALhongjldgJ2vaaWFsRAH0BLpzLFC1vzchtAs4DwVFXyrrQDu2O3xmO14hdWAubpJdy2814opYDJ
Li1F7P2EEBUXbT932pjqFQAQTeRoKcMtgrFk1zb9i0c2tguCKUkkwrtmtK/eih6EkD1aeooMuAJE
zUiTE7G9SRTKvXSCR+KWeyQGv/+7QIinsm5xyx13+VHbt/2Oj4EgwWaPn5Z50SvNB+XBxVBH4Qj1
QAgDcN0TL43hoU8XcoHRHyNSWVGp5III/+Ju0lpy21+CVDPHbcvVPkm1XEf8+Pw1/vDnF2uZ6TPM
HcZv96udWlnt/NPtcUJfmt3JsZ3ElHCXJ9QdlpDWEz1ujLtFwy4vEE/QMASZ4s/Mo7hCGxhHZJO1
xndmpTMRjoY6VvQ5MhX9WHOV9TiFl2ZLe0I8C42pcT+zhmAEO5vSdolpZsXNePdeJLsLIX8sgevB
xTge+TDI/E94SVBcpNyWCSt/XcUSbjDyNV5uLCf7WJAQhx4J+DVreknVHxK3HxLs314iwErajDCa
hLxS7YdPtm/fOQf83H4rEE26eMwIaQMEIAljFUqfdyDyYQTqHbTA5/PJe5vCemPc5/13DACnm1ZB
lWkdnqq9TKfa0OTAUazNdXlIdDZ1La/wOD91EscQaUW+KnRT2pl3uzSKfwFExbe5f/Zw46N/GpK+
x4ubvCk/V2JqdXBfagcWZkxAU2JlOEdrDLvukGM5SpOE3K9jw/cZhbLh4QBGTNmM1dtnBoJxThLj
8rfc8v6LiJygJeeKS4cBlxnMS3683OtK/pBAa39WYpojKFZBp6SVAPXDT/42nTkDbCzcW3J2tAOI
jSa9VsQBCbkcZ2gUDPZmpGZ5mZ/NxJ0eppTcbTTE6xS8m72IZt+vBxdcoSspVaQgV4ccEDinneh1
AvoQsroJCojVppN2Lyqm/VLqdRIfakD1fCJjAW+pq0kY1qOkfTkM96S+KqKyLdXcXAei8qNyHxIK
AqGkBGN9kQGlaMhFWXQ9i7GuTYzzucDM3wIymqI9P3YpOInNKs92tXeQ/ntslHl+6Jg2ppX3S4+U
lq5FVbiKQDuPalpb5DqggE+dlfHLeyzK/tIeFqh9TnWZTrHfXA0durOtzDcwZCWW51E7RdqQ+MFZ
MO8xV6s3EtCD5nP6lmmfzcnHEJ5UcqREBg8RDuv4nYtshF9RhmBc45Pe56FXgmGQ2VA4PhDciuPD
Pr6LMbAMFzjX7v9XSTRl11Q98a4n2VRkwbuQv3z8P+xPzh4Rn+ffHwCrPK4GpB1sFYAbU7OWHYXX
Gwfj+20T6AzJs3Ja59VlO05GGqwgv0Bmm88R7twcgtRJA+o/zdV8/22/cQmH71IVJ8KYgT79sOB3
FtcBw9EGKiZ8UFHIr54mmy2YFlAGPEivTMJ1SzRDSfddK/BYp3SmaM3eVDoIW/n6JFpldc3DS8FU
w8E2ly9mCPuc1hUCwxA9M4s2Cfxgx1D1H/W1EedkRJHUrnHdoNTz/kvUjS9BD5+fAOsoKn748yhE
mheSB3mtusYht+8mKalZdEraLWS1mXyZV9iZEUlgxYa2COE9vAosyid1g3QBGxtK/hOA2cmBUzlr
rnZLyMybR4MdyVvFli9+kgUmPurRE7M0BZHEemTwmQlnhvoLaKjMS/BxQKKnRHwnAs/VDbEDDXtL
CkL+zVwOkZXjr4K20e1t5oN0NtgHpQXDHN+/DsnoWiCe4mL1GS3raMu6vF9AJkXiqUOnVXMni715
EaIIfnFhCuQ6whXk9Ns38fR8sOkiA0jysf/cR/Shbrf6K1WwZ5a0yJHYLtOkwTEh4kelk702d3tU
IDbsSXTzE8WPcWvGy47+RqQdLfycGF7XpwDn/kbQ2TrW7neXcDtWKcda/S3tsfDQLFPpTZgvG/Nb
398mtoxEIlLwsDc2+sJC23nXwLGFQvBmVTYLj12AqVQIl5GrAqRorHZ2/RGZfAHfcLGHnNCBIfOc
+JL5Q9W/QW7q8Be5KhhQ4nAMI6stt0wqlv7QC8dkVQa0Rir3ZObmZ7wmeoND1eZH0+kDvhOcLuJg
JSZWms6TecXzlaBOZmks4h1Hb45wI6AYjh2UWBRBeRqZEhTR6vXBfBAo+duiV8NxyCrfVVx4bSxH
5lrbjtnRxhXQVJEap7FuLP4s4z94IqQNP1yHdppw1f/pB25L5FqihmFMmAY/yg/lt4WiBivBN96m
VkCE7BcxoF2p+XsbAzce/xH0/e6FOHpDaaVAJCLTYIU7NpHU+YooNP6zfiqDsie5DrzKT7bNJHdk
Qq/v2jpl7VmK9D17pEDfeuZ5ctOEGSGpCcxJlkXE0t2Njy5/D8VLXhW6F+KKMPU2echyhjA8buCS
GYtyrVe/XM73LUDID7WAIroLVNaXiEKYdPsTvbCtfoHeGxCvhLcwRybxbcYP4vi7uuzQXrdZguGL
bJQ1htyZ82Q0rmPw5yxevdOVrZFuwpWQSkSf4FYLEW5gng5UwQRzNlelBse7wf8SkpkO8AX2+D/h
RtSwTWo8T21wG+BCMzGog5nGhF3bfDQESTiIstNQYQDxJor75XEY4l+ek6bJ2rIWOOsnPFv7FjpP
bFCsMkjo00sTdXAJXQqHH7L863oRdSCTuZPlRM8UZLCQXD3aOnhsR58Aec81QqLn0bjjqDBzm5Wp
Qa+wTvoEG9Yzp+dJVwnWvE/UULTUQA0tBJD39pFZI5zUwcnDHZwou/KzL+/iBr2xvaJIJyRXpYqj
cGzGuAdWSinoJTrsuUOoDjBtNlkckDKJvGw2Q0oyNAvVlpPDsCTndRLfYzss2YeAkrA+KqklViua
wo/FZ9605tj4X6hNVm4AmiSdlerkO+gO/FRyNimCAOID+5rqmxfwDEh4BF7mmDfAInSfZD720864
1z4yqnny7wuL/ilscBVDhU9nMBRPZotvjHNwuZ3/yei99LEoPLTyfv8f+CBiL5QcylmVGmtvTew6
0TAFbGwWJQznwK7HlndffyjXOvvDo5/KgVItgLSGaDA5529kXjWKBDnBRpkVUBZ1mm3T3wPCT7UJ
Jr+V8+0x2jpf8Bq/0zEzUI+WIaOTTy8mzX8ea80xjBsTcmhHLrHvcChR4p1d3qxtSr12RLxXlzP+
72Vqy3dCv59QU5U9LWb3pPVOhLE6vJViPULZ03eXD899nYNw9T1TPPFZQMgTGHRiFr8LTF6Pz9VU
uIxOMktFqEj1aKogwZDnPHjHNj/sIQ6lpklldmhnPgxuVvBqSxvDeBx1NWvptahtXnumfRhUxb8p
UJVAxrKMtddlpjNg4N9s9YVaSzsMWunQ/7mu1gs79IiOV9PILGkqRLd/TCsGvDIedKK6clQkdhb0
Z8Rqguer/5m+QE5W5dfQ3mmGAY6QTfHD8PAdFyXBrM8LmY9KjpXwDIdpc/3/ybNbFrzNz7ikZkZb
s0WOwnAbFuognrfrk2049NZT8hNbcabi9U9p7kv/IqDbmU/cRsCeg6JJk3qgqkVbcpyxS9ZHTNae
HglsqiVydA/WJXdckgGOoHXHxKIEgwKl65MAOLGARhXpLZU9iVJ+KyFuxUzVwVcWpAL5gkL0ffRh
0CbuzPQdErNZw7md26ywSrNWDDP1b6LN8HhyTD5Puyj+jlgej+ocrdqFtTn1mVk3MaqKMMyz3+5E
5eNzdOMW+zkYw5VZRBvNnV7J16HiRpoy3HnyQ5dUX7lRKdY3Gj0t7IxPzHb7iFEHR6FSIlOHJZg2
k8Zgb9nVz6oz8Vw3HuvLJvOrJMSqkV/vQ64g4MMFp+67oVeti40xIRA89jFef7x9CglxltHP1IHA
yd5GS4+ob64nHVsXo6nwNBeKar6FrJQ6XzVRz7StQYRQ7/OIoMAo6RSvoSVTNwOY6kpA9UDPrtOY
DeNlcvNk0ZcDJE/fgsGd3CEa9V5Uh0dj9ijRW9+h/0JdaEslmyxd4aXSn88YicgMfp2yGZaiCvOu
D6ZXfFDggcVp0GKsy8LItxnwrr1WqdKK1PxQ0nxPj3Qzn1gpVjM4548qV9QQzxWPgFLRconRsRAi
TK1gek9FfWUYE5YoCzD5a3INqDUlaZomEA4ENe3Pw6d6lEa37BUfPl38KiOSs+izHWQ1UngSFeBd
PT+o4zACiKcSsz3/V1mPZQL/niNesjP3nkicMxeWY5VF/FcsLt1nkja/NirIxxlNBECdxzoAXhnj
T12lNRJ54oXswM/pd8GV+oabWKZ5GFqxrvWpSi2b4sDoGwg8rg0T2TaqifAUUj7EQqPgtsoTxj3Y
WVI03SjyVxXOszoOkpsSOOvXw/AXORz//a1RgPcgWNgx+zZ074Q5jar8FgZvQkr3BFwKCUmQngvv
omexH33qlFfzUC2Yu6Do6OsLq5hwvtGWPLW8X6B8I8JcEVIkunq/cqpKShRgas+roe6aQ3fjqJnK
z0dmP72dyNCnVrwUi6hrr3TArdr2LENxwxVy+gPmxnn8UMBtk++qmI5w9TVUK73wwl/eM3jxJBqE
DU1JXlH/3YXjHNHS+w0Ed7Ht44d9zFR1Ta6jcDwN1CIO6aFca1MRPzVR/g75HDZBVOzuGs6W2z0s
a4r+F0wmi3o5iIx+McSF44ROwvn/TRna+ZZrGbdN/uBZRrJOO/2n2QlVt3vBRpctkJ705OXcEy2j
3lpyPUSi/ZfUd6wX2HYPI/yFk4fOEaSS4Xjs1FtgEwnESmtJcLjgTHRaueON5Qi+XRnlU2v4eqjf
+y/km0WmFuFndWFhVp6Pca6NpvO8KrdvX8Z4UOS7kw9HqpZFh3Fe60ik3GZovy13nJiR+9bs3FGd
1XWvIx2jEqQ7hHklpVtQRAEu1CnNsojZvZh8K1Yq/IZgQSPFmMoNY5nnqyZp1gx5P/EMvPAvoe9H
GYi6riKsDu52AHPWMnQOLoohUklu2p0MPrc8xAKeYniLa55Gga/1a5w/HRQftaSP4Z9ubcjqVA1x
ZO/kYbqd/nATwUNGncFXqA6slwz+HYlobuHzfLOaRsxsLFq3llGlrQTaQNdwjdJ/otdn6vXP37JG
iZQ+L4jD54Fc9Ig/Old3TxoCF2fOjsmRTzDncpiUnogggNcwJsn1UhHQq1wMHIo3PevAIQiTUnpr
yog0q9bmZ+fA+GsAWX4rnkSXY31O3EhLDm2ySXQAmRbnSn2DrJovfD165VjXXIRFbEOpsKv81+mz
Pguw+D55sQRdLVfUekKtIBK2SxqyJt2czlXWBOnGClAJnTEcGJnyK2Gvi5lDQ7WNqBsA4kIGuLi5
7CiNi7R2VbkQilhMw2bgWW2KQ++jM5XaK8vNuKHw5LZgh8Nngm+yvXI8aAiDwcBzrUnazikkfoVJ
8b4z9WKEl8xbaa3I//MY4Tag/hbhG34BAtHznSAG8UxpFPnhIQgwHIC4iqUxuoWNLtNkrkXb3lTh
ionb0xJftf3M4SPf8o/Ixt8jWTSrAFndbc33yhXkcweJbSyCIhUnbWiN7rdiJTGau5pOc6QHQO5v
ZLC/BA/b7D8K308x/M1jpnUGOBGxf04hHHSMU3rEuKmbrjRHoSePFXE5DyvpOKh/tCsMvkeoRVcz
SlqGWcMBqrDUBIjn61trA5nudyJNrieLK3goEyV+1Ns7v0ixvt0CnsfYC/W6Ov1pUXufIdoez7W4
pB4LKy1/GSdAx3uzONhEQFZNaGmt4RbxHP9n/R4bhH4GMNrJKOp3HRmdesP3fgN1p5uUyNHacWPv
qxNJyMth5dFRUX0E7//eaIvwey3XjdJudYEwRPvsRiBUAE/10FbBWa5D/t0Uo/J+HVuyVuZR6Z5W
hzHGBMQHhiLA25AERpA6yppd39ohqzVWBwVXxRtl/Asff3RvM2HXGUpgbFE1gn1FcUs/1j0rfUeG
5fjdHTrVX76tsXw4Y5jr3zmD8/lDUJ9by8UgE9mtG2VFe5n0vVoc7hTRtFGqRrPgS1AyActezQMK
OJH3in9ic8Pn1hRuZJRIG2Ar1SI6CAZGDjZAVBCo/M3pYto2ShUJMS7bwLQY2M8p0Qzn+aw5BeTW
fhLz4AWc+v/Z7RUyDQjz6GY92XOTIRKZKtatOQn+loYNhA8C3Y+qsGF6E6HIEYHIeXUO/cCWfGbx
9qoMsMolxEPMqCls6uLKvwFxOSbb1uCSPXd6Xf86FNA2GwKGfHOthLsXQu7CsKScAzni0Fh1p0Rr
kZ5Z3dwmK2v2VftXGxiKjnXjazatyRNPBfuTdo0cZLICYxbNgCpGjCDNImeL1lN4SGnaXSKf18ZL
7rtnoIUgn0dgkGX0MGXB+vvaE8+zJBz3ZfyP02HAlX9SpgAQiXAAtVDtXZeWHl1cvM8bjNNPG7+c
yt0zBywOAY7y0Fz/y99Z5jNokPLeEATKglqJ9CLpfZDVyc/HIU45VoqOkc/NMY8cMddk0AJjkJNC
8y+GWwAKSg9UtN/6efL9BCkB9OvCwri+SQO1B3ZqHen10A45k6KvYyYVxC1zhuvKxl+tJAKEGbZy
2HcYJ7P8FfTE2JRkbYdohSRASl0iNU1JJfOAuKBPBAeDV8tY7DskLPPmOaALECoU93Kn++s5GAVc
6cbZqrIsILvFTtpZyyiwAyOu1VKp2gRYQQrYCpc6pxcz3PVtTFysWbt5ANP/EaN21I3KLTqbLlNi
ZvZokfbJB7vj145K3xjvW8JhyUzAppzoR3oA7jQz9o3EmCOgOWDCbKp2YNYG7WrNIE3So4PRBPcd
bL0yuffyLrtIB+rGgQhbVibvqP/uaC5d9d7NLD1QwY+aM2M46mFtxIXgVj0xsWBsFUVTJwi3n9gb
W3cesoK9vnxNkl3G7b07vlSJGKKGxBWcO+wOclWlwkMkDecB4nUCc7FHGUedTpTFXFgTHoxhr6vL
u4pg3zUhOKQAdXVqznqxfRsNJL30OQzemKMl4PxfH+xyrf2tbkPIZpUWmcoJSEW3e4abP3P94m6U
UijEOivlTiKWFyAhbS5zEMy7Qy37M1ixkUQlnxJbullvgXWRfDdLisG0K0teRJJL6nSN6ltU8qk0
nAT+LOvPKKqcjkw3GtDO9Lhyu1aR0oc1i/1zn8OzfficyyJfm5duTl+d6H1SZnazXY/m1aApmDLN
mmi/RQIOC1g9XxxlrK+orzGhIpgcnisVegzjjOPAGdqxtBXcMkAbPsmF3v5Qfwfjwsn4DMGnjT2S
PytQa8PDT/ogcOfWTjJcGo3FuA7hy33QlbLMUplYv7ZMGH2QS+l0PUAR9kd/zVJ5ZJfyBapT/Y2A
61NlvECcSdsp4un1jyebhU7QPmBqLvxYUn0zb+cM7q7Yw/LEaBo5nB3dIZs3H0XdtTOkH4pNVv6l
4TU9GMF8bupE5BMmc8Ne2KRZKYHq6ToqlnNE69potM1WPA2omdEZNUE+ZqDEtiLnbzmef2UFkQRB
LFyuMCx/CeSQa1qPUjjWnabNk6dTx+zH/jWfXL8GrFZ+/63US6WHHBmaQKFyktq88vRP5339hXdP
OUXaXlV1UE3BpG0Nw+7D39Ke49NK7svDI+0b7QPUJeqrirWHelqs5Qh3qaVgXUZq3+pgLTZzknEi
eHxhf/SqL1LYXrsEIU8M1LO7DVwM7+3lQlOOTKIuTSHcru6AvkugV+pY2XBFY3eK1VwdHC0y/aca
fLKZ86f5B0Hfhlk14eVEqTISNbZQ+wEPAUPoUmM0VnxS9TWzQeMZ2rtMNNzOF+PtzpzG6eS7fAyl
lVatoBOMD7Clw1vh7GwdOmbD3YFwxZqJDZ6zVZw8SDvc/GrqVCSWZH/r2/vvK9o42fxk9Aih5VmJ
n+ViFGX2cLBlrjHdDqvj3RoM+Sq+2hXAgfHUZmojc3MB0AsLTliuRnzj1PfvKhYGaDF0XgIqAqTh
I6mbyujz5la6VSkYwZ18RMyUzE/xw1AtabfrGL5XVSWMT5eIlrYID3Nba7f9W19o4sUlHkTAEpHD
//tnOgX3+sjMKe8rL5HR7xz22DibSmK1duEfNSer/dV8+3+le89ajRVPcIb4iDIz3oM87c4OGJzH
nj2lMho2IlrbxRYKbipW0qHZqgy2zeygQ7wVT+s0KQCSqS3zHhLAZLGgRje9E4XGDT5QoMdP5eHy
sMB2y6/xJotffw//2iLecigGusxJdLu2dsDeY87LCrZxyPUJrCGvMfB5IE9JOAgCIYvYnQD3iI5j
XPUeBXLmxWDRZTThND4v6lnMSsxtWXuJMqG/b+/pamNzZcv5xCTIguB4/g+I6zPGBq0Lm5SQhYIz
wJnVi/FHRv1c/ucGhesZpIiUI4gR2HI0wC6kftpJaG74qw9HsU7Mnt5RpYsvYt1r+vkdDZ9i7dbX
ea7OlQ+CJ8Xe4vG3Qcs8JODilXAhEIQ3jqfMaNGH5wJhzDVlyoYVDUhKQH8TTnAMn1mGQe1gjUjH
SCvjImp0EgVpuErDfgvLVSsNQ5s52NRpIBUCW/4Cbsa1k04z021ICig2ZSaEv1Ud87dI1f0Kd4e6
ams5UUghMwHZ4oMCz4Q4gV4ExscgnEfWryUtBteBdgUPHW7Oe1etmXqmsz5SR2labkAPnwy11swM
KE7e6zHe76rUB4jOx/3V09nwPcj708R4HZ/C/966EEm2S5R79KpJZ46AJzKhzvxG716BCnn6k/o4
87BjaT5B1Jg9lNukp6/6QV/wE+J23Max1xGOurFGJQQIkdsnBcLeL8esw8PXsgRxZf9IC/CLv+nh
7BB8KiZ9FyXMfM5Q49TpyY3dIqyprZ/bzzgowIsK3/L2HFV+Fat4JzXvDpxbWy5og7GeH8uvhiWK
trWAK/3sJFxQN0fqldgXIipN6iMRhPVovORUI4GzfLfa0uC/fTv9ZaBtiC0N0nDUYLAFvctKYj25
z5IeHuHGfC5fSoEQCrE/4UoFpgd+apf7pYUXz5Nn0Yv2V9kgDIKgVhrgFxZXamSaLz5jRg2yepJp
sRQ3O5+rowPfbtE0PdpauF8KrA0eqJj498BLI34UNh95oYZ0bS91WI0G6hBbIPohCtHkChuZddzR
70bqzF08y5fjxdrAvX09sSlfwTr9j5cfeX5ZGbC42oFFN7LRZu552cUi9vqXes6sep4CGDYnJKDK
JwdkRS0WkeII3hvyN/qMaje9nVgQ8HNE2nc9X6BNK8bWj1/HE3ERpD6sIW4obS1df4ANAhf0WLCT
Y8pC4JTXiVEQoDtSuSWb+K2BcUHcftg309JRcUUGl+duUBbBIDD3waVt86IGLenzAkZL6gEepT2d
Euiehtg03NMjbjnrjzMmulK/nKNvL1LW56k2pV5QeRosqbgUC0SY9AHXE4Toy0qH390Efg1gX3km
dQeepAgwGYeqNaHaLF68AmxtyYTWNqVfarOeuj6doYDOgsOdBvm0eNDtS6oGUUWq6ux4PfrEpMhO
zCR74mPnsoC/dkafx3g+pRoNpfJphqtAUrp+JDYiEDDbS8w1LWnfT7zMZCYRfQG63PD+hgzP/A4N
w43LknzZ8z8nULvD1Yoidfe9SvJq8yhLl+gNNdW8kELV28kKZCj/7letoosC+31mqpfQfT+NsoHu
TTd/CPk90s1GTd+DDBzVooQ/1zWeqzy3NcYwZn29TrbiPQp27EStiihmONcmxjwVvVKZkYWL/J7f
Sn6PSx6h2dV1AVWuqxnALyfd1ptysBXDH/lN2nMML57WTCsbpzGWa3mOTnDsv3KjwWG9061BNfu/
YpIzevwAPK4PWVWXc4vnAA7JtKdLtbq4tn3A3WoyZWItWYtjHcWwfQePFjgzBmRzk7pyjzUvUPML
LOEm3eMRPoPPKdRoLxUq/jqTDqSnd8Fh82J4Gbbo53wz3B48tydANovbdsFMbvNhqGOhsTHM1Kjo
wTZslwOGR/t5oAizLT/gtwflyPV+NyBbuGAjYdKVw3duH/ifbpY9NnE/r7AfQJiwYijl757xJlVB
aBr7pWpM1ZmV9XhfOjjnCmMfI+Lj3Q+AoaY/xFFlLbZK6Gnta6xnTGr24cU0FtDHh9TvmyrC7wYX
TeP1TFWVWF5GDc0JdHK+Cdcp2JCwIHfe5ZRLZQ5QEOPdQRS/tFwQnZbCzDUW/pNdrr43r6w40vF5
/MLOSTDxpHtNCKaCgSqqCinJYPjL1FAKlylT3guhVZAYggdekglbrvgt6RSxvNpWTnFrRT5JobPC
lC17L5iMPPeaoMkleOJvq8WcuUf6lr3gyq7TGsbqAwLm7yYsaPGS40KPIkJxXwcmgiZPNZURz8u0
eTjJ4kJ/+JHimGNWJE+SpzGyRhSdNnd2nVXcIFbp1HUu+HDZ1c/jPK5e28o5plX7BsPOHNGHpreS
it6PtGc4hdxhgc9EhE8jNIH1sABek7gIO8O+E3j+SrsO62IBoXjJx5lu+QeHGYH/TdsY95LkVnU5
5fF9BsMGStzOhySn8zFd1XRAtXZ7f8jzedMnc/eaccsTX/KrF9x3vVmBGzPO1iPy1W5RflhuYw4+
9VS6mbmdWm7iF6mjzxJ+/7F6CGVCzDbAJLWzb7YjK8U1/2+OsrPQatsRtLlwvRzjpcwj1YOmumVt
YE5LIvtoUoK6109eU+GkiGhIu/AeHCnBxvqWUniEFl27E2GxcI5/jdX6WPW66wUHGfeNQFR6NprY
b7H0k8VgtJqupUDwFkGqrM1p542PWKZzPf5pO3l8nRRbR9uZH8wG7HkAjjpmLExJBK8tcVmwpFnG
DgadOaMGZdLdt2ESxK4WRQt6aD0CqBjzaD+5s++tNvaxJT45adKGm+344dHEkYRwN28jfNUkap1T
m2tD0w5B+KyNdrtAxfFj+IMWlHGUtESppAHtfMVvPNPjvyPxBk1ulLx+FVkE1Iv1KH9l8hS4nAj6
tdgYXGhipD5w0jgaQA2rwE8Jw0xS2zW3MQaEKeN6y7sT3mr/4hRRKssCJRWNQzTSyhcZftjkUYKB
8RNMFZUh7W9KpNbO+0EmspNqf+/uSpfXA85aAYZ4AAcyKE9GnCweG50eisVYYwNwDCAEHj/QfVXC
zwTXgHIoninAYxoGA0FG1etkk3vvpRLwapRoztPpY8YSLId1QV4S7bQKC7PsqPq/51X1pWnXHkzv
QqsDQ42ZK1RdKPgbH+xTkO/r0Hz6GVCAwqxvQ7c36UpA895ziRBxsg/6GlEQMb+8BQyDOpkjvxFS
QJbY9NjIwuzDdMv7Rzamv00t8+f/JsFqeodDbZQCBomhUXnJNFdbSh8npndse+48HmbW3f272pmz
kqddhyudgkVCFTZPHCE4h2IUuT4UaYbAjGjhcd8rhcvKVC63Ni91emTawczdjAzhw+WY4s+s2GAb
ertSGRT+D1aSx7i9Sl/kJeYBDbFL5zNK92UzrBs6nxu8K8fOl6AjPPAL6pJ+oVFRJ7s3qae+ekL9
RDhrz2PstYn+23qYxbYqihH0UYWMrL2nI+vYOS9B8KjtHy0ROr/husxc28yC83NucNcKqTcoWbwD
Xlc42tJpnbGn26D1se3SYNGdgQofU+hSW6COzjep+vkvOOV+XE+IM2SXL1Z0EisysLiEnItOtLyX
jt13AsRHfwmQDKjiLyPPFqMYBSuPm37r0YxlLhyIsbjGmrL1E3sDL4CNXB/ax+pERuNqNArz+I7r
56P+n6xeOb1Fm0nj52ylK9UqLSOBTwvwPLCgvbxvpJagz86b1gKKIQfVbdRuK5ZUzy5k6oMgkGVi
HKSWENa4pX/PvvsDqIXgaVD8bvVuWH+k8jQ9SKj51RdjD+0dsJij1Q9byViuIuZzWRInL61m3H/v
AJTwCSMcRRMX8HsyISZnmNxuxsBHMbmgKieJi0Y04nc7ZQat7ODMKaEPKZg/T7X0iUobIYlG3Fcd
JNhNXQ3MkY0i6riW9SrN8n/+5qsQAKbJ+GWq4yAnNL38WyrjcNVP7iMg49oQj+zRxemSNTsIRmeh
i+5mLiKx6E4oOSisykWn7dgUXbvCUE9/kU/xiGs/mkciUpjRKCTU8D4AC0XN9u/QvwbSHC9CtMBn
3pL6/HCaJtnCR8quSHIxmLaFHGMy9oKdZsJsHfoPUSkqkRlwE2rKPt0Jng0V4BLTE9GFl0Qgqh9z
msUAiQxzkFrN9QfhudxwheEAUCHFaWYWD3tNUXsndgR2jHyRKGUepejmd+2WTLOR8oRpHQqc0pNp
ah34bxBJPpmqiGcc8afm5OkJAhZMCL27M7q0ew8s48P1PyWpshfYMOKL0lld8S6js2JRqvbVMd+i
OVvwfoNOAvolkF2PMJD+7D4xjvwIKCMqqCvPT9mgfz+dPHTUfbSwQ0Hc1hH08vFoPTeQ9xk78aXs
83xpz43iXZfoo7xkzmurbgO4RDo+qWZDIIS9LYOcm1WkQ5VOCNWqh9zzrp3YzoYhZGtFvbdS5wH2
ipxS++ZaTui/QBi5zqCqmTRlxDhDHPHGizOHPATKECZ6dnKmgUv38iNyMweN3bricIbl8W1z37Mb
dtHyHz9uG2JoP/djgBO5Xh158GXFWcK/IIC5rcJvdmlY6ntIzcBSs6HnG6U9h7o9kOtHIsXpRrUA
m8M1tseJ7pX/5uf+qSM2Wl3QTM1tkha59lfcelbAAQA2bFaWKMaZNf0qNJrlcgOpSy9jXkxxqf7m
yjbnymVgkFRboKK0LZtq/2Z/b5E84mW7lW9v2B1wDINDdM5giTv3P/+DG7IqR8sghmIOxlVv/Wdy
taMRMDdp3PPYI4rrmNxb4OheTG7qh3zT7yKsAYNuGtivC4kSK01BZbypTFoL4utU5afa3n8JIxkz
z7BYdBPHB2akgVrchY3M0phUXrUYv/y//OBL71csGBY+tR1MdwZEr8ZUVG+Ds4j2A5W5t2XETSQ+
Vfv0iEBU53Xu6RUfvF6Gk+IDmlojv5t5PsDSoxG4Q8L8PZ/02Jxu/NWLmulekqocrvGnWISuvnQv
MZSOSxY2Lggb8XG1uLD2CZzZ5XT1s9cV4albPBP0HwXn1gt3wXkDTqOUmy83v85/ocKOnVEu6B3X
OQVUgXNMDamhReEfcHRpHZJ4M3maYOeFVo0Iu74m898sxkNWBgsA25MTI3IpgUP/x3DqriJFEq5y
8TEa9dk+72PENBR9ZIQarzCkdA3AE3or3nI3ju5DVXJcjTiQStSAH2lCqmt2mkezbhqgXW4Hjyza
VCBIncbIzleLi3T1xVyZDIBrLulY8fcKpPSL0ijPZ253rmXvpLZd71LeOKtGz5V+xxk+rMLl7KV2
akvhWIn5C3S/KqM04vaQPN5cPyF2nPTzqNfy9yKnZjUVdbiDtyMhSK7MRlTPf55iG3ELgwtCKu/3
uVx2iChES9nF/U9NgDM6KliwrZB922O1I98DLkQvW0m+GK+hxOXLWuSBeOlhsQ6fNTjE0v367ZTM
Tuv4UYs3kypGi9d4WNlw2BX2tjAsumFr5mLB67d4kQRDnmtA4oAFlUAr2xn4PKcmHnM+qVKZ5XNb
npZWUz2WwEatU0qPuMOUiGUmAOGg+QWVSWvP9QNETQUEjVPwBu4A89doUm53XmveCZKdPMQIxrgx
xKkGME2H8hf309Isyd55q7e1TiHc50mkTl+hfk3DtF/jHjoBXHoBGq+tHjykZHIEJcgz4o0WykIf
AxK47FAU7RaRc4HnB6A655C/nlsP5gnWbDW4X3AyNzUS2TS66EX6pzbAr1EHENGwVQXaabG00UAF
ejdtFSq4Gw3jozGUZiETuWMPGYB9yuF4o8qk+sq2MgCY/KY8jcT6Tr9p+KI3TiWsld4DDC8+iiUz
DDmyCt5hs5an/XlbHq9DyXX03Tx3KCwfuygrbsYT+8nuFVFW8VzjCyfzOVEZeUWLRkRvvCwuCr5c
jAGSbt1R+A/LEukcxUTImus085qCHLo4guIR1MYtlCNRqckkoxJh0B9fO3XyJpdAkgoxy4dAt83o
5asrrfnQL5FXBXfYqY0zB6pAhTeVBseO3JEJPe6fJng0qCqvvxLk0ChmKIsxS8kNg/BtC7XEyvsS
b3S96XdN+siQL9Sqxmk6oa7K3W+HnsiIS/C6QL8zp9+IeKrsT2tO7h/0ljS/IP29NE3GQ+Cyquvp
4hlJUZ7pIulyrhCp/A31UTsEDMtGWDZBGbGxX0iV4INuqGrYNSycu7CQBJw+G/UZDlWccise5m0I
VV+i/Ad4RrTEbaUmmeTibHQhuc4DRxhk+LW7nzykKJaQGTrYTW2Wqrx+MS4QzMSFqm951LWxRAaV
1k7ZD4rqV3kPgpkXblImRja6ihf0z0QtMKrB8L7iZ/nzVnKdIwMBoKShh1KdIZ5FtzyAlIus6nKG
z0PbDy/1JvnMxo5O2BCZpF9Q2ObX4kJCVJk1xMUyTgaywAt62FsXg3gqFQM0J5LZ0qVThBRYng30
HqpTV4G0YYurUOFfPgnvfOjmkxzKQK8zIOGc9aUZKoEvqNedjp5TplY2/GPD0Do7LR7vLlZvJXqA
3N7Z78XPXaXHFl/CN4o5AGXYCsll/f2HO598VNb2tzy/Wp6+nFYt5hmeZwxierMHCpQy5Unb62MK
+4qtBvSLPaqY045l9AWM/sS1QiHpWh+UVq59LXQFOoOK9rdUpUtbhMZOsy1xGkbhoNX/a5/nQQV2
xnVbD7Dx7vEVRt6Yx6m4LqHhAiJNX02DiX2e4xP2/Q9fQxvcrOjajvLs1LKkOCsrWZUEK+b3/wge
P/ePuxZ4OQj615OL0Z6mga0bW6OZtl5GDbLj9kDZjrD0OCcnorEiSh1kKAJjvu31yFxfOZVlWijy
CVMvxhDkQA5CW8zwfXdVvqQy3CkNo9n2iGHvSXpOqgsGNTqz2aTr45a4o4N5LV1tK5DrGoMT0Y3k
HRW+1oow4k7DJ7WJ4WYhlrfpkOnionAHK2LBQ2gYMnKR1uT71AtqYmhiUGqSsEsfLTPqODDyIzVH
wgMQnIUNrCTlbfSlD9QvuM0eKxRS4md29ztbRBzE8aJDBiNZRkp7X/HmhgTAXK8d06Xww9rt1Uy9
23/eJJAScBBFCW+6YjD1L9s8xZQwxn9RxQDoBKLrSp4/4lq+MeUWfYeiiHSw25T7ipwqhEcRCk4G
i5ELxzWXl7+RQneC+QalOR9QwEyO7hrn9S5vN6DQ23iZIyxbhbGI8e/P9WfG2VqHUiQOFRFEZwAH
iduNuNXWFxjJYmAZYQKAL3p7WT1fEUpJVC+vvhN3irZ9Mik4HzWp8ZwXygr6JX0igNIUvN4Z47Lt
hMCZoX+q2kbfAHM5AUEgDsLh+0TJC5fmEAt/vqezkMtxEFJM1tdob/8YJu+3EiElrTRfNHJIvZzp
Kiy63+xzG+ZJ9lp+Qeq0sT/5SOCxc4WBEr9x8kyJIZvJE58IcqgMNKMe8LME3/W5NIRq6t/t3i6X
30A1++C0HXKGIb9R3zRBv3jM8iNSLmy70xOCijWsO6Slg+xyR4nigR9K5wa6ZplLasxwYTDIwGuC
hybFd4FzUy1+z7uTFn7cG12U7OHT8X8Bzc+97IIPFuPm0aU4HjlgQHeFV43PxeJPOoYMvsci0PjG
cBArImYA+OsQwFsJyudVH6ojqPe09ix6U9MBxUFz+gfwhmd+HF5YrbemTvmIrjPN6SQrsHjbyjjD
eu5AgGEhy1AA+Pc0NQlcAKzG86deTgSBa6djjgVBJrHNbXApN9+gE/3dQ+qOwIojZ3/StzSNbGQO
6cPXmlnXbn+AdBlsWep29UqSZEr4pSnm/bBaTSIYLhQP4T8chjBDE42ebxqbzRLRIVjkbjHdvOsY
gYXRRby4pzOJUXRZgXau/y/mSAfVG/7AHS5tat9VcSvj1zd54quxI2qCxXlF+j3tbFbXlOhMMyC4
sOoQqOcUaDlIKK49DY5EcO+NZGZse4yhefpm42lFnb9ZJcZboIhTuaXMcd9ed94FCa5EXw/QngmR
ZBIkQ0aBwGnKt8aU/oewQqWtamYxfP6OBI10kWSXR2IjlwcqgmiksANxJzs1ZJvp5INBTCARM2YJ
EVM3PC6rIJOLN1YpFc6L7aZ9zVXvNb9P/HbfNXNzxvfaMvEnDN/2ZcuVtS3Fs4dFtrROXBqxW53Z
+wdXXEV6K+xlsA8Z6uTg74xhiiusEGoQ+S53H35rswlXGNednwuzYT67FpfQ6RMZv9+6DN+JduBF
9ivt6lxlEYWpb8uj2o2ZKMzQNocJab3D4eQv0OZkGpbE11BCpGjYTPyBRTjPCWvek0Ch6EqHPUpN
4CHT+/JCxtHYJX5HatgvL+ulzdQZP7PYltKWwHeuGa11r4B6/Qb+z2u2xEibnK4tIjtDrw70vwQN
LHKeO8KBqxH5aJ/nBX9fBe4GcuMcWdUBtGlnCs+RtF8TOJjN24RM7OI7QYk+FdYM4Tiq/nubhR87
itjaCQKDl8pxyZ07tdPaI7gFjRWhWKT+Qi4D7pWEaEVTyE5XuchHlnmcgO49VyrpcPFcF6Foojuk
OBbE2VImZzm3QZW4xt1APzhB+V3olHepMn5tzdwZeGHpvW6y7TOkbi52Sr5c40dMoezaSbgcRQwG
PvLWwgN55zXkBlN7MhGo20cW98Wk0klzLHxm5FXG6kYm0lzFsiJpgpZGbbXPmbfZhBd560aUgC8l
56avDaal6k0X26tCEVMjMcuXaWNRwxnw6TI0bYfxTXelUAJFdRkYyKGRSWocIuXqnkKDbehTQ8RX
MX1Shic5uFaQj0EBiKTU910uSy/qyMmeNlfIYlx6mdn4vk1xJbfCFcWddZHQpCP2XfjbN4n02Cfb
M7H/MEXErF+CI1ZaPJ1m/uky+c8dGXK4b+8afAFhEoPS90WRQBurJ4TSyXmzvKZ2racxSq1Y01Xy
9uJoqEPspq+aLKrHg+eyoq101J1fGMCYiOaEEiJBHlj+XigxvilzIQA1Iooj+DGXT6d4USzRwAxK
BXpUOEGZWSfAOGCrAa+BFf6Vbg0wlSdDbmgXUEcX4t4BQpvU0ndne03GCZ5zZPJCsbBOypJ8AL89
Pcle6TVsl28zwhsyXkF3ut6H3WraoGBSCJuLdp+OiHC9GNS173nnR0JwRCGLvzEI8OEzBrpkN3xd
LzSV1DJmAysPqPFqqGvSkbnIm/djxhSrZyWu+12cSAzNS4opuDycIbtmeQoaRoO06bL5zWZgMmLp
sXdVvzhcV9+0DxcMlEATmGozdzQgs/zq4m373jbylkUo8ajRt/U26Q8kyonMaWQszxL6/LlShdC5
eto37MmjdRKDCOkHI4cyjG6ra7XynzgIbS4pNd7BzoI5TNdjMRDSoNgDI+wQVoaNwctT5F1hGNDi
mvHMu0rSCzlT84DH+v+3+cXoLQyPXXH7q6hr8tdCAwIch3bVIQPQGDflCUOKp1pc8rhSYLC8dMYV
40SPIH70rkQC+9NTr35aK6lZF5QUp2auV1xmmFcMfu7yYcFP5JTWHYXBrJYdxBCzehjyb0CcPyzX
1r32x1t6UfEehiD2lfk9xNu7hwHWPRc+E8Jzpa6BXeCeR68qa1m2twdcSpeDQBYQEwBhQ+b7cBUd
t7OEALM2puGIWWJFbSaQojzGTgQu/Xi7OEyIaiveIR2aKRU383blqO9KCOrrfTXd+w1g7GoBy+Ur
wvUQY99hxV2ZyldcPENFl8jDrUG+V0fhLtyLwtXMq6VizmvLCA9xGybr04C7mQF1ii+qiqmMqjMX
GLSsZvK1L7Ex4qfv8J/HeavMdvmfvTDZp9c41/AhQnqqb0N27pED2SK4w+kDM8O9zcB3qnWZ5+5P
9P+U+2TdbjGzXVbduRNE+DLzFgY/tjKISnbT1qwXCqWvsYfnDoh1BKrlwWdbHLyGsp+askdu1XLi
hXTF3L4+AVtyUC7Qf8VZCTNKKvtz/IYVQg4pPwbufK6DfmurDD6p/gmHkxfUfnVefRlt791h9BPw
7+4a4524/M6Wl04ocY24Cie7rr8QJvjR+m5k5FZHortdLvcxHemrdOrmd+xooUMwM1x052n5oe5W
RlTR+wXVqN5c0Kb4Rvb5JSmac9/0HisJEFBNTsL9JVpJQVh5Q6CGnK2cSEtpNUSkmZ6L7fMYOhrV
7G6WgF3EaL7a0GOhzPq/6HLKnPfrXhN+Au2RsJtogUMHQ+MrGk07XCHXgxQYTv2ioMjcbjmwCW6G
S/gR1fsT+BU9cao/tZvtdm7tgzSdvbVXUIjnU8zkfBZfrBZL+j0QLHoXlmm0Cg1WMbhlQ1etPFvK
UUYD7NUiTCqBKQqXnBpnQjXVZ5PDK73DnoJqtV1QbH2FMTMcq+MqOnbRuj3tjAp+0jscLo5ln4VB
oWsJR5weVGRmH7znJk7cb5n9eGTCWuuebqSuOQTBeUn31lSVm0r8mwhEyGI+pUaxEDOLaD3DG4F5
OfSDUsB4TBbN4CCcQKwwE8XP4TyThM//hfyMl4/0/3pGIGz4SNxJ1ESiKuM24BPwxY2fsD8kgvft
mQZUgZpULYx+erN5wzl+Yb7BuMJwo/xAi7pLXwtfHvjrpZtyPVkWNZ1EyAlPkwroCAAl7GqVe/d+
KbrLM6SIsjS+GWTFQ9Ni2GGD5mMulAlb3CzAxQi8bdUYMPcGRMr6OcM5YjEMA4nzafHkecOLQuIp
/NbZzy6WG7sqkHWlRpMBB/6QVNUFGn7c3HVjU7DlhfU9dMpZrY+KsDYPQ3FRX5LAPYS7ZRzKWhr1
YzAZCzUdw9gyBljkF7OOgL+EsMAhAWBKSEzqLdXAqiFXjoUes+q4cf52W6Pfro/fwSnOs4ekkAKr
h+eLF0knCpyTUub65kF8O+pILW9+jnOVYovSum0j+FcUx5t+lL8TDppuQ6p/rZqBv7/yl78Jshp+
Nj/eOOpbI+seRkpKdUtQXRIG8y/1vyXRJeduIiAsMwHnj07J+19YHJLRB/nVtG1UAY2Huc6Ei6SG
Xy8Tp10JDcxsusZ+79f/owxadjAs+fs750v/iakCyiTGYvJ3x3dGLsKSLwsRD7Esw3LGm7pDEHDt
GwaAwkkh3mONlzbQRQ7raNcvaSm0kFJ4sKEFREl75JjNEoCYURyppDfJq70BUjZgnA6fOetRn8Et
GM3tNXlG+XUIMReixpaOjMDQV+//vW0PJ2TbFy+RApdkPl+Fj0WMcFj9ARH5X7F2+CNuai679eLR
3ciwRgrpHSsYabjdEavU/YlCfoB4xdmRp2ZQQH1UgfBuYZZQW1mmiNZRzhl6NLLxq/GIPiDMeW6g
+HEtF6WIo4cj4EcBscYgirwPCssR0VAaJc1Rk8LiJ0G/2HGKUFOF6KxwyGehcihQ9q23nIvHYSuw
eEQ/o/L2jQmOa1GtCJof0Zmyo8LKJLNWs76sJMFTSSGU1eblqrFzzgbf5SH5+IQ5xfAWEV5Rm7lt
byJzFSvHBY/ESyDhWgk/VPx7wgYTOIufK7BBsf/u4yRsMBZFJPR2gxkwgJhM7uEVSdRp508p3tfe
ox1PWIsnRrZx/BXme5G35Puj7oPT2NWo95DEkhB1WTND8dNkGKJ03BzlSnZfEZgXzUTSAE5E4w2J
YYd4Zhvg8h3HmeAqN9Uh48NGngl/6bTbrrfARt/wMaR6+lhFJ78usp9RyCfP8Lzfs7epZzIJFsP/
XigOy4qo+g9ksXwo4/L3IDsOBbi/YROwUMBhnb5DdIC0IwgZoFcoIe9nhpCGNDL7QhGZTb00S8+0
rPkyGv9LylloUv86PyU+t0i5dR8/mEEIl+N7ZPui5hzQsQPhXPls7R+lWnxGg9KulUMsIJ7IWcMR
qYvZwSg09V/tppv9brsqFXEoaRoUyv+KKgLgqUEKZZ9M5KDG5qAx9LbHdKXPiU6LWiJkM90MHYHr
Txdd4jw2Cw2PO27aX/wGK6Mb9k8DxX0ARoTI60sAMzwx3AnLb3EfilOwdtAIFaeMBFIyKbBemJYp
YxyjmeaY9sxK9dk/464qUpLj9XeAHf7VACjyE9opo5AsXLXxMaxvoLBxrtAlwxV10Xt4L+d+HjKl
CLKbSWQofaHFvXiP/daQ30HxGBJqCWQVt2xYt1QkSJiogiiXe1s0cy8K+DUO5rFBMs83rolHYe8Z
Lu9KTANyP+0DLwPWqX+cqUD63iP53R1nVJ61yTT8XFYFchXIE6dBQABLtnotQyYzb5YXr+upmLHt
wcz/RjXdH/ryXhs2/Afi96IK3tAWcMzjSST9HgAKmoK0oMeFSOCUCXOyGwSd9Aw98tXRzrFPy2h+
tBJUDbnkh+TDTlqRZyUxJ/dCe9qmWrNkK7gjSzufth/EO82LBpZIGZEhITP9OtHX5OBk+Y8TQMxQ
AJrlj0hBTwaOvVzfQ+yW1tINR34bUDdSwNr2zgrawRKVW5RliCrukSmCgp6UXtcx7cX0zhtdIj4O
rkUtDXTX/GQXfnU94A7iIAWnncitlLMEXVbhk6EZ8oH9POvn0A6oPIHSWKk/2/c5IjDa8773b4LX
ZXlAs+jFRcysoe5KOKjVTlQGlAP0+2quN6HIdV5ooMfu5Z5BK07L406G9OpnAL37FXkBepA7dso+
sqrGnLNt1Scvfmn7PBiWnZLMKYFb92hpnmChWeZFYdvCqjlZENiMNjdVjEeR8IXhU30JwcLpgmHu
5sO3XqPumYb6icA6URzlThMdmEesqvL3XYdHOKPIBHd+QUbWadMdGOWx4Ia/o21ZWysdLCVgOskp
0D9LCcJGUO/PhWfjo6vIisnM4yJDhMfN0x9zAwmXJcEpkvJQVYfzwa4TLuKeg4gnBnrZ7kXqG7Zn
fMRgXW8oG/BfKe209sjuhndY75HICAYUXhUU6UZ3/ki9iLgy42nVFoZU8XECLBN465NYKvwGcCU8
riB2P19Fa3We1h6t+LlpCQKTdUjw5OQctEBa2EBJ1OLyiTsj3eknTf4/7i/eNyGdo6UieLBUE0HA
9uWA/uFvR5p+qbRQrppdHwM9v9TkwsLLyjy87nUHSyb9MmXYlbuBPF8rXJMf86sw4IpWrcNpSho+
lO7MjLlMDgY4i73FlWyLQQZJ6kB9m8LZmVfq8Egkb4+3acJ2F1BljUyY9P7lNz4SJnM1Gs5H3FPV
t8g/gEZmnaaPwcpEezgbwOXczjrojr4JzDJm2SOe0gwMhE1phlqmyGosw7AJj3wpk20VONevzG06
iu7nWoFKqGg4zDf5IhwYPrW8VrsIWGhBQU/mWZMOvwsnjQCKuJMoIkpCnviBA5wzHru3s/hbJiLP
C+DGBXGSqgVl02++IPL2QhwceGQubb0VAVRdJb9dqgTbVA3UUMdiZfCZodHBpcj72DdtdljrkTYk
VVvFii5iOBjRqYBIQpTR5+3Y7yKz9nmFaXUmIXR85CGNvI290Hie8xhmzeITQkXAn0nrMfEQEm/i
O9bsU+tOeKdGnPj4rkfGLNhb2ve9oEVDutoinjGZZ0Y3n9AP0Bc2jj7rWelPadYjlI2G56sA+NM2
nAksxH9eMckKAZJORXlivq0hKEOTU2K/rM5Plme7qPmEGI/bK2vC3q5flMApMGUbwjYjqcEiK2m8
JI+FSl1yX9YNfjX6UiJCc3QVGIa5/5jAFHCf/1gFS47MNjQ54qj7edmbRm+WWY3OHy6Ys6TgyfiW
v9ZEtTze0XjFPldP6U3JfHNexDbhu3I8K4E0dgW7Ie+U1GmcrnHMuaE4YHy1jGjJj9Ko3lFut7v+
hajwMVJbf4zbUmvhuUG1sM5wKH9FxhpD5YtbDZmFi1P2Poo6H8lSLjhy11J/9TWbL4yThYuf8NT1
Q0vAFJPsAlJupaIy5TukpbhyqPI2xz5Flos8n9uow6kPRP8JU/MtwXGBUn009DzvfX2uQrHL+fg5
8gyg7kWRTIu1EB69SGjO+0DcYMvH3ioPUZf1w7ordohmb97R7AuTOD/SFRB3VQd9J4ut+Hb9hM3b
82EXhztH9Z5bRmaGORvrvO9N17lovZmItE5fbnxx3cCtz96larVrstFlzJlZYkDA1NWHOIZ/YSwS
eQ/wL1bRb2CjJHUlNII9CWzgcRogKtVW8Aa2pIQL8A9WTiyPDGVtF91ZKrStApjBHQX7DtoGhd4L
LuiUGIhgNTrxB2hLuM//x/swbkXvYHmoFQZNa6CJkJfhnfcX68d0vrFY0cKJ/jKsSK//sY5Uwr9K
Oqw+FiwU9anLtXxtkIaCc6CO0O2e7bdSSxVagcMOAnl+boTHP9P60nf32ByRvTaKCFVywv87nEUe
6Fz3L7xf03h2ANh8qEJ5w+cacgG1aqTNnSwwvj3YXMY1Gue/0aS1IE73QEVRfx+3d6KvU7+XVQDU
HET2mel1R8UnoYFgMw73tKNL8bpQFvPMQRVONlwikQ2NltXmb0SgvhPYlQ7Y/4Rbt330cim1ORe2
+putPxgGI6lu76KlySmzD6J4/btXWh1mTZoyoPmWu3xWttNDc93/iIRW38vFjSeg+T8K0cLNqe2H
ZqGAZb8S5qj9thZ+QgAauch43VoHhpSRuPVEwvimDF71SPxXGft1EIfapnlZsF4zWPMQlByYERBi
/jlbkkbqfQ1+9uD82zrXrqgUQFSnmGFs81SBSajFC9zTRdZd+T3MrVlz7Dh3uiQhm2hU9SPoBu6i
pYXezVs8F4YEsACZTXzuQ8DsTh4YfK8KA+5St5iD0swR7ok2RTIxWAyCVPCt+u58yp2Cll8172Ys
ZkYdi7DhApBEOxo/SoDw4/Dy+nZ+P2204Dmb9dFESO6UXcNAuvlh8q2gb5V84lODBJm1MvNvZ64r
VPLi++ELzq8K4dJdh2yqXHkbMKwy4kA6mmW7kC/lEvXUsjFCDoSW2OZdGOkxWlESd0z7XzTjs4CC
eosK56NLyp2Xtz1Genp2kmcwiqyUCK+cA/0NaCc4gu1oK7rqzvzlvsDsQN5JJes/BkpQBA64nyfa
vRC+1nOA/UwGQpGXx55sjlTbc9K+YOO3QjQSDNf+Qxv+JMmB6lU24JbiNhFblcpOmG02ZA3HpkQy
WPNuklYHQzNLVM162FgR0H2SBBn1dMGFTpO/lhE60COG7NFP0AiOwbvvk3If8aHe98+ot85PbMPx
T0UT0grqnbu3sAvUuNjgR7uzuIvJ84zjV8/qY+yw/DWTBJHroQ9hnbll8t0xJ5tk0emSr3dSVUjw
PLDdEsdrwBQ/Wsyau3jhPJSXU5mMiv4J35UZgDQqV3uVsKkSdjC6WCnSdJpfg/VdunRZfg+E/Tz/
/7gNLskcGfPx+hjbZKfL2fnCF0VB311Tav32VO3C3Cf2VTIbtKV4u7jwq4JXhaAE0B1LDx2dC8GJ
lwZFHpjv81CQr/0fQpm9MctsY+3F1S5Iydfocqb04BWqv1rmn+Fpb1eS1V8raUX2Hnz6V/7i3wEA
yGQ48HbqyjRFs7ZadAqu46buOle4jO8mJBxPNPLLbrmlL/CWpO+RxXIwtiKaRUvOMTulm/8Z8XeE
0/l3QlTqzKIrqGD8FhPXRUGDeLD+Q71APjjoG/dKyGL0BS6363tQNW9+B4MmxXEEvfkjLZsbd0IJ
NjuLBRS/RVdJjFg/GhnSnt/4Sb1IJrFy0Fe8pBE2vmdRjJZdDoONoSNxDt9OW13dNamDLd6cbyIW
8lUisTBA1/hGZepMKs6WAU8ZoY45PBU5Ya1oyjVNpXtjX3vDuNF0izBoWHErP4FcFEoGc6l9kLOZ
u39DrGk1T1GMAvMQKDzeGhOFnjlVeNtJJuwhl1bMOJLLu6ThDp8dYVCpG2QVfQVR0ScGGGZvbjLj
M32PsaVrJeQoDRX2OLQy4JoT5R68CKdn98Vife5sg8EFXV8sq9jDGm0KhpPTD7cRMsieYJPDRf0m
pC2gi8rXhXVjVL9Nk9kp4RiGQFk87nq/V6f0ug4qIXClfyywLEoTKUsPyHaf5zdqR3i8x4DNhaVN
UpqqwVX9sCPB/51VVRgb0ruECJ8d0F3n2DPJsQtTtck0i/SarRoLgKdWx1Mu29YFXMpJh2BTNPMI
GnaFbajEMLq490k7aiBkEvWBusvguH2y+IuodQ6bLH8eQ58t9CrmG+22COFWFnU6Cw8g74BXnTbH
/mmjnTphMlkkU5VehpW+xSoYmH743+G+uEwpNETLgf9+A1yUHozuYu+ISTtuExj0fWvBchoZu0Bf
bB4u29SzufLY3wxRGjfklomxR42BRWNTeqcV6A7XyKrGFnFcTEkbSd06BXv/sSprXNASnqix4xgc
Rkkc1iJn3XmsUEUmY0fHgEaoMIRd/8YBwJ+hLw2rZ5gAQE1bq2IEIVEKxgNymxnJco2dbIkRWoP8
nTMEqzLeqsgXJTNmWqiIBTzeWwn30vnvYKlu2NoOPF1HePk1dak1In1PWD69dT6MtD3ZR2RgGqOb
Xj+VVMOxlf95uoDNgjVcE7J6ztJCZE2cLb4JX0hOFG2umagXeXtbjnPmGwtqZ3HuzAiSc7QISeD/
ru/Pu+Rvw6a5IXEEOBaw9IAo8+P9iJ5c0eDv3IgNqbvIu8FlXFUc0Z/+c9++HxH/SSRvyqh9yfLc
dXu2HGBGlo+jy3WDPf0ZhlA7ztwolGu3b8invrgJlUF48HoCdDN00sAQYgcBdMIFXGKCT7lkAExt
7txojahyAzTYd+27Buz2Z4PKGA5N81xh5yi9o1CU9WFflR/5steekI5M59yDUeMllWSS4mxg1oKy
A1V5AyuDf3PJA95aepSWMx/GtmUaWE11OBI/mFgTaCNmfP9AvGz+2WrVvxHEc0z1WkcgYtWDnXgN
E2/ZKK1OMYbY00DFHb8KuLOmPRVINFJGJkF9lt9S2kXvX9eWAFbunJOCaJvVguPSWiIU0QPrU3iC
/mkKiHA+bm77xerLdYpduhbNbDzrZSIJ+fC4UUun7yJl05hsvHotj++uW3Ks0MFhgIJYqk2NN3Gv
QEKAiXmXhZ3O5Tl0s8s7FHwhIhUqDePntA2KN9rZtptayZTwxFHHgSIHbaEFTKvfH7ZrQlZ6Jz+B
S1vvahV+ha/YaR2E6ocDbqTZHbLw/mfZxYx8h8uq3lZgkaAqZkgjns+DqEgrOMxWA8KeMETXV+8C
E1U7j6d/bNsqHSlQ1wi8/XRRzILNC80yGZonE8Wyybn4QaoASmGNeV/vhxe8jOAhiJScODBwFMbB
MLRyUMRyFz5/W2JEI1xljDkv7ApWzK+rMdpm13AkTHp3ItolYiPhWjn0E+ZsbjFfm4zGImhzJvA6
dmfEyHsN1gIzgk+1iyExr/UJg+dXAzz3LHf4g/ACmp3pDJLGCq+/s5SmS5ZCwJkV/oYoQwGTYrmh
pvKDxF+nWujEZBHwJnJ6tC6YMpqOEVidcRtzma/6toITcQLqq9CiD/6nfAwZxMMwgKSUHgcm//NM
y3yHN2ecfkSU7NlKPdrf3YMWtDumRHOe4+MYuh/HadAjGvOYUR30IVKwPP30wn/HRw7PnnIa3J9p
4uI4GMDzmqkTerBe0OireqpYGrBLu2eOZ1Ext2djwAZh3I9aslIDaYOBHgi0MoZpVtfH0Gcbn/pa
2gJ7iV+NkyVmPa9ox2wGnTHkw+7FU+M8CyyIuGv01JHX1kifVBL00qbW1A1k/8b9cbo94L6RC5V+
dUbgu0EhXcdqtqDNVtR/xbvMsa2qCDj7lNN/eWa/2iJSFaR0d+D/MJ8z4lKGargjfPJRdxETrdDD
fYP7gxDKNEVjJPqTO8py5JnOB9XehiFQOaUb9ytrjKvZBWogiAP+5p6XW42JJ8JdBJtgv4porQOb
x7nRDn5t/X6jjAotOB2J4AA5aJ1RN/3isfC6i93aJvAOPd06mHeWKaCCQ6zGwDfK0KzXVL4Yci1N
nTXbSsfyRu2MH2xwciELqZR3JiKFq7cXaFIJXXbE728o4e/DxDEw8P1+K7J7l7Bjg+hWfSpcz0ek
PCLlCmRWKr7kNtQqROe/zE01C/ILF5ymjH5xV3ALvUmAbuBQcFyBP3MVQGXmbCko53bkcmYTlISm
JnhwlYkCRVhDV71o0OzeoN7rjYpvwsuszsFvf1oLDTJgN6ctEdqH6tLVON5PknZYUoAyqAjra8BT
1uMvjNIqsDztRhg0yyT+lbe3N095V0vJ3XvfOkJIj3EWlwD3/eHHPxudl8T9Wzk81YeGAoq4aBJB
3ZHkZ/XYASaVKUGXLVpxdJxWR4DXXfG4tbfe5s/qUBr83Ai7zIjrIm6TiOKSq18O9PJ38t0646IU
7bLz4iA9rpbL5gAmhHAse4hlPqPNK5EEk25pD/vCgy8OTLwT1P7J4aPeTC7afsLzVoEP+rmC13XS
PI8toxFeJ543QJdiXeWr8T6kFegftplCOVom8kx4DuOr/dHHz1kiQCUIqdi9mf1gaZHZemCYEUaP
+wUXoZqbz8obbCROYfqHbDJdaDY12xk0yhMXgW1ZIxBDsl1qjCQhIUIILNJv90pOSm6K1CRh6HtG
S5hea29Z+cvbT5FiBjiHTW/n0Kf2eVBQzDGTivphfgO6QTKAo8JG3305+C3cPGNcpIzN3buKx4ES
7u+OQvW4jbwYzMMZKTcGtZ+RCqocN/DYxC0Y7goCS/+9ymcFyHY22D/cadBXFmCW9n35pJuVB3VP
ks2ct/qW08Moquws+BD+a4GJXQtMaZtVriPok+1zo3R+rDQOxFi20nvBEdJ+XfbmONB3pQX+ytBc
3jDinvw5wheKQfeM2h33QPnx5uG+peeso8cVbW2MViutwmSRLenb5RbKX/w8ONsnJbPlpV0NPhBa
pHYub6D/f06wuT3W/KJhsAkJe4mBG4JxBQ5Xfn2BDvOUh8Jlub4XK/5L7bLrDaxix9ksWcherqXV
UpFsU1D7BMzfCLvlczEfCnDp5YExc1SnbzkUihZYP3urvze5VwUHVL7C1m5k24fxpA59QXB0z8J/
oc67vVYqB7stqykdN5Dlkhs1u5coM9iNU7eO5M+HOmOhP5i1XSb11+3MdcUvyHgpAaEm69fzfdSf
hPnhY+X0pyi6FBs63nKoGqb074NgLJKUBQ7pMJ18AfBs03w6TzP0z5GTtmY4GjKE2PWLfuiorWbD
w4KRYI5IjdaqC6aBWKBjeMyA9XVfUjphKmo1x0hs1snw9x+esdc77WxLYDpvKwAMwqOtPcE15pby
0hGtzxxcWHOSPtJbV4hJcNmvnwjwENPMyvyLsUSSdPQ9sFvdBTMhN7NJOxqmnor/ZIBz5s7SDWLN
VVhqyTm5fpZAuXul8AZN+5IPQlSIez3A/+4QGctfwYRnawZ4NU4pmPQYvGpI5W9n84ZSo49HNNMq
CX7g+VWcQqSC6xSgzrZ1hk8HqxEJXPSDIavXMuNwzFNKsYPRrFSDGUTeMb/DQNwONvLumZCz113Y
P7q3Gat7kFcDNu4QenDMMWobbnG4DZlcfprvS9RyeID23GKjHDfKEwAsa9PST2yJ6ibI13UMjDbr
tOKP+tbAGUQ9juFph94KGyaAY4edt1qzk0JE1wPZzQ/8bcmcwQfEYxLPlBz6QViFYJw/FXcZUn3T
ZuNndQMYmfBRWrFaivAUlycD7Y+0qcz4fff65Nz5Wt/JPVMCE2hGC0VRTOPJCsjGXv8GfXR2ZbYy
mjJpC/4iXUJhkrCyKJcKfomsWPVF4I73p3shjFHtxhKV97//4oexZFFhKarX1nwIkDEVDF0FDmt8
RthA0Wd+H4RElvToiPTRrZbFIYkPrYtPa6jdYXB86oJnBfB30Rdx1E486hCpw06f1fFVi6l9NHTp
hxhuMy4awbDmjNSZEDeT3WcNTpedxmnGGKvS9Rr7zMtzMaWju49xIG5+S8N1B3riXBmRYwAaqrwK
R1+3U4qDDNVuHduNSxn80f2aA1yn2CFSPYUPUG4ItEXjJln1wdoSa/37Q3vA5yullynSEiV74k1D
KGeWMF7/bb3gsfRKumimQr7oo4gWRkXYMYqRC+hviNfRtSLQYWyrV6ICuJ8BP1Elvci53ORDNUQS
FuPyfp1tNc2DId1M6NDZ8Z1cF8r8Be7JiLUJvhK7AgdoqlK6A8WCkXt82PxDirTPm7hcstBhLn0/
L+t8cFzsCEeGESsCzG0wjoPjlMyoS8onkd12hnAh94VhT8qkwPc2frITQbee0qBgiHJ7Hw0VaVOr
rlG2LQtqhTYODbCIfgjwb1FdqTSJal5Wc71QnbFROO2B5BuIoJjSEtjc0X0XXSiFybM9jlycHvb8
h9kQB8XeYp5g28X+D60e3TZPqyBm/Q/k82T9OyG4ZU+UzDVD7NyLbD9nwcZx1z7boc+s/oTE49IQ
rcIoiJLB7oHqoCfuHYqoWrNuT3VJmvOdGM2pjyu+cYjAbc+N6gnI0XZaZ6dDdhCTb4DBbdUyKVTP
Y6EPS0hh0nRsFrMXNQpwBhD5ckFwdYkjYq+NSQjePdU4EWyiZKE6bk6Klzi6/SLGOw0/dIB8TgCr
UlgUJnb3+aHsMp2c6a+S+ds7GbTqGUr3UJVwlqx0/uLyZAOHWgmcGszPVjaFoPmR9rrLwcBsIfzo
HD1C+gJ1w/9IP+glHXiwHYv6mfgcnW/0OfsFKk0lO7YZvWBVW5/B76FdR6qVaB8oZZ9YLFx9sG3f
h+OFO388wxJ9HeI4SPudIe1nu/2oleLdy/fUGHpsJG9GmsUhejGawQbQR5hm4DLsJm5QqLBaM8Ol
2Svr0WAKWZ1cLf/P6F9f1YAO2YLYofSxb4m8ciVgPOXbwA4qeZGHsBSDk02FJI3/Adz2Dl8Dccwx
H0sauVr2D8HIDTwv0gsYhx2D6u5CPp3/sMHdR4/6y7pD0oau4aQVxUMoRcWBRx7MN44BQfM6navF
AMNz1QSI4pZZbfDcRpVPQQAPFMGFp7VSi4vexIJPOgUhKVmvvVcc3jphenukwRI1AaJwAb+D+RqS
6WMcFxzNJDS3ZDY9SGRmR0OcsgZsS4yKn0VzUcMF4DLpSoZWA5FPtyhQpK4IcjGiHUjydAHGn3+M
1802dW1H354aAw/CXi/wNPh+vMbcdLSPZV0M4OyhZRSvDKd6TSslRKuni2EJoz/wJWEybQaX51Mv
O5qVfM9UifrGWb185r0DocxvueU1H32JmT0Sc10y2bEMDx6ICdEmX6bhwGYDCCluJvnSwHF2wt+7
1Le/cGWckgPC2R7wRW46rZX+Atk9gZwbaZBmYlQck4A/bETvsy/RU9o4jfTBI/WEcsppbzW2DU2X
ELNIPgYULzf71dqMPrISONFjiG0w+dW6x0kcDZwFXXyQ4LiKe8DfNsXk7iw6ej8Ow2YPW9eEi6zl
I3PWB2yNiTOHopgNaGJ63z7yeKGiko2Y/S1T8aZ0ZrXwvd9EAdJLeEKpJSON5MwPVi3s3GYOOwXa
H1sECOmQ/W2wHwDsx+QpPFE4EKzesh6V3iEz9vf6r+yz7+NZD7EX8F4ouiVV4qU1dB1hkBQjWZws
2rfCJEVizZgqgPwwX0nBcBa142Zdt1Lw/MV0OU/g15fYrSccJCizF+bTWm7P7PXh0tvXGhCyXxac
ddX55INkiR3Hf2PdqnYcUKk5eM9Ri3iPU2XR6ramYUXEtdGmexFO5EXYtE7g2hlW6kskyJdoksIi
9FxKB6BIlWwf8NY7B/bamyMDp1sHlsEsNiD7d6pYhkYaHe1TW2qkBAIKbr0afjr1aOT0f14YBLhU
BLs/6Psi+heZv56ohxyzm+Lr/U80Or05BSdLOvv78EmBhgPTwP1DnWc/gFgrqJ4RKUjVJxOD3l72
W1XwYVGkNoV0OL6m8w9MaK22b6At+BDcWIYZDJUugVUT9F5B9PuplAPldiEuwD2j4yFSQUp2FFVy
xxeSdmWN/SmkT8+zWuTsmyChLbY4YefqfRRR0pCsBy3AZuJWao0p52o5ODJwsFu9adnE2ekQQ7oV
+YX2KSGDkalgomxdHFcOwP8l9aq0td6nU2Q7sckL9WEJRmz63y2dG7LixIRdkeCG1jSK9wkFuGOj
gvysC3Sd93UsTP3oNN5csjYe1iKmbYbkKrr1F+kT7ayxseGrgpn4ASsr5xbVUzt2Anp6bb5zS6iD
5sdZSyjNFnlkOWqt2L4zQ1FY4WJO78PmjB96FsiHO3lS88e+ljadYd3iyyRBfbKKowix6kJmIYiz
NuBRYeK8/8NzQpp1XulvOSosyv0HpygN8c4dtPTipFTT4+mkG4WW8du+XTTcLMLsrBkcPOL86TTY
d6IakPyJs9QxxQG3p8G7KSKcAWD4hiXvnq5W/+ESh1f7tFaRyHQnaeuNg2f7IbevNYJga5VHSvgM
B1t5hFHL7u1ET1+fVHbDrfM4R2ZatkOeAhNMgE6/z5WI7+cIPJkqZqCVqdFDdVtmciTPoR9C+hKL
6D/d44Rz/cDFwffTnqHrH+WbE1fHEfm/2ZNIaingV7w+7vGZ83X72ufOmz6iP8FYFU5kMIVJL3+W
VBH80p25jCJbeEnNp4CNX3JHPwJMcc4skyb6BbMWsQz/hyBQuJBRvURWAS/6D8fP0spHh0CzuRAG
rkxQG5NXTmvm9xICxrpJGWnhruxmH8xz5ujPL+70BTvMPipdo85j/bAfXHRXBiaeV/SqLLc/w/Zg
KkbFkinnC/lF/Frp2vQyCIoHJWhd2gVTcDMnJ+jQDHVSvvl1RC1k+QVvCNlxARgKfJ/P7jPrctil
CMhXHKal855xhhiK/brY3aHFTKMC8M5l5gdxJOZEAVxWLcvYyEKXIg/ebUpi4CXUaInO2i5xQuX5
cKhtLOMG8PN1dpktrOrmJx4+nOZRyWCgInYx2M5GGA64Xbs4OkHewGf6afcq6w9Kr0rxv6+2qcqh
xjmxZ5km20JJOfk3epq/retpyh+Ms/AXP8HCamD4GZtWD246odCUOA4nm/DSutsh/xKcyG0bnsZq
am60f2lx1+HswBgfeQChHASvV/K7Ljz6Xl7aaO/lEHZNIuep7SBJE1jJc5nxkxQUTfeaL9nT6RbM
nB3/e05FUYta5AiMLkBrP+dJyuVWsPjeh5Dkqawuld2axpl8gAS1vuwFs31wQkuXMBvGIJTwUORI
Q3K5GHp2vhcjWmFpVQLl401tlzMnvjdxp/7LFJS9g17VhgF6MsBdt0Gu7tjWJEoA15Gr0ZtPijhZ
uik52HWZfUB6qMPD94yL0WBViHXlLbUBVCQhyqm+uQ06EBzpO+TyAjWR+O+7hJ4QSCjaIwb+QSMW
GBJum4OAFmUvEiTgWPHaWdAWCTYcD4k36egURG8lit6yOlBJwwJZVXDSCFuugBwEFoO08fPWIC9n
+3ZR4nag+TX5pt1hLN0hxM3ImYjJdyPYtY3U7J8Mk6TCs57syGeaIV5VsRiBdQXdq34Fu0MHUMkq
dOFt3fWTdy0Co0u9OkVsxThEO04XX3aQlIL5Tgtx5Aw2wuUbvp0xwbNBylNFlrXqupYQVVYV3F4D
wInUMVQygQXNtRzzHyZ/aVYk7gOwi/6+D+57Vv0D4mxcj2tTNbcq2uXtBcEVRr+VcVAqhYJU/i34
CER2nD5TBFb2u4O02uHUYwGBh8g25QwiDhjqnWE+AhOfMr0KnHLCAKB7LEXmOrqSFyM2ELrg9Gq/
MNfu+b5SZ8i7ZqDkPTEFSGvCvJ/lYjF/8brU8HBU2vblR7WgrCVw0p2AoV2X+nTevJRYlwS6Mh9P
CsGRrKDda05D1qlE3vZlM0MbOz2OIMBsWGEiwgMcNJf/zJpPw6+bZIKeKAse+rnqM6nAzejkdo9w
VaYVuAgsYaegU5YsfFKUzsvhySRPtSdglhPJl6PQQXGNpkNDLwDLvpMoqRv/be7BnAtQM7WRvlfG
WRMmLLddtDU62H6HCaPSYaNSCuXodXfTB+AZwVKF2Q8crq9Lbgm4BV/Gdm0hVE5EOLzMfNdci+Rn
pcfaToPrEzKiH+6iOnl9dD8QMXDKm6tiHkd3PuHTKdatxqECINjYr0H91D91ttuAt3GiyxERMLk6
8uZx5GfxRERbMC5ye2KuXFyge5bdLvA9r/hlSHkghFjEVWi55IcQ4QofI9nXFL5dgSoCi2Cs2vFO
to+tJXUtSF3MPnebiq9FSM7jELRn/dQGhJOhZKNzzOJRQvp5tzzaJVw1wrvaTY/EDaZAIKExmmy6
NRRAp5uAbfpyOspel8Adkvbu6O4D8hZ8eQmkfWZkmNFmSzXDQ3KgMn69ttPoIPwsLJtdf5/op0CI
tKngkP0AXvaWhaSDyLLJCWdZGPVJ5a23iEdW9ujB1kutsi+Gp0Lks0s6F1h8mU3PbDdve3TZaOKL
6v2/z+El547WhrfiVOVJuMQ6BAiT5pnTCnb196oYkk8Yl9czsYnoCviIV58c+1EIvQfES3MQUKk0
b0dszjboiHG66maU9pOt2wX4qGorJOfAqKUnqMXEi8Q7fitaWEJCyyCxS4vHc7pWWCoSThR249ur
irKVQuXsI3f+jnfX1c7e8ax8l4hW/kiPz+6LjB+w8Z9c32McIB8JhRCH66OZPTIv8jDvD5yuaEhC
cxQwTiRjILgo1M1PQrEtfTm9qdSnkgYuORFCPSdNBv/OJSr4yUWlQW8W8EHsWH5UzhzNz5dccnlf
IWx/TMKFJAThsc7tB4jxF6G/DRG1VkyhOvrQzM4HJY4rgXrnfMKHMX3lb6OYI4wGy/ZAcmLwsCdN
VnW8/ySZX1iGNb3XQRQXGtnN5WYAtDmTlm+8WtyNRz3RqEfZjB0oUzDIcstK/FuwjokQdQ6vpB96
6dalScK+9mzEvgChB8uaUwtXtKbIj54sjJSxMMCALXK1mQMw24vlfvZXPp5yWQg/b83JZRkYZOkt
mMR1YjemwMGL4Pk4H5yiOyZqMOlwoPLXgWJAJx82oIc9YFGgET6I/ewzKUCUItXLdt0qy4AEl9Ob
A5Oj9hzsLjIb+CWbW8K3RI2KXnjaSxS4rn1iWAwa/H2FuORA76F7yflxpxOuM7zowMcaH1O6/uY3
t44gQ/LN6QpkVUQ2X2qlE8wyu2LoB5HWWr+TPrUXm7KiFEIcRpV56L6ZmyZEmMMmiFovcxXg0Df6
KB2VeQWFhRWdV4fdt4VU+xTdD3eJsEvTLKfo1ah8doh+fzewi8lCH5oDL6RBWydhh/HIh03qp9Dh
v2IASqpAsBNdLnFecMtOlupMFES2i+ag8b+D8C36QMG4gox8lEGrs8KJ4A2q3d2WcS9DdB94EC2z
NlqtMIb8TsgdzCGssm9XkVwJIhgiEjh65LaT3mr8uitABt3tw5MZn1v9hdiLKYLvtQJ8IFiVGQlC
RQTLkPOwSAv5SSi1JgXsUP+O7czVssclHfPlMHOGTzx3r1N9CVP4HtZZw0PjfPE9V4tteihk7bOU
U32fzS/KbCLKQV9vHJIO66919nf7SFj4YkrM3W9G9lpR0TBIwm3T1RhgkPXiT8xyOW+O8quWYqnA
7eRe2LpVGxkLCroG91m1otigQy0bCPqjCgLbqWH+PBwQab5nOS2Dwn+KYyq7cngKdwG8VR2XEcIC
j8uHdcqWxAmhXtlEOjpkntfdK+qFEbWpNFowOCfRhTUP+Ee2PPz67aE/QjVi/FV9lV3Sg75lM0kZ
JMB9BQEURbXARvrDAQfLDVzy0ZIBdqBpOomu8jQ677Hmc5iHkNAXj4R9Wjt1ELXdv2SkyMennF5T
aW99qD9WwDyYcym250W85UmoS/9zsWkTbhWLQl1Jip29gQdKo/r3ZP0A5S+hhMcXu5PlUIznpo7b
mU55uGVJ5OA7l0yFygdkC3HF+pjtdI49n5Fq5WL255DpffpWKK0/BGeYLaMRv25hELbjOR9+WJUu
Go/9jdZzaLUxOk0DParmeI3Hd5v6lQKKVCf+2fwloI5lAp5FlEGfIRplsd8MJ0ZXHY4tIERWvkFE
ctWqHHeLHWtUZ1e80hFtGcVtBNthv0YJ5DLvXRTyRfh9p7rMdS3E0vSrfCienlhfl2/b1KHgtgLE
Zm+LVayXLWdrBXPiljaGlqja/eHgr05CHBQ+rp4RTwodDqBdrHcQiUwrHplaMBjZFRiRIbBITB4q
FFmLNCaBOP+04J1omv7hFV0CnqPgmLClvmbkv65vfXq2zL8W+g93tE+5eLVIFCKx7Z/ixeW1X2Oc
hm5FJMyQvJ6DLDU/NMEyUszd3MTPxmXIEoNN95iY8p4iOfK6YhqLez0Q/w/YOQPvotiU1sLcmccg
Ga5tG6Mb2yc5qTidFOy4YFZyAntT4BBGS5uHbe9cNCQIFQPh78/m5F5NU93Udxrsjwwzw6NZX6Ri
3NttQZQQxndH7pmH0ZA9ju4MZ0Xc/e8vn+5SVv0A4+hQzN8K6bzkVQwlujEqqQuoAIuyAM3lC3SE
2Kz/+jm+5zd1iCefKD2rcTp5f410VMJ6WqXyD/nilzDMYe/QwoBt+4zI3xWGXxyblHEscD0a13QM
mS33cR/DMarYhww9rSktlyeUNzcc0NQIFkM8LH3WjSjOtechYZCPfnNyAVngU8+SSUJE6UOXd2Lq
g0m0vMN9r/z9dlRNErDhIOdeugxrQHS8pFfRwimNiGhMOnTdvD/ABjggDxaGbzlMWFIs0QWqMnxr
oGGb/4KYwvaXakPvaOilrdrphILYqE+PVhKyCelEgRrNPxxETS2tdAzEBahwCQsyKoyXReyR59qv
5d0T2+iJWBoul0t6DWUSmqNCcmKcWca7qkfRj/VUSPURLuL95Hy0eA4oGMa4KY0wGrzWmSABxHdc
3uJJc2rfc4m0iTA6Z35BUxJlYD5O2+Fpu7l5JPC1PevHIJGjEwHgnGSAsykEaCgg9FW3ntRL23fm
uohwNYqPH1d5yF/TRPyUfMnjb5PHa0lmEBrw8TrPgDzfnFqYzZvkqVUoMRj9wiIP9v1TWJ5gSar+
stF3BCQhYnk3igrHA5wLOe7iAq/tHycxagaxYCYufVhPj/uWdMq2stDy1lxifPN/j8UAMJN2RWWX
6pIWIFc2L8nomvV4v7+6HEadxKlUxDu+MpitQI928WYfE6jxN1K9yNwRJcYAu8USAmSZE1Qg2NPi
RL6qSkKxEvu4a6bQlTVyo8zG9dFqPqTAidqBwjMQ0iRT7I1ktqqvevlwWanK5WCU1G8RwUEPCMNG
eaZz4mG6QLeWlu8k8EPVPhztCqDFzIIn6/JleNl75MG1+hRt9Sz0ZO86EGdGhQ6BWek1Eji9L7jb
MwKWKZhswPGvYP8adbesv883z07p+hKoraGxX9mcGVqluN1d0XqUSQv628nwSLlrQU5ZSpuzkKoa
ZzQQ4ltLSaLSSNKgGEkvIh6paWT1yS1cldN9Li3zVVLro56rBNiAbHTUNmDXe6OOiw2IPhN3xDlI
FKAhbq/clDHjc1W1t2cW2cz0kgkLBUJNYWkuOthFS/TIq3IEvk9NNi8Pxsnl087TdsG662ayrQct
iA7AfYbm7KNst2l7Tg8B1xniifzToqAMcYdRtWZwnTsuvxWhQgMyRzQT2fUamJYQ9Ojr+fXqAsqP
mj//HlgA3Uze/HL1TRAIXtDTENxdaDmrnm61b8IZ0ecgBYuiD7rXfPMJNaGrqMWYwcjiFpD+wGvW
SUI+Ba0LBaXVxYDheqLS7dToXIzLQUDp06YCTUhREDRt7JJhQvrMmOJ35nzbHw8j8hjSM9z1r1j9
FXTUrnoeXbbGXRBTUh+4QYKD1MXe5eVAZWMf0Ej0KN2CqySHQVz8g0szwXIcHIDhM0RlwByrXG9X
A2QehucPYR/vFtt8i0J6QKCO4/jnWYbMvMpEcM/Y9Vjfk5P0XQ/DLjIFXFCvr1AM+cJPcf4td9lh
/JfonDRNX/4zEXd8nnQkin+DOxCdvMCxyEwjZOrq7al7nLYuKwAxbdNl4YzIQsl1cc3+igIPK7qd
WqBhQoBHHXH1ZUFShVe3uCRlHfcruf3lXSh4OoGJp5Ir50th0lS4Frk4IZoIu++nnh05Qli1NNiC
xT2FNJkqj77jrgkdS4VlQM9VcO/AHKoxr9WLm+niS9lhFAwPubzHQaJrACvlPJO3227HgLKwcBPA
1XiCVM7ZNtkZhm8Prs9ihNEpDvkrTdlm9ETcEdqYH3puEliklvv61l+zC+l2Wz9+RmfcwMjUe6ra
d0KT8A8W2Mr0NB8MGB048muueHeRG3TyZiiLKckc0lCOidtuleXm6i5+mY0IfcjbEIdKmyzOLhlL
IScV2U4FQ9VcIAWhlnJvDdXuubbRld9ey0ZwhTUTYvwDUj789dCJVsDZ6q9u/7NymLQuu8a7rqzG
qOsaoP1+UU2Wa7k2swWrIygZc//eGimvEF4kFmNEwh4Vhql7qOBc6Uvue1dNm1izfIHNtyekfbX9
j12S+mwOVN9N1CG8Be6rkeIR9natDiC8ey1MLANWZl7zWRi0rbPLhY6D5BcJHmNZ3hYGPVg+SyzL
FqpSS5u2njx5INVCYZX8cUJHD8zrZEtDZ6VbansjC18aj1TYUczKhg7aKnlfHUdZGVAenvWbFRb8
ynUSA0RaMG0LUYNfvLM/Xp2BzVCwxRf8ywJ6/xEDbmoLJT//mdo5bdUr5V1s1a2/3foFneQPM8Cy
B5bqExdU4EgdlkeqXXVf6NXksAJ68o/O9cUOYmZBUh4QDorxOnfuELe7KMeGxaKDDGaDLx4yu3iL
B5Te83QGOeGSXp8XWLYMdhueoT6WpCinxB0oMitb+fQh3OZ5KjBQBbNOMVvLtJBUXlAm3Ie/rsRg
WK8ykUSstEBpWeNbT+YMsRdh5KoNeC0IGZWibLhsEcUH3+evRiqL4wTA+LlSPVxuXgYIp1u72lhR
K/yfRYFrk+yuU4S8LSGKL9232DLfwiKdMIJix+C1tHq09p7TPh973nwt0vvmu7Ws5y6101Se1RyA
0MOc25hi+WPQDXK+0hhQqjSsIVM+zqvXgqnFPzDH12kPInWKGIx3kO5zWK2hXiZjgHUCAsHZ/jU9
5YlbDc2n1X+FsgMoNx+EBgOpEwuuQh6FBP2lh/VdI36pmsih9bu9rlsl/dBzqaxhUaoQ4ErQPdP4
EOUL4nCSZiRZQylqXnBJYE/Jlr6N2CNCBWycNYqYu4xyJtT5i+lryVpUw1hFpGTSWUOLQBoHqQyn
ffQq4FMmd/pQc0FGJl7aqRCHA2dFKGWGG1cLRFDMwYYfVphmuNUrwkmIJgkvGvOU9t4dtdEX4PvT
KhqUufKUMx4j/NEbxgii7jHiF8n5HhuFd/VC/pVPD5w/jRd6UxVIoC0fZB16rQFvE2azG5g1cwjQ
6LtcC+S/WpBPk4hV+kCi/1bmn21/8iyDqOuG0pWwXD0eJEbohfJguMOtgdelPH6b/0b/5cc3RUAF
XAjmEsuqXLBhS06bFsBBrGyjpXjpO/FvfcXOn+RV8wqRWNpNfE7KrtQ6EO+e2b8u7sKzwQz75g+D
6KEHFucP6IxFZjWOQ+zqAn2Iy10jKyTQ01ccqfCASJc8eptNkse1ATCFkSMnIFwkZizJkdQT8xKM
umaoCM/DhsS90clQs9zOmccz8eEqRiZxr/kWR2VSEobUzJHh8KT48aLp6CGxMNKhPtYXpGTSM/+p
A72DIGTWG+uegM6HJ7VMC4YDi8uS2LGage0oeCobS02RxmYUZ+BunGV71akZanfUd9ZgWa+vwzuw
rhp6vJZ1h5lYKgAWPwDWfr6zHaWbKg7uoGbqTt2zvfgoIRspFVESfXc0l3IeTQpMI+/RccJSbOlZ
bY8uLuUB6+TMS9h8jEnOWMGGXAkpP9t6gGZgjKlwIVs7BWC2jyLSElRW0BeAZmRejJJCogrSm0nD
/zUPv2MXfsZeU+96+6EbU5dgB4MS2ssxXxg+2GOnCqia9WUckQR8Rs6x3dXqUV6x+yRhI4wkQ6po
JbbjO+DuwMKqRsiXNmDU/KBfjK1vfHVzTVT2D5HPKZldE+zkQ5/0j7sxl26VmD5ddX8ZoO9IMir1
eosW6gI+VHFvX+ddv35XR5BUl9Dw2aTvTW3FHv7+fUT3ZPsIaeyNlBlF5yiImjoV1y3bMQBS8Eg7
dsdwOM6tlE0IHQ1BHRQ8QM69DqLRy3uhey7Rjp/FHhQbwBpprYZ/lu/EwGbdF/yhTQHDAl7Ncid8
nhYxpY3w4c8OP8KfybIlK1bTjAbGQGt9qV156BdyUHOboXIOhiHrzCPBsZ5lU7xKMp3JSp8HiGEN
30DDOKa97xn9uj+zChWNezIGf7TCBz2LdWKs1AIkWI9nfkuOYVFqY6fkTcW0gxXfKY1KSQsoslFT
3lXKNCiMIePEwoZoY7kUHOI0mq6LV4X3kAwuMjHDC1JRKxxyK8m7omp+YE9w6TVIGpASvqBQkIKk
sypKJltP4a0jak4ksGyjnZv0ALteWnblt23MyQIqkWhsLVaN1vmfYSNJjJ3XLFFM+bnSgEDwjI9/
X06ZwmL56Odm80sD0E7b9LmpfhYIH3w0pAAiOPqCvLwFonC7AnJntWSCHTPm0QzVDs29abeIIz2O
wmA0El0PiUP2xFqZqMlRpZRb0P9aIJLm41QiKZpEOhm6dgj0JbAAbIvw1IgtUn+FgjbADZWi4YKu
UBxoPGf5PR8ql3qwuf6FUX14WwTPQLT7YWfKQ/Kri+rvPHuyGsYX7HNESsNcSxlA+dRRIyBpy/XG
7IGfWSfj8F02LYaJoA5FuMbrXri8YMugvR5vu1jLk8Jd4zu8l7WLnEtX0mQoQDbV2vGTBdsvSrno
qhHUrQCgjrhYx2+YRzeGpZOUdjdi0B+kIUd/yvyuO34PaoWXvsvp+lMhF8i0VTAb5c4RUCDFyqTJ
bijwB4o8fdMY9Mnrlba+S3xl2RTaveZvwMCgP5VrePC2bfjbbcOISQQYGVUtictOJpEwhNlnxBx3
WXDlyl5WVpYrV9bs3tMphUPK5KareaDS4fh3Li//yUH0sLqggDEruiIUrNvO/uJ1c+/3O1nUGP37
wY7DJersGnDQVgY/ClSy9vwK+P4z5VY/b/D2lOjt5j2qUCWMz5BmMMVAWmu3aKzY80FPFBPmUZhx
QDQuCYkv/22oam1Q2fwY75kG9pstZ/prhK0a0P1ZyXjokKkPqzerFXytt+xEY1QiL/kr2frmK/Oc
8n6k+sYt2A8iKJnvk/e+khMjifhK1X98N/p4vFz8jp5Ad8fpXnHX3kIXxZU0uqfkw91QKXPG4bQC
zskfW6rxtZ8EZ/d68PmNxOoiYLtt7hF4Ju1BZ1iUy0G3pzcaW3rDFNY/GfXuPA//i0dtrpSng34M
3Ej5yrn3gxJCrl/ARimN+wzXIaVccb3QC44YVvz6a3uFOKVfYaKS7rTv8fmygxHT+WvE0QF7cTSo
3cUV2ey9pfk0fWsX6yQPFry3Vq4VSVmgYWU1cWojnghoD46qrKOkcbJ+ayh1QP/27brZBNt8lBe2
XCJTQcGRNqSmqKoFL44bv4qqp6dp5EOXTvZM8sgEywG129NbMNvDBf4aFeMPAjZozpTeDbEnd98Y
6CpBdaCuwxH5LYSIphS/9LsJeAx6mi8tqhC3XAoqECyqC5SRzKJe3lay2ti6QYgUwU+WyhMEWvCG
v54BQ9WtHjYMhBfmS7hw5Jtkt5ahWlQW9pwIyF11uxYtmC/hsoqYbqD9RvVolnneL8DMrx27ON3+
mOve1E3cDhhL2q4UAWjDEjWHEwmcmCMisP2+nVZKN+HYCQytAAgngbJkM9HJr5uM2DmG0B8S0wGL
inmo+NT9lwpFc+yEgHWT4PVrbwPna+ZuA8QPZnX4YI4y6CC/igyEszaOcw0iYEwqtFgAatXNhfH0
CKLGrFF6IYaXan6NgNoFkIrdb7yfRM0tsZOiZaBneCjo3EwrucfKopK2Z577uFmENU0CSU8G96Tv
A6QEJDOtjPZ8C3MSBKPumllPOPma/waHRLNE6dCQzhm65lsqn06z/pOanmeZb+4EIkyAE9ArtW5n
j10JoUxLc/2TElKUDeiaAiFGnQgGU0TMtaVXZH8PGfKee1BvMFnEVLe2qS2FKa8uHR69v9riDKrm
+0NTZQtZH4euCjN4bdgx19dGT6ftWnkN6Cn6tUUTH+b22Jo4LyxHASSu7wFsE09YTqACHOEZKk0R
jI8CpxaQzBhWOcS+q2cqsuSGQsJYSupAtv2+sdhemWnQSFq3oThms0/ajRuxPQ6IXJfamQSQGgcZ
vcFfPZ6YyBu/ZSU8tQZHg7T8p+UWEnyTW+eH8sddheY/HTAI40nmlfIWz7kxWZJ9OwHZd1ccwkez
RWQffK8ZkY3w4+4S2nqQf1nO6R15AvRej8dB/13RpLPkqDJwqMGJyJQwIMokGVz2sycDVjyjS8NV
porpF2NZFbqUyBNonpZOg25MaY9Mq4y01HU3jS5IbCGcwcJ6bmy3qyt4B0P723FrIvlyeELgHUBF
yHGDL6bCDLtG/Nspt0ftEg0Tr8Xx5YHsK6ac7O3YmLtps+jiwr8hnuZ1FOIyp651zkbHFVp1eV9L
xFCHQSbpi2vRCb6gtx+n9dP25hB0yFeFKBxEQ5S8ZXJ/jNEnME6/AhIcMFYpYicvVlb5zTYceJrM
zEatWk4ySXQUCX6AovoRPbGsSNh3iUliVFtadOHqBHM0XdyOPGrsfdLYefbZEF1B5nWmRz+ga6dd
8MybghNm5KdEdvQrrWvjZHXpSYG3R+emYwQYXY0zo2ei0YX/In4Z53Zc3RbaHLLAaIlnEDhK5Cow
5M/vTXLHePY18Lq65dqtxgK7khGZGLQtJZF5I/gluNQcrfNr2xWZoF2zxBWVSHoUlP4tya2Cku0U
5hFLyLmxeHpE1VrzbhsyaqEh87SC+C7kTvRkkWCJy3P80yBtIor1Klzus/JBL2a5GUnIT60T+e4e
aDkHfMUL0POTqlPfAbNd0Us6dkKeoPsAspn+4YNd7EPbpnbgTanoYrtzXNcY7u3Lbjjxq4MO7S13
OQKuIT14k7LnWCtll85Vm4zXoJzxlrKV2uGBwdDRSQaqaT29zhn1gotm2Tef3bk9VNTkUfvfDJnZ
GPnT59ymkTxq99LPuVB60Pmdw18vQLnMDj5z6ea1B7GzJk5J8ih96/f1azW4hfBVcbxqYzPfuQ+J
yhuFG6EMie8X0ilOcamwjg7IR1CT8lPkLV5qJot/uSUMfPZ9GXdscMjQ9k+jqf/uZkMyh07Wq3rM
+4V+IlTF9QSot+Kh/AZnAa5dFOmdjFj2tFyXnpzpk7UE4KjsueHACcD0u5q9e5ftI0flwUhJWA9f
kGfw/Tv3W5Mf6aBd4G4d6W44v5MxUsxFFIJXEIEY3+iE2pt3256LjSzSkj6PVE+TH7sXKiJLLsLt
5AGhYkLo7SmXZSYs6OJcSEWTHK0YM9k23zaaiHl3+3dQ8ykoJ75hcPWDhGq6hroJ0g97ZogqTXKf
3eLDyFUwfrO6Mp9blc1Dp9LdqvuRYU/TM53BpSTkFB8aLvTHKZqW8vp+jKDogd/zpI2HvMtjUHp1
kuI9eCnXuobNf7ip+d96tk2f0802oP0svNCH1SBlnao9gwLJdmZN1EktZrK8BXjzkJSzUZBpd0or
DhG18+lx2dlG8KXSje7IoHjDMids6CIm4J2xqC0WBeU2j48sWGgT72aV2fp2VlUwz7P7XFXKMlwc
facrjpGJfvhNoBzhtpAnXcAGjN1OfgLLRbyqcQ+8e7bLdINvboIXQd1bQ7TNgFT5IgjHCvTcx/HL
ocJACSnnMDeIyWKyPGIz0a+kmbHRGGAL6Tmo0X/OYNjlosSezI8E9JarrH0Z9DgNUaWlG8gfA7AM
Zq3zGuqvRSGlT+YxE5R7u+aqpStGmfO55XwczNue+w8Y/2U0p+PvVCbd3VCFVNljpO3nnskOIRMR
+0RV7AwnzXXMqfBiXwmXUiZqHcoN7eAwRRgJkRjbSe4IKPvGscS8R2eVRadOaV4CXk6CM8SPuZhu
8034vMhtLuyCD4Kk5jhjKTv3XwVaMBXc/bFyQxyNjg4mHYH54VA6M7ySh2kDb0FoRPQpnyVjiElr
sL4r9irGpePSsZXsJtOy7kgUQ0A18B4C4loTAZTfFI0JKA9Yt8c+RiPQHb3GMfTrx9WW3k+daMZN
DbHkrCbDMkBA0eOWTiVu7TrkloNPMExq5jja2JqMu/kX76Bkpv5cmxmgU3Tr8DYFVFR88jG7sa4H
oQCVPPY/iZBfcHJwX3MlC2lvIKse9rJ04egbXtcJza/A7hkXghk7B11daBcafGpq6tDHOuyDWYJ9
yWqV3FmbS+2a8E1hFm3VFagSFLhge9XtZtQMRpF4O6TdvCMUaZ5kRR0HipKHxfLwQO726iu2r14P
GLHlJB0pgJMS91OdyLI9xdrIdFrWEl5JDKGW/yVyPEet2vY1wtqjgq09gmJEeKSkJkNmmMOAfMeS
bR+B/vnzD2XxdprACe9NxH7u92GadVmg8JYAkuJS2Tar5QmpRUmR1UuZD8ip9WVmQiU6X4SDycqI
LdD0isiN4SU53mUA3aqXN04Kc1rpKxmQdtl5wiPIC45i7/kdrI3elofsI7IPF/1k8DYbiA0kvPkT
ugFXUFpoHMvfReTao7wJuKZRrMTbMDCbU78dqZTkrVVEU+uyLAsBjvi9xxcjtqlXVY7YfXh+ApYw
xiQHS0Jiyw45ayd0w4GXz/tPj9oahCQG809y9d9XiWM65I7amylTNTO4aHBg5Ore4rn7DSLIWPkY
I5z7slSmQR3mtMyZDidelEr+L+L5UhFkiGfG/ZA2bdC76w8qLyr4mAkmrJGMG0tap0h8UK5Y11e3
91GjZk+KN/OZENTspT+/fVR+EM+5SO14GHyCzXbkB9m6hV++Z01YlvjAsyYSHulhaunvsiG0b3zQ
p4eBoBK+wWzQ+86vAlGvIbKYPJHNiEt1LOTuoUb1MvhgtjsxPd7DZ8n5ClLxYaKf1Z+dcwHDREaK
itaJGuA9TJzLOttBTrY2mS/HNXl8FZ81IvOqCOD5C2cPynUnajonjX8+L1mPQAIhnfqbUjmaStnY
MLhkWRZr/OOQjkgkzPaihRi3Fn+uXcalsKsbBJTfOkEf52CQTijPlIjfglR6AikgeG8QL9wL0sn7
zMqtpCAa+g+y70R8SZ7dzquH9bxGXQXrw6IjS0GXhEX3Jbl+m4GBosn8Qpv+GGE7JhnBRgVayW8n
kI+xsCXzMelSolaLBRvQ5+5wT7qc0mQ5Cmqw22PQFe/7zP08bfHhThyS87BeCE8n3JQ22mcwQwyS
mka4XGsNYip0+wgO+vzSr9ZuqWswGB5oacxtOpWn+BTQx95yvziKzG2vuN0xum+NGQ57JO5SF5Al
x0J5cB0ltQLAgzT9pfQfQGBbLMQEyE7FLcIr+wOFWI5Ja33zf2RZCmXHT4G0QKh4x79SUwIWGmtz
RX83c1ksZD9/gtWJo4JIsspIFhfdDUnv8hWPqqALJMlOGkX/M4nz9mqWhcRTZ2xWjRjDjnK3ZT9E
AIv0NQPuV8xA2xDapvAKzwW17B/w9VW+jrbfbfbu+f5jv55NPVNz1S+4Cdq6EbIDW/xo9FTxskKO
iRC59zXAkrni+F0EHcLyQpMpn65CnJ7Ct4bfB214Df+30pB2Wbivqo3D6nfYvYyAy4FPjZYFiUfw
A+9gVtB3ziugjkmzhgQaQxljuQq+fN/rGCHSVs34Huf0pm9x59GCkFN8OjNQhquYvwRXCz6A/ijR
l2BhAjdWbAeiUv25uL7YdNJV1OhZLUievngi2q3aHVWT7nEI/nkgTdSxQnRyFj9Q1OazboaJpp+G
7PX9B3TReHEgpqn4uiDJz4GaEmXqh92cOJIy8ieLnu5bbBjCcSHacCa3DJnbDxjYP53q3bjkDsRe
Kj5kfOfwuBiRf3jB6jxWXcxw/FmJDhqA6SC7TTZuYlzOLv3Pduz6S+P7DdNM5W7FFOL2kT0540jg
v91IeUYwuehitH0TL8aI6Uo1V63mCuv/hUGlry1+K8kkV/zqhwHZFLjoqobgJTfyio9vSwSkaLPu
WsmN9UdhdKpTerfGJt76QcWf15j0YM+1VGfA356iLJo92pmUGjQybKrLNUaDUCu+V6oJKMwfMnre
kv1Dwx/KR2YA8b7HGHz9XkTQ03RItQ/qE3JgW4n9v8DyI/Q1r3xRfq5DAvuQfL8VnyKbqec/lBi3
D1J31dLdpG3tX6/y8TMD05i2KjpwwZiiVfidhCxeXtwCBuPWp9yRVSpZa36Igh6PHgbju+JX2u9D
cqNvuDhoLcOgpeTCSYltLlkxGRJW2Z3p6gjonCVznbCefW6iqGDkUt3+BUH5vODVNxdrO254g3ov
w4OuhJnU7+28IwiCXr4Z3xLrm/5Lb8LlUkIc8lei5C1sIKD8qA/KT3clk5HwLXWi57wGaT6+Nfb0
9IEKuCffr3Hl+PcTk337Tz9FLh/HtfP+csZ8A1xLSUmEDnCO5NoMaOd00zzAGPLn3Frdr9dSOR4f
aLl/jIOor93p0xlGzT0mwdb6lrDjcJATtqUMTbssXKPsdvACs4wRCB48ZXlK7t8cvSdtrfJit+lh
vaydg6dor+dflSrATvwhBvzZ12rydJ2wu1aOZ+OcALyD40H/PqSybuwhAdCSuxrtvpRlSHdE11Ms
xGMhyMqO48m07iqLeBT/lsDbnp8slSnH/HdB578M0k7poSh7S/iTmXFnyN9J/VhbN6vB6axB86sW
AaS1sL383DXUlGjIdbRB50A008k9gAKeoM1zHC+tcTBt+JXUEYNWjJrHkcEMJaGyJ35r/RKntBCO
uKAaMEuw9OWG0UFrgZThpWzdG6O30B0uSRNlyFzcMCeu73VzWYqo1wh0KoYM7v7wnP8CFtIPiGsC
rskj6po/T+kLF+eDObypXnrcpzVv/SL61aIG3+Go2FVa2lDAcvyxuUFSLZH8ifX6gxvTk4JFGMJA
yNRusevVPS1kw/kzkPoaO8lX1GqWkBe4xyaswy5OTBjWXec+ZnAuin6Q0EiVF0iYavMl5Qqysle+
WuQOFqYP0mZYFKvwb1GmJ9r4DdpuLsmdJqKCSIOHIyD8RjSHqgLNe2r0TiiMVMigX6fqs5Kkm4wR
bCWkSZXXKjN7QwAbkpSlBvGMc7J5iPG3PxbH9MQunGiBY4Lo7pDISHusQY4mUopq4uNM3YT8DQdM
yfVwoHjSiB7gvghE9KsFsRLhF5RZI7tyu32NdWEZf2BuzVfa5kXC1B5OmUMNj7SPNoO1BZcLGEfz
oQoxvZ9C53LD2pI9OcQ9AWJeqt/3HqA6ptm0mzNvGHBZEwQMtz/V0HujDBGFj9Yok1yy/6yhLcq+
psPnqk6TIOcSyLOZwhAGufdybs9x0O1eoSeKtgc/ISh9Z8lKnUTO6DgQhebisT1F++eRnQLTw8af
dXB29Ge1XdquCGsM6tMNotu3w3atXL1+PXxxISV6e3JIenPEHlrT9+MSnydo7t1hHdq8s7C+btwG
B1NF7HaGp80E/Dz5x9YVZpkLzMXk+NH4eJhQJBpeT5dl7QONHvTkkOxQzO8HdLE3i3YMu5wWgd6+
05ZKYoBlHZ6xEoIECopJUve68+mfdtba2yETNnYgCcWPIhR2hPjxBI5oRtA9/Ip180JCR8xJkbxZ
iErxmrcLdAiiR6PIX0uQE+YO4akY+LpZcQGHBitsnDNYRSfBXU1JpyskQ+MbMO3GFvbwi8dZD3Dv
ab5iQaHGMLxR3SAPdtkuUdGdMcIayStwbMP0y8/VYst9qB0P3RhBGVacuvVhYtl63ECdd93N716/
keXIMwjxPl0w6Hw0wtJPFVXepjBbtJEjof3D/nRVak1PD3rOwbzBPP/ck7FVJqHZs8YSJrkUPMrw
0YY2mYn/SpVedjhcz+YzGiBfPf8k38slxRRl70TDXjPQKfFRGBlksvjhw7ldX3bEtStV+8SDfy1F
Krrkt9qogJvKWvtkdYuJlM4K0x5MtFQ64F33hQ+U5Z1UXMjtHhsjz2SZy4YNlZYmRYmRB9EK93Cu
l7lajTtkb87AsOZ9eZWp/GcUBIxRVNvmHN4xEv7QvM6NoOcPodbjzrjn0TTscAq5wGUbs+egGaN8
f//EtuJZfVqkELqy5/91oooCHPpynvd3IJ+tuRL2HiHIqsWcctYKs6VW6QMNwjqUOHA0JmZslKIE
yaHQx02SZpJzrzC7PI7e2XfJ2aUm9mjy2bh50LuVo7y7gsCcErMqstvAtLr9x53OiVWDOP2LU3OP
8cJGCzPWAigldqwP8NnQ6mKsRIVnfT7qt7hdedMDRlTeAbU8ZQC1P0yBm6nkB66sqSyJu1meXc/s
JApQze6Hl6PwPZFAI9dGxjO7a6aZogtv7UIL9FDrtxKOLNwVcyVuGWK7mzBvGskp0jahpgXTjSqX
eaSyYtUpjv//XEsy4+d9aJ9cyZFFMcw3IQdYNS90NXFj8lpCbRDZ8Lm1Qual1lzSe+vlsWGQaDDo
0e5PVNIXZgG36qcRz9zeS5sTNqVv1ku2+7sKwn9NfNjKZq6UG5jXi6HXT1kEJb6Z+pp9BhbqM5jq
IdXipWcp+EvOXowsSAB+qSJeRbFxQIJFiJpnFc7dR0VejflaY9rBLlM9irrPFv4bkHGjCWk9Dp+r
Cc/LQMcCFiaykhw74wOVwL6rwjXNTtacWp+ETQH1abN3M107o7ax3USMMIv8pTWr8m7CUIBmWDV9
COjnXQFt/Qq2CD8z6Ymj1CG0bkmkk/zpHTOt8uUhOha4JtK7Jen8FgQqVa5kuTx67qcj2di/V4sY
ih8g/INqoTs8OrwVUpUCt8JQS8wakue53FXYz0r4RusIDfI6H/OIIiY629/fjwzpXpgIWerRJ9te
AvFKHHwuMa79Ec6amGj1SJC+4C8EJxjQQHhGj1Rdgy6bzA04twuWeGyNzToz9RORyJaGNK2AfWYK
oM/jlPS33s0BkpFspK7/j1JZxqh/RDIrVx7f0uRtxmc3qTxuVbYL6WFMuZNN3xOKiw6l0CxvuvAd
diuhvY2iDkP5cC8i96tdt244F7mvrQxljuNUIs2XlOdEjNmMt9nqoNVCgx7fcAZW8CrcMVsXJ0lO
kTISwcMnqtaWQpy7sX4F3UjKQTQJ1wZakJaIS28YIk5RCcPO+zEz8w9dk6DTjhwcFaOy5xKsbFwi
6lEs/f0i4cNy8CBCtP8Qx9RGcCYqmH+hX9LW4cOS6qlaBxAvdOMxKlIeXKBZNKdwsbLEVKxSKRKt
bc044PoC3mkI2agvk9AFQtMrLh7bT39LeJlJC74eC6DOJi0vsf/PaQb6NoVK1RU8fHG5p+/moZHU
mG40bQA0HU3zvu5M2w0kOYWR1ZNtyXB+NLmA4JVP/6XBtqlSJHf/z9CsHbFhUlH51xQXhxNLkU93
X8yXq8rxev/0jINWGwkTFSEVYUQrT+rWZMqyhh+gDg4GEXBLP+lS+wdOpxl/N7rtab5jdkpEgZPY
VaZ8ZhaCVv7sHUAjV/qMoMPHMBVyBt6JUCmLAIcq+3hJLerdEWtOyETwZwqa3rsoUjehLUzurLud
Wbo59SZj1fRthFDbLdNhQP84lJBPtqQA6swvZG8R9n5YA2r28ZnHFxG7YrWsuPXRdzfCNfnNpYzf
DRgVEQlfDY/pSv5AFPnhhEZJjkk5Sp7ggcz4GFISx9TxcSqzmMu60n59js1MIdf+qg0DJkHgNwdp
CZKaJ8TaqCNKKwS0QLabEqSRtrMEBJEk6mtL4Z0kt7MKIxcziWFxKAWdK4FNw66xeAFDvZEPczJE
W13gsQ7y7fLSqnSm5Y7Y2jOUd76ALOs+nPor0/2yrTutDn2sm+MXjYVGXNwUdeUa5uq+V7xSRiW9
ToFPxG/mEelyKS8X8Yd+mv7B66YQcgvHqi7HtyahVG4Rdm6uMLwjzdEmckiQFRWRel94waj91Tls
tkVN+P6/aTLbGYYKK1jZ2jW6TvfLC96xmk60/Lk1QsdMtHKGNtlPMRUa01dJ8jJ7zw+O8QyA9c3f
7eE+J8CeSTL3HcAg16yUDcgG8gPs9fgSgl1GfSqWOY8VvOZ6l6Tk/SMG3Yp53EmMbZrBAibRHzuf
Hn/zkaUA7R4tarWscExevV1CW1XT3J4PN4UeDahNDhn4w3w/ljh6E0AcoHV17xkFOCNVhwSJ115e
G4sQ2XqqkCqjRN6rmKFwPdq1qk0BTNMhgNpebj4gW1wrAjzdUA4/PQrb7pioXf/f6xEw7KVZKACs
zb9IpHMBzrdleWKF6MaE/qcstCZsDrAXRkdt/thjgTwfiBkz0jMYETbbb9f3snqLVxGC7T9TuLbX
8owRkZ4DQLTJ8ujShrUY8DhH8I/WrwHkmThX4LjP1yoD4PrjIYdprQ1e6vVRCuP+51AKm+wPt2vF
kbMWWAygd9+stFdczr06rVVjAtw+lq5CdPEaNiQNX/PMsCTKCV5XBklPglFweR/YgPOtVstWx4CW
Lsl7JIRVemrbxdupFYEfHfyTzoMAEyM9JLnxvJCcCIjmbdPkYJbVNR7W3gGDolobKY+p6xrTvT4o
RWJeKsY5kSOB77jSC9ZqDVcVPAvuInVc4YB5aIAjn0huA9zB+dmRmgdfJYNg0IG2k2HyFp83sns1
LSABiFcJVTf3wDZO02TL7xVAc7kkfX0ZLymhzc8KQXgekERuTwNY5BPn8EUZn9OBhogVZ85ecVE+
ihWJnrDD/3HO1ivV8hck+aqunRPoAgyHK7qPqVxrpR5EIHphmBHexgfNpXy8Wg8PJRv3YoBOtgRh
PePQAvpixVtkHPNyQLWOKCyHC9q/44S+FJpFKZVMe/wjnxQr+A9lzDgZ+Yzz70p9naTMIcfKkHJf
AgylEln4huZoI3qggNex2Z79DpAnOWvEFdHsCxPYCejjZrrHFflmIcQ1qFecrE+moHPieGRFX2dS
n9OfB9AeMKl4kaaOgX9cpFrYLI13jUuecZPZoDdesNXvm+QBZnowXi1v1TwtalWTfwEQnvgKxHQm
XQXzh4WxME6IYv0n9Vt8tSiyie86sU9KUh9MWs1i/XOrXyFjCEQiPN5BE5hHFCvldPRlPGbutASZ
LarKNhFQdtJdFV4VUqyyMp9s+nc2sZJFX/JShpQyDpyN5cCsuvcQJGy4fLHumhwzCLYCDqS5U2Pe
04TL4Es8I3U8VwL6nSGJBnHTnZupEDj0Jea/jwIx2l902FKB+QSwDjWXaj6R26CDRMzOR62ooYZd
Z/ZQ8YXM+cFUjq4T3nFfCLlIpssgJkz2K7apD+GSX6GbRaH6dywLU68LTdOKpLiOmdfZjLtdpyJa
avtGiAxazFbiecsXc4xdk1Uaq/+AVryApdtXguNxV1u1+EZ9k0OKSbedRxKZ6qhLwNujZCSOljLz
+U/9bdzy+nZqCboIC0vo37Y+ayWUFElSfuzktp6wZH9di4IqkZU5+Uw0W5xnMuOYuW5m6pUbxFmb
W0/E9HGvkwCjg7JtigmICajWBoxXlM3wi5v2kg1ZTdSKYTBqf9OCTttERktBzNFDskqcWLgfxMO/
zb9ET2w7J5lFUOFSQolvb/QP8gYZA4RrcwhQVxYym29+DV1YiBsiBxtTxidTnSTPK2b/rLJRY7LQ
kfFHBBVBGOwCvGusSOSRlW5LUFgW9Oat1IcvjkMk66j4VaEygJh0vi11e1d1aUsaJWQxNwSlwyWd
T/sZumn/dJXvc85XUJ7zrqMcMEi7ZL2AFzkaUF6l5DFb7GUjhyIbY9pGjYVPYQs1v2CF1EzBBqkf
d+NUvlJpZe8gNvoVyQkOSYFWr6yWSYX2SG0D5N42vpfSv/mRls3JFAfZxDyF8iyhaXPN/9ylTUmP
Bv/LU47D0SEh1QTXHcyLMjfrzrh/mfw/fgS5lWhv7TeP99MWfSxP3LkQ993+oSLaSsGvhrrfLxei
m44QKbXaLjoe5HoYbc5HB52VP0ksSAeVWxZ2zH851phRH0VFNjtY5J+OdweciaoBygDs3m9Ckq9u
BLocbn7FK9JD/dJfilWP8Nbd4vk77eXMsrxY/3RJArFnJ6RFxld1rpdGM1USMaXDMR8z8gGON3T4
jQ1KhDPmWzb3wsAEhbub2TCw1qayflpPGQxODr5YGloARVlk33U+OZoZtI/hCuuYOOdFmaBERITS
lOc2r8AcpXwUEkcLsWm5QxDn1SJCFUCHHAOEp7nRVM4MW3uSVjZt+meJkO9tJ27nOzRbmduUMX3h
w2yfqfqQd1yDK754t/O9yol2NLOfhB7Si3FyuSHFku4P+uHK8XZdV8A4QltcDr5fCRaI+4+qY48x
Rcp+LGgOawKoZmLi0bRKF2pN/iu5TQ4yh7T6ZrWW1ZlwweSHNNDO+asoKrD5XgH+X7HpaY0ywIW1
DKGYWjZbm3Mod2A62DFdMd48lLEoEBj8QDvKDyF/+90AfId9+Dq44B90orkfQod6U3RePO8e+qqQ
7Zean8GqJ18Spqa0SjoVbDWlZ67epopDnukG7t9aAVZh5UWyX+eqPp52WuS4Kdfqgy3m7p0H734u
iS00MaImUAhwC+OiQyfyeyvQx41V8+W75rTf7Jx6G9/eFvlKSrrX7an8srMfhxxF42QYgPvx51Vv
OnpnLl+QWZmhbuhYh6wuzI/kygS61ze81H6tBfrsTFxx2MX4Q7ELFF82weWHMVUms2xFfJQ8fYKZ
vwxKJ6bWgXjzTrHnvYttb0jrl/nGST1xrtitRAhPlybu6jWRnxhEjuIT8KcQRwNbslVB6OwpPOsa
ZzipPHKjwHcaE3B9esbAAl5rKiwGGJPof6TeSMjbLiJMlLzh0iIFc4WN2QUsIu9xpG6hTV3c7tKf
JNq7DTi72rrspLsBm6wcxETnHMCvsJAZJOT5c459wC0MMJRCrNWVPc2+FPTAE1zvPZ9z94UWLKLt
KdH4C8OnDDm2M0e2lk2RQTTJJbjXgDhHeVl5kremS0FDhAty4ftSvBdpA9C7HWzrTxh7Es4/HSaL
HwJ5mJ0fCMHUiH6xogd9o2ufCJFo9kCa4flBwYNwwNVd+kePdNebQqwHOebne5tzYJDpblr4dVEu
/g7R/lscGwGSJfzshwTDxe6rCGwZUX/fIkkptA1JDeK0wyj8fcGOdnVNu3EHl6HPCOfTO0uctioL
3utcBLuxCKmK/hnXt2pczUAaGIei3FV2vV3VmOtFXviZhscwSSfReiEbYXyj6tZh0+HuxsCELW17
kQZRIGcP0Tqj3/1bCkKgmzubQRX2prNdtqcsJj9um+ZBUDHZAcTM5yAgl3Fc1ZMtVgOSnjfQFWjQ
x47B/qn54EfPfAdYl3YS7ukGxLbVW1P3gMG1MGrI0bpkugFDcBiAZYwmmyJlrhVJxslIQKe82Bbl
UxF12eT94YVbkhRKywfiVmVpmGycaLVAxqUflgJjFhWAV3s/yYdVlAx3bK9NCzvZzPKejq110PyY
6h9Uea0EMYCSYPWauZh3UALK/1TDDNWVJeSdfyWAnV0lXmNjO8FJUIIAFohdfM5yW6LUv2Y74C+A
/gBlu+uLL8buAhviIknqKuodefpqerfozsfY7Vm/DdW4BRJD+XYBJCongzEiscp9HLF1pVc9hmdF
KGt+PLoyipEH3R6EPM50Rep0eq2zsCYR52sqOa9bzg6hBFOX/EPImCx45CisrYxwkDP+fGg5On0V
V9bAvcYiMlhjNasF9d+YN0CmA9F0AW1QjOMMygdMDT0TUrXsOnXLyV2ZYVO9etryUfWon5SN6po8
UvRvoCuVBuhM3Rbi1k8oo/0zw0gSvTexY668K3GRJBKBggV7D2A8mKQTiSvOrspp1A9V1qyLbvhT
+PZCW+e6yMPCLjqXbJccwFcGDQfSXbPWrPF79d+UKg2KwRCo2fQE8dlZq2/1W/s4TiNBqpt6gE65
yVXD0qZ4taJCRNwyvzpbUPe7oL0nSwIhgHYguB6R56HWrT3ma4XKcvkNejYqtQORDEqnsP/dyxsI
BQLzhJCgdaLLtRcCXVNbxA2hs3b9HcgOaEUVqlY4Tmrk4agCsyZc4/MsKFIzqZ3nZlkVtliGVNqr
lgeHExXtkPEFOncerOMrgwy/usb0nx1PZVTXhMsOzb3L57S4+Vm4Ad4eWp1Bf1GzRmRReMslnFjv
MAFq4Ayp8IrKZbnoUfE4VBqwnre/ciZ8dvbh
`protect end_protected

