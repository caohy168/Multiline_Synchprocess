

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NS0UzMRfd15c96SOZUCS1fp6CRs8wjCMJONa5Nnv9aEx79OUbnyoXsYSo4CLFDR8jsi3YC4gTGTd
MyvJDWUn1Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hZnsHcJwARteBAJ9FOgdrtMNGawTGbjcJtHea5OVEQLpN/1E3UZeJQvMM5mnBKjJlNnIIddV8i9M
joJgNubZ4x/J+5MH3hTdxxm7F4LSVBkzCDCdKpy8cg6sRALdJlGCLBd5W3fL/N1Vm2mvnpWYOTAK
o/bvQTpb6ITD77LnrhY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R5vX6KxpkN/slhDNucavw1UjzKwMJVO51VdByoN947hhTDMG4hIQ816kJsxI8/j9YOe47a6kVgQX
KY5bGd+cKmc7Sj/0vw0+AaRUi0BUjWSzIKXTRnPH+tW2WtD0kJSh+7VgTuQBcqSoKv4d1hTuP5JL
M95KyED97q8kA8W6/tEFUdFDODI3RK1AjVcoiYvmLp1JHE6N+4xV9DMw8xy7xHVPnxKUVydXS9ZI
5Kpm5nLDhGrx0aFmATRDTNL/Iz8QjDkpAArYSnHBguJuoeYzuJ0J1ZlDWpswin87gylwAFb44HxZ
nqHKf/UUdwFz42xC+ufZ21dbt3dIGLJZuW/J3Q==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kkium7vGgI4mIKVYu5AQtLq7e+Mob05Zqln0+g6ZaWnlPFJRayAUb2TGgpLHS5PtaVScG6fp7jAK
hR3jUq/6kPviQVKWL2u/4LhcA4kKyI9Zdi+ehWy6Tnh028+egFThp5uoINPpEng8RwwI+6IV9naC
FSuUifTc2tuuLl762gUP/eM/n8VGC0/A2mW/JvUel9ur+8u3BftctCYCVxa4bDpRr5qOXJGA4o6c
E4X6LDHXzpiVoyMS5t2r3OL/9fPqkK0nufzJdd4SZTXUqjb/RszVSlGWdW+08kPsxUY8m1oqS2K5
TalFYT3jg5Mp+kYfDfW3qlQmAC3mJl2SAKU53g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CkQIlfatrQuDsmTnRTe2/gzxK2zxoe5Evnu6XsZZXur5sC8gZMQaMz//gFgUkCSJi6IZG2S72YwZ
/DWOIKI3TWXxND32Nx/hdK6B+9GNQNAe73NLPLq84cJZY++JigrKxnm4um/tNdK3g7KtL3maNF+M
YJxE5p+FssMep7I1eFA=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EmZX2JV5yuh7StMKg1MKBA95BI+QbntliTbj9Ha7iFw6mcWRe5/6CGQ4XD+IIBUvXHSt9N3dYoIo
PmKyvOD4ATYMfvlrtSTiU0NkY1vMMBoIgaVMYc4MWiOOqkLX5QCr1y4tP/2tYFT0XqOadBl7mSkX
zlFIafpoH/LOglrVSIoDeBEC6MfVsaj2w++XvX1XfB4Q+0amZMXDTJWJMAh/IXT47EhyGLO/yis9
ZfieIq6d9JNguG3rVoKcxXkthdipGLh78LhCJkQ8FEwwGSvTbhQ4zgHstrRwdAASUDa6gwXxPpIJ
qqbHLfsfv3nb3kTfiGn3wbY3N0IOKggKgCcBWg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AboF/gdXw5XFu8Y69yIdoJn8uAobuhjjThXr2RSoL7EztRuvDZOCvet+2p1rluDW2+roz8+34B1T
nJYCZlru6Io6ivyh9RLqrWtjUfgNAh5bdGa3criaFYVKBbO5WYESngDLA4l1SKsY/ml7jdn559js
3PXOVkZ5okByUMAkBY9xgMS74kRNZbbWOs56xv4nvKv9udRIBNg9MIWZs33CMGZ6na7v3KN5Epq2
xwDAxNEyc/aoA5g51oYouiXbJQ1Nb2HoUlG1XOtMFCdrUfxuR2W3ymUPchBgVYx0ewk6YjTKjYY0
kbo74o6VcLrA4RehB/+i6DYbsVtsYPvY8u+VhA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cHkeoE7Sw1d0LekbvMrcrlfDu0GfJ9HoUw8fLhpsruaH0GbjCq3dlMBTPam2ODYxDCkoL5KkHnCy
Flu1mhCehzsjfkPpA1Bys07dlEsLcToR1mbANOUTbGzOUIoxpQY/N59lhLSnhvL4bqEb4ULGmsMg
tL3bvdV1qKnitWWmXgHqMeP3UEX52+2ODqtxSE+9LvBE/H0u+tpADs1/2g0UDOWfjx6qgqWpxcE1
nIcDsMEzJaatCD0P8lIqpMMXPTupi6XX6Jd8cXWliFXKHXevMkzZ66K/E5YBzCuv6OKuPSXVAjmf
wZJsjo1WqZ3g1O7+v5Eqc+ekE52N3vpm+ZqqMQ==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z7DnkfqlpbYa10n4bpu9gzVCQdqPQvlWpZyyy52R1KXRRDMK3xAnodeq9EtR6ZOsmm5PN9SkQqQO
l/gjwQOcIVAi4fVzDz8+IKXpDCqkqUS9w/NOg/0X3cTIKaih76PLBtiilbrPCaQggu4V92QkzQZZ
Yi+k/NGNjn8AoxTCOPlc8dFEeQxWTPkno4pRRRAxB6EQGemCa3RxC7USFhUJwDWozHilTW9mQ1sU
Vbuqq0D8vs8lzgHCrzvSriyzzI7Ar30bNUJ6xjfWiDaBEkoY4lQuo15QVyvXbvhwZNz9EXXXNec9
GB7pUSwj/cmVIDuz7ortZFaKgl4hP9NzontE1g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71392)
`protect data_block
1POjI9mkFfbkpiOOxGskTy8VWpLPbe/tfU+/vmVb/njBNae+6Zo0RF0kNcuvK0/FOIbrbt/sIKjS
NNoJJBC0S7fuhzWqi8bWiZOsYg0ebXeZTUsqdiMN478OMPM6njGb4pfkftg80cEDrO9eKuGFoC/p
7oLZSeckwm5cwhDmAHkCXdNMLrM90JNLvpL/dOAUEaT6T7SMRpLOdvluA5qXpIkXdXJ6SUc+o9fZ
l6BcoAx3tTZJ8+krD2qKbe+CgCoZgpDlz/3GmBMvJhfKug4HO+iGmDkv7LeAoSe1Ydjc1Z3ImnU1
mXT4IeJTv4sd2IOwnoOWyTaZ2kRpXliTAvh/vgpuFR0oAlX4w/RSqnL2My8R1WtQj1kdrTqIyRMm
NT8XurS9T9pYJ02pzrL4lMN9j/Kt2yfKglv/lNVYkjcjJYtkefJgsndceJFuI5iVY/kBde0ltg4Y
6N5EAdCnLePypU4+TL8faZlJy6SXKXXj0PSTJZDEP33RTa/u71LqM5GrbCfzX5hiRSdPv4LSNpKj
83qf7p9JO1li8qxH7fHmr+BXa6phlovoWMZ/OyxCpoIVeHVsj53SNSJSNbJaQk+B5s+WCCr8EW7s
jLndI9n8KzmZjcb7XQI1T8ul/pUGO4mtxjPcKtAHwwYOA2K4GQIw1w+lfknMjEy49dh693cWIAG7
36Y/Jqv1KV/W3fNjDM4Cf9VTOJrK1x9raKyYAir2kFooyuXldwGepZGhzReQJocMJUfHqPDKOiA4
uSOtpbpwwNJqaP0WHugz4F95kPMQnZSd8qoD4QA1Catw7KVOE/Z11d5sG5GCvMCJVG8r4iBdsWj4
RtBE5AAXNmb9voQ9kOspRSK1An6LvVKXn3/3Kb5FiulCxXhLz7lX2MMGD02LaOi1Zu5pTwHRGq+t
LIBE1QJI9NIKIAuykJaTyH7zkXtPZA5BJhKnh4ywcB9gWG1gaFAg7/iCQg/awaY+0GrboamVNNwG
zp6iDy6Wr5j27Au8lDGj3JbPRtjzf/0JGCkCtPeBECNkfMk7G9avXH8gNsNtp/THFtwnXsyM3w0L
E4bI9RPIU+M+o3FpSOzbphLaUSzzDvSU2q3foS8fmyO4mxuHSuYbyqp13zaSdHwG2Hts47+1ffwq
i2hPfJqBlx4B1d2G/lMgtY4PPGucxbB6OhrqbOJisvpT77lEcVMwiKucp0mPaJq5lB+dAu5KBJL3
iTs7Z9qdEgadt8Pe9nyQNZlDvK3DQn9SclydWSL5PPqTBsBSMB4Dq0T3VS/XalLVpmmpsg2xfFQf
ud2+nnF84x8PoQXmXmqGKoa1SMwFln4fasvU98O12h6SlPsQVz+G2U8LUbvua/A0p/B3Yt0rXEn/
ZHww8oaLIdavHcjAKDXa0J//LKdI8NUDFhwXLJeFUI2MK7DjXL5jExJ3teifMFablWjyobH5tDgZ
yUvMEK/DrXcGEuDcf7K7XXaXGu7e6b9B92MTWWdXykFYCY2QL/C/CcfygMHXwnjp2Zsiopn1i7Vv
39w1Mx4HDuVGg6vvlXF1bUhYph9xFLguOpaH5QFIDbZiLQNnKyCgUDLyNHCuFC2KzqOwC/xOBNOE
Rj6zP3293wmBHRO/Iih5smqBzJZM1KdxRKyawaihA+HxtbgGSv7yamYp9ULxds4q3stBe86qFVBX
2sJMfuz+G6jXazMOgX9koD1iSUD2yjFrQR1LRULUhX1/vHF8jqCcaEEoggdWrDwDYoqIqnJCv4HD
C6uieDxRnfND+ivgjUQGXgicaNHkqD5gkvJY9DO+NbwKIt41PNLGkpirq+PI3PRT3ZWyqbGVfuhu
090uK3TwYfR0hoPKeTNYA80LgOKKJ4YCcr8xs9U7NGGuZ1kVWIpGwxD77VbIs6iT6JvZ6Kcs4uVp
Q2x00AiXYdc1z0wV5AsFFzReR/ZNe8T9bqd13N2MoWzkb+lRlZpD35TDqDFJx4IAS0P+BX0F/mj0
vM+BAJ7jNxC8DME4rC05oGSA5Ti6honURxbOHpScGiMz983qbp1nigPR39X1GbA+sIpfMrXB7ujo
CjsIvEO45j9dbNCjijqnwAoQ3qguiQvBWzkGGQU7G3m6N2y4VC4qxcA16WntB0InrVdaTlfp6N+B
KOxziqgMdrZZrwASQpJJcS+RUZw/sqQd7MobhgBBqRniHqhPqQBvBluMQsQmZzJlWT7NEgtujTyt
OMNR9X/A9roUq5Hodfrk26euBh2T9MbHf3uKVbsgh3wDMvaeEDI9vlTb8mDS+sObkY4zUp2qI4+8
I7G6PC3IsIaiSNBSASW+pYDUi/xgKUE3LkNu7xM3aGE1oatLV2xQrEvGzcQkbP3gUSKw+a49EkaT
PId7jV6arhjhmU8C8l84PhTmHvfq4LXLvL8NTPlYa4Aj4O/YSZAKlzVSlKA8bzXdPzHJYNAKrkKO
ev1YlmePCkv3T8gEPt30UMWLLoyUE0WIWz43YdH7LFb2HbFCPj3cU+nqm+x7pSNPDFw0stCqxkop
2oZwo13/WnldDesF1k/HEyAh3PiH77N73aC1EV8BGGm57GE2JBmg6GbN1a/iLF5DtNgG/3YyELiG
jmO8Ikax9Z+q1QVcm5GkyK1u4mZ2/6GJwPRdK7ZcDzUHNpW7EDfP6vRavYw5y/eLLflYZnBKv0c1
jUmUgYyzPBZ5O5huf5KcqqP2lNb6lFaEgnDncpQav9i7j4mNOdr9BfY0yVVeuBANgtXbFkEG0gX+
1NhZClX4MUoQZ4rii/UkoIZ9aAgx7FaVy01y2YKjKHT7C3JNMHcdclhdLRe736hTX9sYLu7cHiKV
c0iy3rot6s1I6ZrOoVy9Z6ixCj3cOEZfe55miQNnBZxJ3OmBxszYms2GKtRcOvrbqDiQPuqvaOAk
bSfEQErjkdsx8S3tjYvJzSeMzJuTMAQ3/+SXvsttlaN98J2Jmky36SBcXg9wbO58aFi3usv4g3Ij
USEZbRscuJpoSo8v6fsXfhd08oosTfR9JqPzAOMmNZgHWDm9Z6xMOC5JG8KXVxpwcDwsOT8JhnFB
GmRx4ewwpw2xUlmsPDeyK8uI+m/q0bMhipNCWew8CHw8WA426lcNwthHcehzSpQFmSdVm0mgqyXP
S12r6XI1cdfUsJ0htKmsFH70vtec+NL7XCvZjIZnx7XqJUIBRgYeakliTHighkTCTPcn5ByZwknT
EPCqs9MNST/gksVc+i0MQ3C1vijINnVyu/z/x1Sw5GYdlkRtcGZHBIjGa7fWflZSrNfVLbfqfDBa
2KtZxaN7JLnNKrFmWSMwc2SS1XiWpw+kNwF+gjbEdPEJkbJohYaaxIg1QxKukHncfjzEXHogz9Ff
mIkXWnIscFPwvgbLZe092Lk/191fZF3voNn/DMhXm4rAgO4oZrhKEOSCJAk2VECxd+j3G+cx7XY2
klk2LdonZr6NdblxbQeaJphgsIirU3c8MQw6QErJNfP+mBYynzsC5N9qlU4s9DL68nbT3Sch9ung
HKOVQ7zMfLJPR9yK/xYVOG2eMiUdvrSI14eiABdAIZf2wM3ep7DIqQaSyXMumPQzcefbfAm4eNB3
fmzOXjnv+L52VmjdJXqWVFiDM3kfQHU50fSuF+Mbzkf8iluRuNvjKxMxuyRaWBcxbbnoNCL2TxK3
hwZ/FLAFT6Th1EbL/1XGfUC+6uEPjsScdEx9x+2V+le+RfQeS+KdGcXwIZGDhvAaqB6bs8OKVnIJ
cZvf1PoHDodFje/ZyqFfa+n2M+d9gDW3L6+VW5ce5L49A4mP+PHev92lNVUOjmHnFQagpOENdLaJ
qf5tvNTsxCujMIxCqzVekkInPN6P0JV6tsUp+XzZkIeGtXmxJPkYWAuU8YaBxcWfOFITFjPlxe3+
gBbEModPQ/EoR3qN1e+g0G99e4NuECZNTmsVal78kME4miWt5g1l6Y/AZfpT8zDgjIPptwzy7TnI
2ljXpmSLqWogNcLyjaeXhai5blCeOS+lqWr8+OWIFEovg0hFf2d9NKYqT67lMYWpP3+9tnLrX6C4
imOjvmQoOPrdSYlBvyhIcDDqaABvGkY8DKJgfCyK3rio+ax78EZbR3p4r/sxlVImcyquReunMxSy
P6hIlOaR/rpnO5Lm/Jvc0DWSv1AQ2U6ZlmXOxHsCFyvURHhU3gHYcNiJt5izgCRvX6zKq0ibs+BP
nqv+na9Rj9YjKV7LIf/lFUhX38f044NYSu+D8zJ7xEDO3F28SraFqIPlblj10FHVCKlEYdXTVfK4
Ftdj/Yh9lJT5wyyDCumpKzFS1vYxuJGNeAkwS+Td0RMQGbKJYrdKLE3fm8lZzFvGBiX5xrYgOCjg
w73JwBnoyuKbb1T0o1pTMm/gPMBasQmrcuqV34VanYgyZLpFCPlUwWcFH7m/J/JJduCsSpwvgXhG
bK9jBw7txAVHs/XZoowoozGUYSipzo7ILNLiplHEAfakuj/gxjU8//n2nbUfujFLUdZshTYlDDOS
rDR7UbSLTChKlZ71Xui0PICFmospItlBApx7ovJF/hMct0luKteHd0gKI8zqTaQDIc/bZE7TNBi8
RDjqg94HQImjELQHLvjBc3djo2I5gocagyvJcmTBVfx/0My8Y9kJ2mJFC1GZZWnEO0vXOPAWVIoz
8qUUivKHfob6meprCEhS70V9Bl+Z3Ilp2wfImAMPQImX8O+wSK30JQ6J4XVS6BeYTHtwuGXSCkZ2
4B5t2B1z1KdZpmWN7dhMuaT/jy2up1cA2xtbrufVsRnlc9v424h6d+KQ8jRWWPl9RT/3N8L4JyuA
yBZA98BOZpZ1VNtO2vMgJ/jeIn0xo2xhvAqyB7dHo4DPtSW5WSDBkKgTSl8r6UTVrHUQIq0sjHXs
tS/KmGL7wyCqExOsUR8+qFBnhposgANYK10Lq3ddR4aPmUC3YR7dA4o/sh3gTuSCBAcVyI+RudPt
D9baOCAA3Qxz8sswrcGM8lx4V5HyBNg+R2Q8B+RfGjGMFVcVx0O9zsQPtEYRWdPZFKcxCp+Mr57c
6pekCbgnlhinIFS8jeMnovakRXSZdmYswlIXNf3WfrD5oG0vXec+c6knPv2Dozlz0ccVksNWIf3Z
aC4wrVn0XVW16TC3067EoCjW2pIaUMtD3V45qProfdUXI5Sb5/+JJObdcx8W0KDM10MfoKgm8ffa
1KzXNtkAH6/P4B6V1KtgmJLGhLZAdZAkXrBEsvH1gzRVSr+UqcF880mkKtfXkUvD1RYTcT3sD3rp
5hkifH+WNgETkj/KI7T90/L0K3Ku7wv+4IAp3Bx2JdFiuNcNy+eDBy79UKDuiDozOTRqunUnRvW3
0KyDTe6wPGWBKJvWQpN/I8sk+7nwxnmzu20jhcC2dZnxs4uvUYIa6u5C+XP/Z1sorCGUYByZf+zL
PJG4B0LPyAncP/geAV9bWAdFKPBEOIWF1EMeFuw7hi8IXyG0od4N+yDmdGtqTDhyHq+szQyEiXWH
A68WJ7xa3lInwH5mJ1zKLMWQwz387a6Jf/Dp0c+i9vFF1GfT3Hl7nOH9e31HXezlsEIudbE8hNa/
N1On4gUxkGvICCX4onVwhiuq3eyDUq5rpOKYjzipKxKuU0JXggd4Sj4Qt2WHpFjcWZ6wQxXG6JuV
ktrp7+xDyby3jGneEIeCOXPeIDRxUx46Im3TZAwEDvUz6cS6WlBlQ/JsN13/Z4G3QFF+CwtrQTWH
MBAN+DETZ613t/aEhNUOmttseSS0v2acYclzdpJKjQibscRUw1P7YOU2jT4jWknZ2uCT/p4nv7In
czhDUYfEC/CnXXEV0WE+sfRi0PC98WDTKsiY5QqFxNlASrdD2WR1jZFzTmoWNYV6dsj+9LQk9sVC
wovQz7NrlUnJq/pL7pDWhBs3d7gk6Hnb1LciHlNfDr+FRv+H6+4Kj4LnIEeyrqSyAGzvNHRNCBcu
/KyIuoGDN9MxYtw3+/08r8rr1Q5e/k/OkzFND3GR6p9N0bU333RrTx+Qe8KnjVZeerFYHLaGI6rS
x945t0bsWak4n/QnQfMg6RXShci54rg3LmN3TObhP/5YlkWF/tmqirc/+8J0PyHt51PXFky3+Ao3
7pZawX88KK2lLNnw+HiSj3kMA4cG1EyhPGvWJGM8F7TNO2Sz5DHNGzWg29lhcatK0+QwowkQZEuW
KrByAwTP3VlKnYs6TSAbNBHlWbpKbu1hmXWlfELSNmsVxwmLiXsbHlxtmCfJS0zUDStKFRYfFfoI
SQ0Jk/7jZKBITfXn0/V/AUd0HU/I/v0cjZ6pd7F1YbUGNuqy9fPwecxFMG1AYZp81nT/TXal3ZNd
Sw7VTXiLj678J4GaVs1riyoHqxOCEfBcwFXkL+Eqly5qS3e3h13zx/nvx8zpuzec7Fd6BAeSmsIJ
3Ii9Gxeww1uu63+42dD+RiCX5noabxJ142zMDhbTej46XdgiABNTwpMLnhkcBykHfuTWk7oZIm3+
pVTRd7ZM47HY0WGgcECluJvLREjOuC5laXA5qGm8TI+K870qBlh77ZHrqNw3SsvVGuyKxGsczJ8a
86DgP/vDU60o3fJDcfhWh247/SgGUAjpj+AtWPMIB3MSWbJWhsWQ2ITPuWtxQ0QiuO1IegodivGc
sMRrBGKUxXbhCoznmSRciIjDhD64VCAyjwO/hA++OD2IgyV2AstP2lI3z2cwwB2nb7GoRCZL3VYB
yJHXjTeo29Om0mU9pNWQgg9jn0MFyhfj8JmSgJyxqWZXzv1swz87OVfv3OzJxRY0tld8i3HLhP6B
fvZvndEXntziCiUOfwQPiguaC9azkRdu87D+ur4Vd+7Mm+9Aw785g4j/TZnZitQaZBGbkWcUBn+M
cs/2YHwDg75H+1QRx0+70dxBdwby23cVsqqua4ioy6j0T4D4FO57StJoutQ3aWvfgdMo6USYYxpC
MUhLG5h+kuOjbRQf8G3kX5gLcamU1DkMdWs0G+i7sbBoacAcIsKL/UeZF5CcTflJG8AynQ8JUFq5
mB7sLaIo1p4884Bw9/kC/fjqEJs7hk5qPt5n+53CoZcIxG0NYieO5iXAVl1Qui+Te6rfiPb7ER3a
T7F3qPGHBNv2UerfUP4xv4ToDF7VjzCpzzFTomgVyxm/jdHwd5ckIi+JgnTHgnWWWzDTQe4YPWl1
tZuKSrEj7342pXV1D7+h9r2if9o/voMoPbwiyIihMNyOpb9flucKcqmsXUa78CfgQseop9AR/I0B
6p4OLWUvGsEAb59edtaSpzI0QWa0/reks4+BX7Ffq0KtkCum9DSpS004LRK/iFB/I8Sy6NrgM9+y
NEbaia8W5Botwgwm4h9mpCUHcYyRSb9dciVSs2HTTs7rhqIOK+xjfGCrgXOh/jE+9JSlUtg9+Bdy
M6+Y666sdMMQOpykcIcmtomJ6vUQth1xaKe8GRW21ARmWuiL6NTZBDhzU7IukMmzSgVwvMMNEB/B
9FOKM4ipNM71QStCvlxMm4oTi8ulBb53+GPVWr7zvFRhT4K4CyhQ4Xa31VX65xaocdJTBkX2KigA
jvqXaiyGjr6E2mpL/P/RmqPdS9s3Amuv3PQ/5Tel7ofqo0ndZ9ZxR4B7On0Az2gcSMUYL3D2OOqt
Tr5aGvOXLsA77c/wN8PAIo2yUD+dKpNnXMJQQIBj/cTrK3Vzop7wTevuPUjL93NdjpA+99TtHOyL
lHQs6xLLOVCY/C9cabo4cwZjGY7/LOoruvWvPWTu7qtvMS10V5+Z3MTXd/w1CIMp3iYjGn6BtMVI
jq0zQhd/jZYE6gubfvq727KNxLHBAXV6Hv6Br8LXZ7VgdI5RK5FyS6fesoFSF9RAl0xfiPOiJwGh
bqmJM8Oroa1hjdOoi/ULKq5lb4m+Psc/+sK2iPsboW7JMBaR6Y/H9qYqAiWZv3S9rtVYgDIN2Fr4
hKbvMHufUQp7XIwi6Kb0GdpX1p6PpQmX6w6tpqhIodK9Z7YctaKMBpIt2w0x2JhPvsMxcKSzes6j
pO+4Xpy/TagBW0AOru93bsjLnq06GtPsvXcwyoV6mP+vK1bbJUE7xzM6YKyuRCRnqHF2TIfOL/DD
tQT4dqj7XuNLHJ7a8Vu5yIsfqqTXkVADdMZ5bEVoJMN5F4HZ4i97qrIIbtFoSz7Jii3v/lhzMmh2
d+ewWb3caAK+NXXB4Ex1ZCIVZ1wj2va78oTii/sGP6pMt1XuLjUqJ0iqkEo4itbiQV7mFUJymARZ
7zl1c2XD9CETRoS7/mpXnRC39WFa8nOmlB3FIpyDeEUlb6F8MteDGOkg23Arsg9NTaxEqmRH38cK
6SMz+qR1hCVj+/4tl7VewasZetRyVWQ6ir/5/ubRo4eyXJ5ngqNGg82Z1j9laRbNjDaj6JnSen/4
ftvPe9P8hfEBPgA/YVMlHkF1ESt6N1gAGPbbQXXZIu4eX6zL79En+jlBh/TvC0S8Yze4mJL3pPpX
2rwuEuCy2EHnSxX34BUuDwb1yky+TSnNREOq6XYsqnXPz3PQqE9y+59T0rUEjNQE0a7JGL9u4yUS
kWXxJxhpYnq5Cc5TgA2rAHITZGCdiFUL/Ax/reyntBF4ysRZXLVB3EFwYPBYyBhkO1nRpw1XRorA
mAL2xPRPRnR+zkqaudS8IsmzB0G5QCdhBc48NwoqeBUnN+S2p5TQCWdZzlgL3U9yMAFAwaRbzJYI
bS/HUw1+yYbF6egESir+2DMx02Iz79ce0yew3jP04AgGr8YSbHTCQGz28bZRFw1MMId8GXTv5t6g
f2HkoIk3BO/eLG49jpC0Mf6hZXYmeI/AIpYj4kk2YZN/2dUrQlKaxhBmxQKq3mYyLy2wVn0c6sCn
fPqCiCMfa1r/2Gqb8duaXLWk9Fkt9nsjo6q5vVXLluMQLpOsqBKyw/4kVIQ7U7/e7r3/C+3U2DC4
jbxFjQFUhlSAbRr7ELI8Fqg5A+IWO3+SmoW1roXk+2YjmL/YaGpnMJo3xCZ8MJQYx5Vcbh/uJf2j
ZcB4mftQZWd+6Lh3Jhg3O97cJTxF3OpvgBNObUqr8t/a0C48ug8FNkK3YjDsmDeEdZSFSOPCVyl1
P2Tw7ORHq/9SM9mZWl0lKlQZuYFWaRWuwOuWxCHvOb8HgN8GIIgM7Fpsa6vhhDsrdkOj2lWJDPX0
JFVYcUi/Z+ijYlaqDeMt+0AKQAGNfC92CfgOxjn8Dx1jnTtIHGmqjSH5g8OajicGISERvKnQGmuT
yVuDci4+8cuXAb4x2eiPHdO00aMuzAGLGUfYaRGyW7nCgDgqtZOnej0Yiwr7DIyLYmg5Hho1GRIw
2dWSaxgiaNWUwD7OzG7NGcti6ToMbJtKmIy3azjuKiqAAAohde/yeUQHZYRE+ufk6r1q1cO0ABpE
wienceg6ASOwiyNXyXrZ9RDvWSQWF9X8TVIEOskdOoqPr1MYsCF22s/RqXAldZAXu/hMhaISHDIt
jZZ57FcZOntoT0rJFvZ3WiOHMu55puKrE2KvKOzL7FFUmVU/ZcmTEIFEoPkOYJhOoRTtyyLBwCeA
QAroOsbRPnuBKTHRAhSxhAZ5+1dVLRdFZSM3dRjmZ8PRaI63a3x9L66RyXxeu7mck+nLU/nTwHK4
ZoAy+xbULdtC5UTm6HIYBelLy1yMVMBBGyWaiWTX412DsakEKJxgZQ8UVJLWV7CmBiZv/JIKen2H
lCJtBE1JaZ+C79vY6UmTiSncQVh/HQgwt44F4ECXGKxkFYDv1tjJsFNpx9V50t1ySUT6HeyEFBLC
8/i1FaD5oCOvDMT9gPdpFhZrMpmf6XqNeoLeqGHl7j1ghjttjLhm/6DZ7+KcosUWPaWMzr5Uii4p
fXlcYCYoKhtyL4SZf5hOcDeqHSnFvphXiaieOLcdjAPomIT5DS6JFZqXajWldSc9BhiqywHUwx9K
OGum0EUSKKPtQ9F28iZIDmLMfFmjHNs9Dton+1NgJMi4nCmBtR2IyJ9hkuSz9E7umer0emJkOEDQ
oYltncwMo9QIdI96rfoBPq5qRt9we8C+YCZizpCCS90ehdgOFpTw8ApKFHpPw52aBbtzwtbRnrf7
2mG9UH5jF8+UsEI51/0D0WEh2bn6Tv7P4vZOqvd1l3hAJtTb7t6qD0E2T3YTbCECVkBrLB49n0AU
2Ydze+GLJOOAe0U/A08NodkjNdd+fYErj9G+p8LpXGxzGy1+KCvewWNOuV3ElOQIvB6aLg+buOO1
Ia2t2S0EPap8mFuy0kW0u41OSVnVMQrlU3DOHXqXzJXJZXA0kTcfNOFoSU8TmH8wpXQisc7R6hUu
JnR2m4PoLxVGKVH+g4PXRz+pg53OwTxp5avHaulEGICm3Obe4pW0YURKyqD7xhbtUn3PjwxqsgIe
mn++luUTRwpss3TLt9nBsh/LSUR7nzsiKADqEdGoWR6nt+5WzdEJGUZ5L2/yCgonq+WtfSu5Yj7g
AtgnrwpSZdCV5el3yL00aNGY0XEpxPjqFULIihrS1kYW+s+z7HusxGfE7vU44W90j6qIVhJFl0pE
vYIBNPeeag48ecgqXRekeZPYI1/chGt2ZL6lxl/nct709XqjqE5iKH3UtPQDc798mi04r/hegE2X
zS+bTp9J7sRWtSvDNEKfgL+MfKG2waaLf7ia/ZuQTLChnnyP160qRrcSTDiHpwx9KGysa+GzRD0D
M87OIwQSo4pvZ049IPF2Cp9TVeEdD9TvzHXccAcu5QCetP3vqA8fIbwsK+wCnQx/PJQabJBTk+Nw
o7ml4ni9jOu03YEhm0jyrJ2WNthWACBYjjYoMikC0NHS6QpmA4t5MkC7OxAUxw/wSaAo7+w4zeKn
cTQuYHXt1b29bXEKyAghzMnqGqwRJ+mEOqi0IHc2UlMhBLA7aJjVo15KztKnZprtAhskDwmFjFXU
41e6GNnQXZ91LTmg8MlVI0roPVHYYyTKaXB8UEYVSi2bTHrj8QV8QM69VqWsgyaQQ/Mu07HCgYXS
AddYW2PBVt9tp5a/Xch0tdWRHVaDjkNS6AFnsnyEezfzhgmIaesTLaMU7pOBbvMOEx3pDBLZH4aa
6AIZarTD+U9nLYnmp0Njmt3iSwhYCkF80ODFTHNHp2A3DDgtirRpH9fe5Nbv/ke1VHySIQN4S5dK
NRMCikoLrm7UAo4IS3gcwnDvcmTPwp1xjlu4b7BHN/W8yXfqnArVKTjPEXnbS6m1Z2UQJU51r5rE
m6R1D58Xjf36nnRq1XPGaN1lnoohIWtXft92M6pptTrDgHmCbEC9mV4NoEEgRmiRZYW5DLYcI6kQ
FgRQ7YYjlqmYJdTSlBUyATAyI4sY4eS7ZrnYqelwp7c80oVeS/bAqEvqhOjcwugSmFNn1QfR0MQF
9nx9GwDvdtOjG4pKg4O8xnLAmovmoqPxLbLHE2qEXAKg63+SkVfpbeWzKgdjYqRQzKTVUCjMnjqJ
aI1EztV7lBigHNdB2sSaTNHBC00H3yzHaqZ8slTzKSSk8RmMf/dHg/skA3kEWBffg9ChA7WteDXv
xrgA9rtDdWGUPzG5QBOjlPEgZ90LrjMhUZJmUCAm6gQ9HMkCJsr4wAHb+JzKITaaHoDYTldHgxpB
OfYbO7AdJMwa0Wd7tilZZqdTcpjbedtgv23w/ne4tm3OhhK6lQFlPi+nTl93YoRbbwinEXubhCxX
TK/sBIpF+KuGoq6O2DnktBsgwkmKqGb78BlGsbcqzHOSOxyjtP2pt6hbWPNO240E6Z3h/DR6kV0C
8puMC0PKHJEJAiuGY7ySgFDo+NBE5JB2EAKsAKrkH4aJMxxhiBroy+I4D7EW8xTsOzY1BC/bZggy
KPMjlHI/Gt3x2CAtkfWok2Wjly+RCzdGC0CQWUN2BkxHA3Xx2VeXJLPSR3wCEaR4HyyR9Pir4/mi
TH7h9VQN3mv0UCP6/gkMZ5bzH9S8xQjdUIeXPNfXyMdkz0XUmwfA244X1wSe6FJBR2Rt+aPh3nPH
dT1hllPuF4f3D7k47kgkxy8TCc4G8MZUn15bLPwhrtZFoVqGjlDuYSDtaF7o3zjK1IdA4pKgFk/D
6MWT+aW0YM9gTqV6Yzoxkhqnw7Ii5GnNmcc5pzNGqEJ6aMSiRThTbcis1FHHi1jdes8NJGLlfVV0
l0biWNv5S4UD8QelTy87T65xoqcwE3R67x+IedCTtYhfE8fAKRfBmozRlzRHEwQ3PXRCqd05xhxh
yKB+bqkwCN/afy1NNokmcrbB/UEVMxNIUNzSWvMJvIaFNeC9E5t006CvMAR0SPT/n60QQ3f1aGan
pZ8PiyXTm+2v+27lFNKPcwcFCF+K4w3A5/RpiXquuswhFw5XGSk48sBTeDLWv5fAqYsekh/fWyaG
CpmRxuOZlkBcgyOahwX2G0O82Aja1/Swz9Dfxg6A5XhCJw+XaYOHZFeAj3TlYhuE7GcUmR4U0Q0v
GKLy4/WYbHVB3gJMTZe4sqR4AlWeMdsuuj1fOya7bTw/cspIQ1FbZTsVT6NDaz9y6PQZ2O+7t4N7
4yUMImcOoUGJR70lnAm9gI5GJRCW/yGZiH8U/NQwweA+HqrW5PF5hVuUcRbnCH+m69dwgsye4oSd
MnVnHhEeJEgUR5oblqAYE0hX4c8uosSCggs7g8EcX6LSkD8/QdUAZ4jp3DcM16t2HOIknHd13F/4
h7cuHrVXvMzWvs+1iJyjpBLrcbFs5PP+oJnaipGqUK7xBNkK7HjSxr2nkegmWCTIdRKfYjkB683e
aSVBNRNGxlQWo1StjTStPslzedjycJPSk3bz/rtEVb8V/6L2+lJQkL4f1pKC9kAHB48H3Yv3sDeJ
Uv+dYAmX/g8OZopMUxj1FnePIZDYb4RqncXFCi8FXqRZuxbnotEYv5MEtsLYu5obpwdg3kMPR7L9
1fjkYfV+u/FPCZt6hE5IVkxU/ecbf9PF5zgk102/e2r3t/GK1diADEbtVOYX1CrseyGu73k99U1m
KsKz71LjWbR5DlisfG/rCoxBt2DgUFiXPFUJD5vO6PEShnDAb37Fp91LCSKPha/EaJVhAJvFCPGJ
S/e3fE3utTsuuTxQJDRTAXkgZAH/1U3JMmYe+H4p3/jAJ4mO3cyrCY8GwIHaLMryt8hkSBYdeHZm
rhBF6NRGQfXEzidQOZFaPnfvb/c8U2BzBXBWtH+69oyPnvEm8ETnrt4CFVWmOkh7GN/ctnHmgpfc
PQsHBbCyrVEI2vMtHFj1r+QA6KMWA0JlCiRAvNjzIz94HBjIeM0ujxmgWkOciKfXNcNPsrHCzkFf
0YhiybJhZZ+k2VCzjl22t/7Sg83ZhJSULR7esKAuPG6mkUQ5QGFHAxk3rDEWJ+9lO5N53kb8kwjd
jtJbsK1QnviSQ1V4pdY+s+FnnwO8uGqT4T4fMboCJUVppo9gBzY0UugyuU7kkL4JtSQRZiVv3ulC
Lx5hs8/Tf73WCSvYfnLdeyNVzsMhSiQmhbYg5t6QwtNZFbMXzO1HBO1Zzuhh/sECyp93Ga+tN8y/
DPyCohHGngFc9h0zOvqdaOiBM4rlxIc/B31cwlSaZJ+sIcmn3hH2H9TNtrPvDY3p1cFKfZdE/rVg
iCjppSq6T7yurOExywzONwZiQQNRLi5FFEHjf431DnmEZuFj+MEH/wWVJiew/QxAQ6hEI+mZwUu7
Gm9Tqkluy1YY0baA9p2AejKyNlpwP+LKicdPRR6Ys5VC/v80fSRb256jQmQMXcZsaIgeS1JuENNn
cDUgqtwRVAJARq2UJpR6vUhp7+MRAob2wAhyvVQXbk3COuyFXTWm9Bv7/RuTmwt14g2BHYKaOkya
xBs6AADOPPnsduDDFYeVS5sPOKDCQJlgAh6shGmaJC6g6eHSMFZWxTnFJlSZUQ57O/+Q7QJUGwcN
DmpRyktTMl/gS4k2+Gu3J57TLC0VBwrs0oYmcjiQWa6cf9s7yHLZwshIl7fNPjvO4Uq8K2pirLgK
IBdNt/n9x69ZBGGjBGdjDIOJ0yYxXFWuISjkkLE/jRoUX9/9FLGNgZnQA8QdeTXDaRecIUUy9aGr
8stvhj3f1IJMxDoNrDqaogXxyfWTbhZf4m4bcg63eS0VltzaA/kHpNNlVEUTVPL+vC+j9+08AeST
jzSEbTenZgWCEkSE7EiJag4bVMYzi1t8PcOOvyEc3XjV0PRePYZltUjb/ykufnU6mU97S2J1hG4E
R8I7dMM0/8sCTIsrh1/BsNtRrnvD0ey7spwduM6ZICFSm8SrywPBRPYsYJU4l1X54UGhp8u/50Gv
Y6haFYv2Aik9bMehvU5lW+9OIg2EuCwdr0umJ5EhPAJ7IXEK554TzRkYOPTylZOG+ueA0oA7POTI
/08MMqDsmzPd1lv8kkwIXXtRUhQSs+1ojnJxbM2ymxMRfgKNdeMKd//FW53kbD8vE0W4xpCPcC2Q
/s3wtExXk/gwu8rOVyz2u3NeADO9bd3DXP/3zs7a3qaKnohACuaOm6CfM0AM3zuQKg6NzVZxODZ3
OYl3rG3vuInWIpkX/BF4boiVhJ3EyuQ6jReoMfd5vIWBqCjxrvq5WdEV+Ya6W+6AexIEFmqOw9n+
fh1IRVswl6ri5XbBqNBGDNqrDjoRcyLV+QtaYTCZ649XY5Yq5/Ro/96VVGpGKIotA6s/f+NgzxsQ
W3SG5EAZyQpwkUxUot5wotpLVM+ljMaqussKFprHVIIg7aXsRWsTIHaaERbeiAZpRjPGmLX+HiSv
uNgnNsvphEaa1CPy8iutsfY/jIVlYR+AHJ1Do4iCHFL2hGBRlrEEep70GYC42Y4eaIesVUkH38ni
lEER4Zwwd0HbeC5+Iiqr+VvbVUJTA42hWcwxK+bLcpTZEDQuNeAPtRpAcn0psaC9xRknjF3CV4Ol
8+dMi05NXprmx6iLPVoToufinZUk5ZgKapaoQDatr9mK0PIjodI4ND+bUSkybbmgWG2q9pMwptoa
xUwwATkYW/a/ZSjvzX4S2L8CWdDgRmM+i972/dObSZqguFoHbVErhYqZa7+058WPDIj0oG6QZbli
8cDzCIADzN8iSWUZxKRViiUG7poo8QMR+GbmtjlBf4fQQG3ZjSPJGC5SuF8ZHYLZiytCBoRLcUch
TO+fpVx2iEFJ9JU3P2DBpWxcC/vzyK5BxhvlfCw60jR0gGU3KeyGSIgyPglUWo2/9+/pIybCLo75
WKlP2PnAITIcNTWl67UuiG9Eqw1JBWwWgNY32vlmFnmRzrb4U4fsXXOSnr99hz7CDf7wzAYd8I2o
mzldxOGgvHHb6cbLoTvQeJHS8tT85mEYjT+l6UPPxSgSBOdNiH1RYoS58BdXu42edYpeZTjQHu9s
UD2jKErXzFus4KCOMZWRM1jDBXf4pFom48u2bcFm5WB1AfEcXC9NucfXl1z48c/9Jb+WbOQeM7Gv
rnIliM4Clerid5YDq+WZnVjECsuUWEtLE7RRq5nC2sOmGLOFRIZMa0AaB+rQkANTBbNv2a1NYcAl
5IE29RzmfopigEegzUCGkmN4s9Hd81Bi9jbu3p3Fq7PJY2W9e6wHEiogxKSc88Q80C3Cc3hcfwSe
mer5jW51/m74Cvw0d38IYFvfGJX72eZY7wCumpXvnANBUhbY1PEOh/6hQFbbiXQkBXoBO7U3eEmP
lo84jml/Gs1kld3YfMjVr9GvxRcaQFnjVv/xs216EEfq3+nJEb3JDZD/NDzpxh7Km9WFgytoBiq5
ZMKJyARgPtp981JQSN9PFau2ZuxVwtSOe/eHP2j/da/Ja+G/7I3NRyxbYA5CZQwkzBbscrqm4Hw9
AqWtlVGG1+kzJjkk7ZzuLCh4+S/xE44yeXSxmANiqpJW8Lqa1V1HuW2zdbtJG6ISbm+nP5IVViWO
NCzC+iYFZgwSMGn26dHCav+s6pfZD1v1BP9N93TUFNYSadt0isaw7+IWxiFMnziB8tO2fTePyDJy
dd/GwPEQTqrFCHh7yEhb8Klh2B3IlqwQVZaFSQ9pKtidm4GcYlpauM6wByfXCvLjWcAn6Tl2EpDf
jIfbsKrjmflVzYkFkUDlMEopAYUrQF/jX7sr3M9zWIngV5GCvdTfZ34T49pALDcghWurLGB5R53I
VwTr0O1qcJvAdBWPSPV31lsRmOEqOOPma/C/WKP5KLXgugQcbse0XgYWZAbuURiu8M5lZEM1oCY3
JNhFzhFr2N6mCBZOtzqbeghI9BQAVxdAiFEGu/pkag6lUrMOu+jHZimB6md/JY32Fxwvn6534DXO
HsvB4WMyoNmrX81hoFza2/zOjF85w7K6+raAkgSti1h4MeP/lRuegv30ilsnDZNYGLRSqGzaktj/
2gFxb0AeVUXvwY8HbRA0RLeQ1VWyzplGOsyds8bvEparXvF3g0nwSkk+iwCrRmXc7DUf+zE1MKlo
9J1K/Sjl/kb61iJO3M7TowInljRu4+jpxSR887hGDs0RIqPG/H+/2fjlJDUKtNR0IOHPSCfv/4fa
5bEObwgN70NMlTRY1WXaaPeIwYSxz8YVWcT+8yle7pm9/H9pwZ5paUt7G43cT6Bgv585oAzJ2NCp
0aNbv/zh73xrRczoXd9XDjuqlj+bSacXhEAj9rH09X3JGAP5WvU+OyqkIk4mC696p+yz5cJQcq+T
LL0a6xm8Vd0/NLA3QRmujyPi2zVrGxi6wmefm+Xo0Cv+yYwuu2+OknOIAtnl0q0VKuatoiVV+z3X
xCxQhXPsrhK8vlQYN5oS3/WsOi4X0HElqMKXAqKumTbrnwkslzXlvdYdMv2dcYItozLfq+pI5GYH
5t4FypeelsOanimvJkgjrhWjcKNQfSgIB8/7EuiD2HXmA34J9419bwlSZLE2OgTV5m59+hMBc5z+
I8rrDQMlVDFDhN5nH82B/Vai69kr9FMlLgTBZGRrV5MtNIOog8dehetg+klLyiZkWMOu7Byf6cbt
HO3IfSWi3hOw3PLvijzMp93YsV8LR/pXzTNuG/uG/OQpQ3wBc9JJtH5JDQc2udDXlnEzHHbpIeRw
jThPigjRPRvu9LqVcEfpcqjnvD+S41+QMPuVuVX1Sys+U3Ad6T7Sl9pGxTwzTcMfN344p2szNEC1
h/ohW1DxWnAOlbQaqBXE+nuee9EvPY6aC4RBaKREcbTMxYyfkGan1O6/rHmaaj0ybNR+xWUDMUfn
lIXDhHdsuxRA/Rs+H9U7lwX4DnUsXYxJb72rpGsJbFKBl8fl4Gr9b4xDeYc/LKKus9ZbNsCmg7sj
WKbT3dh6+KXotYEjywvDcY75zgdPjQrfHI2EcXJaZT8tP9ygDxAIcdA+Bj/JeH1f64Z7jl8Ja4vC
vMwZM90PM7S7hRpiO20wFvUnewpt5A4LwWbrTfi8XAiolx1SdvwY1v/1WQpS6CO558Ew+NhGvsa+
c1ZBuzmjQsDZvm6sfprSuboUYcUzaGB1NyxaW/i++EoJeAApx+zM2xRcldDv+UMYUaOnyEGNLCyo
vJDNVXhsgk+FMiVaTRX4IolSiGGRUD/rOFSD1tqL7Zqoe5db/L6sEhsRRCbnWfI6BpyiTdyCkBm0
9MGh5OqW6a1d5F8yNalRKR/HvjjZ7kEaXWyhJXRqgDuQwWghW/BA4YEfBx+BBM07i69B0EyZ2hCJ
Oq5ElbNL8zXD0Gnmw5MWLZSRc8x0KKESvWQVtzv2EY5FVdyqDIw5p5j8wicoAe7Q+iASMNMFRxdt
KiLth+LZS5QS2rqpR5kHxc+vjoTE7+SmN7ID/wGVO7mUq7dczON/cNjNl2pKD+70XjFCXtOjRg5p
zn8x3KoBvuLWOaJua0bE1Hpa6kZtfLvP0RHefYvEER6VKhmiLLoWpLNTPZ+6xh3PssbTo+P5SbkZ
RYXJPviUuQPaKGvcWUqzPDH8+vEKL11sn28bdxoYoTAWg1m6CYzgqZ6NORsaxExXRwd0QVugG1n/
eS/leYPLcpAnMLlhNVDtDLHTT4wBJWm5LEyC/dtcZlcYMWIa2/e8IcwBFg/o1q6H1dqpzZgxmTVS
edThAaSw1as7DwuoeS1aaxEC4wm/swn8KQI3xB7XBlmGzkClzgc43MuDrU4MxUzluM9FIPyxRzX/
W1TP91v2J27HC4FEXFprfAakykfT4Y7yQNiq3Uhi6/tXhJMpDg/ZWY6b/tuKG41IfMfthoQCynGr
YCw0Qy2rg8U/oril5cikuD7PmDj8oqJFbePV5XT5VJq0/LdPNXB3tQst5cYmRNCMCfxG9umQo6cR
MPGNLpdS5VsOC5rgIKgLo7MCBPva+Ma8bMZiCieBz7PAZNiSIRxcc54eXw9McRmp31pgeA+0p3E1
nVY/3avh6+AYytJiXCxSmZY6j2rnG+sFJB0dbLyNNyOIUL5SMIR+F3sOiJ5ZjOX/cmmlKlwINQDx
KHQh/k3ZoQSoGAEXwQQdgwB/zljsCB96A/4UI963Kk+T5hqp9Q1syn59VdAXdlDtrAMmnKqOemT8
vQvErR1AxlGoEaTbgxQiZhBwP2tbc/VBclRRV/GP952hI+iO0BPOiwl4LAZ9KdGN0M92Iohz0UpB
PjeSLXoC0bdDZrfaVVh4aaXwClDxX5CcH+wryM9PBaGjQnTtsUbyb6yBxmYuOyO6Rc9FNXB6MYmT
0WQiCqRWnBi9w6iwusLB7B7QZlXX0XwdnRO8z3u3tHtmTq4ysNMNGOZsQB0TtbYOwTlD4pvlhBHX
gm5zE55syT3DZ0jE4BUZ0sxbfMunnmPKtNBZKaTuYIld1SE+oLB2SFbEtdDyxXENFortAzN80V9V
UERLTMqB9O3xixBswTNip+5Q7Dj4ydGaMBfGglnobQ+E7rLk7AFmHCuJoZcl5fzGQos5j1yb/qHa
rHpRWRs2Ep+dgPEksSo5Qq/BPg6jZ2Sn3guD0i5GOzsDzYxJYCp25LS9B+DNdf/p2ACtOn294J3+
4+m8ntFjO7MUlO9ynieOs2WqCptC6ovORSzdRUdDa6Ihkes9ljylB+e0G342XCjI8k15OM2M9HBo
dd74q1gC6zyD6MjV4ZlCO/eKmIy8w987hKFAtBDa5exxEpohBM944/y+dR2szg1KxwHcjEtSWsOm
DiJ7DrwM8OhJ/b/38FJaQkNszYZE+shvWlwndmnea/HIhwcc3ipjQ+qwGmHu01ixsMFslcSFxFfG
oc14dornjNmkOr+6+YI1rX3ldLDdHYYmrwEqG+LkLp3jZdKpnzvha8/C1ufRFUau0lCkWyexjylu
FKfpjatPuYvOiozzJ8tAvk6CpYHjeI8DhwVuCyghpQTKB21ZfeDfB3bo/FmSMr70aJ3RAnfusWSO
1C46dkp8hE7UFmmCE1zFhXePwr1CbMgNaKbVD4pgvBq5vA0n4+W5ol67Yh2Um3EIkdfkYY9/gPo7
Tew6tKiApwZzOBF8aNW7/Qg61CgZzbu5XAsEf2mqxvHG25fH+48qehqiO2171LRtc4u6Z07pNxxo
hNKlz6/huacrVGs30VtxCxRhnaxBsfUSPwGpv7fQqP5mM3RSzVoJxzXx7G8Z3iF+y7Io3jjuPKKZ
rTWoJszXSXNjZAACShx2NYj7s3E5BYkt0RbAaJGqvE3LODMSCrqaFAeLKZCqmfczLGIhUYBoJtCs
k6HxNseevS3jmGzdofOWqcJBmzeHPGNjyyOCViVrzjiM8E8JfCM2kAp8rM7qJt7wL/yeyq+xDzJo
6Rp+PbepaF0ck2buKlafYde0pNRyfh6RaKPNZ5ZsdvkUrGNn2y3GOtFm5mFSi5zlLVvvHHMUcCey
5/KbO2RWFkljPKxyqMAJ+LM3lAlqwg7p/wB6RG/av2AgQhwfa0XquNHVIZdwHe/BCkqx56+Nx+uX
fofa/gW5A1nxA8Ms6Bck+Svp4/J9H9Arn1CyMO+RZMnzxwcHaojILOqPilbMFsvVsF2nROLAUTid
m+wyVI5AnDRm9cv5wEvTVifM2FxLILg/wWaoEvjcte5vvTmsiLDorvbVje1nyjeAgZDPAa7pSiuy
3tsNHGueq53OwPRcCatDuCYsc3u6Uo+pldkO1uEOnAvIjmDBlEQ6DJ3AlJ5k0xlxAFaGXbcsidiA
ld8aqPLuLVHs+GIvxLIVZcVVPznF8gy2dBWWCcAGk6HPwAWNjDQVw3jZI/n1A7IPUmi9bnmuCrqF
GHazeITf6Nsc+Dl51s4ClTncVMgzwUyqnK9Uiq1eoaUvJygG2zl6so3Rezv1Rx3CW5yD4z3G5Ci9
6/6P35aa5td84YSEhcehKtNAF/Atx9/8Kg2xc8kVJKmfuWt23Y0qPihhaeGLUuT/wzEByzy83+2p
x94ACR/s8f5t1Yl1B4XSgstos5qRI1BxDtIQ69IflHdDV/reJ7366JefzEoMy/cB4zb13Ku7xmKm
AvScQ0yh9DfWMWrFEQ46Xjms1LqK2qmIoBuDg9EsSZxN73GDNV++3eeejHxVAUMgnVQ0zwO/saRY
EwLdrhTwnrhl6QhRVmZroyOQAENx3dEmgNi8JXMdAXRVFkyKLrgrtk1SelJrtH15olUKhqMbCoAf
WaQEC5zddAmKIzab2fOh5MUsrK+cF18rtf2aRa0JEbjuhEcAbatlzGvaipT4ecn6bnEZAJG/qzBa
fUXqMhSIddz17czegKaby+/Vztze65YVM54uhQYsVfpo6Fg7CVkebdXdURMBgDGvtujstbqrt/mH
5t9Z//33wTHKkGW0n9skhAAuhJR41emLfDOYV0gjtcb/jeeHian3DsjdNiEmuBM/7r3/CgByttp2
zAw2+j+KPG8Dpw3fgfLrP6NR98qR6442gj9MIsEzzLfAirkRYcCysrWb42WP50Ka/BnMD705A+eS
x2auBma21xfCivbv2Qa/mTkeirgSHj9kdBV3jnqQTG/mB/WhzkSf8IlaKASFv9Bvz4I2BSKwd6p6
2unLcPuNAqN9wQR5z/o2Ul623RZqQ3iEgW/ieUr5z1lRjSqIAeEg5AMiGTgl5L5F+PaQtDDIee2H
MG39+LR/qXFGNi8W6tMFA+fzfcnZSjgH61JJSyhOPlEgQs2oM3BXxIi0HGa4W88Ak1Zi9L8nK0fW
D5JcRR8QMLlc+9juuTORfJPl1EjPhWGb885EExSFQegv57KLGp6JGn+tTRFwnSj840/DsaOaTbO2
J+/AExcjXHv5QjaORc80GAj22zCCeOTouRureSpF0orSOzTkzZLaba/y2kSYzw5ZlDAZR2nlHhgi
/O1I4BJjQwrQPiysmW/QSxCn5L1SmjrmVJ6SNRn7b98m5KAMroWFP+UrCYHUYK/mNlGo1Dwg60VC
R4kmkEXJiLqFikX1lxcoj1yn5clGKMkdzDRJ3v5cFhmaNPvs++aQ6WkG6XN/SszPaA74gOMZQd5E
ozPWDK6OetU9ks0DGCsgZ0x6dYtlY9NIa/+YOj0Hb474RP868IilxE8FAoK1HeRdeAZK9wLz2d0A
lpSFhMOh+MwyN1pQuG4Fr2wrVQV3eRhZ8n0gpBMp51pD92T7Uvpetxf5XYvT4dNKqPhA8YcsiCXG
i6j7bpmBnwjOfxDzzOLyNVdIKDxCmCusfwtrjMyFh/hQpOdVGfjUMftQJQJD6O6iJ8QO5AqugWFI
NwRQDKKe6xNsRLumMa9fV7cZXbWbGq5EPtujDXbziM/NUZiCI1DnuWi4MhKIyqSIcs8+uXc2HISk
fufmzXW/7TJwqGe2EPoPFIi742tQX+DjcAzolKg3AU4xi2h0GgwsAVJVbcDRIfy6bkaY0dplhHyj
FlvyYQXnFyoz+VVjBJGhRFRFjBYUYNLtiJ60FZeELCQ6yCjw0wWRqNv3K43dYa2uNvfwb8Nhu3sb
R71TZtadISlPTMa9LDCH0Fc3PdG1HNXvbsxM838VosAg1riil1/HOlK7OCfRfKRnDWrmm2R/vAJ/
JDHNJOeH+PfPJTpFbBbtohONo4/7o7Qmf2X95YeqkZFcAeBw6QaQZQXOP2AJ4lZruS50PvhbbOaA
QugMzbDtQFQb8qaJDHTx5uewFZiegXBEY23V44x8PNP5nlCfcB+hlS2s1zAJCfbD0aB6RWqxcqNF
ZraG1lWVWkBeVsLuULvMiR7qg2BEts/nVB3SXcc8DQKKV6TgqdMjpQbsxschU2nTdQWEWFIH+k7W
BkKuKTe8/cff1QyM4S0oaTgFZx2DNV2F0r4xqzoPrLXSZmcTRhUjHp+O7DQOwabvyi5EdjUOIQk0
kvS6luDccH3oFX1unbvjWCbmWguKAb7EtZ2OrXkiOxjJBsv52hCPDdhR5hJLFrSikJelYnD7IF/P
/8KyC8oizdiuwhfuEQ52v5YESiNKc6lTxI2jD1EF0p2RXaCUaP66sdWjS0r4Gey71nfwaH7HtIkr
p0vzL42Xx6esOePt39oS23w28QMXbG8hUSKhAWeLJ2ALoCP54iksNevdn+HOnHHdiNOWTWP1P6yB
aqc1JmWkpkpiN6RrEF+KMrHh/pPsI/vwqBQFmEwMgfecQuNsepuPEpFBkgiXEc/OUfrhduMLRIza
LYZMpOF+OGoKXVSfz1wqSR/JVtpGoRFaQl1C6RmyEEb1ij8DlpYUpC+m4MtZ8LdtLM5hCorc+wV8
26IIjJ2lXCT7JFgObb+i4CToaiZxfmDyVSrU7a/BYX/auGVAME3xRR7vwexUHEyJQ0o/bhDFkzsH
0lAIa+/1R/pJeKfRUVv3YIVdrWuh30BJZXJrj+WQw7iJ9pPbG0S3R0Y2A5TL0sZlJBHWdF2Adazs
Y7DoEtn+Hc0vleN9TROF6zFXeUgq3nlJY2ST0GTZMJvLZqPUmNrrnAkfSfyqjfbXjx+mF4WCgtRt
6h4JAWWpzOZHJt0LMof8cixY1qbP0U7AWd+OxR+raxoqc/XmGH39ifRRKz4hR2oswj2OJ0AFqDHE
exeP37D5u3HutwAmHdV4LJmCrZinJ1ji/kT2BM99v9RQ9Gu6tIWVfCWsSqHANd3+MgdWpQW7UR70
IuXgtaP0t+QGGLXxkwtjNEUZqERBJIi1GC2cqe8HHRGoHAyuyzHHAnUoo0/uTYIyqhkmOSJtP3U7
LWyzZcCZx6jaV+jn08c7olbTb6Bh0yarrU39PTIsOsl1X1wZ4p/ajbMxvJKpeMnpj1AU3BoNm83y
XxuR3ECGd5fVnrRq33cJstcu03/tScvDmybYV1e+zUz4ZXE78FUryANNSsmQ5wytLoxNTCC0C60Q
aargRCG3hzL/gENTY3vVysP0XlQH+YNr5cjMelxffpRVSgwPdZWb8sgyJln/HZgaR40+Lo4+yGzT
gbu67z6LvvJ0U7aJeXCpQ3eusS8uEq/xIt2lknAqrWoWu2Wl/917DATuRaNH7UPNIRAV99Wo+NVN
ixVTJb3uuYjSdam++T9ibs1EBZFIngxC0BNV9cd/qjSuzJWizSD1KWFBJo26dgkSh8M0sF1sBMbd
VyjoBO80/AvxtzlDErluGpKqyVZdVwcXe0vS301RmZVQCk5zbw4iHUmCfDM4yJoQ9UmElagCwtoW
JA6U9/V4KLUR0TvlHLW7jBUSEKuhwAE++VUSXxMx4cBA1MNx5I/vt0VPnRNOCYJdaPf6EfOgikrD
8DT0MAgzCN/HoZ4cNTMfv5azU9Lszor5ib4rDWExiB1vlbI/badIltGCLaor/Xqtp/pm5Oo3L4ns
jSsi0GNKMryel5boPY5Z6hR97+JJ3okFk0Xa6GxwXxZQqu8l1Jv73P+vUjxh8asmH/WQoCXXR8Xx
5vMK9q5/WqqIFVG36zsOIHin7xMSD8cZyUMdy0Hl1CrIBk6fDJC+32RZBnu0AWnBkkbP8bI6QbZd
Au+BaUNd2qOuchudOK2dILr+S8DOn8XYh2aNvYvxGQ4ro1D1Eg08mgX0WiKwqFjh/40hyO7//70y
Cm0QmUKQHiNrIBFo59lt0OyOBxZBUYetAsQoMxKMVdIIC/zWdTL+1vWfwGOgWLOOx6O7IDpiFbJS
1CIPv2pvajRgBk9vAg2nI6v/nlPMy4M3lKTmeZ8bzCdvRKH/2gbYSSZKMUBEHOGPelQA1oF2L8lX
iLsEeV+1atRCAHpyRjWuiiguzFc9MoaLuyFir4EZePUjNCdMxVZAgSaTGiaDQNpiScdRvfcvcaHo
auqp2cWTyOMZ+EdK2Csd1O3BRVhHGSnCzTxOXeNcB70Lk2H2VP09XhnE9zBVZ5B9njDm7sRI3uyR
kbyN8w7HdCeDocjzcbwE4lGTUHaYALNsCj2iW/rpa4290nkdHEzw+4neahjGRkFEJLiVkJ/LUmXg
5P6iLROGPTRG6GsuC6Z1In3Gc6ulhI7TCahkriWXTmiLWQg8mf8YWO/faf9T+DtowH75derhZDSk
8DAf3pLVsgV42vSGA7VthnQwphW3YAiHQv6hQuYBaRbnXL8rtGIXLxSi77CfIQSRddnX8B85+YZz
t78t26UwxrNNkcI2AoAiB6yTWYJ34uQGBoEeL5ghnp/+AUrq+wf3HV9Awl4xGeMB77gFwrvZug/i
PZI761qsQIDM8QZolzR22kAsveZuzuWSovOlOxWCqsuzpW6JO7Uu608Wf2bXV6zlHfDuvtUksqs9
P7Hlco/5kEn+dGLtlkjkv9lrTncFizC7JJST3fUDJir+AK+vMHkQ9Z5BWtF8nyAwtcqLnEok+QNj
X6DZ77XAJmOo0fD8uT5WFgGImvUQQ6lKlKCThvFaCvkctHlhNam9Hdt/6gQ1k7EK2riSt45QLyQz
tkDYCHZA5BuuMKsuqFyBfRVl9Y0L0IVz3yJ6nQ7+hvWu5DvyVcznFtxV5DbLmyvQ+zNiNQRGFIT0
QlfdL4guUj5kfcD2poluOf8JoXRlqf+VP9Ud9e/ED+eAxhz1BsQpotWq9pSD6Rf4338Pd5I6VXZT
lgPIk8dLrPyC9jOWxYHeqhm2V9O9aJSbcOnmzTCGq1/d0cnwVRGBWpBXl9vVSX01SGR/j9+oKfrS
eVKaVoP9fAZSeDB71AH5yV6/Te8Eev+MtqBfqDoyloo+XMrd/HhFiYrUXJRPUEO+p8F89TDW6iN+
R4+fnpNiMOGOSQFEWTYQI8SANAcY6Mkv9R3xdwJ/7whCPNNmcWHEWrKR/75FsgyMtX92JAElvGMw
gsJ4RgCINF2Lo0s2tl7TuunjcxLrWf2w5FyySzo3GgApFM7utSw/9uJBcTBW4Ssemv0+veNxiBMt
Ac0OkF2qpNojG7kiq3aZOuJrIjTxajcLR9tDG5qKoNjSU9R6eX8fdoWjsmKDg7MAoMVryJlQHldS
0amEUjxclWd66l8y2ot4Y6NJP0WSlCJsmOuOdS4ktZQHNCPjxOUjnnh6tsoy1thcIp6zM9pz6Iim
na9IWbFe+UTjdi6Z/0ZsJGNTcYUZ/aEgvzMu7o3QzTVxX6Cm10UyDAm58OVJsvgqIqNqiIOvubFH
jwv28aXTMd75G4YKSDr4wTIrIRPLp3cBZYWKxXg5grTQFDVGepfptcwyEehU974z6dEsJENMmOeN
TrTzJvHvxO5m2C5JIueeJDBHk8WN0lp5/4+pwi0n8MfaxsfoFwd3HX15sAtLI25f9cpx+1ct2zx7
uxmWmkelJRqGrVwMsRf38k9NaWSIQURJn3mrpYxOwAemtU0Irn7qBdOOR9yTaHtMDRO0+BAMn4Ss
RmGdKYMrXs7ecbya6Gr5aPkOtgCW8wm/DVv+yotZ5/cMXMvRgEmwYgC7gTYLhVokby72T8uIPEbt
ROHmTEIeAF5ZhgJUPiqSbwNSCvZ9HavY9ZGHDKRUXHGg0AcmIKTnP8lzZTS4JVMZGmFJFi4Yzwf2
drK1cLUJFgunVcjE7jHkLiX+9v2TMf5xM2wBDGSXqmhQSnhC+YGTKPoavgJwweH1Zh2bacNufoh2
xXvcKfwFx//MusC/BHkrljmxMuoVpnGQRuSipP2O7cM/l4gQH8wy078q+zpEhggkRlDVI5YEPdC5
/sfvyrKz/RSc00LMik/978fiv1V7JgaSCauVyfyCZEJ6wdD9fghFvk+BPmtqLH06NxuSLuk1goKU
3avsACg1aQ6Fg9pv0sKWsEGxEthlEi9eQwPDWChKL6BWthqpgMTtKYMPuybdmbNO5YRPpAOSc8qA
LuPdvtXQf+G/aFaZqZMEtsNRJZS49Dr0QtB3AulKkrDSHtzOqM4vWuNBu4H8E7l49+k/e04Ca85f
bmywzBUxSg678KRnxrYtu49ClKBZwSExMO5x5XlvJqQg9oSsgBItj7VLA6IH86hM7dAaQt9nLMXz
T6A41Tt1FjWb5ydAXYco1yMfQaE/21Ih1Jz4F1jY0WAdXlJvuJA/Uh0JEJqmAad/7yBFHGock4Z0
kIS3YsAf4PVj8ynsHYQ9ebZDrVGp6taLLt7jbIBLI+DGDbNRZ+GwEubaMP6WLwQf3IB4QGqT7Yg9
6asAuTXpQc5q9bmtvWKLOkXdsAmAHfNEjVtUAsnm8WilabTsfNarrt6ZUDtIUNGPGSC0OGXptU7U
X6QwZgqYB2nru7Yhml+TUd9HmRa8QP9/8yvIRICVDH0oKsWjgxOvx5WzLY7DHCro4j6yqB7Q4nbN
YWKF2BfEEK27mwb36sm9PPcBdPyq909Kom/WXySt652vOWyKYhRt39xpy45+1n7htRAtaENG27Ou
rGU1X7gwjJ6Iz6shIuc9l2a7IrWwWFgsINZ7DTenJhKu+eozZkDTrefl8wYu8dKIpJ1r8Hn7gSUV
qStDoLZIT7oeMddv+0W1ibDpF3NummqfTsFUqVw2OJflPhRAa+2I5e3n2z2ONK9zUV7zecxmcMm1
NItv4Tigg1XKwUaQmM4VxjXXOA1NfmD4k9AXU2kkYunTHdN/saltz9NU09PbA9Z9IwkUwyNnqWjR
P8PLyjqN5OvMcN7ew66004CB8dolf/w76oV0fXOANuHBZcBL7Kb5ruAge3I8hfF9wFydDIeidGEp
vOEunKFDbzTzMz2anFaDXE0jgUVwLsaQMp/bz7r+LtaBMV8fqO4ORvWiigQTp8AQ+K6hMOok3iyP
mUgnfOA6BQa3kEct/mE70r5VjC2V194Sv/TBvpOo+/ztiYLy2qrgW8NZpeIsdA4JTZlAHny5Egzh
Jf9qTm7GlC/tR8i01qiXYwLUBwWZ2uxAJPeWrC1E6UCBvg/iHXdXh6c4V+vyTcrL2xQ3E6wtCec5
4nWz/3M9gJ307/l2bfVnCXvrZpPRXWhCv4+V3LZxLeNbCUz1fC+XcS5W/D+Ql0n9MaKOCSMS58vO
wlgm2NqSwjIyMXR6NOd/+/audTUHSCJdBinrhda0K2V62R3Oh4juTgRozMCaGyfUYBKRhzoDyhxI
jFopCtMw0viYK4kh8j6ZejkqOCjUKC+SCXdn4mpoLEsTfJxPKGciNhusDTwM0lsJKEXp9go1Gq9d
SKDyy/t1R9LIaXerJ7WscRslGBg/9W/kUWwh/dLJqaR+hSYb5FY6Kwj8bjTHO6/ZUNIcxFuXC+wg
rl7T3BjquFjc3ku6v8yWo6lVlxntbrkv8e9t1lhCnXq6MJjy8Eh9H4PzEl1pyUFEZK30wQ/5jNd9
P7j8X9bpMkdiKiCVjKc4Ons+XBAm6sHF1dpK1X8OGgg/Hgy0ypwtLF83/ov+beRv0jBItn/ldX6m
vV8nZOnykMTb2WKsp3cZxM+YDZNExXQVksHwReiakF7rqEVV2fMa7ggQIxYS8CAT/DAmtUaBtGpH
K7vjJZK+qNYrIHt2PgM+s0jHLNIEY2/NuuaKCYPa/ZRj3pYYVrMgCtKc7A292FeuD/7xPzPN4R3m
3pBcfDZFKfRP9S3oofbhalYlgdaADX6G3+dh8xtt37VXdZ/FvG64vg0cEmqsa0kjTBP18SlKykOr
c50zaT1uVZijPp1nESFz11sX7a9nDa/0Oxi3YWh1o6H04QH+jcvl+KY+8YG0aW65fGWPWX7o6OYs
UhslkDD5jDiA9nTjssR0avXYSMdd02zEmQK4tuBpTODD+O8j+aUqUr2xmZ0uYgAYe9VxXRiJXvks
Tebt7KeeRsKaPOsf0YfoosiVhS9ig0ufST/FxFLLFhFL1vqa1sEr5nGvaBAy/IfFR338G04iNmGo
isX8fhwlt8WjqRS3eFkmnGrztABfPUXSnMEqdNwJW2tAg7nmfsSzH4LOdiC0IyPOPryv7TIqr3bU
r7fpj6RxYSHtvBkPOVGKjZ2wLM8qq+P5wWqUIFaMb2pLY7OxTKVAwDT9OCxARemefYJj6Uky5+kO
4jXc0rE4oqPxXUS0cBHwFW9N1TztAXlkl5Hc6biOutyvvP/DiEEm5ApzPgT2ZHTxDUW5xBU3cgnH
I8AF2rCAWsLeP/EFFTWWzOnZBqUD8JW/JuQX+GA65eBgMan1zUgIsJ020zM1+bNkX88fTVaGDQSj
YdCaeQcD31JeszE1zQ80TJ7ajFASrxnMskGXuvJiT00jk3t697y+jJiNXS4/InMh2r11iJj00U+2
LN9T0F2REsgVu6m4AUHR56L2FeuIONo893v4jeLdbBxc9619HMyALPBKPhY3Dy5/1k2g+AlQJaSf
mS1JwE+tXV7BFn56zsOaQ3ihCIurO16GP0xZvGO/cnlZ60jRZb/jsPUom0lAdmqbISglc+pL/4Xz
XjmgQH8cq4imX94IV9uGCSjFw438A7WqYMJ3j4PHeoXNfA59Ls6/idK7MSy1WxW6LbRFDpRQg9E0
j9jUv4YAejcgoZ6bYtRb2TZ/uZWbHmJWsZNBa/BsqlMzsrkhbDf3rqITvNwgsTWhwP6FlVtOqGy9
YS2vZ3iawxjZ4Fo/e9iIfaV9/F9e/VJdmtuUIVVRKG+ldy3Dpe84QpeGLyqL4lbRm01XZsiYwukH
zv7vVr7ZFBNndz/biY7u6fX8oMcsrSjw69NmdTqtMSgpbmBPViYnqp2iaug6OBKCB8LI8871eMYC
bzqP+V5z6IgcCF9f5GtwS73uXrDfQ9ErBPAyYj2f+gP/Qn7ghGYlYTUQrPMK+W4z77ohjUgssnIx
yEuIce2C2XlYlaB98NwQPJmPlCf9+DMl10PEbM/lAHs2D50oIp4EGMKrCxCeuvSafzO7gUs4YK/c
PxxRTYD67gUvc7wC2KtdxDRGh5VhKCIeEezZy0nALX7hCM+jIHUrPC/L9ZE4D+jpRyfUheKCRfMB
7+l6KpGhMFu/1EaseOFqaoda7WquAUO1ZZ65dGewbyv8YsHFCNWU/EqNHvnDAOkzckRtPYhpHMa1
r4kaK3EiVufOQHAcxtgZQXz09MwPo5l0bBJPLbtqGEYzAukgMFaGqxkuZDK48376awZxoqqk3CWV
rnjomFGQH3rOqbYswDitWSGAQO/CWJrLbHNGsAwEDDt/E3BZBzD1s+BMz5xPe+8/xheaZ33tT9lN
Wo3l/3ul529YibuHVc9JKYv4RaWceSyvqRpZ2r5XyHvMuTVhYFAZ//uKPlu/XO81dmPcydv9DoNO
r7iOwWZR4caVtA6f9P86MxKielRexEkOFqOfTmLWcvb0ndOk/1rQCHBkYWZ/M9fd0RxurHIegh5+
ThkRl9m/KimznM6DHA6+uKR8k58HKlPn1oIFz4TtHtsYl8dqMQ6uG8rPhVYxGCHYFA0pU44b7hUo
xTCLXBWiyL+USrpCF7iNAUNuTAo8K4tG/c/enIR4rdBvgg+8PWj98ola2ASCYMQo1su4+LeVHckR
sed5MHxWoqBCWiKjTDZtiHIMvC4LCkIlIi4ya7Sf1bO7lbVk2hmXTrKmJnnI4kX94bwGkTKYpcdo
tuDme0UTm97KuWrTDapX/3khi6bIw2Z0VwIMXsdC9QWNl10DeU1DDD2SydmoqIxhoJFoajWOaQ2s
yce/jllSuDIHZhcGqqF5yiMPts8q11G+kbg+g6XfZnGU/wCrvW7BuJOkiO84bH7jyx6WS8bXx5GG
E2NnxxyU6etrRquZ8XTEsKSCGZsd+lxxiq/goSm59YILLYpyAHS3elJj+INGLhKTwPXP/YnnYDTb
JVs2ww6kjMl+PUmvJLR5yVH5lynuQ3h7S1sqkN/CIZS5IRjawnN6OHHddBRTjtB8F0lcbn+cYnNS
tfuT59I0zY3u5lxhtKjAem4QpDMjlBsfhJwfL38y2tU/1NFQrGWUbyyFtB90BHe3osquCnHOU39F
DXKyH+deQZV7BARYXzsSYswA1TYHvh8qYv1v1eUzbpbmtKWPI+EmFInYmugsE7NTfH6HdMcHw0kG
V1DPMjVSBUKLDKwxiagvEoMi30HZ5DZh8ozG6BiFi3cEmDlhi+7x+WWb5lkRih77sBBJA0i9WrLl
+XXpXk6bxocpUQtpsbsXhY5RWAEuGVdzujRhkBg8lTa1/7UAdJf+DtFAr6Rio3RBZh+3GeBjRz+x
VUCjNX0Tbx+64dKoGQ/RShG0Mux+DqVZBdx6ql9LQlwhfZF3LxK8h3InuZdqc5Hcj6x7DJ0NJ3QL
yK2J7cAnsONCdYQXal7yrFtzKA2ElxhPtXKYvp9spWwuKnHnOFEG3CsXas4+EUFYOT8AGl4JNF4U
lIoqQz1GtD86z5pdzLuVG/SiKD8SgCGTN00OKhweFCwzAQOR0Rvb3zAE+1EIYxBd183xqXNhHQ/O
7FgQPUqDUFaaVbGbpjZHPNo4k1EoY2QhjCQ9FdbjuMEKEhF9zKwUZEUPARjlhAJPohGAcp0BdCt4
lVv+6om3JpnNXztMoIRO18JZFzahdIGlWyB2E/2KkcMK+qC+go0JCb+3pcTmvQXq2kLpipACVl92
4mN62r0vFqzRO7mdAvqJXl9I7N5Y9HcMiAOfn30vKnVSQx2ZYYvweIP3PipYL8h59VlUeaFRtk9p
CJBlRuLm84ciD9TauS+xP7jARdz0KRaoQZ5zacJG6Xm+kinNrFuDtYxXYIrsH+2vA65fhH7am2SM
p4P7gnx39UhSRpiSym8yW5VFrauLD8N9/TpOrnToy0KS4UjmaNUjF85q11sluryi4jmQNO21cyR3
28jX1EqCbIWsgUkngy/dZUZpT7ERF1lNa+yvOT1YlU+HgxvGF1qQp5PveP9YwGtYKQq/Ingzdecg
DrVueIV5h3ui/ss91W39TzXUoe40CePF7Rax7SN3ktxvCZvB2hChuleUhuGGlCCSsjLLEi6C+gD6
JGlaeM3sOAyWcxv0qL33/dLjs3tFYUh4AzH8CvKm00Kv+ns4zDKx1+p2eNNVYY1YvnAvL4LC4sYU
4KuftoZWTLE7GqSpCXKa61jFEA1Bacbzu3nmNDKaw0r5FZLLc5+y1aq3Pgvxf62viPVvurJxS78X
/2ROjUo9MgkgOr/EFtYTyiRJCua05rzSNIZePO1LWWp6djBEI5qdYiJXBBArfr5ixizClWbk66cx
0/f3x63shMmZEzzxqbrs3lp+ymf6eWx7Da+6txtfKtLyqUlzJmGb7nEQ8xbfrRmWKD2sXCcnkc50
KscwBPhpApVIWvQVx5n8bxBojAdyXVeSnc1G6VPMss0462VDzUToyJjpcSsun7nscTYtWadAN2D2
tHtqyZej8FKSnDuBso3o8k5/cVVXD3h7dPUdKqn4Zd0S8zpCSiJ3AJkbauDmKzXQEXzQWAuK+8YS
Cz+o3o3hS4nOgtebGyn8eDbGEr53qyOmaq9PzGn9wjjTnPYF/S7XRTMuueyOw2f/cUPYLfxvXUty
BpsFQk99KRRQYAvmiVPiV7SyaFGuVGBCPAjoUtX6ZYc5C5blsIfgMAz0nVt8WY8hnpI4U5Vgb3cm
Vb4pYMTFz8pgoxTJrBpc6ErkpEH6HW+2jubV9TAA12PCdX4vx1YGj23w19XCjRkTBv7+4NHBEQ12
Zt2EyuHrG3oLeV7quRm6M8y2nw49P+NMXjwl5MW77/TEU03wFhP0sJvxgvTsL7cfSFPeZxkxhtY9
uXecJfy9UPTfqa5Ou00v6yQ15AYdlb5nY0hexUK1SEqTaiL8QeIRN8NCakNIqdQVBc3nM0kVuC4g
bjfedCQv5Ez898gpimhc53MOu+6trb9AD9RZ1eEeN+6iwrReY6y2nxcDMyq7Z6wRQiRdYfVibmkv
OxEj0o3T0fs9Lgtxj45fBinEy9nJ4QzcyyFaHLlMnV0MMGTERu9RfrFFan6xc3T0oVXXTX0/9Vg3
0Pyx9g3M6dalItuSPrbUqtUwUxPC/6zU3S1PUeQloKo2Q5/M5Z07r24NEgL2nGG5KHE5ZSWY8OSG
sZtawU5gQBGTdDT7zlaY76NNjegaNVjYzn+eaf3VEWif9y6HrnbibvbRhDjG+jUpeNXqcfEmue1e
6vIUhtn/kNxM4tRQNNo0l0bHkokBx70tF3tsi28zw3Di00vFKpNMI2nGc0QW6CC7EfNiW2weOryW
gyoVzTb1rOWbgT49Ef8MOY9Om1Rypr50/vGAOFRV1lbTc4abrmtfHDK4tFY+h3COxFbGOQuAWrxK
IWqt3eS/m+g2GY8X3bM07bMPm4TOcCYz//IDmUH/W+G+4sXpkmUpwGsRwl8dofln7TlCvt7+74h2
4FqcWqs01XfsgyaegIyl5D03SAm8J4BMuM5M/Q4U3VjGNnEs9gQBSNs+jECqcPcZDac/918AGvQQ
GgNa3dAStILR673vCgWgujPoxxvXyNlS16ZrIubPns6SNPflIr5sis08YNcN2kJDkD/0R8672FVg
nG9cZIkJ4zcGBBtEbW6dwSgNR/T8KgxTZZftgrVZT4hpLy9taITu9DzziUFAO8O4tOaATH0WAeOJ
gJfLOVb+gZkDGQsvqz3y02aRxSCw5aRLkQb+PEH0uPXfa3eWEE/Zzx2KKitoolpIwAaypdFHn0lU
viDWYkMpPyOxYDtDA5pK1p5uws2RlKHRe/r62Av5UMETsSJ64Isp81a28sc+YQLfwXFDa9hkiCas
XHkLDEr4nU1GJMzu2+YFBuGJvBJPgBdzzibF2fnL0GzMyudDPQgaYCj6ghSNB0JdYPjkkubIcvbS
hXRsQU5OesNTHQr+/x1kp1Ub3bnvodFxhUYuGJGOI5drMG2kDMHzd/tNnxzu3LM10z/CnIPCwk0w
R+E0tuUs7XuGqxEF//z/VUCSGBXtaCx5hEkAnqXKr1s+MV2SMycG8w5+Y+No3MdriCYDhcs1z1+0
Uk5TIM1GOs7FKK/kkCZlWxT9ZV9LoDagSZ4W1nSzjXHfVf2YkJDJxd6FATI7cshyrpsNF117TCM+
p7HMLs6AD1iR1ABNih+dDoQlIR9cLrA2eHOuBj4PNbi5lXUMiW+Y4dMpix2wYdSpsZIxXLDfO/9C
u9RbyJG0lrYkzXppmVIvn+xUPQR3pmVSr9QxQ8miBNwgVe6+SE3h7HuzPI/CdLcjl6B5Fd/IBZ1e
8kpbOlHbqW9gZL9ISdYna+pIDK+LrS06V9IPiyKnrwZFd3uq0P36gmMlsZLNd8WRLkYeuz/9ZMT9
YUeyuEpVYgq+MFqr24gMEjn2pwMdno26e+UUsuOd6b5fEDDQObo2OM0csA6ZpA/tKNmSJcZAp51r
kCvQGa49ExUu9LcleOC9uw8ORgven7kCKGOwW22wveQEde6cH1i85Md1+hlIgBCJVXsxDgI7NOld
4Gfhu9mmJYfC2ESMs91wucPWkDms+JFqJTgMyxk0n57n6Ihl/4QS4uoSNhFASyjC+ko7dalD8mfl
FctDmNuksXhipA4YhD1+uzTr1kls4vsmT9+b3F8CD9JNIF8zEnqhPVmddpJ2P8SbBqs23YpbfQuh
6RoTGXo/pJPhh4JVU8XW99AmJ8WtEESqDQcqnUzcXdfTCbPDjlFOAvoQcuKoYkOEBuQ1h5z7qXxs
YxEAIuv2u88ne0X0+oJnEd9EwsBsU97jpRlw/M+XSsSiOTRc5+pAvjToC+ZLaF34WeBa2lYVluYj
refIKVHfhknIaIV4GrN00KkDpUYECyLqMMLGMaxVUwRTr66S9axqWY6Zo9xyAg7xEp4PrI8UV7U8
yAigEcDesvRgafvfR93jL6Qhbfs0+aYcugbs4Tj5JmRVZssJL9KVzUvuYPY3ZPOj0MQquhUIIa8u
PJPg8T/00x+OwJBmCIGk39RxL8IXmkkvqWJcAecXkRCU1niNgiQ5lCDbkuUmGGjZSwCcjZqY4jSD
B2vsg8lN/aJQf2VmsrM0SxUXyVAumbBjltlqzvFPE9aww0f6guPfI3y8C2TpuIL6y8eq2I3PvmO3
/i8zuU1zoZjjkGHWvDFbvuPLBnzf0p/sXAp6c9rj+KXy04CG7IXOf1bEexxKAVNpWM5tJeHVNd8c
FghrfhlEl8w++PoDeETdZMI3UhcyOSapKjIzV5HiMapOrGR+y2UVIRZZkDqif+pHnGlViyhqYpSP
7DUWJPcWfHVMvox88RFMEsgdqVP6Xi4oimZxcV+z/pJAEdvVDp4/jJtLMuOWd/FVMP/HEFyB3VbW
kGL+0fxlvbToKuICepRQvcYJ0TxB+7Nx7auJyqAuYBjIRRwmA981yXtjloenB6oGC6QYLQxIX/qL
1f/dX8mjFTf85RQ/xBZko55oUN28+Y0SC/3hvUub052yKumkbEWee58sKyHjSUvx8V+JXaZU0PXb
ScRRdyH6ncJI4SToSF8iF+FvjjTLXktHNjvYltJpBMkqbbFPlEexWvcKE2pyRKF5klq1w7V1XDy0
H2GATeq+jN04MaF5Li75RA/CzVZGA2oFmBe8z9tHkmLNaygcS/s4dUT1g6dbnv9e50svz569jKUz
+44k5Yq4zDAoBMEKcAqsHip2vtMUUvIh51BbJPZlIF1IjuqJpMVeNzfRhRx+KiYskyqOhtuD6NZU
O3KZcUYEgWyusoYDNHYUSJo5adeDyCQ7AY314UfTKuv1gFwULu+Qr4MM/5Sfgh83xxbfjzIqcaQg
EfCSsGTEQhO4Ubah2pamByUF4vgjtusuFhjBv8c0dgFOIk4Lyldhw5H6sgWZk9XbQM00p3RVERve
pK8ZyMM5L/+jGysZLJgLQhs6fxYDCanS9iF1oumWCd4yZGZutefeOe7DOwYwkDd3MFdjQVMf5aVp
ZCMcIe9HzwpxGOESxM8Vn37yyHtopIWRuihWRsQV+kDSvyyCLHhvL2ZAn6zIwyYhuAyCSxoY0Lpm
Auc4rkr/O79Sfhr4q0vomthXqqQ7nUC7CUYovs7dvVV9pj0dlM+56jbBuDqsIXigOynLgE1DlocJ
pLovtumziKR2YRaKVRS7CQCIvCaCCz9AADiTEnN5S+TbZW2mtkUengZGTaKLI2EF2x2QXuC3JcgP
xJ/NI1OeA9B+hIVgj9kJHMvVS707mCrEuLhFx1M5bXn8kWSJcQwuhBz8C2Rm9eYwOBsCcfg6GhM1
iwvxVW4xn6ZbxuLeYzp+WiqUQVpQ2TSTm4WqNBks+I0cTjoQdiIZG8wqDO34LRhoz5QZVF199/yT
wH/NHETCLWhPku2xoHGs/DGK41EKHjQ7VVaZ0AmW+B0X/5N3FYTkBmllGjXuqGV2MVb1lccgXw9R
hvVjLA0MDxv4aU/Mcil/zVXw/k1DFW6m2hmV4lSDnoxOeWiobvSTVv4Vvyq+fAEzqjUQQfAwReGt
YUrwtAFEKDM7La9t3ptfqITGMAXXhvGdx+m1pLZJuJSUAtBpJQxo4Q1K7DJXBWwaES2NFQMBBbdK
4x8VrwMJCo+Ptg5MSQx6Oa2Mvdduwt5JiDqysBu7f/t3Z2lsXDYDcV6HiEc9BGKMGczWqtyU3hwc
ZcGVBwhAt85PofEOOoE7KezAfB40zdx0SkUHJPXTNekZfmLFqfSDvZ8ntVugtbuntFnAoTu1qKFY
uMjzx0SYiTHdaWz8m0+T2AW1Ox+7NMdi8cTqdJ5+CHCGhnjmHBy/4DYQ+TcdaK2vFMdOCBjWp3eW
6aCygYIBwZ+ykULSh5XBtjeHQZH79QTpfYRGrwNO6Ag9Ayj5BUtDwpV/I3sWzt+yIHB16kF0OGrf
er/POteSugpwSSDZJ1APgyvr+n3sT610sPwns3Pn6PyGCj0w1zWwtmcyZrrT2rJP6aqTNG4rbyja
lmNqE65RD4NxeDtQAE4HhJozZIAEkRgGXU1CoMnOjiZUickMVr/h6TS4sDLzKDg3zQgZXem19q/B
dzkihHLnY/0RqRdeQY1rDM+GiAyTyfF/QDHdDvgT6g5haoMAyklCoKAUIE4fPs2Y8D7ndakWlrx2
tSARNDEyiy+IvvQZYEYHd0zf/QpxkgMvnMqaTCiuoHke06Kbus4koq2ANmTI0M2nGAkLLMUrdRJh
OXFt5Fh8iCdUTYiZ8CDO77R59PVKMHaCSOQ1Q+MRe8bmOpDMts9IeoxN4Otx0M37cQPh2ZG3nbph
O8dL1qRf8KWuBogbSU2/Hmi3KpqBdv6T9ZqSjhM4Njiuc4CUmR3UWLlGb/gbASAzwe+ohs3BXZ1F
TEPkrLU+x7yiChWXjn3T+7NgpzzdBMxhk7tS6vlrqbW4PsXoseE+PtTsZOxhHwRvzNSv6QRJlv7u
QU7PQkybHWcJAxXyDR03vVs3lyh0pkQ8/ABou2EOlKv5ZEUlKEMslPl3urgOl4NZ3W8CIj3w7eow
CpoRsIkLIQEifFyGX96gUOMqFOAt0OU18LQYQFoj9fajtjlax3RwSJEjOd5S/ABDVNCUqNUiwVzN
vsO2n5ZUPaTJiQekk194F+y9QRnRtIAVKxim5Km+FiXp0V1WKOz6GKqyMBmuY4pREpeOEL1zYDdU
Xb/NiMNhOigiFXGTahpt//LXkimXAO01ROobs3GivAGOYfLA152kR85yHq+73WRhFQSZYSu1zw4F
ZxZA5DYRsIXfZSKepxBlL6fNQWP+/fzA7Kbr/yfRH83FG99v+WN7NQfr3lgYNGl8pLIB9j7Ir85u
JzTppQXWs82aATIoOKP8eeu6hHQ7P+T8RVkmYssxF4JXEqFjlfKM9Kx4IM79YHtt59u1S9kphtSY
NDjxdQC7uCLHLEWVWuwX0BNYfT9ky+uV0CKt4jj9aND5ch92kM+u4/gU3QIvLK7FXUIQsh9hnXXw
I7pdA42UYfHOXo7AsBRKY5X/t9qOnV4+HirOairuFIzpQNIpG0bJBB+GbW/BN+73T2OjT7jik61g
s0lYtbGTqygOKgcLOtCimS5RlSxO7SInQqEyhkIUcDXUEUCUUUoemAqcyo3XBubOifxyhJeq+lvK
wA4RPzvkXzWEQ968LQm1mpGew/b5dqlIns7A9AuCX1kuFfO0MllEX0orFzxYI0wmQjhfWmW21qea
lhks1dtjASgnkZZ4LTBt/pyBz2+QxRc/SZA3XKpDWaxYN9NWEHD4f+dtwyzldwmSs6jqqRwhRFi9
kvzO9/q0qzr/XIXbJ3dKi3LKsdAHD2E63vCGijy+mTnIoGnT067V/VERl3NE6iPT31S7QqrDWnro
684E+cPer1ALg+NDbI+EMTe+okcG8T82eZqYHrVujeBHVTM+1TRerhvsdwZKYghpOvC/5yh74s/Q
za2JgzMwGbTzm+6ddJ6BJpAnp0hFJgPUD69xs6KnSs3libNNmVY8v04529kEpiZD7l6tXpcc6aGQ
WS2MEtcUQ97NkW4U/EKdyCcG36ZHvj11fqc4l/vDz+YB+uChT7sZ8gfKhojdfOjZnvNzspiLiXpy
4jNeV7H249QBl/f8LX4n9whY6CeZr2rWjPd3eWoIIlvftpyCbaEj/vYspK/ZPgUcQlsUL9IMszSw
voEBsvpykpgRGTopnz+XPqNNIpEG/o/qNPBrx52awNUq0bmdZP88QxFFYGAPE+NcwqjcGd1tZFZG
Y1hGNHn0kQ/JpdPFguFMXNDAgTArpWrk7lcZxP1AMJkltX9jN7U7hiI5GF6Rtg6NYz8spgzLVOGa
WNCRVkRimtOyCUDAaARHQLkoS5ypUgvPyCe2i9vbN9gRCPq/s7liZq9y7qLtOJTJMTSfNDbpEsGj
YuMtjvs++6AyKPERbZMtgEAibF+3ZcEQc0zBXI0StBrjZQBkZx1MbRKciOU9qfAiCxLEK5EHdGDW
VBtfFBSfIegxNK/K9TcbTi/Yum6nXCz9BYSSOPw1xdCh8z4NyUcppzsDogeJDQ8hlsPqXDUQlAi8
rgeqGsKL6cCm52vrVFb0Sq2PNSQANVh9VshXa0plpQ32C5vue24iYZVq86t18CepKs67kUfK3Z1T
6a27XhVMNoRsKyKvmJ2rg1ib/YsFgV2r/OFGu3dTVUMciCH0TZDyGD4xs3gqM/0fAxKDLOsSgTb2
GMCku0uu4btfYTucSbWib4T/lniA2pTg5dOcdjzbsStg0iTQBL0G2x/89IxheLbNCZeYXJvRkG+K
3kiMMTVE9Xds+dZ3bKH+zJUQn1qPIgOsssqFiS5ip+Vs3m1P+xTnmitFevZYJEE3Ab5RcirPibMu
JC5cz4qX2yZI3W7N9doFWSQAW9AxFzv+QLqY18ogBAH8IcB6+Io1onzAPpnyp3ZSHx+rffj0Y80F
74aPyYZnQCOJDXsFiKcdE7d2p1yaMSPUpU6KxUtwzJBcGq8RJ96qgwIPwsUJ4z/haIdii6FUcy+P
isI+6MVjoGUAi0FBvm4ykJtkS0UfWM1+DXWTuiSeGnPV4JyuIXvvBfs6zLFRlYiYH/MdvZdYU6Ef
IX1AMpiPpmT6AG8IpYCE+dovaUOdYr/Mm00DMpHRo2dyeUvupua8N+76xsOGWSmPdKjC4HIgnkbo
NhmODcFxBKjgv55Grk26JZH1995KCD+lPylnZ/hraR443ejnlES8+KTy+ylO4OVtXumJSFlkL8Rz
cYkAoD0HWzLbFPExQhZ1BxoF8syCWr2v6I9huENHxqD//Ur3vVQ6bgeQsbEQRbqNbic3a2CWx99T
LM9UPdJcQQC8K+3oJPGngjOZzhsa+lJV5ULRgX1+OsPUEnTvwjYc935pI8+HQa77JECv+7hp4/Y9
ZykAswC4idHxWpAObQO0p9cuocGY0PAf/G3mCgMpzjcY9sEWDH53G42PGTVk/HpKTU7hpXootwHe
sa752r7jQWElZpLVe1xy7L1bMg+xx/0RTkFVZbVuo7p8W5rtdA6DGS0OXg3ccYm8XmzDgVPX7T1W
828CSGYHIfAREO/hv6wD0gh2ebRwzi7vQQYIKxUudAnFJ0tR42qf8oQqSVFUzAaxgFx7MYBkIgK0
aheAkVysxYn0DvtkiuSZf4pu0OiDGrrkPCV2lsty6904fz4Z/IJ/t5GormK97Cd2Fvw2Y++S4Fnm
wbKwcA7MuPCy98AHVR5Nv8HtFR8WR8T6lM+F9K5Lm8masrjnqLzxCOexjrxhIoFafL8HQxfM9AFt
JoxwIz4NN+aQGTvHRpVoDo4QSdDmLGigkHupQK7Q3OVTQpmHc2pfzAgDDBUCw6Vvd/SE16tkuQ8W
Pb3us41/TuhrUAJBuPL6xKH6qaQp1coEbSQTYnTyG5FD/iByBpWlSg0ug9kHOtfUIRShBMsqLYzM
XMJR2wz28QRr8HC2oRHhhC6Tpw8JiO5MGNn0i4Z6L9Q5bCtVtGgoQwe3NQl0XGRrM/Kws/XqkpXV
EZ4cw8We1BANCjYs+n4cHvP0qkjlvLaCJBr/JAt9qxMOk7fWaklr5yn8wz4T5cFsWUQmigePLxrE
CReVuVJIy/4VU0iJUxvUuzoS6e0MmcKTgRuWZuTf2Pf9RayEL2TnU1FjU3DYuEGtR7PLZtIGfK9J
3eawtH2T6G1HMC5K1m1+v8DP/Z7zbGtO3OXRLvE8OPqoM/AAjLWaQJrIr+q7Xv0+n5txJp6fVRvR
kjYA00VJnrToJ8bC1DvF+1tWrqSmak8NGHU6/XUtD3PeCeSACGpw7JQ3q6tRXPBYgkGl7ifRxrZy
Lt3j/ru8JiHuEkQlhX05V/4gfSA6EKNaloylIDjVY+d+k6iQiw2yvYKxsOkKwwDup/w2EjIhYuud
aHISRCBNkmLM/RObQFX3iKgbCf+yryaQyoe4T4OK+cWiCx2tSM4vDjjqCwKKGoRQig/NGlRh9CgS
G5zk2SF1TSgjjnJFNjwljaHHuZceIVi9LOOXMQMH1njRdoqECZ6/xpNnIQ1QHu/268VhKiVk7py+
BxsW5cpXPbKk1bjDStLqB5ah8ACECEVfUI2s8shPNFoRPokxOu0zO3SQI/VdFeT4PqaZ6cij2x77
rlryZOgW0ARTJY7ZCNRF47pdeXip1n1jQdvSCk8jsx0BpcnTyELMsfSW4Vw35MYBCtiIDmHNVwLp
diLZ9o1UK4fmnHSAdzUTiHHusqV3qTQtEu3TPLPCwK3F9tc/URwCW8tL8ZaF9FIbWorYBN8SJumQ
5Jad1flecKxMa0yjwMI+LrfnyJLLlVLhnqjwnnej3u8tSeCyFy2nR3CLqfN9G6j/cwXdfQ1WQikU
ebny2Wq7p7NccdBqXeZcu7MWyaGRHLTf3YPgV7BkVj97T89rbAAkcERjEN9a1Fml4QXMIWiYokhO
+p9RH273G1I8jB+27ruR21FNermCYz1xtgJgw5FU+nqCFQ6lIhgZulQUUilwlT2Qj9R7gja92/ZC
Q/jIwyPEDYetog68tMweKCw4f0Ad2KWQNhSLwWYHH29MGsnfhlyenC8hUbu4NdkbW+iW1FRQY7CC
6Pp5y+sROSq71C4P8+rYACMbvyASDFFcA+5b0TcIBe9LqYGB92yETAK/P4ii9Qr1vb9lF4VYXy8k
zt2RnVDl2OupJG+LoKFOeaQ4SEK9hgRt5iD8eksMsn5Y0btBTVHmjlnA4Ket8GKX4BZAOqlcxq1H
Q+2OzZMY73YzTCYdoQHYaIcSi4A+EIoodlZVGDUoCJsXQCWU1CoP8hCEPgE1uXO0UR8A9OB0zVD+
ry6MEAv9JDbVXaTLSeqB23p2N/udmdHvtHyUpWE/FdXQlQUjLw4R0ejHSr2koqjpQiR7veby6cx8
9bpfMGUsOaI8dlF7s9+HlRwhWzXDBdCBAZYa3hPq9DoiG9oymKEyU86JhFIMVg1JjiVZ8myQsy8h
dqSCY7hBlgG4JBuDq1H+mhhY/kif8V5TldmUKCaIEIvl+1cQa4VyG2iCfgxqi8yzpNGyJdYAtlJp
Ntpr260JNewiVjP1vpQd4bVAFOn1Ko7Dz6QHz8BNamtsywzOrblk5AYnTdpyFcbaZrOA3o1mrnuo
x253vql4iNi39oO9zY8AqbIwGGx2m7as/HJUotzv6M6jC06gg2C/R6qsfgfTpfS9P7GoCRIq3cX2
m7yL+WwMLxklX6nFagRaQmNF7yLkBVpY3bPdt60QrDSUTe0YAuZUcSB0skNByY8JUk4TO+wk4C/R
vLd87mVpxo6M6irNtAnEn7wqrUzDg1rPp3nf0oowgb9DHxz9UGl1u2hInBwaNoY+FjE82KO6b5ux
HYDuWKkJvsc+ujkR8NOkQvVfIBAI04ENDmuXX7RvWJk9WvJcY3YEbbUlqAA4YXk7JD7EvMwdmx58
Ogjl2sAiRexPXd+/dfu2s4GM3HWacT4YB5fhz7UkQR04momzjKxWBAmwl5sD1OvnFZysFBNpgmWM
nRzin0X+feuvyNBHtCTOqg9bQq7ggcHiaSN0o1ZS9RPQmVW330vIY4oaGMXkz+k4PD//RhPfzZex
7lBhI0KOTmm4SMYiyLOmR2mq+OXy3DD1NAWxrVwmEsQGo7LcfOZTUOA6IVGoWx+2hh958yKH7pPz
claRlRkDJRzni69b6BMFSYyLCkHZXMHh359ktdFaHywA0SvfhFrp+DJSqXTJAPIcsQOwVAsE/ZwA
es/Gb6H3e4G3cbA2wB3cKRaepawM2i+PmHKely7rdV7q2muILdsnTNivXpjIp5GS76osz88nSj6i
9VFeqcraQAfLMOG+Jy3AKiEF84KIyQBVCzN0KVxwhvnrk+2fcFiXJHF2mAMMyXuvB7TFm3KNypta
aU4evCN7fI4FNq43Lpmq8yiaHtp7teC3im/564/QhZHAiIfsN2KOdO7Up4q6HYXqXzqbKoHQBggl
7hqAxyGTnWARzifeo/TcjensjkeKIqNHcAftjE867DdyAFvKjhCyoVUEc9phzeyR7yk+v4Ge34jJ
nLjvZYjVMLpJuaUBy1Cyp/JYFOe2G1krxCU2Wv1UGW7V/Kk0PrK/kFm2YLAYtaJ6r+oLp9ye8LSt
uOZbEQcS+Db3ViHySCLNKs9upcWwSAldkScY86Z1c3AOD0ntUu6tJavmFe5v2JKEPXGbnLr5Lgk3
AySfsP62mJngYs7rIFvUvfKspzZ3ImdG7Av3+NZcvJ/rFphsRml96/NdyooFglcRuxTI7SEGTNev
GBf2zLPWpiHe0qcmVYHcmepNjLHsQ68n2eo4NGUTrq7NkqUReJBK9NaosghGBiJFj7ANBxcc3Ur6
UjjKzV14STZ171P+jcvT4lmKOP6CMFazd4E2QAvsy8G2tYatZ8ZHc1bTAdmb0mAODfpwW5rO9irl
jB2cI5Sj4JCtStwUmqJ85XSaYrs8H+3CeKSpqIqrk9GD/3ASIxqWhvGV4khvPIb+MXvUv9GNvhVr
LpT5iLyT6RtDIr6iB7ZUVEq1c08+bYNG9u78UXo+iOW6/XIVuBNv3qZ8v7GyL90wXLRtG8o2TB3n
6IfqBG9zWuO6lytgEIUNVbi3qUsyG7GZy0P/Lr3jl5qmwnGTv/gXlmIjKmBH4EfsfDW9I0FdJr3W
jxp5lR0+OEAlKpgchU6AFJaZ9F5Wq5irLyiiI4OTmV0wsxoHzAn4EVBkQabTK3W7fgoBGUUGgy5W
CYto1C8TC8Xtkwgr3eSg1nSdUNmHDPMk50Yoh4vI7L21Kq9Qbsb9zXKy3BfDBueyhTfhBdRX2tqe
EFTjoenluj2MV5ku0Y+37PJ0ikFaF9HkXaHf56HiaNOqNRXAr33rczwxriSLWdTbe6orepSPjCPP
HkbV0zyzYqugbeDVOk2PV0V5+EZvyhAtaFTZ1zZglgAV0DyditZ2LrJW9XhtSkP6YblZWNODGBlS
G8S9LhCIdvGRA1Fma7A92vTKRsS/Q7UBJv6WfE7V7yGlsZj+zJnGkOOADN8uZiZZiz3qLfjYt8lS
KLklzHN/jDVIjuWo7UoDjdLrujpvmz3x56uEQJdJqA4Cu1kzqn4ABJevdGC5GYPa1toKlB/6mkni
gZ73ha+cB4eAaUs4IU2iMTvXLq4IVMaVgBbH4omj+hrOz9tiGo4CwtL+3euq3VODCt7shqHCFYBU
cBV1L9iZOQH4WmnsC+uxmujTk50X72KBYNuwI+v2r5fVQb1dc8GxV7xMjjETmYuhz5tzYFrKN+B1
vbgf7+rE8sBg2FGG3w4k3DNELZPc1MUKlxt+cjiLsyMVmeIt8A6nQqlkGH2pGQvsBPmn399chCs2
0zh4ufrYJrNxZYRqT6K6XtJOi3PXhaaZg8VSlrKoMESPgPWE2Fvglr+198QEmhNqmpQopQOEwJoY
sK4lRsyidZcRlfOY+HKzaGAGd0qKej16kTv1YE5IFASzfKxvgQ3OsuGkxF6NGmbOufGEk1dk1n3O
UjeJ1S6/oh5wzBDTyyLSrvtsKsEUrxPq9zAA98iBrrSh5lyHH25uvLx5p2Dg/qEthGPb7XHFgfrn
H1zRugKqkXsh4QTew7hUWlsjDH+zcfG8gD9MzQprhRH33BQTBtCx8X0Wuz5FziwwTPEwpmzy/fcu
MAqmqk+5u1yYzG7BmS4u5YAI+5ElNrTCarZ9Jf0JoKTLWMo5zztqCPbkfxy1X44oUEwjxWSz5cGD
Ph0gVpKXNLHsjabgv1UjnD+LwYo0FXHOavyTwwOkfl6Xbjtldo3DcLLWftWgGH320TTAIiiQwUKV
uEy0ElUlZB+ffWQWndMLCRQ4PH58l7pFRXpejED+gEa6009IDKFTuuXcod283lJLZEGHERrua0qi
Zq5J0ODMGIUfQw9BRQOApyq3eF206oI17x+7rjroJrqFnBMglHlrEe7VXv35XhUaJbENdosSFoLb
dAIrXx57Oy+tIPe5+YfZ1dGMUp3jAjhoO+riA2f+HMVsuk4tJqMmPS/29ZYBTQcZQyoGmoSR1ogT
OnOonxvMyzK9pWH6U8phRtgGQ0eyBq+VgKKeI3egPbNlfnu+KNUla459rvdLlZWVhmyA7N4bKWGt
2ZPVwQ2j3l4JVMqMM4SyAWqe2OU3I+6OHUCbXK56RAqhM8Dynry+biXem7176xj1EXFu0wkqPRoy
oM3LEqTmb/iCEsHgx34js6UzKMvym8+rcjpd2jnmqO4s9shRog8x9AVWIQMmf+p5m6+TZ5skQLaf
is3Zm+41wVUiS9sE9kwy7hxs6eJj0sjKvNYkd8WNPQas2NnBfp7zqNATnyRkPf12/SrOMRLM7U8W
WFuUU5Qg+LOaQ3WJmFvvOLA7sspWTcEnSlm1bNWK4ekIdJrfl45oRVyxPfzhMIgZnabaFiuf5rQ3
42UYKzKVxVaVCyiff5Gs52Az2Xw+VOWj+l2DJ4BhNjGExNDb9CI3fqic0Y7BrBOeWiC//wgV/vaS
CbhMIuXK2kRfZTnQNqke0BQGIor0zANSNRB1hyMGur/CMpfdm/h4sYVABF5ViCnzjLkrvRz1SO7Q
dYtpS1LIpyHO5OYpLFoM6gd1LxQCuqDWTdkwHB+zBGAlOGe8NZ9g05RvdxObho/NYXonEJP81UWQ
VgL+hrrh1v0XRhGUxDn7LUpgZNaPqpNeHKJ+wGaJgl1ZxQffjjPoQ9o1UaEK0K5qNgIy1xqaniBO
A8UallMiH8Yo4/5E5rYJPFw6pzYfVJUurI/k0kkfO86HVZybrVVZDRTchMLcNT1907yHcGZLb86W
7/MjYgyyfBRQtMbckLKQ98v8PvVOjAVfdeNGvBFGt2I1k0xafPr5pCzboaCCxhne37WvlAhVCxxg
eDeeC7Z24r4WLd141HBqGON/KWdAof6ggtQY95sKEU6QKBNeb5apTLXylLF5/Idkjl76LvVgytux
YZL5Xlc5+PV6a+5T8+9alm9WFjsF7Ivi4c+mm4YguvxxJsQjbPKJtwXnemWZIE8H/+okmK1RpY+3
aGjFDBGcABvhEaY+Uc/ccRp5Mhfuki7vi1o99pqhjExNtFjGnvTHQa7A0M4crHAIRNnSMXwsNZtT
t3nVM7xfTSbD+/uyUmB2dSoAQFlmZ0bKCTYb21FCY1Kt1L6zUG4CBY3v4UgeIb9TZxI8l96irgHC
03nXi9QDF/588LEZin/F6+HsJXq0cvqOIhAVHB0NMfvHB2Qexi5BfQ7WK7upS9YG8OelP+uONjIC
c+kgWUc6zFi9PbRcpcoYi8vA2+e0ANjDSksvlSWaDkFCx5TrUVcfiPvNyi2mvCNB2EOGZg1BgKmc
MhOgCKotMjTWVCAwkMWL8KjpwRi2rFJxomKYiNN6BaPMpoi7qqDK2OmI/ELnijpuTW2yT/mqQo8T
ZYlc8LCqEBTLEYh8muOu06QZOUObzOrOgi02P2D7N3YoXHnQ7MnXF0KeqRGksL8afSYWvZIT4vlx
wAoCAsswNPjfj9VfiASthBzpSJOX71RfdIBauf9NWThokhoLYW60e05kk+FlrgyHTBFIDc1aalbg
+gR4oKBHQAMveVkuaUQTPLPdl0KU455XceSV3oIS1vmHqove7/t43zE3eOMcPjO7BCfm7FPQ19XK
Wd+2aqBYCOpndWFQPdVI2/TJNHD1fUXOkT0iIgp0IaP1yLFNd8S8Cw4nEORxgIRCOA9Z2bjoj7FD
WiK8bABG4aLU2WuPA6zIMkfSsuDLwzacYajh409pxdcneq4VOF88dIKotQihP+TsUhvNzmMyGYYe
3LK8E49O9lRJm0cZaqZBJaJyO1XNnkaYjA/UWTREvBbucA6cY2xGCu23+xl7uvP6hdrR7MFiLXoa
6LU5D+pAdJi5KuWGkQTOFPHueH2Qb/AmZ6X3QwQZ3RinvdBQLSjYxez88felqYTG55GvcuHEfcEB
yCxz3WoKKubaEZo+mRIzPNc4zYoVY5f3kQaU3GJ0rALMHkRNDPM/SqRWjxemvsn6Uw1XQXAH1NR7
06KN6GLJGPl2SKm8BNBMbxj/qeApJkCIZg53l+9Q4i9Or6922iBQrEFOAMG7gJaL3ruKxEir0Zn6
CfHahmCSFOpfhk6B58VpsL/jngorJiQsztk262bPkCar1NgIsjCWRIPWq9ABpVb1gXpnjD+WKiHU
9+5vIjb1dP1CzR7C0N3H7zoawl5DCJ0M3pHVH0C7KkwE4Bbz/MaAGSXblVSzuJnm2EZZe6DqoXjS
wxVKge7/s8k2oJjU9sqtJjCpRdEey7rMlQlW44D73BAg4WG0a0Khm+FHZ9hEBPPX1UJZ6iWyQ8gk
WtSRebg/VrmS91jV+S8zbAMH3kUKjuATbQDKbYNzh+XG8oof7kVjv0GaU5YIaDOZmocAly1G5y/X
mczptaKd132uvV9Zi+ziEzOJ7MGwZHTwBS7GVhL4yoWKnepsAj2CI48oI32DlOODu5GIw61NlhPF
agHpAhkM6dBGtTt2BEMqi/AY421Vp7r/WkjIrgfavTN7QHwxvxmYR6O7voqhxRsdbK0W4R8dBHWr
lK9qrW5YTYJCynECn28OqeHunFhTuRLhkmlghyw7YrJdVSJp2QObFm1wp5mL7w8SQVwcaiabCyv4
vQjHHoXa5DfWBhQmnXMFGSqq/4iH4Kz5C4n/ahOVIXosAB8XdI87NcxvQsWNDl5ajbps0l+W476v
KU/nPQoZ90084gtwssunjiY+WDd6Sh2e305TaeCKb2ZvR24VlHXKXA67yOMVYBNhrH4P1vLMcky5
hJKtBb1fRXw1cZZOaN4ZzKXKtiojZ+PqKqMUaYsMeDlvJrxIOUzNCqnjWSHdeRB+bBkwH/heoYMU
pCL2bqSGKfOMLdZs8pq7JRmzkmLQpBpTg7k7PXPnUwbRXgJiIge/1MgOsK2APqRKbFAKV9dYtzjn
MffSMrYrO3ctMBsMDKQDKt9YDfJPUPKD5jpO7c4TcO5oWWljxJuaoGLA83+JUqzI31FaZwas5h+y
S8XYO2CqI8cGF4MrR0voQvZjRoOTSBsieU42rSp3xvAqRSx4Jk4zyzDuKG/yEXQ8m8Ls9KTp00g5
PGozhh0AibjcQAOzgSDlz0szRBvb09bDMRrnwEjFU5M6E1sh6I019hq0JbVXJKR9lStMxZwzv7UV
nv05LbI4ZUNfwHByqQU26RF/7uymw89E6Z0U55hEeGXLSsC+6i75cn9jVIrxNZY7oqludFkPC5oz
vq/Uim1vFEhq4ORPkCKWUaNKmqJgrrT5htuN1k5HEQ8v1flL9FCKq4ZVmU3itywsfZiH2DC+fucI
VgHGnksdbArVRa1OuQMxDFHr93lkqSWekW50jfv6pMVQom5lfsmAfTsUspnXCWeMqSFXS8dblVYF
N4AuSyRiEh1LyLY2E+v6ASOq0cI26+LN9bsMuVQLqRYX9Xn5WVNodE4uqIJRC1V/GAi+uFy6tzCq
/uvHZMIsdzcjfOYP/RZJedQaQy45dbvXEHUWt0BKBoLgk4VVWrAfagFSQdTp2Q+2ISzZ365LOdWv
CgNow7LP8hbBtq6LzfH5GUF6LHAEUkZ1rxlh2kbvxf9Paw+mJIa/uPGD9MhJygL3jibS4IjYqQXc
5ifMc01ReIqLAspA6lrcPwO253Dvi1S202prrdV8l1VMXsEgZ18uwMGFkXCTOwkCgHd5WsZgwFjz
jEndczzigfZqXPsD1yiwM6vnxCgJSDpZkdXI9Bt7ZCk94781R/UtClRPeY454MVM5yass67fgkrD
dLqWYmYm3H5Od220EpcomPX+ccwGMj1/yXVVINlBhaYLzXldwLUj6Nz0826SroU4EVZ1vzU9b99D
9JsS6bat+wDoiKOVWaTLMXH76xtsxsPtnMIrTMnCLAOJWmagfkm1ZSHcYvJwX+0HtCAHui8DbUWp
COkLPm0yEjebnkpWvob6AW98zo1pehoeo4wTMAIcB8R+++nWyJj0f473wW1iCBtG1JmnBQPBXVam
wBgnS630PLrWD6z/Vz3fNIv+6jJu5gy/Q1SkSXhpgpQCkXiaxT5tJETlfkm1EdYQm8nJr+vY4N52
GKbYaKbYkGCs0u/f7Lr+azWOTyBcAzOhUTKh+4OmB37uSgzC39YpYmqBWLkhWuYSju3KyUoN74Bt
qe/pGUt+XpwpZLGOcmKW8ix0Jsj3GWFlPMxS6MKjpZaxKQIXG50q89XPgFXVtN1hgWLgkstVO15Y
ct+Q6DTSSbZim0kj50thV0Gm5jO/qzQUu7KN95aLGkdnMz/2rVsJAPIG5tWNRaXwAdP3K+b2lmAK
xyDSCSQaCocSPm5t8t6ca5v2DSHa5FP12YtvRq/lKGC5TGt3R+93GQ/n+eR/tucf5kHRIpUWtZCD
Y72mCYSJYcABIwtJ7YlcrocmKVrZ9NYt+oLr3o1hekHJYFd4UIf75aXn/pggVveHYGr50VMOupg4
cAo6X0f8reaIxhzs9vqwAK5YFa9lBdSkYZTPKP/GEqx4aTpDrn3TcSk8ExT5uBUnVATZwf/IV+hJ
oRHOpKpytxGDFrNI4yyrxTcpCa1FhDG0sELk1sOFdOXt9X5R45+Zb1UTWGKzvF7qu/bgc3PpxzT6
jE4jMtmi4ZNV9T6gwZkySSVQxfZRSjXgvsQhah2QbKpW4SRORCKWfBsrIvAIchlQFTjPw67/xTAz
lLOH7ABMsEClhJUHVqIeTa1mJdfaESUcbPquYcVP5eiSuMDVvMIXiljm5fHd7NUwXTuJvfL4AGF6
gHCv/YvEOhKDEHJYYy7gHY2RkS4kFKfsC9ldDiIMQVix1v8D6zAnq9lUVV5adc4oY5dU+DfHDtl2
MR8ydYOJDqUJGVdJh7wdajFjSjlDPuKhKddAMDpK76QjEBA7R6dLBGOm0ukWS3tmhEDro61CUtXq
px2DZS6UDfwQi1Sz23QdlNfFk1uYzyqY38xB306J4zljwFH5FeQ0GG0qjQ6J/eolX8+3Ntwh5z+k
PN05Nnmcw5DQ9Waz2QXd6525qD0LaCCXFC46CeXa2gvEbHCcEV7HMke55Otz+g7OtK0qKOfVoS/E
HlgC856iFSe1ctFQHi3cvzwQ0s8PAPTpm/ADewK7kKKUjiHX/HxSxWVRi1xn78ou8SgsYGYuOJ4T
oDad9T8UT2zotz+saIwvz0xITlnpVjn0FueOQv1g0pEko/ACXdjZAR8NA8yy+viS3HiSsuKEk7LU
dNLq+969iFXkwic5qhyBG3lXiM0Hx1JVS1/VcrBaIByQpkBuuo6Z0nPN0Zvh1PGK7OvtPd/qjqg5
1oit0tVmOq0tGUoF1izzOB/8NBwgvgZjPJdYwgZXRxlqSHlAF7dAmsDR7V6MthNh4f1PMxVSP7oK
qHcltkbhbPz8X0aOQ0DHWV/SRK3vwW6B2DlVyj+S1DK3bLbUiai0khNhdFmf9jrQz/IVD16unZCd
Og8XinAzJzaoSs5JLudFYzpUzbFwg796p+hBKYMbWiuLOppdYC3lkddf9ykgHp3BiBAa8VuX6pYH
egbfhOv2DV8sVZW0cg5Dw+Z6oATCmPI7JVRZylvMdTVOAFusdHQkvenUhnJay+vVKaWb2imUrCwo
/43uwE7xM9WPAdfZiaaOG3mZIKTP5TkzaJwbdiEvZnM7eLLruyGIVBf5Oxl4jaf2pbBlYRd4UIhl
vF2NUqaI3pmTaywND9qSk2WDAs7mrFnKB9WPuzmezXCTJUKcBcf8p2716sWeWKK4JqG829kVSrpu
C0iLnNCFQsKgwD+yyCnmR5BJNdhBA1qsjligf9bQlJEaMvo+xvvALE4VPvqIliiNnX2/d6XafJfq
YTbvwwSuYNH0ksUHy5SsZVkZaFTBU+Hd00e9Rl5/uh+k9YajQCLacp1iD2wJHmedWthM41N7HvJ6
fK3Dd1jq90ZILBj+mCny+kevczbRFcbQgkm3HH5Fe0lnbYPMu12amPWZOKTGJBL75kYvSqtKYgcr
MMfHqWiucS2HmKB1ZOu13PKnpbdRq3L+scr+YyptuWJk4mahijezN2PTnzMhZLB873ak4nhlrM6Z
XjlG5h9zVyfsyWsKXwdYBdAjSblY+AyNwdvLoSDtJyI/XYto5bZJZRJzZWRrB3nXc10rZWw98L9i
4zXkrFb6M8xa5vCim+574KY/cV++FKS/Dgyd7tfslSoCha/3bgiRROlhGOADMblYs+5IeJm5Xo8K
ddrlbBvTLYpihyzpnUPOXbhTyHDl+rBDzoR2fe3Xz2pLTpNyhC/0fqZ0kuRgRMlLwS8FjRsywldP
X0afNXPmSfymAqTFAPWZ0hGmO2viKsZ2FNsrzOPLS/sPl6FwIhqghHSnlc7xND0XZjgpxGoBexa/
DusFfAQU8YGfPkoS5BnR76cICXCvB3j0t7N/njDGZqfL3hvJT7i7XhvF4d0aDsB0Ugb8CZZnIWqr
BeE2HjiHwclU75PCo3Dbh7X8Qt6bRSrPdY4n8xK9uhCRjMSLI0v9ajsV5WHkf9WobJSFekZ4h+HP
wZ8fK4DfNJBuh0r7Khj3jeGL7IHHjp7lut8HvuSPubaKF8iH1nf3UbAnvbwtCwq/GWAbv+xy5UoB
i2C8D4YaiA1iIwNlTe6CG11Ef0YfK7uuvBXwVRYI8QFoZfPme5SOZxZvCHv5sTXMsswMb0Nkd22t
Qb2jnzNQ+NummFhyNL35EF61LCOEmpZ2lZTer18ELLXqW3SYGivwG9wP58LPrz/g3F/tyBpUikQ2
hZfjhrwKroTIFsT28xymV2zc40yOTdkvRyp/HtXBiYTmHsJ9KzTI+FxWh3Z6M2fCcuEE6rxhq6Bf
puY45B0F99ISwUTnzxiwAvkWmSzGX7plp1pJ4bl5HJL//umIozGbGTPK0JOoLd7o+Uv+kmV7x8Iv
j+3TnkrEj/XliwDwLzHSLueoUhUUc39L12irVfJm04WqVgL2xl6KakqryqyOg2j1cytgOq1hPUy7
JkvFLGImqkRnJZpCd9i5XIDwRJNakuYdsQC9ZKJbIqE88Vg8VkDk5pS+/mZtiAAmpNQGYs2svjxd
tGi6QgxiAYTu81h6kY33BC3fc3iMNldT4tfQRjy+6vMBSGYIlHn3DyBgpIflDpoeYTBS839y6Eev
akSoD+fgD2Vmc8LC0rteO1ikCEbSD9Ruo3cjDrnaTABDPxeKHOtpKUu+3RB+PJ/qObfjN2EOXV9U
qR2jIXg6BDOsxvwswE39jLjTUOhUaARbUUwxRuPXIbrpxT4fh6cax0nlFgE9Nz6g2mCfGVjIrwjn
sUZ2GiEhd839zV3qvsEv5t4rm8wYxVGT0kj4cQYKrndfjCBtHvwgaIfHwOnGJYbsoHbVboZ+PfXm
sAniuNuJgzPFP6vPuAI3FbxRUupcu3XEEs554+RNJytmN2GM5lF8K0QcqxEj3nYi6D4UtgSRhcNB
dNUoFyOY0HdrwtsJtgvHRzAb2tfVCul7yBsEMQP+xlpms4fJRT4KLpjj0LkAGvnRXeV03YFCafmC
h1Px0jnEK59vP9mv/U/qbbrbGPMYHOgk4PmisBlXTleNgGdvu+A1rO/BWGy0IarPLVSTARPcAWsj
Ds3zvzd2ofiLdcy1/jxj/mKYTE4DOzCWPsQT8bkMTrSjIvON5u10F1wE4dggnwEBOQ6Wck2GB25m
vZ3bLc9dVWKZ14XL5S6LVSh+FHv1VGNZmz91JMZ+xYK6rVRGoF44L5Oh0/KzLe5/CP6kFAgBkGW/
K5xUFYrtwnm4kQieO5xO5NeOtHrGHhpdBFyySSy0BVzQIcdQKGQVoI7FAFlPIGji2rqoKCupnM7l
tI2RisyLV3q8sxr/GDWdR7lvozNDX1FrirtrozyGGM5tpkVJOQyHKoss0hq6jBMlIVlNhMGQi0a6
/0xb5TrpuOoz5GJ16sW2P9ASRZAbza04FWmznAht/jor43sbG/nh2/pLNkj0tIgPTOxi6sX9xVdc
F/dLV3E8PDINTnUnXs3dHBjtQawFuwSRc/kNAFZUooftEv2RLram5du+vA9wAQGKt09iBJRlsetz
IXw0zYHU7xd1LmDb6CX8pcalgwlcUl5CASBjU9xiLNAlwMNzEwJJ3OKQ9BVgfeYjhiTKgDNc2g0S
DKj4VqTCQ2TUNIscoLbs/7Fgqisyp2htl7szV3A3oTL1Xr5X7vFVHstU+m83sXFs4+8Lo+A9k4bz
Tx8RzNwxJ44NydldDwzzT5v1jDJdWV5uCewupntghrtCjIyDVhvBLdFuLIermZ423u1Vbu3acITS
1/Hfbk3+eDTudv1zNA7JGWSMrvsZgAT7ptelO9lCJfwWSNafzivJMn0R/BvGBu02BAXVrtZ+P3Qy
SJcMtDJLISclz4F6ZQX0A2jVSJw8Xf3bV6KhqA/oSf6ly1LRynbX3zZbGEtlte3c3bW+Fub4Zfep
qWc2F9h1W1oXJlzexJ9OKSc4zz2PMlGul8bvQaqqi74IdCiSV4lVUZvWTzfTaEt4n5aakpMULcvw
o1+5n4jxXccdmqiHEcsBUpQ3w5jV5OT4VdJccECaGlMm+uo8thdaiXMTiyPiq7L35nGLjuU+5X14
/JlxcsGJV9ETfyaNxQsKYqYzBAZXW1AAq5pGTnbnlvchXVbPOIiiMhvsb6B7DRHqyhpF7vCJye2m
54rf8pBJr4Kxa2XK7D6ZklbGiDnfLjiwjB2EHIW4d7q8BWtXCIjwZvz6farIvCtW/LSkNLwvOxhh
U7m4xaJd5k30k+LBuXkO1QH21YaAPtp3wDVOubih72CBl1yFl7eSugnVLamJXflELKEvAn0uucKe
Qb3ti94yRpWebKRw5nho+z6Hca3vqqtFWoPccrSNvxWmtOF2/77Pun0oUtpTZubhRTFVIH2/FKfA
5tjzS2AxfxzfLIlj7GNuzwi+XV3714Y25hy29nCJ4SaiCmtxFSPtOjJtQCd0/Az0X0m9hGT0R8OC
g85z+XmifVc4S7wo31V+iAUVkc7flNKRgj4YoyivBgVqL2+sI0qHzG4tjl+9j5gq7l8/9qG9XBjT
UJj4rIUkgiHljLlWvEkwOjRWfCSga7XscRTL6N3CHuiWLKrThW4c+nfrbXzNynK0PEXriQAYPkgF
+jbw3FMy6d1Go/WX3UOpRuiZGDKu5aVFqdfi1jUroOrNot9CfSfNHZge18d5xYV4T1PTyRHHGY5G
wnIm5KFDA1Zv7PVBX/PRK51RRA0U7RxmRE32MOHH8B43XeBx355YGFan3fgxxa8FG+e6LrJSAAyO
mn+fB1YxsDAxP8tUA10VMsCb/bg+CeWSNifzaIp+rHEo+5GXUNMQ9vrCMYC9bRS4WPgeDr0Kw2P7
ULSVZJbeVZt9x/ZNxYPzGSuUddCOv2RgNweNlCY4me6COwRFskjXvFj7c7KtTpVdjXama7rrLmTU
IYZQQ+JJu8hW5wtKItjRx94FogQCFROsnPeWLCzAl1+tzTVAO8OvyEIyXdfE4S87qle8thGfA2s0
qPMNCaJfr2okgyjHzRtr7KYVdlS9Vhg64L4BQ4ITlKqOnqO2X/VRhZr2XGe60Ac2t41ZCRkNUeqi
iutx4qMq1YjYtk5XqMyUAd6INmmELw5KSwstWmewPSny+w1r988MJgZZuC43JewbMb01rbGDzMuH
Jk1FdF7WW3iToAuBQXRfDg0Sg62tLoJdTKf/xYjV/7m2fhplJZzFPYErxvVhv8dAne8yjwDCQRLW
M/g/gLIDKF7d+kbP/7N65f42392bwt+9qouxj7I7kgZhEGQ04UtQZh31dBoEsp0txgTA6VlGz5no
6zNcOObp7GN07wOxv/hszWr4DYPq6A7ajEMtXkyCuv9rM+fUq6ObFFeMiDyIidW4HgacCJJ0jf9Q
dgSA7aE5j2n7VBpVNp0AS5WiAxPOuL5N2ioRMcGdWoKv//gOToeOtcC1dq/eo7sLLBM6zh2h+Qcy
zSSwFHLdK1F927lecDiAzPcya83ePp7Zh2kGjQLOifD/h2rLRNTHyRpZ42GfJGS00ddk7Fml1VfH
nfodzNhjQi4fTozofNxukLJZX9IL+8CR0qPTvOHo6xOkXFYyLDJ7MQKgGK/+VRK7enfgRMojAuYD
mWui68R4JcFDIMJW90DnclpSxAamYmQXSXlcq0rtt3EWOh7mhO3wI09nBfJYR7RsQmTAftDD13hV
5pEj44I2AkEd2MyAtQLolpq16qG3XAdgybVIKwvzziUl9AGBLOXc3d1tNS1aaSGlTzJOMWw+U/Fo
v6FqTYCZqlytYPJOCiw++ivNS1AQVdIhFZkljn/Efg4J35fYXXx053MYYl8JEUWgGaplgersRewr
E/YZChWEgSu/Ss6O/S3T2Aw/FnIZPvcG/zXECJ82dpwwxGuWgi9aYDND6wGqxEbHo6bzzcjJkNHO
SOIkK9tb7s2DCfaq+TBcYawMZdtl3iNeMbSRDxqYV4LQs4dsiMYv2pV4nUmR79nYoA9tMZqpe/hs
skBJEUybztEHnCJt8TgkOZergPXfgNVsHp5pnx+9LMfk01o02tPDw40/0FtquZ2XUoCCBjrC8Tl2
Favq/SbenMCaGs2OzxNi4Z0xLNmiZvSm8A7OvoWWDr/XLU5Bvmboou3j8HlXBJeeg9mkS9WSMe56
lYf5dYxgzZar3G3TmFXjjKScO0rRdILDhGS5089tFCZefT51vcT/KWdGqsMLLSa5yukKyXe0wW1f
GYYXnfCwtZ8uDijzHBaVoAehBM6hYP4FPoiS1LPtYGAYX8kjnNHRPKhk1sMthRZOJVsV7Lba4PqQ
s1Ex7t9HDU+nd3IKBumQiWtoXRITOI6bW6G9K2YOlDAV9i1JytjK+LXkAnXBMoQYCi2Ib5NRAVa9
WgQ0NZ/C9+eRrrlDRenJloD1Dbv5whZxgeffmAzy2FaPpUavqPXfFpyg7g+yGzBkdYsI0KMEJUzT
z7OO6X/+m14wQoN0/2Ovq7nOeGCNCRtxRrbX0G11otoTUWNbkqslmBhu+c2ZQYE9y0jPkHws89eY
/ebZc4PQvPyApe0loWzEjQdzuQN1egBW+vaS7t9Kt3kVQO9QKLcWlOtuO1cn7S42Mk5N8AZRgJwP
tjoTqbVVfCktfitew5ej0ssP01Uk0qROBBWHB0JvPji/rSj4w6a2DzyehvuUEZeoLRqom0awbIed
VNHIf2syY5kvCuylIcQEfokrm1harU93zYydaqo5sV0Zl953no2eUxY4trTlj7iqf/gycMoF853E
d3poWiCAa6Fha7c8P0+kfGJ8nNaBV3VWwGQI4PpBUaoL7ir9MowVrTFfRN7WGizaQwW9aIWn/SQC
/Z5/EucS3htFuD7x/tZ6U7++EYoz+ZRlDw0Kz3A4K8J47Z6ZpOOstNPjqm1vITndoOuL1rOU8jnb
Vco+XPZiuIgkuOmQ6wHs1BaxOLAzXUKYE/q6VTQxljfWjH+s4K4KOZkE9t0A6VdvEXjj7o01XygP
YckMXCtRAhnHZ4lxFdXuqXDDXrK5ucjUTVCv4mHeafmB+CX73Wo67iC+d696m2fKXi03Ur+5zCWy
lyWmCZ4/F4b0+fN66EK5UEHOeRCT/9goINu5WEc12JwGvHKNtsvio4jXIpSQnTfY0Wh2TRrRhskN
kgDqJHcbY5xbyZ5iRk7Cg7uAEXmqySDZKY7M9TCmPAJODfASoN5sdZnVuKJGzIPra02BAesvzhT9
jar1zlOt7EUwLlTLx3sLdCDOBwsWxmiRD4LGs7DwQXJSZoEY9kZYr5wN6hbdtm1Jl75X1qN5evz+
ZrSwEu6OqJp81aXucwXswjl5x9o1qyyLdcdetFAotBwLQYaZpco1k5upCxO6MC+BXFSd232ITFfQ
HpIvcMRSXqzdHAkTKNJECcR9UfcrYq+M/NpTDBVzgbJEcoftykZXClWMMmtzCQT2/YfijGkU71yF
hYNRIdx/PBB+xnyT81lGA9d1VuYpAXD+5wTXQlTM2bU4XuHtDb8pZnHJlNHcsFey9KsGwzt30cs/
ID+8I/ZxGd2ET26zycK2eVBCBeNOwD1kCUtBrCoCnX6Ogcp6dJ15ZCZ9GUdFNf20Y+I1dAVBlzHE
nlDYYmoXiLpucWTr30tB9tVKfp1G/hXNZPbA4XueAYBCMQ2nMQFSs2KUBxEis6ZfB862UOHvji0i
Xnawy5SmLeUKyiBOZJwDStK/DSolIC98+In8pYovSlbwQGp4axPJOTcgmz7PFcGyWM/auOTiWYhC
LV2XUYUUmCtB7uLsbX29P36sLRqm7iItNNqKmaWB4bfdhTPLjnJ5MZHy/j6zeJyekB8i/Px+DWaE
062VdkolD90dGszY8J0sgj11sicKjzFTMBUB7jLf4k6ldxH7d4x5XxGawqZF3fgdaivbjployURq
VGlyzV5m9q4HsSYr8ObAo47ue3ZjNBikZ1d+uXKaBzcHTfNvIsxXYrPY7U2k4SYBul4tqES3sYgd
neiTR1psLsiJpU6UEAv3E3boRzT2FvczawZvGwt7L/FD72v3Aeig6QrqV+ic9IOB7/o1K3OxrVos
7vl2YLFWDyvMXqUvJC1nglM03txmRjh1xO9JKUJGU/M86sDTsAPrjGc47GUtBSQ9eP4sWd900SZp
8Na4Rta9avY6yAOVpS5ivg513Yo1VBLlgHEQNLV5c3v4o3a5iUNG9J98LaMaqU08WURWldlx3sgq
asPs5eIoRHR2pl4qn1J2Dsdcxz7xLVXqq6NgUM9dThlmnlJBCkjjIZpotGuIwJL2rRVAgoRFYsu0
V0Lx0IY+jWXWwmtT5vv9V+722hqMEPYJ8ysJJEQHCLea4aFiEonvTd7nVfg3p3scarUIeIk3WYx+
PV8NFZewUstGa28ZeMNl8Ndsz4AjYHIBA1wb4YuwaowDVrsV2S7wX/weVgL/cpeEZ08a0wHYiaYQ
2NaKacC7XN0Z/LF9wR0YvYl2D3nfwrvcz2CmXc9/2PALtqjuC9mkkf64bTWouxPDbGZDoWOjGQS0
l+JcBtEghqzcY6wUUq8AinW0/usB6qczCiBb6VRHDa4Ul0zPIEMXooY/7V/bLHuUM93h+QJpUwKG
AIIBa4nfM6MFg+nPGluAPEkhx3hgnT5mgaw4S6rBf3+gAieyzV6nKpQLU+JSWfLbW3AxTP8642Zt
EIkWgs13AA3n0frR8Z0ZAUq7FuX0cSOgwWUMp/Fz5gHBzDY4Bs3vmiXPZB6uqXaYarUA2jnks8qY
TnIgT/0MStWbZPPEk8pJ8H6ZdYjcpE3V6sSCLJqlk0Bs1mPSPLjnHOsz9LvS5b2xf1o4TF+dFw+d
5q3Inh9lwteX2Q0PbrN1YujOIW6iat3KvsOX5VreRP9Fz8BMYNRwhKFmWLJcDsOXRMD6wz5jMS37
NBK4XZAaAyHSJPKGOe50xl7mf2NAshWtjEV8vEUkIN9DiYnEgQHAUCDGCLn2qeRrpJ3u4/31jr1k
ROvcRKHfifNhyEuGwBSlCgcs+oiTfHx10iSdPMVnIRidt+xTzez3vQP7yjZP+BL5pPGGkGKplwu/
5SG8Xt1EqQX8hxZdnks9HlHzuiNIm3muu7Oj7SEum7FAH8bXkMxM/9u2pqiRbGkGDV8FvCiTkHj2
C4xHh5CjyQfqt5G3Gl6xojoF2WSdOMJI5LEpgcloZaJPt6T4CIAYI1AxMbA88F+8Zr0XKd8fPyXP
4cr7DFjCZQ8tj1Q6ISkpiY3mPoy8jJxFqADShHM06RrDpRKctgTNf7cviBWJHjVj+suUkUwRYYAs
6x7UTY9qbyWSolt+N0vQne79vCCb0lQZgEgqhnPaT+umZJSSaU+3J+/Cock1ppLeDcj1AyqIu5Ak
QQ8oytEo0x9GBOwTo2dKAsJEubhfCshDV9siMtkLTojmcZ6HiR9VvRtjfGIx8DCLX3uthhA9EviY
OHBXC4k6ZlFEO2LLSkPvgcHYzdOnOdcGolXYV5hHhTPb/7gUsOmNVpPB/H/UCiVsQ4Wi6sAJVepd
2P+AqwuPML+F4r87QkCaZcNf2UcE+res+PhUzIhfgq4RqJwVXs8/nZU+iX/AaPcUWs8DTy4WEHKi
eOhGjfNfzTiG8s9Yj2qIvLkuuLpfFFPE9uO0KBqVtiIGKBrYwA+OTTdQ2cJL+GyAY5EdmcobZeKd
wrS54iWSQyD/oY3qfMw9SD7CJbX6r2jzhhCmc60DeWfQZlmBn+JnjCHamdyJ7cNcLnQ0ns2txPj3
Wbw7AUQwYUUC5NbxvgJP+s+rTXs1Bei1czzG+FfoCOZbmu0EkJnHBNta/U7W+EJng3zPxiaXIgyA
4r6SLuxAGABAnNKveR4Hnmuo60JxSHvvYmQArNTgaHTcib3vkRtfvDC6ac2AN/bcLedFVKyINwKf
KRiUWd+kZok/TAxaBL8INA/WA7E8q4GgLWoz5iJdYITTIU61ke3l5gmLG2q+ZP6VGHAZs7MDiAhY
pOQonIMt8Pt7GyaZWgrq2D12xa0AIfFct6ep7zO5wxHFvx0UYk0AH/XFsoH0NbwMXO779SbgiLaX
ZJyqEGT2KBN+YH4JHrzwYg9+A3TXrUpG04+hfahGUrtIdlGouP340EBUliohHomvEBlUa32rSCXP
JIA2as1FnJICRFBtf9MLcAQV6W1YmnSMOpB7ZGK8E32gD3kXt/S6ijH44ZOCjUr2E71e9TOiVkU+
Cvnb95LNPqVhotmyVy6lsu2usIX4mW3XJ/CQz0rb5Pn/5ygwCOy4PjuLRu4pBaAUg8fJkbg6efo1
2fzYhJkx4IBpyS0wk/CLT3ArLPASsuEl1aJohaIfbKmVjeuckm7YcEIGQzyQrEgmxcnu8cAstvsY
2QAwnkuN5EzPKj6AlJqyGh6Wrkriu7hkof1YP/NETDRQ+CrXcu5ylNYUCQpW0vIgm50PBmJKrc/7
l+1cSk3ER0bRllMz6WhA3vs9V+fCfKhBTDN/TVpZUzQJx4I3dxyTdEup99VzJyLrlYuiguhEpWWK
g60nerU9PlUSSnqVxco+cfWrDgdKV6gUOP6fFwpjGcU2LPqttUlQqguAaSyWShHaN6QcTtrjwFnc
sF7z7w28m9X+26RuNQ6Qk9Io8WlG4ypRM3eKaD1rtzZ8pagm9LdZh2RclDCw7522JL33hwRGr85D
erx668j1S1ArBHTtQhTDOvZKJEfsvu+jwM44/jQLbYj550ydw9afupteknRImfkrfY6ezemNy75o
/V1e9RXagkX+pLU/t3cU0IpiXkwyM1zeS15+//PzxU+NkgUyNISvbdboMXT1I+6YW9ss3ddUrP8m
jm0Hp/zSkCRo6eRde/8LOqItqXWA1L/sVge5hciDsbBaPZ/m0kGiIMBRFbADVSGbF7H6AUVummhu
Ifh91tC2kRLvUHfUuUj/8X8PGK4Lq4kAni9h0jQCDhXkm8ab9V0OJCEZLfRqwXwLgrjJNYv0JYe5
VVvbYcbtgit+iK6L2V7BkE6kV7sWQwudekmZQBxzDkY1AHYRdDZgOngU9GAkjcSCnvap527WQNkl
Ftjxqcwq8NZsDyydm8DylUhUMXkYADYAPJoIiK33n3oiiIyV7nksR8wToieHIU9T6zparX6Y7nLL
5VIcDmUROETyII37WCDj9yMk7+3wt0zx7dfd0ccAV0QWAmk0IH8ZcOL2/EiJp4kOuOsj7E7hrOWy
4wUovqgdgQDxGj2AyLneLy/oNO8XV7Xha6SDmKD/Ioii76Wqfo7fVsd6Vc3xSNcXcGPNmkIVhF4l
HSkwt1BtKCj370eyJZsbDcEcnsywwNxoL0hGbvKGMMXOS9hSjKeVxAGLKn5SeRFQwuzYZ/o69+fP
rpIbMKEB4JJ5YOtV4g6FmYkY8hE1hfHlykadV8zX5gvSsCf5AslMI8R4oG9KpuL1SZgIqw3oM/hj
CrfgzKxoFQgvrC616r8iX5pL6N29SYvvcNGMHvQAk48kTmQB9iewIenYuk4Qmdkp0UHCpd81pSWN
ChcLvrnHog5XyUf+bOxk3N4DBPEDLg6jc3LVnT6g8f5hhqQZYW+n6Mwnj6pJTKI/9DpWilGLjO36
0oFYON79owbLZE7W0Op2yv5afiBH4C41OoVIPfYlazrLBnVJgcfjsRN1qAZHPIgKnenPhQc7njV7
PvVJVR9uw/EIPXO5h/CfafW0QeiqUQov5ND6N6TgXdJS7WWwRCHreggUCwhUqiviG7BHZH5vUCj4
TD0L5qEMBeLw03bRojI45iNdKNaUV1g3YpxpuSnTAR1WzloWGbCobFzuB45QWPpt2xQpY0Tl9yqa
+b0+H13WS8y4hvoy+ejpE8NIKTfdYzCxwsMi3s4R+k5anmwAS9XRH6hNnmjyHKElEbjgaxr3julu
YRvBoBneFonWn8mwaofNQJ9eXy1Hf6W9dGfE/4tRcL/RR2UpQnczS9iHugxwhzHd3pMdgIEpY7gZ
GW9i+jO74Gv6VY6I00+SwKeT4lR2sipDBX/mCMsrJaqyf/XZ2l9JJDNsskaKGwuO2gZXdO8z7jxo
yIpMsSEk5yXHgZam4+BoZYYajwxG2k6uowhIMvGDei9FqMB1eKrOOXATzLbiUd2rzEU7yC5Yolhr
73WL4phaoEIEQ3DyzQkNwIVSyzIofcT4YH59lQv5iW/TVcBkbY0lEahMgNSEXK8Gq3jthjIFafSc
6Yhbhv5I28ebgYOnSj7mPvIWGaUXazTfgxSXIVefk09nYwpF2IxThRWEEgmCDRuGxwvoXJYYy8ak
aXLGA0K23gMFP7Ug8KrP1gj7RVyZGYUkxDvBX/rIO+ROGCde7Teyex8QxuGWRp9Yq4mq/WOlRd8z
A+/LgJ9hbGKc6XnRHdsZvnenCdXPvLCMMv4T3fqhkFfV+TdkffdiYNFl6xlVUwKIWmNTCt1ngAT8
Ja/NKQoLyEV/un5kXQineLl4C24gTUVf1zBiMhdqC0vmHpp83vm07vcq6OSkUNR7URHxAKoeAGiw
00UwAwfS3rBFkarSTnPmaAXTlspJkE9bBMFTWA6qfu1vkBs1lsfLzZ2GSCP/fxQB9cdXMC2my37I
lrTIOwwF73/hdHsgkktOlb+Jdoq3EGCSSm4kctbPM+ZimE7YgYYxvEzOVo0T9TFVO6JZVShPk6Jz
pn3w2CbPYrB1z4Rti/HwdeKas3lmssnR3nIJ+36ANUsE3FeXO64HwoFMn02hbhObLtvWkcbMy36Z
KgR/SO58le00tnNHstSmbDK5mg8ycqq4QTMrCc2AEOHctjVxXZ3t0fqRKWKGtoJSYwkhz2+IPlyV
8JWnry1nIMlgJOQXGhLUqT3mJzJT+R32k6MYWNllxarlgliNMC0Vv9cRJMga1DvZfqa7S/thS00H
CmRj83+HRCsWANM90pW/M+KcBc27Q2z1NQC2kJZgvF0yQt96Psap4eTQQYyAmQOg0KZKQMI6Epwn
tsNMor6Y3EqM4D+mne0QsE3bkT8x2Bp0C7zyRGrET9MD/yKNpGJ8EwU+b+CNTEtgHaxNml9WosXc
ckBD0Q0O/Of7p2lPdnaRt4if0mBl/wVgVd5kJxTo9ZMwh9T5mPWmZh5RSftsojQ1+5ZlKoPpKdNs
CzYglAzWtuHAyhNFBtIkblN1Y+pkjVvOKFjuKwn5parnTPKd0BoH1MSNyY4tQkeaXKO0jDQiMEod
WYAlWdmHz7ksO7lmwXOunNlHKT2uAr1OaNslrbYVMy7NNwUMGtpwCocJi2b2u0QtbIvIGzQbADRR
teQR1iN5camIqlLdG5G4tG191o4ijL4Wp6RCcX+iBAVcabuSCqQMLRD3KWXBsl/qjZEKMAucfxq2
k0gSxOfYSt6HQHD7bXnYRkLNvxQdqWPtMZRPHQIByoc/T6vE0fzxzFnGEA5i8hH/UTht83B8rSXh
Hb/NyGje/Ypj3iKsE0cg60tul8gSzBiCAaOrFGFne9LE7cX/zV1PjV/gS66C+ISeBY7BRIRLW6iQ
luB70gzvZnpLItAv7nfuCuluuF0o8r0YW+K3xTRMTjp7CF1P04AUYI6o2BN3zgJcNjis/d3+sTBA
SSJyg0CS/5u7M94Um/1gDS4kfmZRTwgjXx4edmOEcbMvi6y9tievcQDNulgyvMORzqIWqGkPxNgE
kN5OXnOGQrN9J7ZIINZ9lMBBRYuv0k89atABZJgVLx1PdaPnA//NtR+pzPZ14sOwGmf+6I4nE38j
uBv7HnY1m13ugesARWZjHkVFrERTu9ml57O3d1/7ELTUNUz6jdQ23J+NhHIhafgDlg3dQ2jMKSpe
g1o0zqW1X4Ylgc8eJfWYdl73hsZciDzj8UVB40qz/FfTKbo2l9+B6nps+CzUKhMzYoA6xAwRh6ab
ylKCzH80M90ioaMHY+H51UKmOC9/SFRPvGxuIlgBXOOkNoaShVrz/D/wqNqZ84bLDMifTRM5Mduo
YzOyIHdoW9BfQwh3kGh5m/PdejUANL9NRSWHtjZ4SXIySt5onPoYkcdD3qvpZjdjHL79E9JItQox
fZCeMCyb3CvBT5Mf4yCzT/zJhCOiUQrHXVTxSysLcRs7GN7sN80m8RnrE6wtmQo37DEulOQtfBDa
thTs/yKqw7VGHRn4MIH5opOdeE9J7qhu6IsiYQecw6F6DsokKpkgox7JWaBup4O1Lix+PWBWtprY
vwxxFLkLSp+QqLB+VZrFJsXULbouCjIxqjGBW/ttZl5sWR99a+U+4Dlp3fNYvfyTjx5PlyegV0jt
x+vG2Qshbx4+rhJ3xR9fJlsxTA7DfjrZEn+V6io3pDtuREcqNxuUDsBSiHCZVDGN1TXgdCFY96Y/
Qe/VfQkAYnuy1Ousc2GOu9aSM84XZZtbJkenzxz0Tv5B9ApxquDizSxDxmTWsWbFE5m5Q22KGasN
4BG4HqkDqx2Nnb+SEmMWVt3NSNLwy2m7+su4NbQFjtJfTAvdVN0Z5KRbYrgAw+K14Sl3HcVV3u4p
CB6kwl6e4SbUbkT2U+O8305ESJ2buRkd9qp2bjd8gEsND0rcRt9B/omMJJNRlvthe+130DxZpsYG
jBxv/ADa5+VjXFMnhP4Hli/M1u+BCEBcuD/kflqIpBlOzUDOX15Vcy77yPFx9ORf1agjw6LjECTK
qxB2tl//FYuHd6SCEHeeMXqqS9KXLQBFW/luBY9YqCVlhXzC/7SJ7lsxDgn4UfZwpnYbFX9YsKKV
VT3FLdpycmjhx9f87Pqdhjlla+64t3ViY9DMEWdLR3GYfNCjIMboGR9YyZ1jKizSuVnDKtLlUML/
U0WP8PyjKkzlTVoijUvzCARl2oYZ88GAeL4/WRdxjMjlQMaZQQVgzIyg8fhNS3d6EUTtPyuvRKje
8Le9ESMWUYSqPSryB5o6tUyPFpwLSCCjMkWBbSIH4n3DMrclF+5o6cV0v4sgosPS0pP3hVsW0/Lc
UxtmnA2ugAUtUE/BUJH9JbRZm3uuX1NPHetwWCQ/uQB7/Xq56ApiOhBNKnWA1cX4lADommdNrfvO
HTQM0ZcogDF4GKZkiRPD8a751F86EjjpD08kf8rJ8B1e00guOVxru0m+K3Sjq7cgUwkbsbjmXiUx
VzHvmjODQnLXCvfOt6QerFL3E6fBj+OKbQRlA+Z2yMhv8IXCQgqBTsRB4CDr4a2fzHbDvr3gEnw/
z3QHfZwRqWGqhb4ceQ5Adk8apNHUurgQh4vg+58+aa5orPy8MNaTsl6jPlf4/Z8ka8KG6JIx+ZfC
4zQHs0L4O9+PJF/wwY9YTcRvlTNPWCvW6otW5WKlw0Whrmccq7yX97ZlBJg4tXhqv6uadrTdh7oV
/oaINZsDlAcXj0xV7Hns6NTCui94S7cs0Qp9CKgCXAoTkiS4PA0V8mghc0nfpfRjE10q/bS35IdI
4Jzg/C2cmVGAo1+Ve2Tk0tQs8DlxAi/2mehcTWKUiMgn5kukM3FE7R2JwdnS1T5A9cX5/2UYHukx
Rirj7+mjmgFzQZV1dEPpA/uD3NTpYdZQaWtVEMXG8dGJ5ocLqzhC3lHwpqENMGvwof5ZjDLuW9+w
x4RizURdKgqESyoZvLBpR2k7PErxJUieUKWCI8Lo4/Rm63V3dyj540tu1OH+0EmOVK1xCa6ckPaD
ZeNRuNS8fvGWWURtoME367Sqao4EdVPG9gXqFDHmxXiJNpExS3NdXry8vyiuU0ZKsl3hK/QoC+dx
WV9C3nhpbtqKLun970DYa3M6Duy0HCvTnfn0bm5R8VWBHeSH+HVwuE69BEy6pl+XhysIyzJL3uaM
NigV9LibZtu7vRjzgDH9S+Qn+95wG8qCt+Bm65v+2Vp8gOtMhLj3Eu2G3bmxORtXVUNGnuty1+w4
2+EoeqeS29/1y53BStUvIrpiXGVkn24r0s/321s1JqzqH5dJOnfxA/Wm1srZd+lAG8KEmEcJTX5x
YR5f/lntuXW7wCiOSFSE470Wu0brmLb1rK7EBy6rD+pfBFlCoUnqQKURXzEdMpoA/12QqdyLev5Z
G09c+j6M7osA7/rOX9xh/DrY3pS1PvsXIbDtJUjS7sNDLjDdFuMi1pP0SmEnmoVECD/xY0kHSkWi
Rs2SB4Lrd8JY4Ip1Pi+Zpd6aFRC52EZDxQwQVd32Oh2vB+RxxlEg+0nbVWJ+zpnJxrjjHu83V+1x
VUV1vJv2cpZYQm9UYe9oN0jJaYBqa/2TbR9NLgntJsiuCaWC4CbVU7EPsrrFczk51YEkIEACWQNS
qIDx2H95cG8h/I0JZXFclf9Ycs1wDwG7cnSYk2MJCwVnIpG4/hU+H/0AnF5rx526Jhn+MXPryAQf
pAF7BZsfJq+zyfR6mwLX5fTWynHuW9cf49JJqFAv7yvkHEI4LtkA8tpe1yWTPTPSTv+7dWIg3sSz
6Yp/VNnOyNjto65x2W/3zOdsxtHk96My17uy6rmIMj7fxTu7X7LN92o/V+usRqJ52dCORcVZZ6OF
1wB9vwGCgRCEbWs8JAOu4kE3QiYCGqbUU/YQYY0ABsF95cn+e1qSVKbQfgHwMvm8dmNM4ERlG5yV
7l1RhNoYPYoOUwkZrsha9N3hQoXkmd+V0s1BQvn9/kK46KJlDLmlcFFXifD5NFfidtcstLZ7HI4h
0KiPa+QBUZ1gZcjH9YRWQoHffRPLqVvdmDc7YhDku15Y1fXyEIOBrQxUNb1pJytQXwijWYaRZKih
xuQEp3yUaZVp2QiieZsk48E9jvytH+r5FMqDR/k7BBOzmEzrHXx0pqEfP6sUu0XWM1XZml/f5mQD
lhuENyPuwnYS2tNNWs0FtvxVY61b+JxNQ3MJqWtGwLxZmtu5taNfanv+wcegREBJhAyAGZ5y06NA
wmJKz8iMzcVa0E+pTT4c0Bl1KvETH+fkn9jjtg/WTj+5eX2911dEJGJHSsuk5gGqcbJZ0g3PCku+
cJ8acu2cmGobcA5FnJFzYDGzu+0UXByz3LsWMuC3olVF7tAv7EW4nFMeuM8rMYE9+REoYG9CHQ09
HRzo51G2wIUxo0+QTvS/N5mozCoD6FvVuVMwQX9kx/Wi0pfuMQQMCSTOnEkrJs1SciwHJeAQVcu5
e7kVpsCiorCTW4lKchWhXjy8X7q+gFrxuz6V4/RACeClTsULmv+3bORWuYMraIG0VaRluIVGs6gj
sFnOGVVq+iA2TKE2BHB9yDRu3GCuks2ZU5d23RZywmF3Gs/42UyCsJN/r55zUwzPuubp0J0llWLn
8ryNwwK5rWbr3dzy84sdCKk1gfVzYRzToPMZ98g5fVUXiZr5eUDTpEMyu9GYIaPOlbxJ2ES6TMSf
o8TaA0/CrvFtaAj9uuqq1HDStBEt1M9OqoOBU7t2XXivIfiLuPiL1OohDeAT9DhrVCttrhDTsSmi
Do9+MiGF+ErIxwA2EqUDAHSs4Q5E5bpfuQgtu+quNpP9zr0jAwTZYjbakvI0/b7VszZDMKmGkWpL
Od50b4bfGaXm5jq+gbg/1QqFgoFskD3/4843X95ODnQ7Clez3qWKfrFKfWkIC5jOmeJI0zaD7jUY
kr1XqPP+ubqSAW+miV9xOep+lduGzmcNkUs9K3Y185yelQUZAQfPby7H8lnZF3Pb2Jjfcy5h3VWt
7LQpxVih1IPhgr57lmLPw60njrKkLQubHjBFGr95/tvmofgJRyHGrEgwhxNTG4CuawOVPEcVMC9O
EONzTuEDSresBY/UPcmXeliQhde4V9ng5yQVjZXUxahqgCsSY/GPyftqko4m1yQS5b3bOpK/6Gd2
tGZ115rYHJNnJBl6YTxqhuDoRaz50SkqMP2XSLGCZQVL34j8awMC7hSEsvKbDnD2VKhwTHJSjU5L
IQLhp+ol+7uK+RVWYQWqKXIHQZba3ws1hT8ZgYi/sOutag1Mley+GKxDmtFG0rvm3Cs4V/GKv2CE
rNgiidxHHEpWqScleDQ+xvxUn+TmNNEou6BTSH7aQmWoaiWoSXv2WHLG2/l1lFhelT04rwNGQaT4
dB+M9mCk3nlKjxfhIxMPUJTSM4aklQjfuWiMYyOCThorCNxah0xPbgFkbmDJoKGgXUscnLH0Qzrg
1hofwTUjem4ejnizcDrlG8+JqB4NSbO3gZLExbdI738inU4GVvYCK4MMGhSOj1SAtkPkWqxUnAcX
EZ+tb8xogKDNZbQt3OdHbw7IRdagelcJ74UymtxOsuyIW5ck1TaNKrs8LDvguAjJyWw/OuQ4odHF
JcJHFGWH3tezFgqKkNHhcA9ItdykWcJTEACZ73NSqEUr8j3HpY9jEY/nOLuR/H6nngohf81ulRsD
nEmkBXIt/vAZ3bFECCN4Efn/zDAkuyUlSQDpVPT3bdXosAnNED7JLqzhZDqD+lpPZjpc3G/Qoofu
1ENV0kvwvbFbmIgmZdGTQrTHWpolYCJiQcyhdQ8Q2S34z47W4/393RlIn4o5ctDR1mtY7uI+mCPJ
+eSwzenCrKa6hoFiTSKQBPsT29/SAbZg+Qw2iUG2Pl6uczfS2Pt+H9D7o1E5n2dlZ5eUWMQ0SiUV
oIouUvKLfhrIc5vC8N2AUZ4eFWxTGZnKK2khtfoIlW8lFKS8qHs2NtE7tV7EdmRSqpNMAzeSH5oG
WMUM1jYRW7SzNNPOmPs/RwKCoiosOTAEmOWzki3pboxbUMyrfWqk125zDI40C7tHLcQHHw2ZTZMr
N8ZF1WJqkL9Q5eLdc4rUpLZRJTfyzH+leSxW8ybnJJSOcQJ9cb6jrBDK15NtbYUESlOYqb9eN3up
LRMkCUyu4OfkbCpNf1Nf78Qn223KcxPgix+oWJuKTmLhrTWdq8TwIAme58CNZKyl1BB62M9p4taI
LEiOa7VXmMvpE4VYmOz+HWISEdXMRKox0N4mHL68KsiTnvJefQPAGu+5vxI6bfbXe7Ze/fu7F+gT
JaCh/1w78zwK6aEcjQMRCWoHK6eZu8haAqAijAtwDAALUeI1Oz11J835XcmlUt0CfqHhk/RV13gA
/02WjFmTGcXEAILDQyrIS763I/SoMjyCn2uwQ+dsoxjl3ibg2bJfAF2EmCPChP3e45NFCx3d8Qu4
XwC1MLgskD+oK2l8Rhw/B9jgFrDmuMsik//NZQk4FPho5WdahCY0bxDn3HVOfuAbatYigABIFWTg
aU/YoNvOxlHEOZCBaVvzq6fpweMYGVEA9arIz+34y4BvMZJqhdGVfflixwWThRbZ4FAHJm3rqzXZ
HfNbbMzooWXv0PciQhMSmeBwcQ/Jc8rWVH7NfXaqaQp4EgDK2+Dxj3ykjFujFa+2XRxX5079udcg
GXvj5Yhhfbbtb3RYlvHJDmDnPoiILJ/iYfJhX2L8dyWQytsbuB7YCUDfCvyfGUf3tohmQ37SwAh7
Qi136Jnm4o7yh1pi1qAT3jf6metgSW46L9fbP3T9IiblJ9kS0ey+uuCeVGK0I4DlhDLopD+s6m1J
kKQ84gE3SR0/2s46+b6ifto8QLzv0FW0OkvufVuLL0sS/YZKb7ZxUNNA17BdFEvTVJ2+0ItKD83p
D02dva6EsAnk7vCqYPergbdaAYtUEubY8ktufNLjiAvzD3Tia0ek2rHd3r07SkHVU8yPgsZZxsuL
tOQpS3WFADYtP7NTioAR/2nzZFC5XTMVzthD7j+soKMsO8mMNaP2o6X33HlvEyicmkl0QxFP9eMs
x52i0ta3hlnqm1OxJnAMvnSokr63iwBspIQyGxvBidNqJ9fAZVLJEyx2w6RI2gRs3dmOUjD639nN
jeg+AgrykYsJUoL+o+p1kzJp5Cmbf2XbP0Sa1q2yt5a/KYnDpcHPM0T0hdhGLohCz7EqBpbCPQC1
QGPs4QBeX2VPU1ZX5eTz9HCu/AJduMj6cCPc/MHvLAOzmm9dlWyMpYCI6HxGFhUys4O/VfayXD11
4nUdbNv6m83BD9idTbvuWa53QS2deylZiEa/QZ2hyxCFRs9dZAFE5z9ZriC6kmCU3+7UHiUQs5Az
ve+W1+D0QeELKvtsj5144/kW3cb5fM/E93ETaGUgLI4+ntgx1dEcOHgzmbLNStWCPiXiR9cJwMXN
aND+K67QIpTtJoL3DzCprGltkAXVg+5Y0LZqmxpSPH7a3UuX7kvqfzWnVsP5sK/sibmwF1dSz7Wh
+Ba/AmICy2DW8NmhfVJ4vbbXM5zyOQrG+tEBluE+AnssP9vV6SCg9/KhwYGSgPWSjQ+FQNpwazyW
C6I0vIPzO+skTVd7j6C913uo0bfjdyMQzjf5fqaKz2cxk0Dwtj2A6Vg7R0fFm3ePFQh/Jv+cSrW3
AjncXl79jEgbHliSw1CmdHDJAIbOGi1ox17PYz41BWUmFzOV0H88RzgCWiNaxvmimaCvMgVqHqVA
vkjvC5c2B/iOfHYVd6WW2jmSD4gPRfgq4HDzwNsPkX/RlpHJj2nRgQ12MVJujvUQhDdacHSp9c2j
CdB6ebD3ehAx+BaG3Zs+qNntQLiVHHq8RgfiUdBp5C2vTf7u1NaL6cL6bYRCA40CKI7+K0TOqbfo
BdetndbhC0xjouwoggjZ5AZRs9kz5T8JRGProLgaTr+IkV/FnkSHzWGVCh3wDhdL/mkhyYy9ufoh
kTKF5yLDR264d7O3cCqJMseXR50pnJZ4tbKn2Gjhn0RO4Twia+71N/RmhROAWSgKaLejng+NmdiU
OnICO2cCcB7O7FuO2MQiOtaCsrj9pYrOJES+4M66NdS/ds2ElMvL7X4Jre7hSkZLpUgq99VInteS
MumSN/PdIg/ViRWecUc2xRg/cazhr/0mWG/EQKDHbdMcbMLcOjl4UF2HiNxdoigY8q8UZAWR0AMv
cSw/LD6Ha/wpXGhSMT3Eyxtsy5+QJnSFBXz2ytJTMwMcwJkc/Mzc9nqcjwuikJUPjUYweuOiGrSX
oFj3NJHgWmC46UggHO9O4BvwCO0Z30Wz5YVR9c/XaSbeWoxi91dqByI3gZEwrZxi/2qABAV5GWH5
oyAGjknAyksx3/CgDG8AyGCC/YCN+E4RB2cal6dfvMEwtEkdD+qvXqWtvprJhUeLNyoEVFsD5/Ms
mWcW9YIfCJLDItn/KiSww0OKK47EUM1TDwprxI+TUlVK99YQMr+tWcGIxDmkJrVntkV3Vy4rqSFm
gZALK1ebtMbJcKm9VT3igzvLf4A+3UFCaJprto5GVWDe4WZWRcmBjqtsXu7G6K1zYkQs9RVPegbo
CybtDsUDYEzzse6/fXwh1RbPB18FtjgKhQDY74uSDMQAcFREpflxJjHCPgRIjIldcCm/tDu1fx/1
71q2T4KAQsy72WLrB29EiWzA+dN07bq/zCgGcGi8khgQGMKlP2z0gSZasjZhS8IV1cLjAa89yw3T
9NK55lGOaBhhP6X+840GxNCyUEKWZWJtw6GLvp8SSa3steeltY/fXY8Xd8T/AICDFtUTnvIs6UUU
98GAjwR6n8K8mNnOoVxt5GgQ55DAJBKT1Vbw+ZePpaoYRHNvqI8SMPVB3BBajriLcJG6NxnzMgjj
YnXzFt3ZU2SJ1js5dku0EkPSXKmqzGYrVhInaGiI9uttBpqNf5vBhlhd6dO3QhDTQLsayKCqFms0
8CFey5egArDtpWFp4hNpG1Lc9JhPvIxYJXEzdl69ugleZan7ntLPRs8OnZXEUdnbAaRJbOkW+bVa
fY+dCxFMD52RTbVKPt99MsDnq5yX7adgbr10i21UHteRRg9Ihaf7zupTHu/8v+TJ9prGRzkNsKh5
jArbiJnk6q+ljqrUJ7Xp2jlB6o0tx6BNY53tk3oVO7dxGpnirA9kNgoiNSqu79k8s3K9o8JN//GT
CDqH/rum9LZlnmyFO7+0Vy0SDe75ut4Y0SG43JBBsX/yGueZ6LHeVL/rByMtCu2vS5VZlGIE2HAh
0HfLdRuP56yBjZoxdExsbG/f2VblUPOMdnBdhP3aU+HohMr81qmTfSC1oqnVZNLlM+0u0f/mGh3/
OzvOPTwJWXqnhVuF5pO9bi1KgzK2d0EXG4tTJUpofKxC78DlWip6y6kTQa0Hcdww5nu6wmoA26cj
InD5ufa7xs0+4rZK3VSie/0P6e8XpU9BjQ184fVqcfeZlyj+SUjK+1aI6HgZoEM7Cx3znIbTcgDk
ziE+Y2u1T0BUn//h3pNrSYRjRoN02QNPUexuPKvhLcAyIzIRd5bQCk+ydLPRKRii/MABUbyLme1D
jWPZM9e6Xrk+zLcYqbk/3/izTpRQR0XxVsvmvoQ6eJJCFv8kf+iEG2pJ6s3vTKTQCD4sIGYUxN/s
aFdnTmGN//lbUCz3fPihPh/lkptUoccxYenAVmEOkGSR+YE4Jz5A9pKa10hxJJUBO0NavKqw85EE
mCl4ByPld47lgokJy2qaIeG3jjf3wEs5H4ZTEOnEb0SIYfaZO3t3EhP2XcRvrfa4kENTPxpoFDbL
T7mJ3ThoNTaWbqpSWPAPBkAs7Itwdy+7qN3YC4j6fmRuH8GjlukSgyQzVtuQqCNao/6DW7qRayKl
JMNyULVTIlBxE7iIrXxHidNViVMkh4ViXE9h5Hpx4DXhilsYHZmVWxssEj/NZhY+VG03WXXqYJ+e
pJTPXfN0BGgnBPvBgBgbst+Y4+ZI5Hy3jdan2x3mOF1BzrZC/5gYCDj6UiMrd5ZtD/WAoZ8IF3fX
9jR+0w1cjCtqHAK18XVY8/hOaJOeJ4Jc5OtCmr4DxCOkydh5LbMHxTCFumFcnlCIGL85uOfyhd0u
3qhSiM8NBLSXlwLJTJ/wd/Y7bLM6VblbojuLqrxatHxlXwFhq9E/CN7oAm5AfRPBXs2pitKpkpIu
E/NfbjkTMFpSIFcYT3MIe+kcY4IJzt9kAbZnNpBq9Mw7a3CxMHjpWvD0Nha64gqGNXS7Di3Mb5fQ
GL/2TB3LX52b1QLRbKZaipdZT6EZZF5Eavi0M29vjzIsP+8Xntt3X0yISP5RrOhtt7SqKBvfFajj
s72h9Ga8fJWNofgIQwa7aquRfoS8wdXLRYv+FUIdpte9o2vF4pwYKANFofeqKRhHsxUA9gGYMdwi
sZh6Ac7AlmpdaoZCdyg/cG7wUb67V/3beV+F84BIKF4JQCYYtuHypLOI93Btha0Ngp2/4hsMt80T
8YJq+FN3xahtA4X5doAWp7Z3ijAHZL5y+ErovYfOkRKJksVNhXF6UqCoxHUH4u4YpTBMebN35q8T
PKaVNl/CCRsRFGsT4AOG2JknvNSOlESx9PVmg2TfoZN3yoZjsZ0jqui0IAZ0bICEgUK6Kr8L2EVt
wj82FTcgMaScEwZJpAjZBdQMPUnxkNlONJ/Lg0eZRjSODypqlw+WYLNCCn5AOSh4AV+jRNZ3Osza
EHhqqWcQeE3twL+DN2YeswI+V6rqzARqbo6pyRDQVBTTGPGjX8Dy7BkeepGHk7gAhHAxtq/qvzlD
LvUiwb0m+wZJrj4b9TntXTUVXij6Ae99qEEwc+Pp4Q5+u+57lScqFu+MStZzA9+JgT1o1DzuJU2I
+uGhXUo82cpG5NxgjZCEkwqqLg400+V01yq907Oxsa2HOKl9hBLJHSjdfToOz9oXRMSlxxTL8mYj
lxVjJlXyIcrBH+K69SYnGBfGvp7a6UhKmRZYx6qIdtzx9fHyJ55YMAev8oXITeXLyQ32OIKQuVGE
rlBoPM5bWw25MaPQjzYyeMs95ZPRaRcY8sVwke4YD2fyoZqMugGiCE3wnBc1iKKYa0vziJys/Gh6
fhnQQBwpRrr/+OBYNZ6Lg6CQxPIAxEPrlyWdT3jmMLz6vqKR2Y4F2Nz6S1p1ScHS75rPv349z0Qd
3RUOpiKC5A8yzRjWb17j1BioFpqU9hgE8Fo2vF0UDHoArFOhhZxWLQ0+pMNAgj5ZmkQPhsZpacRC
4cTZn7hZFsaxBWkwdn37nIas7XPTcKQHUyaIu+hogz7aYGcpJuIhM+rGIQUvovRcBm3/5Aw+qCxN
EgNA2WiT7kSHXtkV1B4ViGkS4PNhECX6tp7lbsoYksPqU/X2nqZnKUtr9zt2p6+PqHc+J9fOFuDT
Xa3rCNvfRhLRZ1MsRAyMs1vZ39+CLd82RiUInp7uGGgt6wmvQNC26jPvIySHR2WnqFI7w+NgS5ho
xTqWpDRTKwlzljJwJikHXcI1vxj1cndFQBLqnN/DspdFKvzgdPpUcY9VLWmLK+yudLk4y5pXayLV
RqZVaNnL1IOZz2sWeJelu0PbTKgKZ5LT3wzLE2nqOKi2MLM3AXLVZGEogfKXld5ByCPR4yFNvCiR
enTmRbaZFOrDDlMhUliLVqrS1tRC60Kx8OWLISy5111Dfq6yyjlCsXG+FgTu1GFeOCJPrrcAaRxX
DNtPxHRGOWv6ygeidDE5Sv7stdFXlcxQUfyEpMIu+C+dHjmcX9O1tcKYZubTcdcNo8tLlthq3MBa
MsQAsIFbAwzELjEup2AVPeRGqn9WuDIyjI+cNRWBAS3sm7Fl00l4BB/SJR2XH/Kn33H70UBZ1Tr+
gAO8ZUEUo2Y30omJGjRiLdPh/I/0DOcGX32VX4KazqRWqU0I2BeXeRma/Mu95VnGn6ottZGQUZ3r
Mu6GBmK180T9V61g/Qt47/SQbljso4dUtvQjjkBqwA0e9RYq33eo7GLU7pbZ/nCDWlKcFlwnCHdz
HLJvG7Dku9QqkhrY1zfrbBiC5wv/nDOR1X+2h6Ym8EQZi95l8+hH/fYblJX+41I6p7I9w8D9KDrI
k3TpTFn6N1XdQ6LeUjiUEYx+dqCq+zSIOx1MQrLBDD2gq/KSyiAEjN6fr3/Kam87pPe5uY4tHSof
rxF7UspB6oujKyXVWVXxLfrQ+4AHNOtw/OrVg5OKiwSu5eFmXYSA44b1lHz7oOLMFjhutV+AKfUS
HMlv5oIwaKBrMzA3D/VmoqxAW4aXrQ8pU/jBfgxSz0Uwvb6b13b5Q3NgUp1vuKMglpfKjCqm3aLz
B/6N8DHan4XdP4R7cKWLFQrKVBKGZyUm9J9uyQOUiYb8OYUoFkblxJPBrKFqguwrhQOii2MFLO0h
CzCGTXY+ajZto+rGBECpOmBgudoeDNpT0DCasOwnXghay6Ee+pOjjLXTQNj/Qt6TmZ+pv2bqi9qn
24SHX5cRWQyw0pYn/3/SdvgXXsDBHS2orMjhaHrWZTuz5ujTCq7R4OV1oHig05bMA96z5hGGE1Yj
jYrlv4GxfMXV4tS1m3S7WVQy9Dr9JdH5VX/4IUhNIs25VF6nkI1wjzPkNRlAsKHFRw5H23jUc7UI
SHJs2Ys7GJ/hoqWXGrxbPZYHLuh7ljy0GPMOziEk9uQcrvOWPQqjriF9Rj4PDP2Cf84OsVXaffgI
ftmhUUVohI/p34R3C1b2jOsIYTsJHg1HPDSqqtxghDre0/deTq8dj4gXdknp5zfRlQHTeTMAS8l6
KcM6WN6eJUyLJ/gB1eoYaffHcwTQgeH1JqU39h9BS7PIA/ms+ybGG5825TE1Yw5sOEI6TwTsQflK
CjQWdFh3w9Y+Us6JGAa8a/njTuOGjm/B18evCE14OES5Qmcju5v3rjc1T6ZbRCc3GKyzH6jP5QHp
0+diUh0uiDLPgngQHcaIZyVD4gO8Mm7lvPzMJ9BY6jqDlSLB70hiw55KdEsYZEiPI2xyqnw6jiAr
mjqkGH8LvjFUHjnoa0Miw49OhFo8RPBQYDl1NONkTC9CHUTncuKBY06PxmXAgDg0aaXZPmc4smda
fMUWhY9LSbhVoGoHieN57bPp/jQbiW0h/18zc6rWbqQLm7wylYg2fKlLFVMbCoLYQKisz5AHCpq2
NL5zHqMxJaavisFbROR7QGnSb/JswctqEcfz0tA55cb3o4dCWpRNscbyqkDMcHlO1nr9AEIZavPw
WAEWItwDbbfBLX1dlyyWfxj4e/mW9i9w1gPFeHVmGU1p9PBoE+6XwFLmMPZSSNScheGHNt56Mblo
l/yPoYT+kDcQFBycgY8pFj8shM/XvTWi1Q1puR/0Br1cA1dXR0JmEX3wM+3J8GzzSyJ3GWWvvlNE
AWZjQNvE/rTyuSqmlyZC822syi4HiuRCQC9QtZsN9SCf6Whriwz3iIMtvhGndkdTxfokKNhv4ulT
0i6QETHVNcYiUrj0fVjDqi1QlPeYCXsIN/N/9YDkYzHmwQVlsQcOZjP1PvjBXNN3W35LrIIjUjZi
TzLcVwwWpwh16dd43QTbCAdqzg3QwWptygcNoNtd4rJmKIDy5TSYl3wILM0Xh6R3zBpCoGNpGOc5
1bjmXlvdnjYu4IpIZeGKEo4L/YcXj2ZawhU5zIyB6LnYxIZl7Bm9kRTBSA3ngH+1WeFVBa0eww6f
6AYzdw73wtglxAw4JDbag2TW36bfTes5UmV5m3AulhYITOrS2SlX40Pf0j5j+ijlEPz32Z36Icg+
HoVfqb0sM+wLTXdzrRPTuiXYagIwqDRBe+1lbjMcNa+8CI1jdmGxvejU40ZqA76/TOAW8HEHa46W
zpIwrgNU2ZD5pjOsQH9WVSd81PG5q/EtAATpSi9XiCR/g7bBI5fiNeODoQivwR98sccto+JXGbsz
GgTWnohxaDp/5rjOs8Cr9Q2La0DvA7RfHGgrkw2+N6BFnK1qonrL0Y0qgbvdACirtE5iZfU1O4ge
TnuQBj6/XW6U3A9pyHCKtHnoU8bCopqC035XdKyPOIErvN8X2yJg3kV50xotDfMb54OBEgwE9THp
2sMevz0m7xegprpEloicg7q3kr9MhFSnCiHhPO0WWDf1WUpkiaXB2QH/zlrEAo9RPCTBMnUTBXBe
4XhnZPXvtaKZqEpvoh0ZdGVI8nnKaFeiz6Gw1NC51VGI9afGdyopaxv/aTPGhQYnnnx96uVHF9rF
wIe46es2cBMbhEhP/+14vzDH5+Z0JXYy12DgzgSscApXGl0dZescl5x9tlm2HPgp1Bx3VhTHmKet
nNExHc4xOdRsg5lwungpZ3Q2ElYKMGXqmcUzJoSN3nyDKWKKTN/g6cqDSM826ZenKNCm6Nop17uv
GAUHRU0L9FAv4ZaMh6uPpvTzYBQnYdK++4T4LRGbpvbooDwEnzIM3V+3W0LZ48Cin1qfjsV6bpIc
fUy+Oyr//KQuspDxeKDOjxqhy61TtRVQWdut6iuUhQtXpRxU+HjGf736tjiLu2KLQUUI3DIBJQAt
A3fFSu8g5EZBz67qz4ZBBRXHzJmu50JEI/xkQYa178VEMdas2nEb8L2vdSViDS9SRmCrqXWToL5g
iJUJeyGVhLc6EfknrjCDFlXPcJJMLCFfgHYhabize0i4pB3qnVWFOCyC+A1GeRa3QO/P0xzWTPuo
ij28M00emefCTU8dq9plMnEy52NkGWgLt/nRI//zIDrW5ydvDMBvNjXIEJC72gv2AnZoa5T+eSi9
f7AAFqWYeuc+9z8hELdXnfTeSFG0qrgezL9MNQvseyObKmAb1UfGlczHUbl2inipnVckPg/0Z1Mu
g/mmLWvE8elVWJ2mhfPdBmT4DrJRoSvet2NNVx2XhSpLwnUtA88YWsWjvphEORHwrygIUBGmIXEM
z58Odb0hcmVGGMQbYyAgU3O7UuhDnrkuNaGtW8K6R9PAUOj6WppI6vqr/A9QVMZsKlmW+x8N7xcR
wuttQS42m+V5vnG3+XSon6HavnlBZOdh5erxF4sZK8JSD87ScvPb2muu2Kts+zHh+XkQsRNtzT/n
Ixh8cnEDiGQvaZL15CrqckxjLofw6WrbKWj0u4yJJlOPWTfF0W2it3xQs9cER5sPSU1wnuM776GR
qiaG6rRvL+hnVeIsaU+TxlIpv2qfK9jsRUn0RHej7BDX0/BwGbIICMKaxviUCcBhIUxHBTbvH6pn
xqiAs52i+WhGBHTd28B7LWIgnBCvF7nbbsZEpMMb8UmLS1AX4vON52BhiYWrm4heTUfENgh3Cl9k
e1DGMaOBf9/FGp5zftkUbKT+dN/mqesV4spWUs5S7ESKiThS+VoqQzvpb/8d1DV2e/92FgjMWg1D
yC1mYLUxRKb65fEanHBo3AOx30A3I8OA0FSxQeKDys47+bH10CJeyyR+3pnChkIaRG5y712+Sipz
cMn9Qtbj3p4JbqnGFqNUNkT72J2QmdB6vnK/i/dmsS8YwLSTVxtD06AxZHGB0/c8w4KcTOWbGuKQ
yghqg1Pc3vnwPp+Ckh6RRFXOa3EoS1gsyQhO4t6BgKuukAoikzrRhCxsfCgkXNGQgU18ytJGrY5f
odow3N6w72raXDuNYKloOBnOMkiDbAZazJnLIgn8MqiDhHIBbGIgQrb1zatdyAoIgjaIFO7YH4td
CTpbviYqKuGyr3ny7cLFkpKfxu2azbc0vsePa7NP1noHDEGm9UMDLsAQGopG0mfVXSDIHaBjYMwy
x3T7W5dAMmHt8X1XXHJxr2iYa0HjtP2r1Ps1cIgJgZziagJgTUcVG7akvhPAODIxCtz3OsDjIjWl
qujibyj4ynabeK4dkIv4dI6W6iC6vjp8bF4O+5bhv2Qpz3XLrXoEao/5xMQsNuZhU/MIzfhz38ZF
Y4un5Qt1ITWUvUZ/N8GPHQEczPlbb10q5j4WJQwmKqecwsPNVmoVtKZG/UxBNsZZGksO7XqjYLuW
2/ckyxQldmJ4jjD7s5zY3oH2NnJTAOJBVTfVwHMVjoJed3SF85Wjml8O9ZrhapfXYnHLnaTTf+vv
elIR8sAIWUrx5jsslH38wGwdGjcUexe7R1w187WVRoj+aiA6yL+1NdM0NWsRYACS4nCfH5kKGF04
9Afn8xrWpXqtYul0QyW1/uEocy+MJG28LzvQnjc0A2OdDuwFdroV5obZJho9XvzUkL4w+FT52beB
fseuSECp3DE0+RtApCneDLARSJBrluVwx0jGebvpxNDA97vuY1cMarbCAiXxoYpcoQ5YCGg4M/ni
SBcQoNQ/h0LxLRqSN7FGcqH8zcpxBM0JooARRFMS9RCsHK77GAFDrff+u1nA5VN3Kgqxv+vjsJcS
xzUDkeIkeOtK91ZuZgYDH760Gb6xcd5o5X+mTu2ZKEl33CJrE8r4JJH6YkDPJy8wWqrnEygIYS6+
6OTfp8RJjJQEzrLJOkwTjxjykYRezD4sZOVTcjtpUCAJ30qyk/Oy9GhIQA6YB8Lad+wOSJ8J1jXs
+vAgJBo+oYr510QVOIrSbMGFDahIT/dxD5WmE95J8Z3bndte5/3n69L6epyG/Xb33BS5ULb2898p
MhmZsKlGumkZ6BeEJcmWWHTDhXe3zlqeO78TATtFfKpJUKHlHoPgrGEE41liZEQgT1AA+kff4ab7
Vb3RT65HUXczznXyi9iYWYOcTz1pljLsB9CiMttDZCZnToEC2j4pRRL0MP+kXmtWM2RfSRmU25Lj
yPoLM8x1vGcLK6yBRtwH7aO9UiXQecUQ65haBldSQDM55q56iRQFBTIJPIwXczDoOcImqxO7pOMF
eOEUHW4i1EajUylb/FiiHod1mVKVjyJaQnJsOtVsaIigT/404Nruaywgg5g/FAl9KJGuMqQ5tNVq
CpO+TvAzY9lxZa1IL/ei22YOnEW39TFeU9HuB051y2/YdCVcPsxCCS1dD8C4kIcdJ/XjbDIbLAT5
ni+ov1vtMQOJsPgqUia71R2pBl8TbB81nU2+ai7zOW5dlea6+azFZKO9nDNRMut6vQEfSbaAQT5A
F687euBWGrM6qOkdu3EtajeF6uFWZxMDqm/ymYSJzcArjJCKxqvNWRadp/bJlDykvWD4KsARKhz8
ievr1TVVNEJ27Nkmg1bW46p6Hv1TzCwr2wfb8/emBBUHjjoAiYCZ01gE8cjw6Cy+R+ehQR97ebaB
tH37a24YqHR0Wrgk2ZBLFKebhLLI29AOpC37sOVV8SS3wJGg/383JXhY8+Vd/SEPXrxaOGWjPuvG
S+U6Gr7s87hywxIi3wgobUwlspg5SmiPrjoZCE/4Xbpqv13HVZ923zlaEZtsAw37vyqgAD9CTwrM
G3luXhtGxQT+q5iNsNqL/VEnYV3+0cBK3Ciu2rvZemLD7fgBbDsimeu7VWt4cMz319sIvaaA+Qks
uS4OA0OVrwglIzO5zUC7+FOI25DnH5Tmkho2tb/tXod6sSvs0BG+rGCx8vx5CPndV547YfGTtAd4
1+WVX69kT9YMebrzwdgv6nCdULEvviR+CmJ0BezyPlEiS7Z37cOalTS0YrZgx1nKymHqPQhIvX8O
zS+4pTq2wWVk1OrHD8dx4MRJgKnJ5GkNKkIV30R0SoS+dZIkyQ0ikt8M69q9MExy6UJwqxvieTEZ
RkLz2uZsSuMmEo05J8xZfqq59AbHo7tPCgMlW0QUbHLEoh1athJtznZ+3fS9XZTdvVWfS8dCS3sj
5sCjWq3Xm1JdvJbe8VajjVqrKS3qXbfSyNacm7klw3tHnKozhg540WDAOoHQI1fDPEQb96V2Ygbs
TPLNB+ppzKIsduqWusazYN7t7SZ7DFdpmHOCyXswXMtMjUlrBKfH3YhT6FtmJuJSOjBbl7LAYylj
uptHa5uy3idiRgYYd4agedzUqIRx4GCsO2Z9F7DL8YpprKehmjeU6yNoQ1dekZ5Sa01uqjTaNQ4m
jGhG1Fz/S5B+mkvVU27stVAusYcOKGWNAaTUHY6G2OYWuOgsQLsi7zF2JB0ZuvaUldlmeomAjb58
1NsiEcDuBOM9H+bjWdUa/eg2dVNvDTLO5yZJzbOg2janP2Q6IBCorvJz1pJm7nSPQUU8BKmKEEcO
TtoMKoHPA2v6E8P1QFfp81bsdwL2rvbTw8+UlNv/Rj4COsnj4mKXXJQnqQEWiZ0T/Es8yGNVdB4h
T7yRn4QobYPouzTJ0lwkxL475go1ah9f48QOv1gNho+SZrXFfIQJA8I2blBFVktvhwec08At/79D
3KXBMZ+DEl0MJ3A/Wy/4pmqwR2YRkwjeb09yOyDSVhSqjAzycMbduD51yAzm35CXPvMw/Qgw4zqS
HZVtT7K5CD3ztElGnXU+3F7BN+tz1jYx1KgRd8H2tVyQLM0+EluWK5HtPzcsaJJRjj/me7Am/Q/I
Sl3tAv+GCPfaZK6lbt5XUrTPxPIGgmNT/J1Dr6cPK8uzypFABC5gEE81O2hd0R4binZ6efrSiUbH
OMKYhax5xZYj2XTJsqfljQw/f8TfRQzxMr7sKkq/hlTHH+uCx0wlI5CTFjkGfTbt6Sk202Ds7ZiZ
2s0GWmwlZCecYg9jB9te3LdzxbNOX3RWjBzzdtPvZaIG0nHxvlmcKlAzzJvHI2S66osNVIDRX2u5
vgEaTGorw/YcBgZN7FLqVZhA1W8t+s2TabEnR73e0aXTf3mEF02NSkGyHc1Aas92zyyh4EvyMyHS
KE/JDsTrvaGguec1vQCVK7Uoda2FwvXrz4Ku8mnZXHvhd++lsVkK8n6KvgbiO6HrYJgISwwLIJnc
gkHknCbsLBMZjxWN6pTePp5IKjZ9gFgpzkaJVGVAGoJSb0CrngwmOE5hXxxCEIU7n6FN74Bm0eDH
ziGo5R/khI81uW/2zPGcWQU43tHW6Tsq4A40YGXkkAyiY56qECFvirAQAiSwejnqYNw1csTLf+tj
LXvFxM1d1ZmpYwlEyBh3xcOHbfyoe9nIewdgnKJB9q+xgLryTmgsTLKGzDD69PsZQT7RphVqecAN
3QC+wXVFDfbpkw3RkHiDqY0/p/HNBDdKeEuS1aqZJSMYJk8/F9bJ2tonZeCMH7Ca5qIUBwJJrVN5
9SoVEKqHLcjSpbmeL2lGqQUYaV0xcZJU/BBQ/nKlvPE421auw9rkmY0PIwHEazW16PvJX5dN+HXT
xmURySNL/XGw2am82dvOFxCnKsa4ZoP4zc3oe1bauLIkc9c7WwZyoL3DI8gomMqnf+1r2cWxYBvP
84pK3LmEVYNwnbleAYzQ7qiwPMtnKpUH5kGnFy4HscruDusVuBasItSdE5jhZVI4iZybZAkCNB9i
cckCxQzSdt+FokCltBc1g1PCSMmi37Wf9S0rZKYa7lWoDTR+8/HDOiTEIyPRgJ5mxoz/emfFoHyv
Wpfm/u+yn/2YF7rsOiUf+xz9hyqQZGDmDOfPm+aL6Gs1ifoQJfFU9oKi+RwGVWzLnBNhbVGDDLmV
nPEnj7yw6wk3kmzOlhIthxfSV+Dv4u6QHZrLBHTmcXJ/rxRnOIp5gqnsFkjRZkcQ9L3xUYtRO513
+7Odoacdc+jc/cn/DIK/pCk7QE+d19Zx82+DU6E59yGm5cE6yz1tPrKICQlaUHG0MPHZwEDlGD7C
Je5ZgiQU21e1wumZP7gcB3qTKAXN8P00V4Hu9FBYpzsRcB4f1T+CfWeOeOh0csYN2MxL98lWIG+i
D3/lLJkLxOY+y0ilR0JNPBIUACgsBNHNrqWy7NqWJhJZfo0E1oDUuGCPao66cCw4V+Rydbo7auka
6njcB2v4/jJ9t4m/H6ntXDojGfeysgY0D7aooW4lvh1BO29Fis4OC+WaO02iZr5P0HbcSC8lEXAH
DQZl5NE9NYptxlJ/rj4NQWmLxFChq4Bq8rLeRs8yOxg9Ee4CF2Y/1kLTO4HeUsOZlgwwDeJ9jtRm
azahGEQVB86us5PAeMAmfWV/GcCXBMgjpSnUppjf3taOvWrjOHdm9S5+1eGu7t3p6FPpRduVOWDp
yziOFtSHIj22M0fW913JxhY0ytGd6mC/8dfSS3hTO8Fd8DQoO0TVUcrzYMB8uUaArUedemj+L94R
KB7gmkCPghMQ0aNjk4tUkSFyx5Ww3RSVvw/bfXncEAYrAoXQRTVC9e1AbgLdwkiLZMQcbAtpbm1P
nAGpHSjUnS+t3pEPnZjDAASdRy1jpagGlFWFvYT01kxW7fOEk5utuYpvm66BKNNx62QV3/CSaaWg
MSDVkVaZsLtNDZl1B6vWxBiiplNuMpmGMNIjpQzZ3m3oBzYTON8iDrCijbFnIDYPsSYxKBLa7djT
kuLv/t586TT1Hx5cKzGPhRihBYFFEjCROBOB09Yj0nVLsFHKjEcGSvYo1loZOhyEFQZkO7aFqNnF
w2K9yyVQT1h0WQnRexbaTog7EmXFXXdSfHmnSaA7I+orFFfklm1GS/cW+eN6/pS5vU+LtJHd3mii
3Tbl47vULNyVeIik7dwH6T6DksnTcjnKukgNY7bHEfQrpvF/xmlg9/xcQcyQQHlPyltNWm4gk1jK
CC6ua0egzaLyoLnHmenNEfQMf2OXKLQIZyLwwdaWnBYpktnDJTRvZYkqwgM+7/U3cjexHxJGA/jC
k3uEzRzfXje4MDGjeY8IeefcGkDEXtP3qZIHJNtsLQX244eqCRD+UvW1xRcQw/7NDd5WeWrMgEVz
cfe3ThwOHfMnBhNoCGItG/Wy8bPL9Nxb3QlR6/AVOfcgzGYiF0YqZNec1e/ShBWBMywx8Y2wohA4
8gbnq4XtuqFufjXhJLGRH1b2yYSPC0rZU/G/SHASqy2zBXy99yVVm1IqrwJHS/YAbE/Q3QP4I6tj
np1g6iOEwGgXW3XLpEloanNuxZVGqaEBInGNL7Xd1WjtSTvx1pw7PvnGrcKffhC83LqNZfT43GQg
jzVR38idQWqGLQVfHVsR1TQ8HGIR1r92sr2wO3eUqYC/SG3+3SdMxUd6qG7D4awrO56jj0T2QD6h
65DUGGnb45GMcLIPjDwVSDPIGgMiJ3+D5mOBq8nirHvEIPFq32aMYez9WLnmtyfmhCdPFrxe5n/V
heFDyDMZHQHt/iXzuZ7+m47L2H1r0mqDKv6iP5ARLS9TSTTGsxjX/fonRhyQr0PLjiAIVJbeJe31
MAZUqPB3+WBqEcGXdl9xUgp6l8qv200XhLpR0ymeydklD4jLkUgMZVNAO/Zh+DcBLbc9SZntzE6h
2Lf0cEF+hu/gxBezWOnHUOD6yfJZK3eSqQ3IFtOcKSAwDyFBWH+jY6sxxe0gmYXiJs5AdJi2ZwN1
2BvMobAplOhwfhp+uxkBHgTQ7IcKwnOunHT9aA/AOOSFdeNjsdJcMchFmL54ePXxPMNjBeDf90Q/
Z++/ysu25AhJqtwlfGQOBnCnj8F6LicBVwne8GOUeQNZlMZZhmoMASmLBuL1XUWroi1ehZIOLu32
NJx+njzlH5OUEfG7ZqLluxFgMmrZ+FX6jCG2MjSRa6x5evQW9M3P+JXAXWHtk/EB+601tGHYX1eo
SwEKDwp3nky9z93cCPvGRs2Y4Is90jANFCkXBiHSXUadmPlFGusjW+GklZw/8QETxS1fc/HDOo55
LfsY8JJbIKAg8sOC3KCBykQmHV1/o2PX0PVszNzw8Fmvs5HiG/eao2fhcfhUAjXNvWYLCFt5GQ7E
Mbtx5R5bI20xLPOcKWGE1wNuadfO+msQGU8kMMISJcHNKDfzpemmZVNn/akc+t68N5a0ixnQt7e2
nhQMedmpDticuyzdXqRpsNu2PYIzTf/x5aysJ7sggMZDPlVdztK072YOMuMvY0Onfohey9f8LWqw
WU1MQoQd4cpLTqvIDAs3fB+JpnG2qKeQl83/ZO9/RsEDMxaWYnsID8nBupQqYqGy5RqONbMYmQ5D
ytTAyuEwWN6FdGWIOPbXqcjyl7yTvCAy4vdEkDSVdZ9COgmm+7fh5TgbilwzhREnMyoBBCkqyIaX
b8v6GjiYQURM3WNTLgs/lBhN6ZTV/Y3skuP49EYkPdT3T6+cM1RVxydli04kC6kVY/V7O7ubQtBo
jgoVMxg/6fha3QkUat4v3DIPpKxSaS5ye0lheSTOdoGSJQg19yQzhrdfipQ55eDAKWWgTAYQXjrY
38jWPDWAnXMDyis9IUNeN2Qz2CKi/O8qvzyqdn0ixqkChgk5SggPtp22HEIXlqzyk8PPMaqq3bS8
O6Ai9p5tCz/LS8bW2oVpBo7PH9J8h1LpFsb/muEbCB3YkRaWopk7ItQh6ubbKhQhlQu4MkRoPMhU
v2yif+3LPbUE0IvXKdVxiMkjgXFXf9dympnWZe2kIV2sAAh/qYe9heVa771qn0+GrTSveUSrYzQz
4xd8VELhQELpy2Onm9xTHzCRBtieGYZ1zYvxJwlhininJukW7v6fsS73at8JDXiMNRaRjMQnVONk
za0xnNs8DvM02hOdKBgbyh23DvDQdsfkzUp+N8WH1QL01o2uf+O0VjVASblr8nfuVfsAFyJw0hRa
WYF2Ki+7IBZAyBEe+ZBzHxBbCPtPKGa5usnpoVlyKowiJZS2IFmmaYI7H1/j5Dth/JgWF03O3FqL
ivNlZaNwKkqxdyI3sx9+AgRSzfq5XlKx1ZeKxnQiQ3PAT1dYh7B4xYybeQ5fIMnUO5UpnnfesSWE
qdYTXQBNogX9MtqqHCOXWl6jg0QxlZBfwxRE36144FtiCK4tMgzbz/C1fjvBW+hheQ2Ic5pVre1j
YpNzq/O5iRjgKgSGtM7ex6k9LK7b5TJJu1CPGEQEfFb8333D8ZF6jCEkyh4iTVe2O192Q5p453wy
V/lLM2umH162w4E73J6BhGhZS/X1QBS+0C5v4CmhM2J/wKgugptuGKnwtDqwQRtfgjYPhHESHjHx
xn6h9VXXI94gL5ezskI72kmy51exDIDmH8Up6Do6091g6IBJhTtZsIjjQJXAUc1w6FsAyvqISfwT
hyWbYDPqeJz3VBCavypDCwas0y2bjY6M0Q5xYSmKu/3VzRMLtwvjt7USQnaxnUzlJxNV3l3ZwcIE
DrKftEdu7wsHtBIcyuT+KX9GoVb0CSs5h+3gxBj1PdDgvu9mNAHJ+V/R+2NmQ3hyTtJuYakke0/i
5j3bcRd6W2vCMztNObJ7VR9gdR9vlRgzkTRlSyyLBIFkxQ0u3deFOjDyPR8VD29RirAfbQq/dEqr
mNd2u0moWgHlQT9s2muIoizyvUiy5HSfaAEkWn+3R8sWo9n+fBvYOMh3pDJNjlNlFLRIzYO107j7
p9UbJG6/lM7HgaYWqA1vXVtc+xsrq5VH6sTZ+p/5hmNsuNLg7OvyDw+iJ4Jy6N7fLMPnngksu9qG
13bfo9DSezMT3U3MiDPyRFEq0sKAUcUc5AbqUtfY8uz3WLSJt9nWKCfN9QhE5HIxxKHCW0Pu0EUv
Sr1Ga1y2k9prnuACdQrSgex6onszja51+zzKXGKyaHBRtcYX+cU0pwXTTxGoa62BwNYwRDImt1nh
fz5zsMY0SkZLdgLJs0c7EuFRjphiEkiVCdO+ZJ/CUFaFfl0/wqKUQAMNWDvi1Hh+eL0aFr7k1g8x
iJ87y1ZsPOeV8q+v7+uwRJNIs9FQ30/DjA5GMpcxDAdt4fcnWO9OhqLtMQolvg31vzeepF+26Szc
e9KGurnfGSJF5VJ5t8/na3MUOoRfKaISOvGqvgy96ytIGTOpR0GOEkDmf2v3MrBF/SheUmVz+WMx
fGmVuJ8DXhzmdf6PbJpfifkm/yQcYGOuWMKLCRXgF/pa5qQ/SHUGRBrLux67UNCxsip3ovAf9ZK8
UCwvgd3odT2JR6CZQoo6uh+atseqaIq90CgNbMhUpQsuYbjiujaxdL8HEC4P4mnBZfJCd2d4+/a9
T00gmblWgU3XaP65ZeVmOkue/Ue0719extOuqJVcpMWbpax+8ZXq9ufDA6OnOGAe5/x+4bgHp76z
nHr9Txf4ihAGU64nQYpxUP+tlkZPlpvovxQ47rMBNHdobJeOHfRaJmJpB4XuvpaW7viwwCxY+ruu
k4geSy9xZbjpTUWBBgk6eGx/aaQo4zsjOlFlOW67lqVlIYdqTEdmkmYSAXKFz8lMSQ44K+X0aHL4
AdQ7WEEkvRNkNnyBxqqZWg/6gw0PhjStfZ5YNhxdcWqp1SMsYWpsEgUpuW9qtD7yuAAD18i13qOb
k4bIVnpS3nDIexc6TayvXZndyscfxeiryjtZgsmKt6MyHHqjGhH8F9xCPnPzHIv78tDdFlO6M720
GT1b+k/C5gJ9ojTDucNjf0wzeJzVreiUfbb/jH0BPg+TuD7INNF3vsyvVfZAoc/UblJPXulD5hjx
YUJ82Wa2uiFaboc4wCOB0eA7ORTAZPUOlh0EZVmQUQlmsFUJy+qwedifmUzXNoVtSXx/s7MFi9po
Y1zS0XF6wh/csP8CJjAyHCBE+FGiMenjjHuANDsF6edCguqI3/u/vQxGIR4E9aceFsbt/GKdOYyQ
eOmjk1zgx8fzTXoPaTwjkwxhU1IKGdiRLQq+Bw4wB8EXPDs5byqEiSg0yYMV/avLZOH1qyWyzzHB
Afnz0HlIcWbFnzYYJbmIPSY0QgXj+qAxqDVq7qAWGy84jPL2Ko0dDqldLVyF5I1EUdEkg5UzCar2
/Ka2P+BJSmhMPHPZ1MgqqmUaIhjwMfnKMVsGN2ThwixHVCd/0/9I/ucR1RP1kxw31XThdAk58x/F
bw0EPecy8Pnugee8nzbTfT8IB5xYa5cPxr36hx7FQvXxTQkijeg/hTKSRHr1rRK8ivbw38rlZJO8
XezrxYImLHn6QyxQR9QpJuULCxgdfmZdBm37kPgtWX5lMUCyymxoc2Ib1Lg3uSSZTuGCkv2I3UYu
y2UOSM55bjwRJ8XNdZS1Eb3YvYt4Pp3N/qkoIsemqMZb1VRmAhdiCy1l8efbtVEOKULGCgOsJpeU
01TyDBKu5dgagpAZWT6bnQX98nLoh7tj9EccVB6DFz2B+URq8+wZ7dJC2XkVr+gfivStk5Ipn+Pc
BHHyoR1tCyGTZ4knPeJYxnYBhVUPZ0cjWXlEP46Q9cgFVEsV+uDPcbS4piwohLmdmDw3KgMCgc60
PvwEvC2IdNii9SHEU3BlWmft0KnNMp5CaT15KocxSiQd+Fm+vhnAuW4HR6EY3pEYvCXQiNCXIUcm
6BupnkBvTxdFQ8FdQ8ZigQkpp5/mFx3cHD5tV9je5BWkoJ+GUyXusCCRdVm6rYrWPCBnh16zUQGx
AKT4L3Dw3QjSTEqGFLt/W0FvVI8Hn1MTS5c1h41+TFy2QohhcmOGoH3hQnTctKjyzBg7UjIto5ZY
xfwDu7gq5zJbRpi9ehEqhNTdqv2E/OGT0taGsmjn5pEm7f173lLvPWf9gPlK3whZSvAXm3e+xznf
zYmb5sXYfGMxxBkA+lLUsbSo1NOdTvsJTh+QzBLCnkV1nnPop93N9Dcu0E9h6HzOrp9KV/I1IKeL
mOsoM1Z4m57q9vWdEJK9BDH2gBVtuuW/Fsf/GemGha0aXnAhzerp2GIbmDW7146z8ESrYzSAwQII
MP5AmDC7FUSxwekXbuG7fDmWYozO1IFIFwoCC1lfRyc0mg/wsSS+TvfPy8wzU9sFqy7WNGbTcQBD
J/B0x3xJsndnPb8YZgsJVuIUx5qbkkHXXP+d094grJUxihOVfKNYQfDAb62LbitRQHcAPZLsWZNk
ExmnYizWLL0mYgBgISYPGu6b0rMmUZYV/AZXWza1FpB7OgmKkSX/VFIYCeFZdRvr6iPRVz4ztAH4
wCopAWlZKqJtKZRSgJiqbeEidjXUrH3GcPnsakwYXp5rbnz3wGTlKqx7Wp0WD6qeYkY9jotSTY68
tV2v7Ro1yUDXLhzHpp9xTUxE2my5MDmXk8/4tdqj1mN1L7d8qrlePDlz5+oyQwVgSxK3JybN2iR7
N1RT8M2eaomkzbqUNScaBVOFev7JzRKWqlHjbb/C1QdnykLELfMwABQZO8m+2sLSnEQnaJmNKIzg
TXu8Aq1eCM52RHn+YSni/QvBrYArVzIDvm3ZxWsJ1SyCPJNx4cs0DbTD1oqpmJ5XyiFt1vQsuKPP
PN6XofxuzRXT2DebSbR35hjsJSJFjLJnt4odTRh0rPB5HAXJ1rpeshUeYBkazjcSH4LEihtnhBmZ
y3t1CsOz7BwH9uiv8w1UYW05EhLfKwaXl6eT3o7eMpqZkaqCHW/iiCOaoltz0SSkYiTRvyDLcdFC
f8Qr/Q7WqzCqJBBCSBAPMIr+27+0W79djyszJbaDbTWf0lH51wRxuo5KLgyPBBf0M5XjvmcPZLey
mlpPIlVQ1f/vGziNZaEWhgVV58sXU19P0r0Da1EbqTsuTJPqlbPXuzDXwIccU3rUglEapImWnDI0
WCvkc6I2NYmOTb6uaHzy/UBlQZTgUW6D0+uAZ/xpeMbaoEsBjmNnaIKYM791VpFgVKH5lhselEDQ
T0J9kEByGIW/NgtxJzW2sjeXf/GxxUYMw6FAeEpNy/VCdS8XXeVpCXLCbJlqIUCtO3iqhKep28Xp
6NgQAM+MXBKsEQ+i1VXJhnY7ZvYUp7MIygFRSTqhF1iAg0O9vzSp4GOiTC05W/Z8stxkzjQNIFWD
OiF3E7M4MjqsP2qpVbwxRTtWFVP5xLOpbUZnAxT0EnFd7uOe45uQqzIb/gfHGpO+WP8qnBZwjx8e
jQ5NOMtUdopfAyiDEn3ytjn8vr9bVh2p/zfsdBfb26Od54UnFwDaKVzvdpobu0CGmTfY3qWHyzX4
OczqJara0QCSZVrmiAEPww6cX3FnYShZeIw3kCYK9s2Rtr0nOTBShhJJ1NBU/A3wsUedV71o5Qyc
fl9munEWevY2cls6xP3DzKopVLBtiZUAjDrTvZuPpBfckx3Xvoi4Zt5ALVciBuh/ZZlJ+Yk9ytJy
y9EARiFo/Cyl1BuxCosIJ11zQ+d5ern+nSzrqT6J0NfWwqMWEHkuP2CoPvflgMvOJb4mlCgaXIHe
rfIivdaCQelHWAwDS0Fobh4uhhy3mHSUHfrtkRG6UaeHxbYWBbFQIqTmJw0HoYnn1CpnGkHg8+AF
HNerrA0j6ZfdSvpgkPX4hNFnSoADnOf2VmZXzFTFX+jy5uI3uSel/1jo7/osENlK/E5sqQpuhqSE
EUyrn2BTrVZtt1aK8+hlzN19nhjsOStGDoaMS4Jc3iWbYzNZ6/I1v4FWlR7O6CSv1J7+jG3goMwq
ad1fzHJmfEzRuWI7JrptNtBFx56qAvSt7oqctJ3rsbGmyvEgYS19tBN41wPR8pNMGnnQOaF1BSs0
VPYOHnmxSqDjUs139Bydhdk+u3DbH3kMacEH7FZ3b9QxAVR2IMSEj/Oe+yzSGiIvQJzSbzQHSQij
GARdZz/2P1FsbmZwszJ5uNz2kwx1ShcxMp5Yx81p7YN0AVDUzEoMojWWB8Il18L3vcuOEwNn9bom
Ts1EJ6hPTBznXWChbbYggXjCsMabd5tJAZ6ca0XDu2cKUX1VGQy6mBgGSmP0Wn5OtfN450cBsXJi
cCurL188ZsNRS8Q8++AxKz3c8AfyJQOBeasqiiieA4pjcqm+DAcO7Wh6nrqMWB+MfK22ZTWR3hDO
r7DiI7c2wZv6ERkhPQ2CYTt+NC/iE2PFLOaWbHyIBz8eIYMIrqJLlZkRH4wL9QFefbWIjZ8MYME/
ma3ziKHuw+ka7YJQ2PSS438NVDIQH/nqPQk55MBm7vCNxAm+5VB/DS5tg/xDPBUP4czggu2DMusX
CYXAEEaPC9OWxT2N6HPf2/ySEP5FCexqjMrRtcVeaQVv3WcDyNIzmxh2L1tlS9NisJPL/xt4gugc
vTovd+HAWxWAB+/m3LLRwvF+NHq/QTvwunc+2nZrUjaquMOtg6QZ9Jsh0docmTmwF/+IaSHyb8zH
AS+Saf1Rm1GZNBDhqAQ6UZSdv4XFLMD/bF04jrzga0fjEwk1v9iksYAgWTNN8Y01h6/uyV0/jrbL
LY6UXPEzM8KNJDfeqlsU9u56VdTYOoLUDCOvhTtQK8skCNcW0Q+wcjDh6rGIiJ/ayhAEMxBT1Wkt
+dosc7fZVCemLuuhtCWoaAvUFtCbUpUALI4bzclOAUq4Ph0THPwAOmRV6pRexuPixpCBRusAQKMY
GctZI8U0WjG6SbK37AgTf4QEaTVxG1e03HEwXmOhDAve963wtxpPJ98I0BGwYjLYHtqkKuY79r90
8XuC3jCEv2PCTsfsA3wbqyg7EPVYXFL5lWOepMbWbGHIQbfGCrW8Nh9qHOMvH53gjGn31fJuJ2xM
2H+p9220SU+ZlusnFxAY/nih0/uaxTlHCP6ELI8/BnUJfnXUFe46utvrO1ZZ7n98j7KmwDcjeQrw
nOEv15hdddJ8pIy3FEzIUH8lflAlu99VYNjhYbbnHRNxyeR/kUW4SrmHubYze9l4yGA5X4OavaL6
PHI3jmLDc+wFYosWaWFOXW6OSLcJK3egSCixhpd84alzPmZr8pSN/byv0nP3Z2yva/na1TgfiEvC
987satZBmXo/XBjIaqHCOh0uaIwEgUF4ZsryscVJggeSwTtTiJf0ON3J5fElCgJE4dW6e0QWCK+l
YvE/ycJ1M6mvdRTr/rR+opo8jKM2Qmq3oHKOArpB0hc5KTmnjVxGhEUdfBzjbyw6yc4lJNx73cZe
H9ZmwPGLWSg80AhHrnOCfETbJnCkTrxNua+fbYU1KojECs/J3c+kPYYfmc7JnX9daxcmc5guLe2u
KvHRAB+EfCCA5UXg3lBni28n9XR71+VmPQcC3zU1pIZ2apu4+FR6qtZ4S/DzNWDp+gQWOYTPsT4s
p+NefEXhfCevGeHFZSPw0fSCjlVHpXTQl1DSQyascph0M5w4JQPiNZj8LB1Q+qGUqdkc8eV31I6q
wrh7A0fAC8L+JP/MrapctAdS8KmGn2gDZ59Jom+gNdFZVnvPoLsFlOSzv2JTvalL6b7gY5xKJX14
HgVBDMnjkzWyC+VehlqKXn4tHims3m30mFSj+wzSsj6KKUeulOj5FV+9I5+J1JLI5z6sQiv009z5
gSo95aiYQoC3L97FwiJmKTScsoCRjDh7W4ChTkX1Mm43AegdP1L3DiiSdoF8xFn9IUMyDjvj/tD+
8T+OLld0gTbLiq7mlyBrhioeTeXIP+LLyn/YcigEkhKS0u1AJE8ARZ/D0ZZ4Q6MrgqIBoyUVfh4R
wnJe+Yphk1vAjtn2Z8JXogGfsLr/IPw/Rh434rmYJSHD7/D5rhULZ6RohR0w1Juxb8MTK56f7SI+
WOhjxYn/ZkHrVmoKqqetsmBOdqSbEWavOkUcJFACMOBODNq2Gz3l1TmbEHsGLCOYOOlhaz+m9821
vDTbGf4rSd0xhL7HOFn5E3713dNchlqMQuwK7Sg/yfKPVs8dyrEkZdQ2a81K4rG42hrd8+1bF2UI
SsWgJd7NL5gUs1V9ibE0U4cYZ9NDbZTbSecCtkr26vMihI01JvtbZdvxioP76LJZQFK3ZIjkxvFM
dgdeuKfKjsH9LS8h/CN48gItOBVqQ1h9h/CX8WpbToe66LsilJ3jTtASGL6BF1jpaGWWqN2+tzz/
pnW3rfiaIX/23v8fLTVu+vc1bqmB+MBsImMDr0iIb5AQeB70vBnYR3XRdZbCC65733Eq1Spchyy5
CBlwODOOuIk3t3SJhGsGh3Xj09BH+fjSqIgznACaD2nDpNW0ZKuL3eaT30dNjdk3eO+K0RcOO3NQ
BUu7VPpVVjdKS+acw7W+Mn6brZD2Vg7mySCU/U1dYA3L/Ka18TjEeX2jDJvycrVg7Me1rSk/FXg9
9JwynECCtxgf6ngDSbwm1A+vkIZ/ILbZ2ZarhzI2A9D87WTbDlDj8Zlv4PHMzz8rfwznD/mR0m4O
0ZGwprHUQto5NaFY+TJ75Y+HFXLSGPGbdq2FVDD6uc9O0j7O2uqfnygjVVH9qbbs7wui9Q1kcW2A
r8hriPa8dWHsM34yk1oBVbkvllAXjGe9efr4XaRTik535gINQuZupt9BX+0BTsNZvSkDC/yqPgvG
FEOrV91LpA4eBS/btp1hc9dTHXPcgwqn4dzjZzMxUPxErQra3luTiMvCC1GMVC7WpetmWcut2XuG
T2xeZjdLQyHqpGWB6M80BY+TeQi/XMjWcBccvkfkOAmu4hJU1SL+G6gPQFWLSiexXn3ahPg5EgHG
rkqmbQjHsqMOF5Adl/qHt0ogZkQFOY+WDoE09rzDl048LTPK0tMFSKlY1LMlbuXd3ZT+u0EqQIUd
yUpXalrYWr8Gbff0bSsrSVA5GSPaBPUkNpdOAnvwYINRnm/f66HBkGVjYaaX+9GcsMajolbeRDbA
eJL2Fd01LY9JTFYhcrzIAeeHp+RcJ0oRk3btC2ilXFoT/YuTClBCQ4bLn4SKSguiVJP6P/22qf9c
mEzMzyA5WwqkgTttzgwc2AKlw9nLjLEWXo4f13FU8UPbGFaWMxRNOsW9AlPvid7p5eSA83fRdJvB
arFw6jD9DtV4nerfYvdh7knE9m2i4WYyzRB/rBwiYaTuGDLiYuzsxzt2l4tmHlSEaGHlZZBIYnPx
uFySSru11Yz7ypiSPAary99jqDWtyT+d9qkU6q90a+mZzUtOGeKdAVmbsiwhGeWzj244Md7CajlV
OaQ8mq33dftO7jSG9JGvL/ftsHo6ifvqSk49z26phjsKEL+p44vYZvFhrSEa2JBd8p8mr69/IFzf
inQzt8mCT71gQIDWsvvwqDAl2FxViDjduj/CmB0WbUEYsuF6rXVnV58i4ctxL0Vk7/8W+JtkkMmA
pHzU4bWscDw28hV5OIqwYL0mnkZtMwyWfsa7SWGc3JATyBtX431WGW+MYpuvJE3Gm8aolF02hUjp
LVA0BQ9Qta/VBzvByOn+PpxsDz68JjBL71D9Swsyz0jGFHZ7zic88V59/0VwvA3gUzhr4sfRd0W1
+kWoQBetr6nzXNSI322dCU0Hki6pe7NeKPqJ/Qk89Gb2/JMcsFPEldfez6cFoWBcSr/jGcG1LebC
8A7plUsujiEnHFH8iFI3pu/3X6X1776gPDf5n8bKZH4+Q8B+hqxIEBzU7+7s8BrDiOJQzfg8Slm7
ewlN52CUMI5uMqX8APfT9QHKW+J68AeXmR8gn00gzm7/EXhOOmOjKXOANsMNWv2wUJ2tNR1YPo91
LLOaoTpKHNC5jtfGcr28oBeWaKOCx8zbAxbod9awyWQKiQKS6mzkEAG7b7UUj7aHWPYKMOzxTpJE
jPdC1dRJVNSxxlj14LBANeDjcMtRVbgCUflRhft62+d5iRb967HxZN/T6mejLr7qk3NHXOIO1fkI
3PP4ieMwjX76ts9xeKNslEDOKKwZspjQxv2xcH1gLyrI7B4mk03f5V4yq+oNJOjovOoLnFWQsseo
kgO4zEQkzXQmSTpUXg/rPobEysPb8GWRLg2L7GqWpUI41WXNoCd7C6ACkbyhLRdB7gdqs9dH0sZ7
gE73rvdwbBxIt25ZYSxIsQYd/23KjHASmzyU+H30uHKOvPl8M0I+J3/CMYTcWalS7mFx+PBMbx7Y
KO6uoTOkeMV2wCZOxfMytdGfam4Dvq+1fznwquRTyoXiGVA2B39v2XNLt0bcpxjBZSbRdninMJ/P
btQKF2afg6ykIpxVzWGwLkMXzwBZPdvh2yGZgyzNzWckQpxJYJ8PuDMRd8TUfszd7C2cQJ6Js9SJ
XjqRrq3Dy91KLrT/8uDqDncmRYzgal0XrspXGvUGvvXeVtPqip1nHjcmtDWJZpz5xysqrGGZicrH
pFR43c1a/ntVQ45h9L3JhoJQjbTz5SiIKOJ0gVgu3LKs/poB4WWqlRs4tKmXE/+K4425MUxsOsnx
nxmaJFuSMsbA8TfGd6vy7QBwPKk3ti4NsvtnJWv/rqqJ4FzNQTXXEkHRGYOLYW/s7jcLzJPyIYbv
20K25pzM4gWxU1cYsBw3QQHaH7zao3bbLiBYltEFB3W2RLSL3jvqVFvFxNmSII+CdXiAggzMjx4E
rv37XpHrTgSzS4KVBKLIsiOu+zVlQtPionD52hfFjNygdKtPfW6Jn59YSmOQ2/6dKeEblwZ5nZqK
hVL8niU49Cxe9yzSI5cQ5DPCjrJRvGSrB1TfRoGuNUt59d4JJjsdVzIn6Ky3pji3308YNjlxhcjh
J9WeivfDonAk7rXZg3PPIKB0EXPsUI917qpwkeAaW9rgKczsGksOE9gOcDamMkDdSB1WrLhqjHVt
q1re86cqv7Hj299azMjYNbtXpTKISyN4NV2Qm77VdzDqGCH6xpfl0eSspbiRcwPGof5ZyUn8m/UP
UCYvgLLzmkcIubcji4i3mi03Q/rwWXIklPeSB7WTH1KEILDsgavba+ERyG1WxfRnaYqjyqShACBq
T+UEY6e5FkliWREFcpQa8cO2nP3FQavHTNMAGeHZJdVhxaq0kdnihSS2FwMYMdi2ufSX6YboZs2R
RVxVvX42dLf4rZ3yZrtCvfS0MyGyIxYerLj1NeTwCXvt2apRbTSTQs5P2spaJTfnJ6miFtMyfYFT
kHqw3ADUNeY1zZiLMYB5OsZy5sMhqxakwcWSKRS7PDy+bhodj4nuBCt0EK8DgALeigkUnJHdLDlW
knlniH+EmxRIEj/kvhtTbFeBagf7mZ0/O0tV4Nib2JOfKU2gCgiRmXkXDd24NZM30XxqSvaBCEz0
bPtNFX48O3+FYzRBMFOlngs9r6LHw7k98nFDhxhsijfOR2MlTnwxaadpeNmVt/jJQ65EhM9Fvnq9
MUBpfOS4oEw84SWX+G1NjMFpDUZGtt/3Yzx9TyhnYc7f2tz9vzULKnoSI6L/+KX3kNPh+mUB2Ya/
vVsN8fSXBmMgsppLADE7MKnEyKm3tnI835y4xbMuH3SIllew33sgb7GEMH5axDvx/YMcDoDL6hmO
w2PgLP1YzUcen+JbqM+6x183HeBjvXEsGnT/XwtK/WUyRReKpR6wvH2KPanB2k/XXByMv9pG1Okq
K44Re1hzhCwF+d0oGQexsU7Q1Rit7YMDa0GBaSbviOiQhuEwIJkgXd39UgGE8IsC+yE8j6n6QTHG
Fq5ZJZVQKcgSqD42k8tbUZjBHft4TNJimBH9cmETcfk5AoIiiPx9B6v9v68qNtQx5zOuQMiMapuo
cBvWy08QTzH1dSc4g8pbd7miN28upzRoUVVG4Dk2ZXULZURKFUgbNV2eaGa4uTXGEEeXbCx8hSrd
huPgTSuv9rq4uMU82EQ+YbTgP4Nhle0ktsoAyHRmd3OkbnCo5KBgcoSg64eecy9MOc10GFiQoL6Y
zdoYTK4kQcXtPmoUECggsbdwCT8ic6uzItfyc9t2ubpCLroVNMogjX31E8dCF4rG9GY+zhBVyULD
UeDPPMo+wWXYwhVyl6ILxlpkayy0L99+Go+SXQeaxwlOhyRR8puDnfRozQOakq7r7hIRO4jLV1jU
MLaWI39qOtj/PVbneeYh6hm8zfgnU+J4DRdbjpols3im6vE9QjLp9cuTnRCAUeANkDmBeKRL3O/+
WS16up5fjkQfRsnqojNvGC3jc7PU2FLCQPHDj5RN7t0tZtJqcpdIY2WLii4z1bxmFmHHGLXxTgtR
+d7bf3jaTGk1xMfzkaZFgull/BAS5F39CWuXa41bkD+K+RZ8C6xBv55uUPGoEv5Py4P+L0GpHzjy
dIZ60ty0ozel+vTnVVTnxjW+Q2mLeVCRgKERYgxkZsXTh85WeOkm5G3UZRwkb0kKPbneiu48lwq6
yXlVyEhmS4XfYTaUSarHzrXDab/0/fOZ74kGahZhZKW+XaJ82WwklM9MHx7DIQoyG5Ggy8z9Z12Q
coH92W4VzopN+TLN6WE32GAYmd5J1E2hwj4zj8ht15jZC71eIrzvo6jAzspmg2MVaH8wfEfSiWLG
ky72oOqqVChcJqUS6ySd2JkgX8eJA6qOirGNWvj4yqd0FtbUnf7uU9iYK9Ejj9EZ3SLFzJfLyOdj
Fv40xWgc+g381vNdKgZbZg2mS/I+15t5Tbet7Bl7LBNitPOHrq+S+6HRYjHHNI44UEs2nBWE7AzI
YJKxkA8fZmkHaNiELkVNRyB0NheaT3SKBQ4bjlUH6gLgaNCun3ejjCVv4ECfAS/ovQ/h5treEnTf
cE2DqpHLiwGhImWkfMeIHTbxJfaF44jd5PcUYKtwne2710+dUVM3zLzv4r8ldS45LrJsVpqoQ8xe
Ku4iXCo5a+iYjWcmCMB9ffh3+cwWukua6+fesir0jRIXpYA9+XTG68dersMUSoRRoVZvhKo7ULw2
iI0v7zs2qE6Dd3xxjbj067IsFUu6lHnkmY7JuZptAEz5e/e9KxsJZ1DuX1wifu1sfbCQFCUQSuX9
6grecODpd5t4jfOwEP5nUr7N0wnvCG4SyqLl+A==
`protect end_protected

