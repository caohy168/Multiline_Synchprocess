

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GfYQTAbkK82YBj6Fia7/EiXaKiFR2r1wsSVWKVPbLNCTaHFEiWIqeu5aHiRd+wyP5GXo6B3QEjwq
x+oaQ3SNfg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JzcMeGzt7TTOpJACuOX9MGV6Qpdb6bvnGnDPkVGUDq2yQVhYeY1VQoAjSp5hMEFoj1YVPBENp0T4
0cHbYPe9RLPryarc17U7kLdb5gLOrxk4GNs62ZgiU9/ttEj1YyCwFM1gjTl4vwwTM/5WYHaAicMa
PkpIlB7D9ClIldMf2KE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ip4ujq41Js4GXWtTgLaDiE/1t8E7XHc4xxLZft/5KVnlQ0BB6mfUqweUbhxROrhLa+MvgLTMcl+E
qOW9/xTgQvYzIa7y8sxSLqs2CwAmCoPzZ2mP+alx3rDY5AByEC2IJupvLu/o55I1dTW6QQP5w93F
KM+JTgnnheuUUuwO21gm7rplkpa7yNZiQH2fEeqM9o8BCp2XqiAT2WzNrEgXv06zIZEQREMw8PPw
a7/DUwca2hCRUdZy0Nj0bkhJCsFxFP97HBZc553hBfzzQWjl0bNK5dM7rqHo7qN79VU8gIB/To+S
7KL0NbuC+f7wDe+pxgs3TAaBHEeyJYiHrI8VoA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZdQm4T2CW2eJ55eTzMtQUIOXglfk2cQfvXjpIBGRm65nUy9wX6vifYTHlGerI/TuMZX1x3wosZwu
j7eO0zstKF8z7VxWF4VOInC71/Rnh9I457xwp3eSlC00xV7NRsAC3nB4/njn12NZvExYI/XHPqT6
jhhSiwmMPd/gUeZWisgieGVDJM2yIdhj20K1PghB75XdYZY4Pj0ftdMGFpkuAsVIIn5sQg8SVd1Q
Cw8nGHkRz0cOMnsGkQA7PHkbVp+48SK1muIkzxBaTr29pRLffa3rUgmBI/ugUV6Mbw1Gn6PQr0Y4
t+ZQM6P+FYQhugf1SEx3OiQfK2+Qof9XiIuqiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tClDtHP0F0DdlQrePUJxD5OMZxjXTcO4BxSGrhIDmMuFTs+UD6OELI+gTASuqsMrn8nhMNo7cnGy
b5v23Wzi+fx6INsiCWyJKxRuFYE7W9ROeSCKsJf3fkEVCkpPA95q87mgjT7ImLvZvdGh0CO1QOr4
5M6uyoKpA5RcHrPXTmo=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M7ybBoCpGQpopR1Irfkk5CTkQs9JTEZQyx18IVXY02YWGCynpnaJl1Vi7TRpV/ZmwwLJDrxiHlkk
71Yxme6qsyGN51roTX/nkea2oZnMqAcefuxSmfy6rKgLd3PQdI2GsJfJ0/tk1KOxLNi4L5bxcnI3
FsgxfK7cv8CW5f5rkOFr2DQXS4dTmM0hVaUl4inzjAO7qXpuRJ37st2kfcSthN1V3rFWX8746/Wb
vOKzmSiWNlVVNxtK+wjaTDAE2Lak7aGG7KA1PECQ1nCWPOCL8Su7JWyuK+TbAg+45kfBCXjYHE8I
uJ48WAdfp7E+QSTFUrsmZvS/Bv1uIKS9KKzEvA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vAUuqtlza4lXunBfRH+UTsJLTtMFOxwPMemr09O56a0xDqTUT9iPXvNjy8BLqbIH/Zf6NzzfpJVr
oitiVQtuYAFE2EZNDtslHtVOhr/0BHVJ1aiM+/Wv2BmKqj2U0R3SQYNOBhgufTBS5htfs0SvrbsJ
65khVCZwVHBVkKc1DmbhL+YqsYoK5UF7rbdJJcjEO5hI5H7/32ufxyc4QYfCCS+8XWvItAUiR/Uw
acmDj1C/vy0yY6CAYwm8kfjOKfBVGwkU+vc3KBIczEhowh0eifemjCjHLwvGI9AoIxHZ3j9yBC2D
ieVPbnIA/7VO5hhSY58gZ7M1Dr1xPPFXvlmiqA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b2STEKpxWPPLSvVT2HnQ0J/y2+dMHEoqChpXM7AcDFZ3XI9UEb0ixKs9xMVVzH0tKqOqmwGj1bj0
6DwHVfGYesMEVtjA5+MsTBbFv5XdhtJ/w967NE5OBlRfZ315LEO0bYHytf1zi6CrMxw2527KAwBt
XtIWz+0d7hhw2KLW1GiwZdAXjrziblOy5zwpLJmtbyt2BS1KI3V6SECiTP3Ca3jc618o8Mlb/8WZ
/pO62E1N2qwwBs1s5noZOiHIgxLmECrUjRc/OTKTN9vSIhCicYMtRHtW323LhgGYBtolytTKnvyM
CPkknaI2HZWpUEPvYzu4ujK5LARQmyxrhGnbyg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aRkvCX30h1ro+j8Kbem+YovQTfZqK+gjYvnpJg3ALQePnk7gXiG91jCF5+DK7TjbGmWbOzFR0Fv8
QOXeNuuRzbt5IYHfbZEq9hccOYuH6acpW5YO4vcKMKvxGvITMWCuMQIf8Xbh3a9IVN9c6zFInATU
/4b5K5wFz4zDrGXy1zmFTI+vxNu4pcycAvK4Ts7x8j9nC2cXRtnqm621HOJvQ/7RLb74SpFDKedR
5wWQPWdEVV5KxEo5VFDqC0WYDzXbG4lD1XJlDcaJL/YZQJJWVmJ48OUs7Ni3ICSkeyanQ+yPbLxq
l2XfokHNFVb1I4B8siXsLCt1QSgbE8XuO0EN9A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175312)
`protect data_block
us2dbag/qou0ecG+xb8zmycfyZyLt9GoW2d6KY5NNm9YQWLjaqc0VPXFrNS2NuTGinI/ZHaYVuTV
f1TeQaN6kxag91ViIyWZPf9D2fQof5I73Aprf9QN/5DwQGvqOtOEEA/iXRnK9LqKOB4xdTeSx4NL
4fH17Hu6KwNXUKE4y+iICcWWYAuVI2mA6VLGy5rDDaNCRMlEq862T7myJIHOc5d1L2LWPfyndEr0
JWzhOMJK1+dvPvxdIwZ69OyD0w2BjmGFxNOred/rCa/JrbZAUF6BiHW4owqxMakDJq55TpYn9/V+
/pstv9XhzKM7Qx/AfBh6jMtd1oQLRXneHdbT8VbZaPEn8e0sS5pHxUARQg+5iNMPM3akUAWLdH3d
cpz8hW9mhNwbJy1IBt8Mq+pH89C9hGzPQbWIVMdCrDYgZWeNrYLHd9k/J3c7i0dAfKEVJhWKoNav
YE13qmw3Gfr/1MXKPLKKNrwHWD6uhm9DOZs+nrlDDg3vytqL057N1yAh3Qisaza/W///JUHwAQNs
7xBCcXKtdYx9XbAom7SlGajKS5xvfIpM6JCb5gp97SJP7lE3uMrRhJDb6RaozDEYomfTHnqjlHIh
cesqceMyHdkK7DWkIlkLwCOamkkgWGiuaN/WbJapUiYsEoTfLnO5zBFhB4fspc7fe89RAHMmoRxZ
NAq/8FQgAzvm6tcQyYBWgL4at4owdchLLrajJOAQW+w7f5bha/29TxdG/cNy8bLvDT3MgS9Qz4l2
lCih78U254/7oQJie3rzJSq6B26IVbgAVfqfIdmoBbgLcjxSd9IHRzCAKtG/XDkWr5USgwLucR+4
GxVkKJ9t3/reevlaVgzqz90kX2lxSTk0pipyXdiVAJQayhIB0rzwaz4jwq0rKide59fn35XzliWN
q+DuUfJwuXoI7a0yXMCBKISGDEATjBeeiaggmKBLznShKFnhMKbDXL8aynp5JNNwdMVmS73gljLT
wrMYWVz4tGhcm+zCVqniD18msGmzrEes48DE02qQxTRg9KzyqtiLEh+ds7EhTrEpazbv45MZEmXj
7Zz9UAPUdEIIzESryRbCfGeYA3J0dpNtfibE9yKEC9rWyvUv0qMZwEodAAwgKyPZDUGVWEN0NwDT
Cq3wUBR+odQ59IoxN4xzFdyFlfCLfENkyCYXYasSxZKwGZTULzZSOlD+TM9ohvyKpgmasm3clwPF
+fBdx33J1wk+GvxK94+ig4yyu0hexku7Ao0+iV36+6jrpUGr+FXcbzjxLOg5q+96kqRxfM3xyCBm
sAPgFWnfDa54WBVKVBZq280SADRQE2SC+0P8sZ//XE+LJYDxRCKEoadrOtJXG8PvNAinpWUOGDxQ
HdAlw6SxMaqVb6VwCu0z27dN8uI0XbcPWWwJgpqBG9aGOG5nVB1pdP+554e1jQuHes/tvbuLC/6B
e507FR9mxYTGeE9HwBUfdRAMSnfYuTLzITTZwIcPUOcFI2Ia7MkqG7+1pQS5JhR67dhHYeLScfm3
xMAC3mEWwCc4OWLvxWwApbE5frPrM1z5BxlkzxVNL5dVLc1tB6SsmJewnvrp84pr9gq+ppyxV6a/
gSTj/vwCLD4ztFRZHc08LpnFiUsmZ0dV5YSoT6ugdiT9quBx/AUYHBt2dQTOI9A7KqovLgBRu7ZQ
Xwzgh/pxAd0orjAkB8EP4bM1NuvtwbyYN9CNdxmnuBJw9xTEoTGIaHjxLVit4pszTHSaCuTxlxtK
WAma7xizY8inL2qTXEyK+Aw+xg85a7Qj6tEO0VhbAKNpQPY8pCoBac1xf5XguIoV2+9euzi8ZxWt
tu5QjKM8xJWFxYpdITv/O5nK7wWv9sU9X/5Rpia536O9YPuQWxH3OEIpfhKNx/Ak+xEB29g4HPp2
QPLqHxj8Jste+h+eifSaN1eaR+pAiseOBKctWtFG2QU9mwXrx3V8yGSnWBcj+e06YHxhe2Zcy+uV
PrahUy0I0TDZrPP3i7tBahkGkpmHHXLqzd3uE2FT3TfhoEqt7K6szFagev8hZCm/kMt0OFJL7zN2
LiD3CXSHVhwwTr+IRoTZep7dk/TcBEVIYQ1s4Pcnj+DuBOxQ6jHDfttt0Wg3udnL870NMkIn/ZNL
UjBUdQHkuWymhxcYj4CMRyt4zqwwh+tdnQnRg1M/+t23v0TpEabZEdiJEJ7mhfhufEIIY6UGB7HA
QTYmwM3waVucMfY1KU2KiUYkl8vGGBsxhX/vejM/rzFPbm+ZuuPBGcHIwJO5sOzdO2Rr0KAVJTFJ
Gndn5Mo+Z3nAc3W4+dYUAC5iXPzT99WkbXXaQAJYB3RgavQsViGt1WhpG8g01Nks2ltW6oHEdMcE
lQ+Dz2A+jrC0gRwXWlWun+ILNc1NlI4qF6C+/sD7HqOORtOGyXgQ2cb5wui0Ul6+WF/axKgUfdwI
/TW3EyvNu/IFc9bbvwLWqbnvoYwFLj5V1XzB0KFIsHp6f7rdukTnw5ne/Ke17+KEENmZdWwkKCeA
VvpDFm3Tj1Pj3QxmvhuSdJzTEECYg9Ok3PatRXqpcFGsKv5N5oC43L5jIogKNFSk633FHcpRz8Hm
au1+5Vd4VAIVWVVM6cN/kYrqcoDjCRrx+skKlkG2ytXkM836RvbtuuY0uhdew7krdTR7VYHoIiB6
BofDx5z92E8KNuB8d3rl2zrqYxuiqgnsCCMCdhwt4bhZJdBrnZB9C16Pkkobjlc3QIS26GMDNbB6
D5FbpIbL+XCSXxku7cyw3v1cgqrlqAAskji0MkexVKrLajrq5iONW6b8TCL3BtVFEACOnRqFjv1G
ACQtuD2D1vyQMM841z9CyoQJrqLNv1Do0u+508OFibshHbuZlzgSR4UwiOqKmj8/bPfSu0aRkGmR
0BW5/IgeAc49sLnazJ6OPgAXw9hM733xjv71exW0gWirxxBqMFLAfDsCNiTkxEFPC8kRjmtpfFxW
uFY74pLvrWTR1Dp8wztEBRzvYiGFtYM1zNcSsmzB/ArEDfg7ovIIQaX4UR1tycp0ZkITdRe8Ahpn
Ocp29z87oWipHbcz0mCkke9NJ04AoALKVk9ME67aBY9If6GqDumhVCS2TSQHVM3FtwBkLTiQqm2e
kPLE8CELTWI8mneh7nGdP7mmUBF55CWJlg+cSiwv+Lx8HwkPY/39aqdbjUdUxXHYVhIhkHwwyTLd
79h1jWLL1iBHyijMr7WnCUFneEREc+0UD4MtyzuySqo0lu5YIb7GlYmU1VO0e/5NovjeZVwgt+Y4
qH/qbGHRU4IZgzSTcLBR6kAmZYpMLm2RvMw2P9kFkomZfq3fG2uSFgpkzNtPpoLt+Q6/M1T20yKH
G7w8q5pCGBB7uLC6exSuy8kyoOILY3C2p95WrtewlhJAwEEt7OU8ipr1taFM0wVxoA5ML1y2hO6L
OlYpxs3pCBsDVjMaW4y8Wq4sWNlCvXbhhrIC1AXnpmHtJw38v22G+n2oLHy2/hMS+wvVvAE1ONH8
w8CY89xzVOeKrR0DpFPN1HMEcuRSIvzks/EbCJvf5wPhComb140JDgptOpbxlMyQm2ZhZtuq2jkD
7O6azCRGk7qTcbcg6tnOQuCo9tNK7soDnpfzlISkDNidaFbIt8XgjRzCjq5Foz3mBwebA8sHrv5m
M4hHu909HJaKpOhiVlgN3ET+rS37ciQUFYunsHiP7Q2KkMP0PITzVVQB/XxeYQ9TCHVTaufDclG0
6cvZr/RjWBAmAuX6/HG34NJ0NL9Xa6qlfPlKhBauwD2Hr9WSnGEslEKyc7jvflXIEdVmIetGZfpp
BEgnHWE5H4NxUxIYnySSMaW9VN6VuY2d5YXIlfN/Gb9zxfg6OpBbUiO7m4OsvU8JesRrNjES2+Le
LaDU2lDJ3YEOFWcFcxkow7hw8ng5Xa7hzrn9RYvIwgDg+QtpMzUsj3G3QDRe0PQcqr7zFsbtjQLa
UUFUJU9b55LV1Qd61LxxKYCGUimeMwBSH1lor2T5/5SvBO4UcHif98Uvu1qGDJXSL0fFPFUlTcv2
slsVHVUK/1cqRbt81GsccXaHFVlwlZ0Lq9ELQZZdskfhn49ORNveWYa3p96V7+oPR0sBVoi+HsXH
OkPTD+Ahnhek2XOgt/0JscVmkb92DRhamwkQoQOE+HoyDpTjfOg61r9xPqKtRqGwNV3I4WO6rt94
HXe5gKCqPHpaoN5oO7MIjg8hnyDMbucKfjkNvrPDKJyuEAZsAgT5CekvFx3Abq6VmHw/D1yFe6EK
6Pw+JanaU/5nh2krm/p+coGZFoxyjUjDbAqWLFh91fmstSuR6dRozBFrcVsuGN5fqY4mef5UHQVY
uu+0rkgSxQ6hqtqPcsHs8/iysirPCqGJOpmrjB+sxXkQC72Om5j9QK1veg7llu5m9VFtZ0VLa9xt
zuMdNfL/WTBg4nIjAZ/edyWXrujqkP3VHSuWyzODU/wxfAM+MIqvgyPw9JsJi7AmDkKdR4vpGGjN
8dL6r37znh6HhXLWkUyt5E5tCD0hGc+JiDZ7eMbRq7/U2LmfJCI7i1Y0OFA2S63IK3mNpeEfveCm
0LkEjzsD91VRzqVfl2D36m44ilpQvh73031f/dMrxtCWqGHh8gqV6ZkRniVoZgQCQ7r5EqCCwOn8
A5s5KKiHFwGFvKG90c3qQni7P3hHiVsWtM6HRxebstJ58m/b9IHnbk+sBQ4TnhyziVR0IQUDRjwq
g5Jpp9LlS2I8QR6AxKbbhAh12fVqVWd1ShQ8hK/i5tu4wXcp/H+86JKYpvbwMnSsDqltxqXmhK3X
CI4zY1ce1ORk6pSRv0WYB4bn6few+oqIBOUzRjqSMOsGpr+dkJG91zQoZnTj6tBQliABtjrzFe0L
S4aLVRsv2JaObe166aqqqARkX4O8MdXiHbncES4onNa6GS5erHnAhBqV4jCvpX4XKr3hRyTTuOUs
C89RypuOSdHOAMCyiBY8s7KaomAY/iDM4jVfg6DOPKo072nZsc97ZKDA4/Q35k74gpQmEVwDx7Vp
tKlzFjrJwdd+gp9tf07Nte9CKmClGGMcqfXXMO7lh+l5/kQ78mrpXdyoSmqXi7pq8Cd1lcrVjBso
bl8pKqsm60eEyd0nqgXpknGs20y4mQJHHnZqIHNB3GlbPEMUxajeB2RNz078qfr2AUfbjUSo3YAD
bnQRzs9ZeRmpyW38XRYpv2CIxAuW/h8RXqtmaDwhIYsV/FoRRy6aSTLoZWEKPcm+N3qdhEdkvdc7
VYwDK8wWtuw5FKy1Ij/M6Ex2n3ziLsgvyWXX53Efuq+77M2dnQ4I+PbO/ENGzghpJ2mcKjczksbV
Jbf6u8fWnYaa5EiNwVShYfcLw0u0seObV2/Pd263X4++5FiBi9bhPdYdcKYjMz9lWhDafuvy6QKh
57uWfyo8tRPTgz2jwzaOP81rJoPHfgfwA20Uc7iOs/HdaBchzE8YZfrE2eGtC9eq6bkAqoa8vDoy
P/dru0u9MvdKDsfeq7YdQHGwKoscAYJlJFNHmZhE1CvFUtbSFNgThsCRN2pLksvGqeguFZt8CSvg
SjdDBEXqqaXPYJ//E8uTNblftw+Dqt5WGocUhHmqPUM/rwQGRH4MRmMaq5hshwNJ5n1Ygq7Ikt+7
eaFjc0PexKUQczmxoQjDVZ3fVFNBNc0Z3DoeHUoX1YvdccWaqbtFweMnFH9EjcKZZPn3fY5/Ce8C
avXw9/soEB2Vpdc/eyLE0VGWmR2iFpEKsMcXb7oxPspvFZayFPDElulyIk2/RFp7RfeU85P6jVI6
JR/KeM4Tk0Ccr9kfXCbPkILloE4Saq1DST8fn88ZPpkK3UvCxs9iwNhkvXSS1qziIvIkzsptSCs5
OdnjRxQ9+X8kChGBN1rOm10XMvLn/OcR7OfdBQHF6Jq5HO7RrE/+DRkgqkXSWrPPVLH7zk3tPst3
5v59ZtrFhUY+DcMLvj3dbjCZ+Oh0FnbMU4Bb0LwivNFqx2oNmWDPHDc3OMYRyQLeg7xCiHHuyET/
DduaW0BbAd9P26k8Mp0jZShW5Ekmzyr/MhF9XDFFp8e4k6ybkQFp8n/sjh5xbztoyjUDduqD0k4z
BMYURFSMr+zjEVLiDOlqpOq3fdrLtQ/4b0yvJO/CEBhaJz6hGa70EWjGW3kfDgSpCzYci5hWDoeA
nS19/oh+39x0LNtpfvEesWdzKR1eQwdpeCIUoqQnipOt2Zu2nXbuOfMdYm7A3c1iNFRINi+TzSek
ZySlnqrzfNHjNDVPBlgSJNhIwfPlshI64SL1j+MD+1odLtaPD6o2iCGwIhwWHl3FeW0ISQ04+/yN
8hMTEBOVb14HbKRtX5Y7FN58+pL5fLv0KeyvUvmN6hYKzuLXPsheHTeahZIzv83pnO6QqjsXyDj7
f6WIwRzp7TPY+sN/JfPkHB7LvMx797qdq2Nwi9GItLQ6JBsFmsb1PMplCSp4deKYqkx56uEvZGkL
XVEvHSxIddFZe7AIRRjNswg+YHla/fXxI4HS8255XlbkdzNLie/JZxC1nDmqRACRdAUmf6Tq0J+X
w7KofOGD3Pzh2fzVrsJBAs1iF5+xBG1s0BP2VLdRJFXTLZI+HwMYzXavWlKYj+OW8t+x7ySJn484
PzwmZ3hXFVFz7Vh2iFI7aOVh5f94tM5/OC32s1iIWs/E/7VcFw9ZlfIUXL6C2TJuklm9gKgtHRiJ
G4hCjDCfwvstYo34HWRo19gdcq/0sdg7/lhcBNRHTaKQ/ZyNV+RwPGwPuGcv4KL38Xt8UgANZMNO
1oweufoQeSFI49l1fVbyWsEtPLpFpdoYk091291IY98P92H/wlpQ5otqmJc+HoObkZYUWhZgW8Z/
Cd6DBaFegWr0xB1fE7fWr4LI3RJWTGRzxNNlGSdUhNlgpJnFi3gJtVTeYgxx9D/Icvfxdm4EfRw8
fPXFdprwXXv2n77MaxSCYNLqyuu+gBBWY5ZXaaSpuqtBQxGOAFOR0HI2J+nqyNZ8AaCdvpSk+L13
LHAZr3VeBolw7p3ipe/ZM+jz+ST20675U14Fb2W/+ORifMFysAXDoUGKjcx8qhVG8LzD2auARGav
sW32xSltoxEmbTrArtIdgrxUbXVbED/fteT/QR/dNSkjpGU74fp7gyX2Z5USeByt8o7OplcKytzq
WMVJDv8VV5+a65yOaJrK+wgmwnM+WK15NfTrapxwNLWhvzgGxXctPIq2q6x7eaW0GkwWlvhTsZuZ
aGQ3dx6vsWa79s2aO+Yd8vR/Ley8jHaz0IXMHH9j5IRBIVTiK2+SnhqusSAai8wDmJom4X7jhoy9
GXYOdMwYLPyCfJxnVf2RCQKMts0agWmPB6Fh+ewHqco81QTEVp2rliOFRIZXg3NwiPx/zpsxgw35
7S+kEKsS0wS0llN0GBOtn9Yee13DAx5sXg3Vn5r5LvkQGQW3nDtcrWrNBtxDYbZTPL6OxJCVmXVh
2O+O5IeQ6SmZN529xwd6xnCJyI9HKOXYj1ppiV2BMXQ9ibvM1v0YOwR8Q16DHymjJ6/CBSCzS8jK
aMu0hjduf6CHVhPmCHPo/ZRGSFrsub53p1NBYkyyYIbm/LOH55QpfoZ+RuFeQu0izQyFeXye6WPk
kHQVqdwOU1qyI+wExkPZRmPO7KVBfHIM0rPTQm2WUm4rtj80Z4mP73N4vbGJzJJktmb+3DWLYTjz
RzV0danxLSqFw4SnCNiu93GwYsHuS2tSQ65gPFJbxxZeUBC+tVR5oOnDiTUi+ZRIf0xTabLP+Kxn
p5iRnazzJvb/CFHVao8lgDVJcUD3yWf8+Es4oSbeu8501QF9k16JkE3BGPQJVj1FJy6nwYf2EU71
FF5ud5gIIFBym0mLk90jCm0nLQ90ZwrYr0uUuA3MOAsVaOEEb5eWD+8sIfWrBArlr/Aua02WgJka
lJ3yculako1QqLcK+xNiyt4++P8pbP7LK6j0k821Gbvr0QKJpFOb7W9ENEZmlDYNH9tj4TqDo2Al
wGhCZ3ryACO0v8BACLvGOoPY89nxHJmeJdHreJE7US9F5yxM+ZJMHSHb6EPOi/XC4sgS4l2fNDbt
x4a26RQudkN/FH7QfM8BHzY/PxjTIcX/fK6Z/k3cDypC8DfOGCKgKPYwG/al4qEWNaRy/CJ5Vzbw
upYPNnYieHlTXZAaIcMGzDFyKEH+IVbtWj4mockPDTbZI3WGlraYouT/iqVh5X+4Mp35oSbcLlo3
uKfrGtfGK6u+wvCCne2VL51hlyw47YA/IFSmLW1OYsLxe3nhbGKlMMhlsVq4u3f6KslSe6CUWFka
khci3PmYR5fovOOTjaUoZu+F5aSbJ+NzSoV62VfQL+iT9nbAJ3kR6pg/wsooq5mcFhhQ+b8g5LoS
NpDk5E5scopMfJ5gSg3oq8WXVzgqJmGbWd9OBVoZY6lJz1/YV8eG3b9NkYfr5BBy9gU2utrgiD14
9sorbiZxM4RB0hKLYIDQEqq6lBe615FNecznaUgUW/SuuqnIUm8KtJJR1WaalXt5PYKkU8G1a99t
yxiElL8dGQBULVmkU29onEP9unyOLudZ9A+Sixhfmx24L0aaUnj7l/hOg8iPiydP4ssYXDQ6BJRo
6vt0OthFMKQbiiF/hvLdkC8T5Dd3ARhgjYEEOKn7YJS4TsPbAOp2t5u9JSbkvYqvl/nD8xy7sh5b
MvRalWxOzELcN5uLfbY2GDJTrbEBoI2lDieYhtjsMLZsb22CFLKNM/piSiscarBl/UbfW0f8rc4S
D16eqYayKL4ohHjhchQpBXSrY/wifEfPh7vnvZplDjOWzlxSqCSyzXQBF0SrxdhHCR/OsprRxj47
5vYkhaDV6YNPkdaRvRROhn+Meia8HWI9J1T8brgHjekBqtDPnRzMD4PRnjvV8lYduNNm6DHX+XK2
giZUQmEkos8xWnxMxv9gV1AK6URFQXT8YjePF11bqlhgOizBFzs0ZpEuigPo6fUrViXliMmIZNGP
6zMClYG+53eNL1+cc6q2P25J3YL8whE6gP17G+143j7gxlkuCrOcN0eezQtq9+wvaxQrNzRHABsl
ncywxt3iPeSx7udIdsgWSVwdkgrWaSFyWPUaeK4mFfte8ag94UOPrDeCszWQOtTC9BkUIVlZF07F
pxuYZP9gjsGOGsNCwZIUu+H0M9pX1HPAew2nzPc+aY0jTCBR3MWkewVTA/STh0M6T6nPw2wPj4T7
KwV+NGBwMyRofi8KLJqnUnB7SLs7mf8u6+YkWA5drq9ZtyrzmNWifv5RzLYlzR38wGeLpR57syzy
gVL5f0Po9VFHpfCrBiw5Bst2mMpii5Ab+tCG061yrkGXWLc4+XAye+r07oCAJAaLTD89HSgh7VUB
GHZNSn/Wz5VukGUSswtON3jWBTGq5ylHU0WbZ3MqF3DDeSvtCvafCkkOtyFVoyK3OPfDeMl4BvyU
aNAkrg1Rjm5YLzTvKD+bwT4NRV3n7KfLb/GztR1/to44B4tyLrV9i8cQHcjCBK3w1Lmmu+sW9izJ
0/R398V9HJ6aokpk7o57E4fxDIbim5JTGro1yHHrwpjt94SodNRdJ+P/RvoyVuqGSz9XCbYM2Fxl
9s9lGDTV98CPXiIfImpDTBn5gSFDX9egOYsEZSUkN8TC8x5MSppKmQW5kh6awujUsJYqok0kYbYu
7Ls9ruq/LSNEsZxlKxvTBRMMPgzOGtnVw2aEIuCw1Ll37NcMR36yVJXklXglB8RkfVWCvHc1gOOl
AXE2AbbWWNDuos71X2x13G3+qJjFo/sVCY1EgrDxcK7e3DVYPm8qFWh3YVjmRNfr6U2T3IBvPmox
DUPnM+/e7dQIBuOksxtE3IV/JZkgluVxdumsdGtP75HXAcycJQ7RDZ+D1qUSMBwSb/pqtGIKvYz7
UYSZxuDHU04pQn9Cg8nD3QQXkcg11jNzILRB1Ip7QAw8lBNfB48q4AfMxsy/eOWiA05/r5pQckww
vuggxyJTedMrTUPBpZmosfiv4uulQeBakQqi1k09UW8Zrwz9lb12dA9RPK2PxV3d0mZgKEt9z/Q2
v4d9ZyypGAvX2wiNrvmFFEefn9Pjdzs8yV8lI2eCRhuBH3HrfetspMt4UeoX3T+hDO6eLuLW6rhu
wAjv2GLk+Sa2c+IoliI09R1fgNy/W06H1eHD6PrhVFj9EYLQTWkG3e4cZl25as6cgEuG9ug0j3ic
d6SZr6rta6+4HCdz9tEZBg6kxP6z7BNuS8jqVsYP2nufwaO4R4cWKYqpwLVNW4hr5UWvK+a6JAxT
QSaYktUDGnDZ7luDBE/OH93I3gYDlbYbAn1HuDuZsDWSjVEoVefLNJFRz7eTIiLnO0U2PRWPOXEq
ZlMQn3lUSrb1o8Uia6Nr8sVn0h5lKu4/Ik4Zar12us22iOrN359eYdVITp65zlAo7p97srE2JSEa
uPtGOGF7ZEQh3An6sDYa/kGI65SUVMx3qKON84KBT6GwgB/gJHsEU/w2Bhjt7TP3slQbYt3B5png
479xhEmguQMkB7q9/+nlNzLZtgcEvFCFfOx+HJpIp1Lfh2n2sakD6muXdmYDy7TBAW/ublxz1Okr
WOAQkXq+w4WblQMJAROCC8hNoXOUYb5e7B6U2K2ycW529bemwZdyIiRyeiNn7AjWfdZX+ru0PItZ
mtbSpPjAkgJChkclgfSVKYS9VN3WjJLeXm+2LN1W+0EbKRLwRKTFdDiAcGSAfARg5kfWVEeQ8x9D
SWobT1Vz7p1eaylSzxd9LRme4ZOFHJQPv/FvwnDPg/oss8ashtGiN1dO4OVrXiim0IfB9YTbDGyw
VrkYZVTtRIR/9qECBDQqhWtpHSQ/oP5i6FTcrLT2gtbSz1bHIsB7jjd7CdaF+7tIc0NetsRoWB4p
7LbhwmB54hw8tfENZiWkAYQNZZ0cvn71Tkq5fMWewGuDRPPMGl7Ftf9bx1sPJ1d2U/7v4kotpHBC
7Bp4RM0p6enJJ4sGtsKCwJpdXKIVSH0+0+IXkwoJyD2jiNniN4tdSop7qIgqq4MmNfzAS/fjtl6k
IC/DJQAPDgL1gP3gbiHu2JXVEPZOOI4hgCVXiLa4VieRb1gbALsu9k+ZZbvYGxt92+YACMwlkhW0
DGDl5LVsqDExe8m/DvYYq6SMv5E6fWGwNLhJEfdFSrwA8E/1LkdxHyB0WOZBN0fjNupEwr/jJ4Sw
QR4hu/BksBocqaSoaYvAlLOzVW233h3GBXo59Ogk0ziOuij2OBZ7yPFoyTjWvlRBX/xhMe/xFRUn
h2RZ9M9UeoG2j8LY8XIPgT7xPk9mOH/DDbO6wrVe8oCuZFCUHeN+nvMKV+isHW0JFHHxnro9NayE
AohlGKdeEU3O63DlQx5sUF58074p7rEDGu+WZYqy2iU48KN3gsZ4lu2rvjYWu504whlz+IyE0lwG
PN1D4BvE19IoZlv+X+YZQ/tl1ddw1PnTNz1mALD1rWduKSjzQFAPeBywqKzd3S43H3C73/OGT/b2
U31inaW+mXzRLazyyEHn86vWZVwij5e2/p4frTDTNzcX16b18/OUbWAMLwaeKRAtAgKuX8MWM5Ep
1/XZno5Lg5FNuEmVStok+PZWV27tPsvmaZF1en3rlErHmCQrZ8YIu5suoT/o0hxv0kp2HvHd9OEL
WNJeT8M74kZvttAQ2GkbU5L6L3P+NSyu6lw+d7gbdFPEWmYw6WOQotriTGUA39L6a7S7oid4T21d
XY/3tkaUXVp7M/sYqUs92K8mNwErGELp1ruwMoW28mtPKqVgey1D24085df9+8PHlyZGKdiXXX9o
KOEz+7ZhbLKdG//w2gCsPBYIl0LzsYD8fkIabiqCKs1e80zlvRMM5yEZk8SONMCSEJ25jgB/H3Oi
DgVCpSTLKTh1d3IpsaY1s0O+nNEf5a1av0gHwBayPlF0bGH53EzcdxLDy+A//BBAOaljtemAHmt+
IhS0o7zEE3k6XdxKCNokMBsxPXBdy4NNR89i4sb+bmDpY4/qzltFD0nWT/+YaTCSpbzUekn5pGCV
n5vj2v1U0ZVc0g1L5k0SO6zOSAAiXf/5g59otkkviHMZea3NfgGudLSD7yiAus5JfzqqAZcanaeM
MVLUkyrUurNR4bneDtvaFWv49bNtGrwKNwJG10+NhmhHCx/4+TFHGpN8SqYYkE18W4vd7JqA6aDY
va8PMszH5GLYL0DmVYDDVpJSWzzCuU2Wg93zGbGZXSKTMhtu4HxDcFJaR1HjDh9n0MAkUMV2k7rp
iURq7CroGefmHKY1N1uEsEk+MXx5q3T/2neX3+k5/X7tVYZE3esfgSu7OUvr3gJFmDCF0jVQT2Ut
Z7TkLj6OVtbZKJum6merbzRODf3fXM4CbB4ln7uQfc6dDgr2nkKymVSpkmNuYA235IpXe0Ov+Cge
f+Ejnz176LT7YEbQ5/8jos8gq4NIYK+LBQiBZs3aZY18+LTXfDXqGq4ZYJi6gpNh77o7mjiaVP4E
IDxqkV+0iQZFLJ25FtyzkeK1UpLYEnLkWzAOHkBi8FldO00irslzsEikpAfD1vCSp/ldYLnVs+5U
ZylZ5WExv3042so81h6h74Dn4ZAAsV/ZD7fFfRUuTjoQt76ZLyRLA2s52AYf/Cp30POHlwawNv5g
FNW4LsR2LaBCRUaOmwkbPpyFb/paRfPPSayVHNz+rm+frDH5bi3c3wKMkEyUpHdxOnYc3ZiYhTEC
BUKb1Il63gv/ApZLQjHjlPIZb3rNY1fXZsklzH11CBOAoMJJNRX7hXkgT/5YVfJZ1tqLJf/lZlW8
Zj76e54ALmdk2oC+Qc8kZL4jj5pRSVKFWdmisATDGsJwq1BYHLDAE/gqnfc8l/TtcYb35ElToHaZ
TPAAYiioI7ZeQesKmhNanoW4o6iHB4+e8P7cgRKodNjVTCx20jbarUNoHfc2oMghJ6o33rKsNiV1
5klgSeumOKGkPx/kQCYtK++srdi1yo5P6ldqlggKM5Ss+XPfw6BNpT/SPysZgY58q9pCX77Vdexi
iibN1cDEUddlgEn0ciLsPW9wk+3U8X5d7oanCPvNk4vWf35QuIICcx/vRYsjjqc0pU2uMFiP06FP
Ex/mNGObaYJg4ewWeIehm2DJsJL+MXOttgcU4E1EJ08bc+XyBYaXk3sKOmdMAy/vNCXaHLi7kTNe
o3gFZXkARz5/JA/2mfntK8/SnALlEHYqzL2OISzLnyYl1qHIWvlrOdeeqZ55Bf5Rb8w9DfCUorAD
ucQ6b0jNO0BFZ6XzmMiqJZo7PQOoKffTAH4umB1CKqyZhvLg8HzjItqlipPJvBJppIsWvpVAVgyc
eGyWsnKT0Z0YYJvWyFQEuTAiEikaFfM2DKZV8fVUJcmeVbB5B7XIk4VLWoPO6aSVtMmjucSdE3Pv
5gBGxg2fLfpFX9VK6WGhLODXeXfJ4KztI8lbkJULbqM6iJepcQZ8XpAkLIG29CRD0EwJQ27YU/bb
k9coxDQ646WsQRkMtenJ2twbisvQl0nbd5ljKOxP1kULWYHEET6tMlyps8xTAL3LR26+trEPsjj0
3azBZhCDUdCZUfFjUWst82dIUJ/AVRWI1KR0FAarIWmqjWieGLE47+ewuXxI2DTRswmHsZ7taZag
KDi6XOMtNkZzNFaf8tepSKyRTOoH1o0ns1jbmyRp74in+27YiVlcNogImclZXxYLMwU1fdwHBvHK
H8MZjwyw9miQun+uLFMDqA3Z6wiOUhnIcP0dAMjDkwy/19PxuUCTGgZZ/hJ8et0IArzE6g3KXwuC
ATiG5oY88xMXgDUquNCIGBDwFm7PX213nXWL9tLfPLohb6UZcLZAOAHidJvOgwN9fbl2XwYt30Hz
6W0wQtA4HJoEHuv2+vemXwyLFlA7EAg0858ArBlu0Lpn3BjJFBVHBN5iz4l3qqCMAFWK06P4Q+dD
vdsaK3sm4j40aNoGnqbGcPz+2aX6ARzXxMSKCX/Kes9kSvdgaInNVGqtFtO3JxBv4sNn0vaYAG4c
id7NcgV79RR+ctmiDz1BZ6UzkS6CS6gljgXPbqJ0iU1eByD5SUdvGrtO43HijJR2tvn59di09GQ0
GrccsPeq/pmu0jHZKOCzv0pMKzCmq9TUew6VqB3YeN34TUiVgE/AYqGbhahngzW5HooLGjOTfYrv
ldX2IX8hqyBTkWCMg8Ng5liDODw31XSeVmk270SFsPghZmYXN97LQ/XZR31LlHDEIrPYqkYAD2Mu
zmeU5cSXb6We3+in1smf4QtvmzdZr/jBAcSdh74EOv9JR+aAxU2fFmlRCpT8UdQ5zIvklZx6GIrT
UnEu+kxVrQOYOgam3FqhOwRJ75jgs+Pi8RiDSkauSS0CymF9xkOBgCmYGT4SY4wa4vxBfOPe0aLs
tPPSy9a1tZrybw1YxIVByxWUqFv4Bzc5ipQUyElceCZB+uY3ezh7yCRw+ql+o7rPhHELa4l99MzL
sUtS0kemVD/x92z4aDgxrWqSn4Fs/wNr9pMENofcXElOHI8Z+uDM70PWX3ZN2uLeSgcZNjxToMzs
C8eXBX76JV07ocy0OtCx7lZ2U8Ogy5FqnQT77rPMJX7I+2xh6GBhqSQPfqHi854FfKZfXeOSF2uf
Jz9gS1vD6+9479UPSZkL1BElYZHVn16gFZSYstpIhisLvcqrICG46F6WwXcwyIbyBC9JNZ3Q322a
PJ058y7k4eAfMv1oTuVMmSBWHr79gz/Ydzvdebt5T2dJJsJCRKk/ZIjByvyPnhgrgQ5hQJZ7scgK
9Pce12mfGAay1DRxGDw0EsGYuInin1G1CEM4W33eYq0yPhd88U3Ye8MfX8TQFaikaAD4qkz8B9dE
69h6RirH0OaiWz247nGyg6gEtXTq2fHUML1r94oGdhX1dshZ1KUe89ptaNWmdXVbkAOMp2QhOsOV
khe8YRb9Ze/rokNmOTgCWW8UQwInDSfOSRjn1M3xlAhTmA5tHRkfDg3hdPag9V5dl+ZIhBQd2tPK
sAvrGdbdY2xLVy+tFjkz+ZVEnVeS8jwrGCms1FAzy/kCkYPbBq1xGNsaJlHPvnJ73V7ri16HqLuT
wxPuwm68INJJxlXjlBN7uE3m38tE0paOPVMN3MEAGntO4okT50oOUIEahRiUr5oUOG96ytp1WPdT
Hcq7fllC5AxiJLEg12dKdjWqRj0ecfaecXYM6qKNPK49Fjv4u5ObLHSzP7VL2HAZs97r+yQn6OVS
MC6/wK7DU3GLvRTc0Y4ys/bNKlPXO45hYdjuAsX+WclmS6E1sspWATGfBT/6BYHFiIHCufVxXjQ5
uOjpxquj/rd+FCseFtt6QxXN8RTWISfUQhwJcW2QZr4gRnSG0gbltfJ4R6K7HE1gsXm+QD5kROmq
sFr6aZdOqm6zaDpZeUqda4+j3hDAZdm243I69j+1c5e+7lr3nzVxAck7Xu76DAZFCp+PRtN4Akm+
uO/Vb4TtFv1dNz4APTroNzEdqqEFHOT6q3+zAE405DYuZZx9HVXgsQ0UY8vS3uHqXg0Pl7z/fVK+
P4JiYZIZxqBLAzGxf0612QyQ1rQvwYakPlIJaq1zpfOt8ye3PPQVjE67o6rPWL/CCHg/e3mrfoTR
cfVAdV3hRLs+RJ4tbvV6RMHGLtoiujNIvZaXd52kZVg3pLlkmZgtyA1KzJTPdDBxiMRqFJocQkJH
YOYFkSeyNKRid2IEQZZfGTlKXZ7gXJMIwZOnBtGuKvEkLxctulZZGglyUQMlU41dnWjH9adsC2/E
OXsB13krAKkQCpll/G53c92w8cffAIQ4v/MNfCG8C5v/HDENv1/Q8AY/BMesKmWyspB/Q2jMGQO0
9DihBNuPU41cGUzgDhNoPtAYRNgOOxAdFu+9lkju7ZGKlycJPiAEGSB8V+Hvk/W3x05//tgbIh0v
PtwvKhk+s6VytzPQkYMbher0YkqxFI/Z/rfZXK80N9YvWBsYI6BpU3BHyNeouXe5X2rjukwyZyMn
1OHPjHuOfk6+u3GHeaua3R9+tXA9sXKb+OV8iPQknAs0lGsUhgF4+wSlnLziSMk5PpgJYuTrdJCB
ytytF75SeXx7biN3m8D/QDBv3ZM79kmSCQN1tTxf0AIZ+DJ5hnzHaJ2josUVAsMi6DN86LTm+ykR
1/7el7roZYNQGcEklBDaxqJ/kiUlbpcGhzTde5VesmoxReEhKWcQhZTPM5aqZcbBYgTgKnUrYL2K
u8pwzigwqVNKxCyNj866p8e7tLBo57kUAxqc4bBIo+QBIBNLBD/Xzt8WO0p0eNU2nol2Iqb+qSwC
EbPo1Ej6X7LczlojzOAN8TDw48p+qRi7oMaG4gd51noclg2N3m+cY852MQJ71n9WaivtieD/QXcM
P8V84E/MRu+sJRcMRdwxuJFuUxp+wep4eBhEzqN4T6U2RcOGk9e8n53L3j2zza1RwdySBZzkJycJ
bnp25+4CXp5TP32BQ5TqRy/2XXTkWx/SknKGh0jEVZWHanjQqzuqc6OkzT8mlwKzgzGf+/flRn3o
QV4rfb2dN8eJx7049m3Ad6Hkd85V/+WYYtdpKZ1HfkwGsakj/mhRuK07JPCv7ojL3mF7yHf9iz3S
Q0jN4+cIXHQlv1NSdZiHOdv+vciFpoN5bGm5LE3U1rR6NQm+9o263oE1tgO0DPjWej9h8Hm5EQ+J
IR/GndJY5EfVRmm1POKBqq/d5jF4IvnrWMjbugGmYcnMQS/Jyv0EdupAiJZj0sJPRsECxMnlBdnx
sMoxQ1zIpL1E5gip1Dd4h/FRY1b4QdkT36uf8SSf1Y+DryxHFMKM53VKvI2WsMtI0exXLgORz7nn
SNcIgD1MXh7II7AINNCZP79r6B/7cLoGayADNadfh3Cy9kOZ667OYNYc8GnimffKDEWzAzQCpp+m
pae10dr4N91PF5kfuaT7xrV7tDfRB75UJJ7BYzFM5J9QB5vvgD13Hos7+b6Q4Aqi2rqiqh+3YD3Q
lZxrzMCh39xU/HcPx16W3Azf/47jC5EVEjksfHu45MiMzrQ9qs+YJpT5hbqlyi6JCMx81dHRWxah
rADgHA3oGbwNVqurpUts4wDy8I+KfTH/1wLqXg7y5afL6V+wDpy5oXgfMXQOt544X/UTh0zLbZh8
Sj+0NElapUlZftfLfAl3x5oBT4DR8fdEV3Wra3kkP1Ayk2gQncREFqEDcpD1Hx+1RlECkdBc7P0Q
MDbPaLsdWXkbLKPPqBbRdAMm7PgDdqOYHZHJ4+RtshQwNKd4vfdSLS0/xFF1Xi2x4KQUklChnCRx
aBGwliJuOWfMTwdjcBxYv3caSYx9C/tMoqeW4/MLC1wLCKPjuIFx+XaR0O9ryQfackuF4/em1RRx
dbOet5+bUF36E/w9w8K9LohMM7jymuALzglwz0Byt5eDkSHC78xH/rR+PxDWt8f2j0VWnJvdq+JN
usZ7+DnVvAebQxqWcfX3U4WQN2qO+5k0UYrmwqi4vuWRxqXlgJuGFKUm0w2VOznjTftNql82viUs
AIjfSW04tGllQe5QUp/FZ1MLjizBARi57OwbYc34nl16ILk4eJMgCE23K0797LwJqHcHfVrLXIq3
xShy/fqW0Rb7W+PYYkr5VffNaO0Fwpx52ILLv0L1+ZQDe7CDqWzREXzlqrlvwSBczEt0TXVijdo9
Fu9P5P27ljfdnjF/V69Rgckfk82u903iCLl0qBN10iRLD4FGTev8Z2JYxz0s8hGSIQymEEPMKTCW
IpcfSy4Sq0o6tGPx4zgKh+kAC4eK9hNFr+4LVtGMr7wESsgYoMKqlPfxRc9NDA8nd9BloytoIaNN
GUdV+ZQrVv3Fw76tRS2kN+CWSRorc08daTEZKW9SOwq2yQhNU7SuzUhDuQ+Nh8ekiOqc61a6Ibu+
5RtG/0xl5HTgVM4dToHliqpWtm4TFSbUjLBN2VDSTWI88w2liiBeSV8w17RxwQ1FJ415TJaNsKMR
7Otzh7V9SqacjKgq2nrsS1ps4LNwgcJ4smLFqLXIG636vMY6ziNrKLtllhnr7zaVqcLXT8sOxLEL
cCV0paCw8WrRP513vPxPOIR9/ZVFmIS1hhqKRn/g/HKJFGF4LBBwZ4P5zaJ+uL//bfYvKBCiWl2I
31C+rXKN8y6q4BlOcATKx2p7itOSfocZajsUpGnohX1OMD12uZn1rmJpGxAWZqPkzwLWEuuN/rYi
tkouyrPmkPiyRbI7fEr0W3xrCTv/WDeov75MuvgQJrZ7/mdkCuW6VaAqgUaxMEF8StAHNb8Q/0Tq
dmgE5ZT3PcnWu/llOHeL+Pg464qAWSKY4J6k1/VcO7umY0JdIYAgKuOEhQTdci1t1snSjyOtKIQ2
utM4szxhQ47dSJppaFNuMxOwJ0gEiU+n9VNRsgjGpmK48Z8HC5TygbR+YfEmLTWutb5v2L2FACBo
UYYPH5lkw5D9qfiDU35PVQgBPJBK82ToFyGQC3BGKFlCQVBtCo4/xR59l0YPRjLUmNlFfo1wugl1
a1xdShCIJ2ewyISBr0dQJV9qPhx/S5VdUmPOU9RojLwqZXfXbTO3vOQdBLlErTJjGbS6M07D+6H5
G/rXO8J0TR30P5wxVcL299/NIoy+VxwsMzEd93wm5jD82TIBz3GWn2Dk0joxikKiBvKSt2rv3T1z
swclnN58q3dacz/7wIbQjimher0qtavYf3PYMyErdYTUcMnxEqVSpCog01QXhgT8PNmijGrAGRyV
+IiYeoGbTDDgD0Eg2Oy5qwkitpJ9XE4E7lCaq/E04UO6WGM2M0PvIGYVQj3Vdmj0TLOwVMLeywty
c+p0L6lFJVKyDOHUZOjyGYTpXSwti2oYd0c/Wyrm9jSRwYjxYcYNebPJ5eUQNVx4hoaNRf/3kP/d
vb6PEJEhJ/O4FRKhaeMSeY5edfrC2gl+qmoNGTJ+pCWCdj1uhPRKvjKn1DZ/kbv6/5Ys/onkJuAl
mHAzt01WmB+M15HsdTnvbGywYcMETEzDcG2eyujgrjziyWDW7XFT09qAm1SQmSNAGcyJJjD6uKvN
SvOtv38EJ5GcNIfQ+z4rqUB4ss1QWoGmW0mSLY95LeX4ac4+83h+f/hn4vos8eK/sGoIIjsvxSUO
z+G/vgl9WFFgFbnzGw6L/Ervv4VBPEuTaRzRupkqdbfSPQg8F/HE13RjN7fMIMO5phrnIO0KxisF
j7seJVlEBaNLvUi0wCOpXVZWf6Ghk5Rq5wX62lS95nbfXBqcVW32fM2ZIOScKW/7+uZtLFbzgc3Z
qR4oNzWRewDoutK7k/Lgib+9ncPHv0J37rL+3SkoBqJ39vHRA+pvhpPECbKpOucEmTHXAXPryE6+
VkbA8tTsNv86qe7PZnPQxByIjgpHFnm+6hulUInm7O2DVf/jyOrdvRpl2YrBZN6z61J+xmyZF6kc
z9FqTN3wfA6NS7nk8IZgYPYj9NbmKOXytEAroBMON0iKg52g0ldcdNcEnUmmLgL9pedd7xHVHX6S
lV15tDI+ZSrdIrpee21tQj4ft0lHyff4L1a3axuabqTgP3DUmO/b2Nr+OvC65arQxwvZNyFA6SSR
wN83+MeBih8WBW26SIc8m5tB8x4nHuq+5mSZ7II7Oa6MHAP4n+v2u0iVfxe9xt4/WErcm5srV4Fc
ATjYYIFwxFLfEX5AerKKPW+yvOI2ty6l9Bbpfsc2/ik7HwcmQ1uZ1l/oOoCEyUgjCjnQxBKdYAM2
+29e85XW5CmLlOgczb2WeMk95w1Zl3IIi18DrKa+YVc9lCp+0Id//jPoYRInYlCwVttt8RAmgbQ2
85qD/ZJ2VyJ0dSvBLX4JftgHxH1m2xa2C3jcCBXyFMjslSjiUmahQfolpfylL6f6n03cHDjMx3kl
anXno8CNOtJg9NeVPw80hUaThMZaCE1rZpdK3LFSCO+CwMxiqiRXk2D1t9wdoCGfB7N1REsXGdOF
tRmctdvSLnYU5hMOpaatyVY8ZdP0C2vwyEPCBIF/2vR2/K7kWxJ5BNGoiKZp37UzzzDPSunEyhtT
KacVJAnESZkZCtfwx9iN45uVotazrhZbO5P1bn/ZeJbQsZXFmMs6pm9i+T6XqcoQlQtVAWsVCCHK
TbqVtvEOTkKpKrhcS9TD7Jb/BvT3bdCU55Ih5Ga0fSa/MYzw2o0ov5cqrP/8o6+fu3nUIrBDnzVG
kMru6YxvEEa5zEz+xJ3W0dHDYOBxrRryqBcGRyEQVSl4kxhAQjpmxwY2fi/rt5ac/sAPGC6P4VRj
5mx5+s+YUXxwRAx8+IxjvJlODFVAPB8YV3enr6aluIESgrnMvhuoWnVT8iQmwxOSyCpsxC9DVdU6
ZhzXZhJkOofg84u/V6dDQgnp5PHPNKzUoAFR5CkP3d9r00pmY9UJ44RjXXm0wvWgWlUfBTwQZw6c
O6Bufqd5Q/4blNfNdd0iI6aeN6HQBrNPN2fZgM7TG8TnsPY+/iRgWaDUdsploqJSgm9J2qDoUc6V
bLKqdnoVYsT+m5opy1umwzLg+vLGK9OnZTx9vZ4STDGfHRmSdR144ZrbMsbNM9NqvhONcb1oc3eQ
h+n5xjDWo3bLlLB3LyId5395VR5beL84XwRK10EyMSqxHXHEvb+Am2kozyf6r3HojDeUkra6Of/R
ca2R2CZLW/Da+oRSctSUz+Z87ZOG86a9ZCGWjhyvjkuAYFVsEa2UjcDyiPBbf1Bngu4yuJqY4+j3
R9Lu8nRe8k0htv7UlD/5P8P/dG3OnN+r16mRPsZey3Hy2zfeyXA1VQj0D24FJweRYBXMmTiVe6zh
N57RYf91PAVWVOMyif18ro+zk75A+btUhTKuspvClPthvNhhgJml7Y+OOxzBnGH+74gqJdFlUXDP
MzAO+0tt5Tq32P81x8TtGROIch3RVZCi4gnLjTthAozl7XxpGrUcAVRFXsXFW5puLmClrhL/h8Gs
HgAGesD6zbiMmZ0Wl22tzI+LtbdehnrAY+vmBIDPpRTZ0D1wy8ipQP5qYo31qP0b+bxGWXZTVKeX
O3chd1vr0xjcr/3CiO0kHN2qiXSfbUc8/xfXko8yadUvgNwVxb+AdNQGRxFALW6bZUTk7zT/P3+3
3pQ2jS0bm36UQPqq7EGID3F4TIrRZbfyeDNsHargYMOGbrwXMVadMmEWG+FX2eEkKcIPAGC89NA3
mTo8M5EhyS252gCrZ3oXpTv6tEZV8BhabRFp+rgEb+VQU6IsPMaOpOF86Re/iHwDT4DQWoOre16/
D4gVC38v3nYytZI9buvBJMJDZB8Ogk8M9H/wAjCmpHLP/zPyoqzuOLmAoCrnFYsvcQ9TrfCzdUbD
UZgU0Ky4/2f8Y+wThYU3oO8iuzk4IGEWEGdu+3JIA490Yn7A8TQ9/qyXbDqnQAWvg2q28fk8VD8Y
TXm4xL12hxr0TUJOmJSZSizamuZt672mBfMiSDlb0Wz2VrMTIY9ZqmFLpvwo6hF9ijyIZpaGmbjm
u3Q/1ILJvNvPB6CaSW/tS1Ms0F2hru+HxyHnK3zLohYHD4yMkyGV66ExLIoSDtLtDGthZotY2zbT
KMNsbMi/UEhEtBKqF4XBpzS9zzfDMDjinY41BlNkYq0I2LsM8QRFbm2LN2BCW2gfGRYInoI5YS5a
gUrDqtieAyJ/L4w16L9vIDsoeV16GPq+FsCt7+8YQzCAuCQTyROs1r1tW0LugjKhNZOKDPmZBHsr
OLBCMwgIRd8fQ3ffXzTkQiAp/6Y8lWwNGqOYbHlVlSo0FGw+8Udw56Jl7Q10TGY2W3Tt7ADLmZqg
C8+CGU2R6i1YTopljdpvcN0T/PRxxbc1cwiYXB+6fDqkQdV6QNXa/Ua2XKcY9XqOIETDccwoR3RR
GNMnD2ctpkEeJowTvaJNyzzR1W1ZsIHBMUuesEpwe8/ritfu4YZJpkbbFssrDWmBYAn85GYPCCK0
SBAUjExYNpsjSUsDVouHn6AjJ1dYQod/gKH3c/qldFO/qfmo54P5k7yqcDSWDO0kPBEmJPlMlwyG
H3c2bQYoRdSFifPVn0NHGaBK59vUjV96JbPb9OHhFuMhpFsIwShBm7BfTPw6BuTj3F4ZExL1bM2p
J9/limJHHIrITCdlCB8ExLSdonKKfA9Gotkz/Xtk0Fr+pUpRlvgtiyWF4wg0TPXEjKQOnJ6XmTl3
mQri3nab8aIz5Xo0sT6C2axixGLgrmYDXH+5ItrlqIxR2SFSaXCnvYpWYdW6gJt3UXyICQ2NQ8LI
JG2A8deGGPeunWEoqfUJzZkR8d3O++7k2YxtINQJ1PeeU3h0xbs6R2YhuySn1dH3Ksqa9y0Wcg/O
UiOFv/uVQlvDT8wCqlIq8av4mMJHslLY77sTZN1kpy7vAw4Z93SEPh5CSvzmoWhEHY9+vYUSjGeg
Bopp7A/WHSiGEakgjtYH0MBcRbQxnRgyp3ljnAj5etrW+NzL9b7snrnzsdGO6gOl5HxrSrCPdsl/
7mYXo8Iu9mX3M1gsLyorB/fmHD7WR8Aw4zPPIdjKGu1q7CD1ovjzrk6aXA6mGM7dbUiUPS0WqfNF
9KfjpqwxQK52AAzHuLhqGXK68ez/F1ht46RbwHPfsffZymACTU5nc3r6wupXWwGsx15jkr3SdIvP
ed00pkDa3NlqPFIkvJ9RxImEXhMqURzGiVC1u1d4EAUj3sUDCVdghvquwLEUbeQOsUjP7ywStrXJ
Y/kWaccuui/xZE1UnIA30h5B57cPIO8Qte3lXxxd2HGvWO4IfRfDsXmzlV7J/P/wSmFEhhplaL+P
KDLpr6xY6f/gGGIl2S1Z0OYQ8xZZCPHiKXK9xhbzoHGxDo2Xh/tYQRO2tFfVUYXn2OcW+f3yNfqW
6/eBx1iruGk/hpwVuP+cje9OjzBtpumeZQQKR7GbTh1ZGLElr+q6BZf28xsmSs9w3Kr7ogfuLCX1
KhqcXkp9Pqai0PTPS+116FnD4S0H5PCjq0Bk/JYfDMqM6lp1nWM0ffTVC6O2CLaXHHAbcY6bZaPf
RyE7QZbG3tfGrLnr0qcuyBtjJzPbcUysAmDxITuWDLUqdXp7jsQGQpkATtIjlwfj3ki0+Yt60D8D
KdWCppPMn+emCyD0UMcWaHlksVFatjGCvSZB61uiWpC98Br/wGDyMjPVuVrm0g9sWHi0dxDGRGd6
DqyqzhsSWL7V10Iay+yJaJGx2REjkk5/OZ09DmRf+nBndSIkjIfCrpwT9ocQX6Ac4HBGw75Ijg3q
Pk69p4dl5NZdHRe1Nn96fuDAkM1/SICyPy5XoC8syThL3hURCa28mOmZvrKHd+hQPeFmEeod5h1S
clqD24Qy3k2FqXcsCAUudLc2SNV+wNxfQLDy6la3gZK+Qrdz2CXO0ig7dKaiIh9LZQab/sdGqk1o
YRtmWR98Jkj0JEiLmHTKgzjMDdeea6kUTSn58PX1JYHgn09vEFZtDDWaA3WKC2GvI0lNmB0y3120
/q+kWzMK/wOqtqDTRQ5DoJWi9Oe2iAQUphMarXlqEXEhsLOZtDdkbQnPOL+pJ7St3brY5kMt5/HU
SqGFZoJa2bKFnLwW+tbOhI/pQX724MJngjJ87Jk7DnmLU+zjuG6r2dtbi3KfodW6XFUAR+y/uT1i
RKDUJ8S5SJhxhglC+4fSqtjM7rG8nOQnO1LFtu9UCYVntZ3cSJDIXYusEEjJeFQdQKBB4LMqqS6E
RW8DdcxAaypzCh6QbstaZRqZ7hZy7ztMOAqV7MTpyvF0mNXO+oMFxL1BZkdSkROgGTbR59P+rtJt
FvJk4b3NWTeYA1NIzpp8kBdHxY4D0ZwyjTzqPGoZ6mrsU5qNYTB11kQuicNN1LB0u/DWTXu53m49
YkFPtJPj5v5U4vKDO5H7t+1J0LORzXzfAaD272kJhBxSNoHO+eaTwiTdrl/KbT1WaOur/hstgnp7
peKEiMz47hP/hUPZBnZO/603Z0j62S8cFiN0aP563VHOkVbODpXCnjmnhnqejtm7/KsJ7GsBAOeE
EWgxAz6hTVfAPL2oupHOPZZ/V22JZa+LPqMTykWn+Wk9op0uZ9G8fz6o6XQdniylJJPdL7Nh5dLz
wyXY22mHqoK8lbv9ApY9pE3wNdWaxGKN69HO/HMFumbl3YgWCT3CU70wDB9tezZCkufh56M/0Jx3
ZMbUxasYs+d5XUwgvXe1uCzcAhfvYIPANmyIIFu1TFDOIdaOWvaY51NMsPT5sMtZGsxiSHlt+wPU
UxJkje/TGDrXwP3ixT7/bzc8aov1tWaftxnyEeZVF/rjorL8ASQZDdMAdqFRgZQikDF+jpeSEPAd
00tSGpTHi598QhAaG5sxgTrDl2GehjJgmm5AyDINC7EoHsODjuuoa679hFUWoncJ1LQhomy+TSQd
tE+fdzAaalkEI7at7qgIdr2FORDtHYZYWj43x/VTWv9BXHcRElBYfD05Qbs7v3boIzTJNTcJjLPh
aNezW+kTayFF6EB2uTiLYgl7VO382pdz9IaiJ/HJn4M6Ev5cSvBoOzTduVtcgi8+ncqN1LRz4awT
mE6JcHdd61XBknLLQ4x6dw8qS44l3+l6Ye8N4ANHp1PkauR9yidhr3ROn4+1R0lu5HFw+NIyrbNw
5CEPpCW9l7ntTaTlYbShyzLn2WRpo6B9PKvR5lJivcuSX5HjF088IerLFL6di+RS7I4iexE2WTwp
8OxGubC/V072lLpQzQXz/CWPE8UaY3EKSkQlA4wcOCMSpmTlL/N8INGUoq9znDUEvW8ELtgE35J9
dOEn/q4Bk//RTiEDqUSDKEToxDjt3RMuMueJ1QKEC5r51/1Ji8pAZZYtQfCgLhuJJuC6b7qvKxHN
oC+wBEGM5+nHsrIE/lmL4zROqeecd284daagJ+oYBcKuaDg13P3doCpTDS66Y6m4FtO3BAMP0eVm
pLrt3J70wB805GG/D6TNQdxN8tbbGNEGvJdvPB0Yi6m8d3C+PEreIjUxxgeYFV96TZWE4fXtzcwO
3vzYE+dgqZRpA/dmkE4RQpLQwDBLoMM6ScfTfKYbtejxrD8zcLWgVyGVMbvC0rf0txlgt/3R1RG+
1jpLxjfBiWMAr7We7G7pVQCsVFCHPgIJgqE/L7twJBMdDJKEt4F+nWE+lpWUYMFSIOkvGXF0i2S5
TGbk/BlGKHEKGWHZazGu4xoyqPv6MMcHqngkfyADz7EhFEnE7Pf7HdV5hMDjnEkf9ZbQKZKXVmeO
WxMbIvEp/qVyMUL98Z94TXj6h84DrFxNWFbjn1FSM8SOYKhD5cLrmHACK8wYi0IvllKbDRZp16me
I4+qN7TSRIzC8qmRp4H6CVUh7jWEtoiMZtD21LyNfz9sCDL281I5B+laws2k8b6KgOU90mACNg/3
ZjaLHPRPuPAcNReI9eGv5CAfQOJKvzdwvLZMo+YYKDj2HGr/gq7RaIVGBR9MRXzmiaO2kKLxho92
q7nFpw4tGb84KY+SzIwffg05IyylbAn74yW0NvKY60BNfpZMka1CmMAuvQTHpnYhhukvjqzBvfCi
7hL/ZW77NZBTAVBO7zi9LbWnYYKCpNf1I208rl3Y/9yczzTwrlwG0dK+d5F5B5a38njNx61AmnVO
lYmHgpQ9zPJBdtHpfxmXWolzPQUaXWu0Hqpnz4BwXg70ePe+dkLux8Ced7onJIA1txrEKqm1v09P
OE8BmxsDts/zlICouezvb1OvheHTqLpnF6XPsnHLv++lod6H1IYbxWvdQZjGkyJ8oBeajrFDrL3L
ZUPbAn1xE9Th38CUu9luulDUa2/2EkvzNWDAS/FZfTLKgktHkEakC9HPAV9e7BhvIOPvUVWcPj6j
iy0S2Bqs8ooEXdIdYhtV0Iwkb5R6yGc3DyXgDncY39YkweZ5XjtkeZu+3yN2Zoz0Wekan7ERlB/i
LXavzNr7iay19r+nkLCqMv47rJJVcazCYtg+H3epsn6qCjTzElWhWUuIoXi967rkLz9VUMSErtJN
b+CgP7KHsGXHwTWQVTCvPeyCtIEwqP8jHwJFrB1fROJ7ZyYJgqvKgEWujfyIB8iGns5MTwB41s+q
+3K/HqG9Vf0zWwEEwpS1ebV3YAR47PWrHaXc7ogB9i7/ObM6BAhhda9D3jKuTO2bcJ85BojHxR6N
wgmow0jq6AFUs7+ZwJb2RCcG1DoKsZ2V+JivfCxSE85GOjqlAcCjbEpPnY83jsGLkN/u2zO1EQHe
N5kLwzLQjwFZ9w3J5CEyJfPW+pL5AoTK/bP0I19VFtePlf5/8DyKZ/7aed/EUw0jFh7Y1Kvn4Uc1
8waJb1pxoGiXV1h7bb2YRuwwtnQ6q9tv3Xo9PHOqotIZJsCnSQA4ijomZXarfQx4tnLgF/SBlmUB
Q21LXuK3uwz6IutEbMFYzeON+WB7lCVue/lQcs9h2ZamdyZyaPJ/izMGkxvxonOWDdqXwhxYaVZ4
dua+DNjlFB6Vk4GeuqftqEcJbXDghEDM2DEnHJiyFQEFO1ewOEsOuBtvwfaqyZfSxbnsiBSyGypP
Gr6mZLuxiIsv0novrwqJfvdg4AVW4VXiZ/dy9KqfJHyFXulZpRXg4i/4t2j9BfxX6FqpddUbL7Fz
G7Welgw3UMfOOrk9hEMNHnCZTqIQbPe6wZ6MIfYQt9kuyB4YZrK/9nG8lp7+aPXEMKntan85aOTe
cEwDcihGPbIG+7SVf4dm+4RsBmissvfh5Eoc48Enajp+03PN/o+SOX+dQbi77j0W+iC2eb0qvFOx
uX0wx2GiYniWO4oSLb4D2UofFQVsFpjhT25/9c/uLJPuVYWcQy4uruE6PbuAcBU5YPxrTnHy6ndb
DT/TroPzeycU0A6RLoYDW/1AZ1Wwe8XUm3ftuomRCtpe4iv7fmVzSrwndEdtA466Lu/9dixSUKFh
IKO3MN07XrmlSlyKFIfPPPQ79ZYcc7fKYD1srDd3QpbbANQP3W5y6AHcV9YhDb0OnnfEtWBEyiY/
4D8lV7auDyANRCrjYGwdLQBH+Byz+e+OKsMdOntvp+YlC4/+kV3c1a67+fxg7oovKCBTFcqJnw8W
AgtBkMRY1oQloGUfCoh0QH0/cTOwzcJ6FqIasSU3IVG5CK0o5BvCy79JTSf4tFmIutjS6772zVZI
EWdnZTd3YF+lZ+V7WGnJGuf0m7Oq0QWCQeTW7VdgrxW2t2k0hNqXy11OnyxEtqNiVsE4ZOtbnbxO
+GP9ADW1/88xCGra2nQRd1544ZqA94nqKGe9LhrS9A3dnMjojWsowG0PlnzWeDL0yxYkNb+T7w1O
oPu36JfJhucnGB9nTOsUQz+IT2r0kwq6n21yEDSS0dHPXpVfAVN7uZ0piwbR6n/kj+k50owMqI8b
l4tPSrx62Bl3D5hTNuxXBwtgc1E/eC0avmLm9MIjHCa/bU+TJ/zi4VK6i+E+qZ9e86cX+0RSpHQD
tlQBDkespDt1wfn/89ectGgwCWt9Y/KWKxhHd7j9GWK5yk5C7dmROzR3qontgzOQ9Os84KjPZFWx
tVW0Lv5ykCzaAwue++cBDKiUBxPZ7jvv58euovVYocrBkKg7YpID3fANsFY7lj64XHKVeMnV1EP4
KB1+fcBAVKzWRfVeAQbJ4nfsIYiBKiQgJJ1fhr+xkahVQuKTYokwU1taDBpemcUjFUdvjydoT/bL
VGEBbvngqoYFnZKzmcNiHd2OB7PDRA1dZ8comd/g9eQmGOHouOjmmXdVUM91SpoTWhAQF1QIlKSR
etykjlAy6ozMIFL0kNKerLUFKt4goumXFejxkSIWnsiNfDF0w0V4kPGcDptE0QuXwl+C8GHgwZ5T
2NYSuxKzE7yX20lYMluSRC0Jze5T9ZfEA9hUHFdoiEJz9Rbo4JrGsXDT2zT0KJCP0Yy0ae0jyNC2
VH1EQWTDxubnBvxKkfQQnW2AhynBBp3DPq1etJQJBNstIUVqVJSSeYpZPl27u9TAs6kvf2QmajA1
EChZ0s56wYMC0Spr3N0ASWAvbvPqyCco7UzjsQo2/3BU5dtkxSIloYVzBYXZSc8K+fgnIraouHvW
qKtWupknzdQjpkaO9zywpZmdlzwrdC56nZ/bbDGf43yj8I4lO5kebz3J3yB7m5QeFOz98tpZUJev
DI4DPr9voS7EuZOvoND8xT+Oey3wQJ8PE18ws0mT9sqpdeC2mEWLuEk8eKfwOyheZNEL0JJEHb1i
yxBCZEM/psIRxqwn2JmCATEjSN5mPhwRzDFzWM9OgaH5Vf6j9IIuP70BKe2thmyGKWxTEgXWG5P/
1xjHfddv6RHWWpLoqjxMlO5OWczSys0fFUbSr3A0QXFbQDqwlZT53oTrMReZ73pyfn5Cjw431MXH
mRYmqJ8nPQ7R2mLy5MdNVR4Ki8Ei1KvVxWA5EpZTVOFkL88wNH6OgzJLXw9UGSsjRdg/rGm+EaI6
83aAn1aYZdSKRpPxgWBjqNtFUIFmECUZ+06wBegVXKLqYfnqrNdfMBrQec1NLiL5QaHX3KxwZC8N
Jr/tdlG3XrmmJ/WbSwGCCO9lFPJfo52r0WEJRQHC8CsGftdmaqWtneaRwNK23OcjQEdwRVNVBafD
d/Cm4EFVooz8zm15nE7xIu4dmaTlB3v2d8EWBxqgc6Ts4fHG73KgjytDYOttMlWkxchjFo6lAaCT
QbJCnAHtfU3znAQjJxtiEWk31QI6SRg6QhiGFFs/HtlyTQK8ODpN8gbVlk7PmB0msdiQ/Y6K2U8l
RB16K3YkhitrSU/GW46uYM9jE8UG+9Xt1Pj3vj5W7L2yiyyE3fa3j1CrVGrHq307L8kkGjDdbIc+
uxWUFlsD1rBYpFwjw0jh2vRfKYBqyIu9l1/BC9m+wO+LEVrnTVmR9c4+dA7jxkvaYn3Of+9RdYn6
7/8bU0KTe0yQ6Db2rPLNdiZeLOg7QFLb/DxO8RsUEU382lOF5iTbzOQHx7vUuWx9GSO5SPZmWueT
NasL5CN1vn7ItkTkNew0cODGPARCgv0dqcLoyHGrdRF1fJLk8TDxIwEWVyb8DGYXqusGZ2YdVVyh
yBXGOZ9NrNtqUH0SeqG6W5lH5zEd3cmyto+NHLzTG0GJGdbIyfAMaH6sD1oUGNOhomMMQbW+MJ59
h2Y+G+waG8cWroVFFspUk48MO0p8Y4EcBFTv98P7goRNCF9hjSvWfvQwZj2/qvzx98ABulIrKdvL
J3oPL6yAUUeC/1AlQMEoh7UVKgLxIatUSxYSGxoi1a1IJ3L2wR3xi4u/owzvOtgz2HFiy4Fc854X
K3+/ylFaS5njTU3i/8cdc8b6HfsW27mpFMRXbEXtuDNaelInYvOoS/uHucOaygxBuX07IvpmoRSF
g2K8DRfjX/8HchaBu2bZIUB/eg4FiJuLcbojmqhZBe9kVuARysrmwDvwPcpWRTqT1Qc7qiyBk8i9
/Oyfu196QMer7POn6fhWg7mUc3r6/gna/ey21XI653q3yeeKp1vnG38oNJwOITZcsD/y0gJ4KBEi
illDQmBPYsWQt5v9QEZDs51fSndOQMPyaxclGmFBnEG7+R1RYP2esjQtZOForCX3lHgshjdPlQ5Y
JScPbfjIrOgM2c1TITkDj3XFxWeLfVwnyi4NLwMWk8OhUoI8pHlZAOHcRn1Ge234QOoOOUnDpNKQ
0dERNsrH8teFXq/pHxWa07QZLi0JAAW+rRXL50fY147Jg7SZcrd4IHf20keRrZIQCqd+HujhbTCK
pRayj12x9y8I1tjErR5ZVemTLXoQ9+Z9Q3Y/wcoMW8tFRUqCtEFTPVZPy9C9ncQZaVir+RguPjdp
pik8ufuGVdZVNZIt6VdJMJfxefLnlHRdKCKxS8ELf5wdpvwMRnZTpAxVhzUXynwPobWVLiu2bhwn
AvrkOv3pbpxQT3sIrqxvQ1cCICfFQQH6I1YZTMnzLGHwYAy31n5/T2i6vj1dSNvLCMratFPhLpRM
/PrjD7CleKta/whWuzTvJuQc5sC+g06sSlnTk+kJlASO4Qej3TNzIm8vX721ED/F2MkONmc7uvgL
S8pBYAfSIHOHTihayrpchCy1um3qh8KXJwHJCc+4yIPZdyRCWlpsgyTVi5F47630pcAvVa21qj2a
V1JfBUsSkStj7hCd/MC9ApmTf3aD37ZIiXs7dBXzWCThyDRVxw4hNYOUtm5qY4JPcP6PPKL7r5GX
fYNP6tb4xQRhoVWIrhaEemWTcINiyq8oZtz+xjRHY1hWxtIVA/iHGwxH8imADfulA1J8v2uizMPs
M/YZsLvM2NWt3fcDxEJyUQrtX6F5hPzLBVOEjCU+I/y2680mYcbiYu9tjD+PQ4kHJNoSuug4A5zn
1I/St9+3e4AZfIUunLS7+JHf2ONJI0a+zZlSozgsF7gxvTojLBQzL61WqV0H9HTAknuTXpdIjB7i
TYNy9Y27Gkr2uK2FIcspHdU5gdO47x+dT033Cc1pZRz9piSoVxr1PseqHR4Gj4g9Uj+IaKnA7m1t
7mSSJbTQ8inJzZ2ykdncMYYPMABP8rig4CrCTnuP4B/Gb6ksI4yv947xbI3oBzuBIOlwqv5cFj/a
EBQuFFpHAvC9DMsCnlFcGspEOXpHYuZe00bpMnEPNTSy+og83PU5Xboxm843x54XQZEb/J09b7e/
a5Xk2W+LxPIB+1jU327Kb1J1hQx9y+4PB+nagTF8TsfYtR1etp11z01ND4Ej4ii8++ad6Y5jRVhk
+QZVZKkQirYVGATDCb2Xq18vVUqdq7MdbbEWaQgUXPcpElP3gfk4j1aHIPGJFQLggI2TO1oT/T8A
7vCFKYWTt5vx8bWs9tU/sJ8rGY+QWVDsH5BkSTHFoGdzq/1AkbDrwm5iwm3VJJOjk9w0gm2B/bJd
l0Q4FgR3WnWGo8DEGSi+zKyvOrfsAKX67gBXVJ9Q3/8A15+Ke2AmQ2ejH9QDpC/R3RfTjfiwUDjJ
QfhF9GQp2aRy6nJf+1mq+36Lajem5u5NA1cTWNSulEO39nRqsDiZHzKW7Q0skaegDOIqetrQDA5K
qh2PbFdDQkM/bI/JEZk5K7S+AT/21A5984wI/OhRK4uyslfZZfT/xMsk5Hd0BKMopGpf0kr+ORcL
Gwkj/1tzN9xCiqe5pvCpUlt/jedJWEOHoDt/M0R69wJrU8TrRuL5XOeHwduN/3EYP2KizL97f1C0
8WqPuARE61ESiE3/AM+9aqmuH0eSBNldO4Y6wNKQ1kWRWr/0ptME/aXvK/jiDrY2ZK8rtCBBD64t
vG1I2W75dgfkzl3CvTythdfKn/hqvrbPMu/DXCH+EJCN/LIk6RzSX4708+5LTiDSero/4338I+4V
bPUDaGnaffcxd1tFI5DRbMxZSakUQVf/v7yJaApYIQDFOd8o9/8PF+wS5KW6gVAtFS5436h0A3Ga
Rtw1Pkdn92AOI7VXBCjdW4d64cHIIL/hN2eJ33CBcoBrbYAyBCZpH6+6eyJIwofNyEGpCrJ6wegP
pxZSEuZOPEFD4KqLNvg1Df3QIWtGdvLcP7GP5GRfe9PQ5zBuhULe9vYMhccNiFWvc1Bz9V+Ry+wP
dxuusFa83p3LvBDHT0Kis0qdNQLaCahotFmhYEHZnITCBV92ONKn+tSR7wQLU7SEoAEvJsh1GTAf
DYQpnyMrH8mx09qAl/YERrJKzSgXDx6cp1R/LnbkYtRYZSh6NnbgpC4OaglOf4h0CjV9wZlOHp+i
+Us9FmX7JMN8VL37qEgCViSe0Mqqc9fpEol+HVM1rKdXtxfpR3jI7Y0u4wcao1k5uIPnoD3PZB8C
vtIOB+pLXpuTnlqkndW/icswLN2gYbaOwl06oNOZHxeDQGqC/MkHpihsbPFCVhgZmwtgf/CKUQHi
8IeA7kNC/DqdKEyBisYFRSW/Rx8FTaltx30WoHuHuqCqIxfJp0+tVQ9E+YIAKGYzoiR/9BZvpWzz
y61eBUJ8oe+XcunVeLKWdMP83iLtkDA9vEtF9mfX0+W44eim7Rz8JFin/dbfUDaKfgnsZrTSCaqF
HNw2Em0LZVr5NzDYxQm9pPNscQi/cKfsj4dABm8dUQEHfr12xyoYYXHcJmWEBwhIFNLcFt5/wTyp
AQ5905q49adYl5ZfNthM2EvID+gDZa2d+qirh79P0UYntLwGyrMutuhf8+W0CBo+uplitjaOM63n
086Anxpew2CCaOzTMESTRdPZbrvpquVUWBYLH3aZVDMyuEcTviMooaZi8oj0akXCxMpkMFVxVbcG
5FUU5N3Gc+61tINHoMwlHPCumVIAkHEJq268uvKUBMQetNAcchEGgT44DW+Qd5zgQp0EswGdVVSA
CDDBqudlCp9/EMyVKuOtkKhhlWNqtSS6miMLiHZu4uCyLNKSXMcssoiprtav9ofGT0ivIzUVz9Ae
ot/6zWFej/r7BfFJHIX10QCLMENK/RrJbdqYtluIy64bxernT38JS94/JlHbTrXKgNzEWwoBHRR0
2i9BMG3tuFwsi9c3ZtJ/dYiRGQFrpC30+fEMHln+b3UOMRuCVDBcWjI/AYabrzl0Qbbc1IhmQJF2
mkuxW+trhoOruL7VAcK00cXPrK18jJI8k6XGS4HgPbOwQAi760j6U4S+IhbSm7IOXP8D4hA5JsS3
0qxlKGjgYil5gRxHGGeR4mRdEdN3U+GEp/gCJY1y6IHbwdZ4oF9L2ka3Orqz+ytzSrwXhNsmOH+h
aPWV1ImdY3z6YUjnJ7mPayViiw7csUIyLJLZKbbt8tc/0+VoHZTrhVeLWAJqCMY1cIpqHZTxpuG6
og9pN/5ABmY8/aOwd00AhQClw8OepYWUxu2tOWfYGG/QojnpqDBGCvEzwyFJAiyHFjr6XtJRbBAU
PDysztU1s1BptKSLUktQ99+3U57CwFqQIRcmAUl+ubllbLZf9Bi1pGMyepPEGDO94GLi4OpxIFtu
bg7BWSYOfoLIjjatbrwH1tIuoM8ipXwetE2dO2AeQus91wo7mdGXCov/5CqpZCImJhsb9pe29Jcy
xikPTNhAVJ694ggVboANuMjjABZhce46IxaYnUsz7KA3/Q6bGP3QR4GBThd3tVgKRF6ielflzlnM
F1Uhq2zn1aL5geTj16wsxGa6aFggSttY4Bm7nBRDGAHHLDD4JWo6eFiwMrDqe90XJpwuj4xngLdR
/eDC/aBNMb7sRKoTUL+bXgn3OHrDyRtDJlVI6iw4c+sXLXFt85FeLU1iiTMP1kjj92yXQ/eSbNem
kl4SXKiMQJrF5Laao5bBTI/NQ52yjrnN3Ssh21PCpBXrOlJgDcPuqtQhuNe3rfY0dstzzlTw0Nu/
dg1Ag0kzykpJ7E17z6beWtdO8WSXSfoklukGeKtQ+4xuUxOi53xelnVSxhhkrfKUbB/xl92xIopG
+Aidkj+FHJiHvuAgpiyUu36qvUXFQX8PS47JW7MGxWyTYM6feltooyU2Q19iLTujtcxNplw5mpcD
yyW+PS8glrAsz3sgHgivURsSH6MEb3czJH1vos8LMIb1GeVxZgy8Ckrj5MuQFLh4gCARFfWXxTsR
6EC+x12eGd3ZT4DyWCMaaT2NZ9lwD2V9mgNMNg7fCbs102tTJn0spL7vk3jx+bR5yM1DS1uuMqKK
d0wXeHBZmg13xzERhwuTKmj71EjbsmV21Hq47HiUEzlgg5Y6Jue52l9DRsrxEWQT1ANUakW6nzKM
H91kqSAySuVAu2vVOFllmRLvZAJvEvshl1D7Kt94crTDvMSwSS7dAUCwIQmiwJS+tbOZoHZaO/rS
QTB9fmzNQt7PB7s+IFjvhVSfrIHF3izg6++NjH+LcglJ4hSCfeyF+Ly3BPvOSp3hGvPjkiZIhcnG
b1WIt/rpIAhI52wVhneWuOZzVv3RNJsLIEWntp+2lEgIWmnsZr8b5o75+MJEkO2w3+iXn83g1Fxm
2Rgle+nErP9ZTk4Labbt+yI8l5IGacQrc34YS4DkWYWYoYCMHZGkRXwgiaGRrhF03Bt2D8BTrL4P
c3lKuefMq0mXOqAbybywFyYhq9RG0FkC4sJ6SuJRWlrGDC6IulG/Aj4ek/wtOb2HVDq0tm9ntUvO
3mouAFKvSXUTN1Dnui02rjP1A8qHqJoyoJXFM/OpR1YVOPwcWP6u8uYaFExS/YrSFXNen18EGW01
WKeKGrkDFy0HxrN2WDyVsOUErHrXo4Pfo9rtddk8uXGmGwrY8odT3i4NT+soTwNqjh/SMgPSsg0I
rft5wVhbsc5fxLak+GOBLhNr8/K7hJau3Fc+O6Cy15kprFCFRNXXnuO8revzYlYWoyWmweQX/GNN
2QEHYyrQmrpb5q39Y5st0WtcDxLXyuxnnHoBBTROPdFklAmmRwRd311jnH2pG3l8MV9uqc9RSinA
WbUQuvI0sqZ610UOGGcyCeQ/WbxRF+uDfagrjtY8X8OjEEI2yTGlB0fWyP5GvZcvDhwRrEXFArf+
vpWZRN1DBBU/cNOo3y/+IoFAfUZDmnD2hwlWiDHLEZ95vKHvMGXB7T5VK50dbO3+mu6LsO0bvxWF
KOn5QraPAE+l9DzmmNhrfjdlp1d7drjAGCywqmyLqs+75TOXzGXQH9dHMotdmCAYmjSI938hZwq/
/tx7nsxBZl+WrWQfqqlahQ565cE28apcZH0mFnRBBM7WRB8qkmUnTmSWXfLImciAt6JHm8Cd2BBl
zn2JhCFGeODfz6TJ/8OSqOL+eRDghB2zLD814pWevKaCSdAc13cpM+HWQkNTR9NB0SJi5iXL/rRc
sRr5nxB5WfP5pZCcdhREYW0Ol5piqHVmWS4GshxgQ6EdeXOvhNfJuBsmc6P2AMi9GE1m3YKT/g6E
wxmLSmwH+AFSJLZZ4liovBnm1LfLB9vlPr+UomOYdkUZ0mnBOfzBh5ZWr4D9aNugqgxVhAN9Ss3c
X9WU5cXFcwMSTmfudcYJlnUJrJ3bcephMSaWfl9ph9GdMdrtZzmeygKAppa81Vx3vXq28G6T3Upw
QDtyam1k/2iOS5sXcLTTcFiG0DhWTFDWYJoXiaUHmTGR4BV10v3Yb2Dj193r0JuCC5V3cgr8bfyy
oSFF3FHhe4q/8xP5mYsWJGKoY9GPMVeXboCSNFvfj93UVCnBsmBAxrBoK77FpQzdApVtplxSoTO+
jvPZIWuS4YNrjkG8sL6PCvqNN8SolJJE0ZZnsi09s8x4g/xaxd+LEYZHlD17T1MBnbhlkChXspYs
0t3UnopVG5NR84NhaYuWqFIYrUhgu952rGv0YglUAKHL4KkUBCpEYSymaqKfUg6nxcQ8UGTkHCZ4
qw6kWO+bbUDB11WrrMFSxNbl8pqS/mAmS9QAh91ITe+RM+jjOfaSJD16HEfmDMkEZDpSSw1fBLrw
7bYWoA+M2+qFE+kpKrnZhEyTEd5Qm+5PgeAtI6lVkU5eWNMOcnFo3Abdf6tPccAl6LZh5NNcJC7L
0RzHx3Hg5eotEAnTaprPctHVtPncxGv5ScBiKd2RvODvM56LQh2HjbM57TahGt+6Qy5IDQgwCxhR
Ir5tg5LLcsuYUTFDp/+rt6zMfQmuseHxmSST4PqdhfAzNenljz0sI7PyD1zZqiddvKAZ6WB4YOy2
yjXjAHQJIRS4n7+wOPBSoRsQgDfimqO5aMs8AfoPWxp+WZfhvDy9j8DRa7v30gcG+2lQ7DaiFdCg
6hYVRu6JDftKzM3nm/nKEd+V7KyCdD8epFw36pNcE7L4Mvk/a3GEFLxXPe+4nPy/N2uix7TxzSnz
kdyIbRqHe2NpOQw7qiKp4DdKKb0CNgq/edwUkBZOn9ZaoLPbvc8cj/52SbR1IpzQY2uHpyeh0EvC
knpUAWaLO+zfHcV46b/OS9UEjUUX6n22q+X6KLK/hco4Ac0gNybwE8ibY5j5jnE0jxVfHMCZsNSR
YMUzNBn1PuDSV43n5QvjY6FxWGJKpYxy/3crWyov8ygyxQYWcuc4AYKMXlSM5u0vg6Nad0K78D9W
1IHYmj3gO8RNQK9AuBp2g+V77Ke+NPXJBuDqe4Hd6N7cy1D/OVu4ChgALWtBHiKcErlyKvne67tH
STghoux9UWmyVsrVrDWD6+AOLkgMmCr/pZA6Cf6XJNnmMG3oIE/GPU2LvCEb5hYEmkf2TvAPJbTT
Zz9CIMFYBBKia4snmE4vwkpUdzIP5ymiqbsZPg0lfKoFN/8uN9pbYt2adEEnep5ix3z4Y1uM6W0z
O1nJ8tPNFVL+VMKQzTIxkYF7+N59WPSZzd+9KKnnojnyHdYhWFKXs91Vh5mgQilxXEdW56dZRznb
dTnAReLN+KIKwQ3epKW1FqjxvAvCzwxgV+4mM7ElHzORxmLYyox1o1xjedB3QC1W/lLXUCRKXyoc
R++OMG+dCJFZ1EtYRiwIluHGo5smOOzqd1fJ2exOv3Sjk3+QvkYuo4fk2JTRJOVBZ5ldNUk99QS0
so9wd7ghuQFZRU9rwkrA4C8z9N2KZWBivK3/Db3BaDUH1wjeljxzsnAZGxxCfYASrM1NnvjYvDDk
rAYV54EWpp0Up4bz7d2XDK3nWmGcyJWBuLdxQEz7rxI6aAyMLw5hIYl9g2BxBKZjJMMhcO0Kl4KQ
ESqZCnXcgfo7qI4HhR9xI95tGE4sI2BJCi18nQH+AlkVFO52UvG8sPguYM9/yXCI6nZdkiuWhpA1
JsRazmeXUZtzV7K9kOdAmND5OUwKlTvwO5G5R+tPe7SSEwFEpO/4JOs+gbg22yykM4prGMKeSnfK
KuLzbf+YXn60TB2PBSGum2oisiR5+3QONXO+u74MYPrOmtzJ+QqOGbojIUhftf8INv3rR/6P5V6K
tFiXEzz7PLaME/0ZBf7yOYWVJFMabdJjsspq0Q+3+2LqezSvIeyJpwMk2n8OXWIAkRQ9dYK5P9IO
ju+bDg+ULep/E5/ic1ucKYRa9XxGKXMV+UqJEOzxWS0P/uLRCJLniZcfWVwF7G52Nr+4lj+gCSug
c/PxwGsetRxuEuHeaBXMPrvXmr7zgnkEJ5Fxyt4r+nkGke9l4ebrM4KbbFGz2gqhRhRtT3u3TEb+
0cda9CyGfWYq0zZbzniEAp+PjqdAedw8FX+B8irUHjkzteHxNHCyyM+Ycy4vYs2N5mOqOlGqbQrU
9TcWCOdSX/FOAEuwjEvUEqFOkRZRS6HQsMHbGIxlXoxTIGy/eTJPjLYxUHXMKMZ7mY2qRvjvFApk
S5gcLCllFpJaIxPewzkaQ1/OAV8IZrtb6vi55XaQnDL86JXCEb4iW3Q//uwAWLEP5HfJEOEMfya5
0CHLFq7XxdxwVZJvpFY5fGpxKzkg97dUXQDRjDdOxopaGU8wuTVVeclP7xQN3NKSivpKz9Aoaz5F
MXhEFEp0wSulLVn9Sqq86bTlipis37lG3ZoNYIBSioG31WXEh9pKDhC8xX8FW6yfxFZectWsJ6cD
QPJWysbrKBuvW0pq8cmpoa0Wb1NmwUiTS7yGJvdKoGVDw7RoodC0WU1GTz7EpkOwfQwGfY8qG/pD
0Sc5eECUdhokUTPMC9garCIt8Fq5xAZKF5UEx/FJ3hnsk2P75cWyi51iNLg0W9s1EP+MgaIbZC7G
2o5O0zzZKdfZfi2gO3/vwpwQWnFtVhPcxiHoCVUzbHmeaxBToU9c2dGN0k4TvTxzZe9umMYXr2DY
4ewnC430ao4P6/LeA8vwwmrVb99E4rrZlORsoIiJmIU8riiUZufm/+alnCtGDkqz8ImqHSEmAzYX
/+6m20NPxT1gyZo4hDjb0IMV4hoX4kb7xkz0MvUtUpQM265U3rIq5E874BM3pU6uDvPjXf3B4l7I
xJHVDEaoOb2glWZsaz8Di4dVoPVmXDvq0EQu7W6UHQpqqOZKx9GFZiWVjGN3bWQLreh4cKAm8MLr
tQqp3NWBofTrKZPFH8ETIXjPGBo9R9aVxwXzThv6Dgxcqdm4NKugxOfCI1qIEwoc15tWTXKyvY7V
13nsl3u83YI4vqUHfAmfEgrPtcj76vofIe7sL6vJ6qRUmDJogj5cDM6SgIeHTpWmHbGStidXG2qF
amfgOwFxz+RmkfCwf6ec3MN65R8ZHRzGYX5TpFV4cX/K9dvoUDDnz9B+t1ueLGfSSPYiqk79htVk
GTRKzjNI/nu/dzkh1Es0KsnJ+d9G8KLd351nUx8l6M4HOI19KTYImL5wae1MgGestS2paadUpl+7
r21sOZagfABBWefjUOn/BG+hkN3A0XLg4oWvJouwH1eocmMyP634rhPp/Xlh9BDnpMIvFnNb3hwE
BqwR1OEGIw1P9yN9p9jdZKVLvBCQQXgCcknZmgDlIl2e6r472+1zU+RT8zDp8QNHmbL6cDsp3O91
6CPkGOsDQC29PMyAZjBXFb945D/4Ev524DHF4pnYtwzMTdcDsPq+doe+8QjAjfPcHiK6ZwMQIIzz
2b7+9gbaIvqtUJ/Ozd0mncuasL3yXWTpeJAxmEWQU/LsBxldpBGZYXnGtdOJ7mGViZ3lkTC2sA+m
DVfdKWluYRUKpJq4x6QGEbjcinJvT/DLID1bfl30WtPAEpJJomv3CKK9j6BSvbt0ar4rsV/cWzKK
6Zo4bqp3lox2k9AhhV8BSDltYK1c1joHPzQuauBq70Uf5XfBz1vgeG39R0WnDgvUIZfa9LzYIhr0
dqF+D+fho8BkFnYGeK/MmcQh2Wvikr+khbQlKOCTT0ReYZrFu4xbEbQLi+uwiqegRkVSsJ8rSgSl
x4+v3st8D/kWlmXJJR2wmeouIy4g4CctTHpsc4cohSE07OzLvSrUsf0pFh207ZcVFf/o8MsGT0lW
S/Y/OWhsLDfVDpf37G5cngOJtWWFa0j3RtPhhQspyEXxGA1aQAF8M81dTe9zgE0s5pyveCsoWROo
N7p86kstkYIATss8F7WexYIupO5Xt1Bw5ngCiZ8JQsiVseGnPm4QCYyDLe3LXGCYCIeL6ZoDLtEx
XLffIRFEZZ4Y7E8BOT4JmWkQu8UZr8LDkeSV4SfdD8wK0tj4r8wgdJNoWAHEFZr7+iKuzk1Jn+Oz
b0OwjAN5cGa3BdaLsWr4IbvpL8M/F+RRvAntlyoae+K6+YwidS51BMQ3Pf5tyiV7melnPE+JU3cG
84rjndOxfpQ1QJtyp3HGWUA6NWL1UBTeXOz9YoPjpC4d+cN/Ne0pBSWCgt1NDjHZrQvqBztNhbWb
Lg0nJr/N8NOIUCbSgD4mostqWQzbjSs3D94nx3s71G2LO9aiXm0pNtA5eFYCO5ZcR60jEqLO14ZF
O6rDRId3fJ9OgRsSpvwgkMCiGwzUXT+Oxt7Qc6kHvh1ESt0qNUDS+9KJCX5b1FQp8ZXK6F9AiVXr
rIIWOEXbsBvpFwz0laGZAnZj7RI7fRkaOnBCyifczQkY/MWhiXjzh0eXH/igvseNhw9ksfpwdvCx
Dcjw+U+dAoKn2qP4W8VeafZJKgAyMMQF4/9ZCjngCpiPX6stlGU2f7SsSEONFqObqb/DevzbpI9D
DS+TfEKk7HlSyhnE+s56wB+HN50L3ZJTvyIwWSfBY2b8w8Tr7CJ8f6OgDMz5Bleaux3OVioYFsMk
c00O8odQmw+ZRrE9Dyc2oypVN7wtQiqXrzTknW5PilM8zptRIkDwAtWB5zpSTgCRpoXhRU1N7p76
O90wITreGSUJ+EuhATsX/0Oz40X6Zw4PozQow823XfiQ+dMa0JdCMmjSlN8ZXap4rUitKA767zjK
LQS4JLPexEdUvwtq5xXmhpLYVMAlv+L+ODd+BdpEZloUrdgKvq8/w3SMIQ5ml4u3kCHlf14lDO7l
aK9uT+jA3amMUnslyXhsvG9s4vrJYUed9s4oJdjqi3roFdrivhri6DMPQbnJRbxR7IWiiVGUTSzl
r7ztVbvMB22THufN6Af+ceFff6AvNjJuOi+DqV/96WXjOONaNOhruNlHW3BmBjkTqdKSXi78vbTf
IQtQjBejVw0EpCJ6It8WXDuSZqO840DVSY70TKDb2hvD63ppKLnQ/sJFqkQ916lmqzGEgMh6zWsP
9flByc8XxpuDaDY/KE7OqmOn7+LCIrIritqHrKPBwhIiQYtdgSOlUDsRAHPAuaoZZYXsROx6yo+u
mnLrwAFmdtWxs9Z+135M/p3LF4wWdQGUR3P9+NUCu7rd5Ccajmwkbu4IxrU2KQ7gAxeVtq2wB+m7
QLDSQhbqfrPDOHOCtAqTeqygPc/T4xIEwqa2IvjBPfCB33mhfsYPPkDS1lsl3HGd6CmBnHOvqLvb
YOwsd4aoxJUpxCYIa6pUYv7/9CjutCvM3qbXYuNk2D1Stk6XWfHiUBsRys1BdsYSvX1EbQ3kCNCg
b1B9SB1HXhLKAX3VeY+2sj3gl+milq0Ma/QFr/SZbuoJ+n5BeZjykYt10eqjP0c2A6XJLeUanmnQ
7oQMXSn9t6vdzCbDE6rFZYXs5Q6A0zlF0j3qnpL1b6W5EePSxQbZfPPX++qwa+kuYb8ZDBx4UY9Y
9ozQHIjhrgClCeOe2wPSk+JPvrvFHKBlviV+tFdxQ1pV5V7Z7TM3+oxOWXaOQEuzDtghNHCqftKv
EDR+NOP8JuzGiSlgwvsKaXu6CpT+mooHn2Cu+yFffEEL6w/2GMNyNYQdeowAR8te63SeLQ3ZI/PE
YRAdEsq4IKKwxUufN98pV/1of0yoNHbljneMD/okMY1cjdkS4QQPSe7H/UMRwAw0P83uwV6X0zez
FHhuDCRyCApnzU3jSXUInEAM9CA3S2/R9VPDt0tFoHdJrWJJwPZyN4R0whX5gMhiO54j2NVa+0UU
70wecqKyMy8RtGF1ej7XaGL7Jnf2Q0YOELP9qkLpldt8fF4PaSZGXvNuyLqp635eetB/ZLJC8Ang
WQPV/hmVhv0v7BXEJotf7KaHEXQSkMuJ8FzHMB4Cjd+ccXLaO+Sd+VmmpAcX+iq2Bwnhk7c/jK54
02VwrUPE2EiVaks+5E/EikY545RK5qkDiap1y9qiURrOwRRiRKs3yr7aUtqvFP3AfX3kmAuxiEtX
+BPXv/xbU6edPlkLps9MGzbeibur9hoY1SApM5gBM5NaBvf8zPXMW0DA8Df+jZEGtx6kUl/w60uU
7Q2FL1tJsC1kEL6c7XMqyF86skU92xNeFo3bLwTaxmQdIwNKooeJvd+TTF6PlnF6i32lFxVjswF9
UHxyAKHF5CZ0uOrbMN4WIblv3QDEfjo9bT7AgHAGKr6jK3L9jW/88/WSurfGneQ4X0vJBCH5Sc+h
QYE7IUwMeql+hO7a9MkQ38WU82xYZI0mUWQt/3TaRNbXVk8BOBWxifCmxkmMml3ezoXlMX7Ld3kP
xCmHRnSX2JMz755B12pwDKkTAOZOHGIOxVK7taJ3FWA1okKIcANe5vYwCw8DhOfionqY0fiMBpwV
Wouc/0s/aCs96H0jHhnZ0V5VsvUjl2bJNJvJFTG+0aIeCGX2nh8IlBZ3I160337nhfNs1deOet72
jcTybS0ofgpB9KxA6Q9oZkJ58maq3AWxANSc6wwVSzn3tMaKBc6eiRAJ08rbR3OTIvB8ZtHkqWA/
H2hPZXrPYeR66JnpQlIPylnM3V+vE2MOWYsB+GyVdV2DM10OJxh8yt+vfJtT1jVgB5FcRpBDRVIM
swqXnkifNfMq5ptvE+5dwX+3LwDDTMVxptK5sZivGpTxl8OP9C28ftDd+KNtVmqt7C5C9TYl4tKa
ibVbMSScyo6+a3wVv+Lqj34fESWS3va3St1lmBnhHG8zZAnxn9uPSpkdLVtqv/h+iAdpmgF56z2Z
jLTeuhwfZd8YmnUNLinCCW7yeUGCERe1/MqvXumTEMUb7hY7+MM/Sabtzg2M2+GbZkGJGZNO6AOH
Q0+Io+uC0ijWVzfGWkUVRL1N0KgdJu2DeVxOyP2QSiyFBhqdba2NLnnMKEJV+9DTZ07NQRr6f3bL
NNnZW7Lp2Gpjwp9IV4/z12QatIXBXIi1sp2+gaBSG1eq8y/KyKNDvj0axlvA0ERIJgcKy+QDzDg7
AYldsJscdXgNnhHJEHnXwArTbI5r/qJGYHDge4EsF84mIWfYyAcvUY+rcuCJ4Z0f3ShuQ8zH6pw9
/iMPt6n0TDkI4e3BTbeZ2Gpzr6Cc1Vu/XxlSX1/za5V77qiDmiXJqwXTuyjLh807QR9ooJOCl5bd
5PXfAvj8ZbLQeQ4yGfaHEql2y9QSHH8yfyqxLVOR/EAOhNvzCe3B8MxoUsV5M8flmjzaqIq9euhu
2KtnzBFV/yIbSXldABz1+dxlbc8uCt9GjeF3vWxT+zCKH9pjCGvxYMXSE7TdmqBJka5VqDu3Q+wC
FnOi41vkpqbJpYxWuFtmOzPdcx48k1/Hep2SUirGVkNT6F4yMVD+pfnB4Y8mswcVkjnZHREKZaZ3
znMHKz4PNSjoLT5JuBVXpS/75Uigme+tr4cTVse1ntyNuVIhrqQjhc81EGJyd1Vn2iLn0PuUnBHb
mTQELXt+Ruyu80hcSNzwmxOiSUT/qMOv4maqE1M1Lw6+cJHzBNUkfqvAVfDxydYiLqammFZHW/3o
nYpqrmpdJm1/cmpThA6Ow9D2QdecmHH/lOk+X8tqVnUj+SCUeAne86aDfBmeOh6Cese+tN4KjzWu
68blraheI5KJ9Q5SPZoauuBuEM6QWvrJ9M3ch/fGSXO7HlnHYnJLBFCQBARMcLqc5w33sZwHEMBG
PuPPHpp6CjlyhZgxfz6JGRGBzf5Nj0nBTnt6Hm/3npYsZMS7D2DQZ98sYT30gORYlSo9ktfWJYNd
rHQZJh+iGRuogeRs6PVGbEjwr3fpi5SVaUoJrEIoGfI213jjbEhhV0u1VftMvB9nzU7C5JzSaU0D
jmy4bLO6x9zGD/GOdzHUktmaRJR6vG6aQtiZhKMCLOl58M4DZucz9bZhpIPzYt5kEo/CBkS0A+OV
zIch6iEroLqqPSIA70CVWZfdziHqV7+ZEVmg8WtBHL7FPLyUwwbRHZRnxzwoDrOk+sSWXDKIIYON
GgDNDRurMllkoxmgGaP6XATaL3q0YMaaeEkujmBU9OzDnL1Hu/oKvUsGRMaLcQLjGCcajJ8Pnc6B
2BnH0qI7CdUL0U2GADU5iGTrblNwpDhYYrzc3qUpyus3PhwGKc2rTsYJONVpYrwSCZO8ju81LZmA
Iuonw2z3Ou+udAj4epUCnvqBI3M+peeZmewMoD8nzbtj4rZJlVlkxJ3H2N6fBk7crvoFwDvryW7d
EmfJbevQad4Q7rEjm+kfmmEQLzswCh2S5EPqgJtxP8ub4GMWKI8vrVmSzgAERn6DRgDIw68lOM+o
nY7lMYLGMzFbmQSzErP0zrMEHn3G3k0b6r7+W7dlr6Iufk3pdeLBMCNHZDQ/yffzdhQVimfO8SOH
v6ttcJkJkfGf2/Rx04jvU9q10dLbFOOOu82t5oygEGl57nK5xhYqOAgJ7SK9LWRYgSfyut+o4B57
I8RVZRuQYfi/mIYjLZWWIYBoVyFxylSNUiJ/NTwIZq2SEtJE2URaIHJ7h5Ou+3a/zudLfqMTZ+Tz
yI2r61OS9Q+wsekaiESlhavHZ2maff8Rv6fsfhSxcolM10tKqw4ec1JBWMxRJwV8q6fxaUOVOTdv
fhRbqysbkOxj0O8ltxOTKg/H9xiIPNUR2R/QcG8SqerqKSQHBzhbnnr1G9cg7qNtRMvB5PkH1Q6E
ZxAwHSyOOrywfi4oeDMXuVmL5rmB0zym3AGMWvlBz39QNgV2SI/6eSQlBfHxE2Lpw48LG/rUm+5v
voPnnvGWjxqVUOV0LNV9wIiiA71Aow78xXScCYXqsWCLV11xY4za35RwHJPlR/jagdCG8t6Y8ZWp
ZrjzI+VsF2YFujxMJlvTJ6YDIf6rfbvqAhZbSuXblvixQBEk+vydwlQlCgsbNf9Em0K4EKrUUWWb
/QVkkOgYlVJc9dnXP2VzEEwj48HIfbq2KotxHRg+I381Bu5eif03nESCCMaRLXvL4WhmF7fRnvF/
R3mbYIKhGlt15dhKL0bS8oTQwNUoyjmZtVLijNmp82vXPStcT2DGn8EihO+f4933MC8aQqXyEMdv
aP53KXLkMkpSPo8AhPwlBkPqXg3Zt/T/LEFt7ifIW8i2BBt5x9T190uxl6J/2JOOuMfNQNiPHGXp
W1D0QvhJrgQV4laILhtI2/Q4N7zmaRHu7pmWGNjAmcpHGGyhJ7iWpSjIelBkzS0BQRfpxMFwDNXz
yKkfjkvEf66rp4XhiPh8NQMFFk5UQ4wexOO5ql1fytcsuNI4Y9KXMF25I3ZjJ+hy8CQgf+7jgVOe
tDp8ZyG5xG4PJUy9gA+z3i2VfD2NiD/COIXZ9zO6o0krjV22oj6wJGG8bmN/iMLOPu9ACat/v098
9X1a8KJULhBe6cMxe4tJaBQuiQW2HsMYamQHJ0OsJrp6FcTbFS6G3jUuOlVwEsoRt/Z4ufL8uBx4
40chccQBKAjcc+QQFRgLTZZOzi+4q4nX9kab8YuOxb9APGZsergYTNoVExFnCS7rifkcRjddAvUP
PLqRWx/cnuWOr7/5pSi8uYc+2Hh8UjrW9KxgBp+sDJ9I5ctCAziF3TH6HZueQxuNenvRtG6Q0NmZ
fUcMlJU0NXfsK2QAnBAjJqx5KEPv/007cIRsaksUWZI2s4NaJgsRm5gxX/xMEoyoUJOkoQDB+Hmw
9MTLLWPZDoey13eKPLkIoFr0Q4DAdZKH+B2kIduaw4JWAOc10hg3Nd80ZxSH9m61jDOKYFW9Q5EU
cFp/oFYOdVrsNcrW8Ci+YscaoWMVOh325z/0dC+OFwrB/BoMMkMQ7+Mu1skO9XWbztAmIbWbbYMq
pECcCNduHTk4efWSS/G875usJvPV+TSZh/aP8LC3iO62NoOaMbfzA4TJZsVsm2TAZsuZJNsz3JmM
TlMyzL6OyIj9UUcTOCphzrbVL8OmUU1ZH6eLw3/dlZJ0iT1iP1c/IM10eGhCKmcVOUmyx/s4fXko
fWGzrazk4Lu3gWpi+iQK1vcYCMw7FHzmrgjzklK17SEgEwqa9w0t28yTy7kBOz6c+2ezKLQayk9N
2oZcWi320eaq94neqr4DIexRXymR7SkobWQe85OCqrxbTX37ge8bhsklae8CKL2J95PZNcdwjRGb
jsl32Q09M9YKa+x8Y9sfJJir7JIAgSkCYbSQfaQAeX7ucjmO8IvP9qObu0QioNwOsDshCMzEvO5s
nn9CMVY+aQfc/qV3sJixQiJJdJqpB8nHAsU8TDWoYoCwkPXC1FcGx3ymhGlr1OEkxyu++skBUoGK
dZuTbNo1tnieTYR1KAkj7LGAec7qMTfxkG2mlFmCwFqysSgfF6jZz2NFUDO+KZ3HZF2iKAg0bp/K
rW2wYBd8LGsWLKxNMxjztv68Qzdvj49sgDNfjnU52AgpidtPJfv6tH5AuLHej8obsS7TzVNj/KOi
+duT95+zaVYLQMSS2+U1qeCCDK+BPBAiyB8LmH8ifBl0cFTvaEwthtzb6Xrhy4ERqzEGS9zKoQeG
NxDD7Q5GZBa5Fz8sydwqw8r3r+FdDsNh0Q7GYbJJZpClJ2iQjCIdd0hIYS0zxxpUvXX+WpVQvhcA
dE3qzkE4iqrx6qgcu0s7C0J5FDQAg0J47V8uKI29g+6fWT/n2zfalIranpdPbJ51uG7lc+uiu/7C
Q2WMBNJVkLxd/YWxtkBrd7TBx03Dohmfn5cB3jFDqMq8x2VcopNrARnDjyaIxts5K9aWiKuqrVpB
shzdye07D5v94YhNGHj2opdlkEeni824gz2VrGvkq0J98GXwI26d+z8aB9r1hcZm9fqlZ59ZV89k
+YiLifeNcCt63xfvxT9VbEicicf8vJmgwjNYwxvOUpc9NSygNypaH7irkGccefoKlodBrhXdW8tZ
2I+soxZ5KpSyjh12H68FFVLZOBcejvsdmHlshsdJgLhZMSiL8nHwgOj7UdfKshAlvEKRoQfwwJOK
CRvUk8tlE0bNEBtgRwDtcNPhFDKYJ/1DoZCNiQhcOfDByuYvfzyD0Ow0XH8e1S5yieZxB0l1QXFo
VvzDX37rva1c2SPwFIvNl65P17waYIbhnrciuPRlnIL/boVMXwXujbhxvLQXrr3I1lmYlbhXseUQ
zRMzQZgIHfd/yDm24rBsLg1AM0Q5CECEH149mFnl3kn0t1p0Em4iavmaYqIxL+N5Mo3kuIColtkZ
uYZ5gih7C2Xr0fmTqRI+FI49i8TVPW2kD2LeI1N4NQRv2pB2Q2xRfjrz55uCoQyqurZk/cobkjCm
iE9D+7rJ0pfX+29q2fN+/st7WP3lLvYxU2mF4tmLPILJalDs0FwjdDi9LNhoxyFDOMCHJ6cC5OY0
1xPbWrYZ3lX1+WSl6kPJ4mKGgAY6OvmDCB8Y8/NNvyK3VMSYPwzuAjXcIU1zzF02SHN9U5knHYSY
4T0pboUlZQCTXX3SJgnBTCh63pOZD7mqZjI5KN9og+1yCWpTrSdWQV3IjA7zfrqrOtFXSAPubmIU
wEw4uzZa2pn9T8/SxkwyUSCgLZTr7NZxy7G1GXs5+Gas9qAmILFfDmSFgBzWRQjOAgqu7P95IFFu
9It314yatR904KEJ3zURfAKNvhcnlAEA1FB/SQUdwSW+V0T++w37zHlc/ntOYF12memsI+HZQxH+
XVdIrT/e9vLONHpVnuJWSOMnUadxjt5mItBhwT0ZDM2ZdqXBvXiCNCktNDui/54ue1WbwGSqGu3L
tNc+aZt2GTJk3gtMXxNZQPoXTYUvlHn5C3pdeefNaHoTngIEXNxcC5xLLqarMOnPh31AXWfV2sUW
dIPxnzt8mO2dOtfHHuCOctVCFFSOUcQcztvt7z5n0KRdROhCVTTpahFUrcMDgq5abEpOaCiDOZi4
OMHypx5pnqrkn7W3Ky4ie4dJbAyWP/804Sz2Ahc+Awr8/H6ggJUPlIC70oOgCUnTdonby6DEE6MN
83PKYUtMHYuYsz0PrhyPcbakdEZYj0OfCCnYDlEuNSlJHi5Ru4BP6C9nF9u0pxzAix8p/EypuDto
HZpkacYOaBElpBoOZ/X/kipjjPZicNxTaCOugMHnka0b3Cd//VJ6XcDnfFz9GXgVKKr90oTqkcRm
55oel6/rYCgaau2F6lvQu7aET6fru5E1GRhM2CGCAMzMQyhBIENDWlYTmLXLJbKyKoO8JnTly8hU
1srgbs3voFFhkHKqsbUpmeYYpfvIOl6K9FjqZxYzMIupp85KXunQfZjTuoNj9CKTtYDqMACgsn7C
UJ7Ik6xbf6B8vUxDoV27rWqJbFCrV+VFhKMXWaHixENfAB8JTXJxeCEcBcrPfx/VqxEnI1HJhW5k
9JhYI0sKQOoDC4N/ecPPXgqnkIppulRen4MZVaKwoxGv2VX9BBRA4/7mFDTfGmOOI11EP+buNmvB
yzpxz8UsBpfNsg/VRfa8GxmndlH88jKCl6Q5DifhKd+de2hH1n8wpSyl/AK4zJgd8I/6H9290CWa
eX6nDhPypjEuPzhGrWpOGlZCSF5VhS0e1QK4Vu5AaFYlYUBvQCfP1VMx3Hzpo4q4ckl4OzN+IzAZ
KYuL6CYdljFRnX3PNKXBe8SYYPb8zaDK3fbEtohgWhO8/LyC+9LEIjffjY26MT7+Dck2SJOD8qPi
l/nAQG0gyDoVvevHUDYAYQbtyTCj8Z9DEH9ItcoVa6dh17bc+ytrMMbb/oMrKxbqRzDYa0KTKpXK
gkfOdi7xeOUdsz9+o+J1pmHffCMmVB3Q0QEs5w+8Nu1mdiYbLrQl/RdPfLEetNJDOFeOEwo1eCVe
Ei04XIUbsvDV0PyW1sJSD+vXOSWZ1CXdoCb4RHfkTtYscNyvtOuokYUezR5J4/6zgX7LfR3Z3jtU
QqYlHmydn00cEWmcGQRq+2uWJB56CwbXAI0miWfUoXCSgSiCOSPMs3iiAgYLZO05w9iOux/QQ6BF
nBZVvCZXOzmLfNBOJSyu8rlZYhlt8yJXSqSIKRdYILexcgZvBFFvehNVA72UX/bWneVWlDO22oR6
yg90BcqQPNBjqV7R9B1+2R/JeCCyVZFSdJ6HDaWVoWg2GBKaj1dAWiwnjWRKiobdN2GxV+HAMv+v
xYO8kwAJ906TmhEr7LTjEyHf3DMcQao+lq1Q0ZzF0HQGSEoIdG4uaUwAD6y/jheO/UqLTSwKxRUd
4yG0vumVKwIz5rJxo4DHUrqapPGluzJTufagKtH1loT3iEZSff2pqE/4ZFQCgs+CNEwQYRDhKFob
7fv7bVBtGb1HgsoyJIy8kPTIT3hxxak0nUboIt5ro7/X9SqW7zGU3w1zWZWnAIDXtXT3WY6x1ND9
KPugWgiazYGJZf7Z+ssBDCGaIiaVoxqZy9PBDAxiDdb0oVHu/NfKtLhADJCG/SGyn9vo5scU3eaJ
yh6xziApM9beoeyenySbTewEIsf15JznCgfU3KS/+AHk9GPRZOv7hpV0A4DRdUenXn8PIT5AeveH
gQ7EReScgbCFPZEEvPky1Lv2esg6XgSo3er0oaRVHv86XTMAUuf7kYGk85AL5efI+JmzzJpx62CC
LiaM0itn8eJT1SdxUuv8WSfb3jlBqQ9DWqaLq+jOq75pleuJZ9CedDHj2EKVnVY1+cLsASGm8Eh8
Em1jMTYhwVm+F97T4OomYoYLqZBNC5QkvQxvQVUBgS4vi0G8LSQZKhkIQ4ElWlPLL0DWjRNefGNx
JngtTIve17NZWY7Nre0y2/cR11W/3ehKooASbgEIzsuU3ndqykPo3D3WXVbVJnNgzD3dL3+3n13H
usLLLTk3epYJTayE5/dpMxqG+ohaSpyDzGyqFNnXfx31SsKNfNF1cfMpQhIwqjDEz3Pz8D1KKZJw
JKBbytNBeF5Hh0Le9SIfYRVbeuilodnw4jx+X+m1hp6F4dOE3NMIf7uwztSEXwnkW/tflYBsPBJm
FdfVTsEzSd9wNMjrzJSrGrtvVTk+lcBIcCmJ7o/gXTvpYvy/szsHMT2JBZdVOexIGW5I1yNJy72S
2+l+ibG6hH2P1hRl6OtzdjP+jR53ugrYKBBSoLe7D4vmz7W7OYDQ+Ax62OpIP7ygehJm1R57KAoJ
9NRQOkN0dPjxIK7xiJzlP2L0xj4JsDSiNp0TtVFIm2NPvnRy226eSdh+D8/6AnVhwgDuFVNNTjvu
rrtvx1Nlc2wBmfzm36Axc9S9Sy4Yvs3BAJZwNxPJQ1huMpCX8KSRuRLSpWXG9sXCsuyG7+uwSLnp
9LGEcgoeXnDZ4ZmulHVVflQPFQsegbpPlU4rimn3GtyAvj8RDaigmZ63Bs4oXrZzRuyFi1TZYpGb
UxE0LbS3FQ3hK876uvAYBNIQZf5WXcwus5GdJUYxZjLiXSVOqfsKi5nWKgqGdgGIX1JihY1EREsl
iwjsCIQPXos3MdbVWhbOktwPW3cc68ooystpbJZJQA6MncpczcfCy2CsiI7jNN10XJWZ5kZQGUvR
l/xqcK/rACSefycpaQBsaC0IrvAQ8IHeNdU/bW0KkkxT2CNZ3UckXfI/42NdFJMdqQlsTYeRTj0F
vwIjoz0BO6YXLGfeKlxTtdLMOOFgO/7zIiAtBJFoHnFBUuh2+ml6zXPacClTvksvuaElweH2jxNH
7vdjCayOcXOJVkG9t1gLTCSXxew35O9blysThYLbSVyVp33A1CF6km6P3IGgcJF1SW56SYNelNe3
+rX1Xh2UZ/UKt1n9rxw7+MjoZyAr8v0CIfd+s9oFyQU8JnYVXrrxTfiptIFpVJoCuAgoujp0FaP2
sKmiNUX80SQ/8pioODKpyps6VfDehr70qyzpe3HO98aYT8p2O58FZ9FuFy2oOyG9h6nEPb4r2hap
13zlOL2m5naNhOcK/yLkhuIRkIT4VVnZdrMrhPag+MKPTdjVhRGxy0M97HQbVkZFHDCPVYcBkEL9
bvwm+/w91AXMKPEYQBRPg/oryDVssZ1RzaQwN0RBjsj0z4TFyxlQeC5ENqrMwPc9xBBql7ncLw37
ZhnuHKjeMjglc7M/3o5NtZMwUmOuAK3rlaeBQ3I11ca1WRS3YPm3lwfyB3gx+oBynh0Olf0v3Ehb
9ifd9rrtr+8TrdYGnYjYjrdJXCLf6rXlfVSVF5ecOdraClj2A4RKroqRyLu5pZq/VQk/aryYLHWN
YJ/R2pntByzPvwJEgZVaTbwWB8F4S70A/PTF7neTVLVWZvFGClujXsQhTWnTQOPHwD1TOpiHCVQn
34Tr+TsZY5KSZU+xD4ucwHCmlrbXe+s4MrAmVkERYclKYzqE1we4KlG37GTgcRI6EtdUltPRN+6A
LEIlaA29uvXf+fBHu+bSGYcV2kgsz3Yb8xUcVO+ZEIRTfTO4WqQHWgvGwbxh2ECljmiW7OuTlUNY
HkswRXuN0jdeN1/SsZ2sfDEOEM8ywPvXOvbyZjEvjudrPeFOAa8fjmqLcMZAsnzfCbvGS7YcFyfb
0rRURiAEChXh7LqvULySNBUsNAi57jkYEn4WM3NCtDszn/jKENkdwL1ZjdiNqiqMis72pPMcBKZm
Q4Uu5avUdm5MemY8hOPDKXyPlSChz9i0LcYckgTq2pqRDXN6XkluFeIxBSfZW85Uut2DSsWbs3Nk
N0IL29qYOi+0cADUMp52jgY0xi6Unbc+9Nwz0D+4L4adt8V7iQWlGJjdb8JOCY/wPS8zX9csWUA8
StjhngrwU+DirED9t55ksMzhkK6FLp+ZMOaqYAGw1kcBNdXiuMKtiAiGIplRNe+D7+m8/XzmayUm
Yih8cdfeVa9O6+veWH2CmbHgUUa/157A7Qt+fmYai7QCryKYtb9+hEeZyduRdpBT0Q0iYB+0M5KN
Bd/PCJJmv8J8shriQcrxLCwR6CN33wqoPPRmI1wuvtg+ZpU9opv5cuDuLrnVg4VqGhRMXr8F/Ih7
n6ETNOu47CZWyGjknndv1L2MdzMIH6/PClLBfO83h9bTfLcb7AdVhuQkENU7dVlG/ZK4xAOrtBGk
Ch6q7uVltaXObBcObi63sNcbJBjnMyOw/8eW1+JMp4hunt8gTZVuxaw0Bxr2ShDMflhV6gYHa4zA
X2Ak0x7pDG/sWsY6ymlukOWvJp+rV1cw40qND5aonvu1MD8yVUtDqQ8RMEmeWkko3dl+SD4pzWO9
+2eLP91k6O4Akv2GEvgamozYcCtFtTkR03bPqvnhhMA/MqwGfjwxLYIydObZAUWdF72C3w25irIl
uQmFD6alVRQuvrhIfEujKBMcB3VncJGLcxPdbi/ZPMl4aC9ClT0BydQqfAHOWF+dDZvS28uY/+xl
ICKlKdU7rIhEirMkspBD+yM4C3si4GEXTS1BmYuDMKdP38AUtsu3eRLwHvxc3X01hIQ18Twmc6sA
wo1hr59JJ9gxcFBWRR9YZ6Koqpts1C4INDCWjzN4iUNTIq02Yf1Ee3Yl4jEoSNIF0RbWJNqfrXlW
dg3N62LJ8hjCAK0UN7lJlPy0NflltHUyp3F3v9PmLo/Yri0tvEnJjnzd5qZDZ0B9J1C+qdgW/GR8
xY2YsbAbp2jxMLPT+E3lXY3FqwmzGV51V7pwiSqvoTYs9QVpZIe6QWGT1uFF38rdH9HqJoVSe/nk
N3jCZ5gGEcMPbKMTBCML39aa+APftuvkmiBfymIM+/oZaKln3XlSxX8s3rzwGXyEwITj0TpdjEO1
QEKyBoFn6oD9DNBhskTrv1iPIxBVquHSOpvlHGEKnxZBHHOl3UnZhFe9y11OGjaVTntDTiWVpP68
c3LDCWYPfpYKm0MMtxdtcbL8IxUkZ9pzqCumoWOixbZpF92WPa5VoAOebwH+G3IyOLzgj8wc6pal
C9Kg385sWmLrp6nF5frI5sLlQtrg1RKxCX64jLLlLpEfdTswz+B7b9UNYwyYV9pgQQCVfdVEIoG/
zOCDrsevS0Eta9bcdlouINZHOlkpwXCBQETt4fmdlC9ozTfBsFoGL1bW4Nihs97zsxvU231Juquu
XZ+n+Q2C9cFaJ0gXYIWiX698Z2+RWwJ3JCOtuCHj9C6T0VkL9zCLfVGJKtwSjNT6SXNRUrDWaQYV
PJBHkTXqxgm43zu5wyH+r3SKIyN1819vBiOVUVQXXQYY/FFPa7Kzfelvmhs0GE6wIj3QVVKC4ibR
2o4Gm4qdMeQzAMmHG6QFtzNQyJuCxhvNkIQFA1HGTOe+mDxuAmAyVPViMN5Qpr+KOynWX0BaTb8Q
5gPMJH01HLUoWSTRpfg8RlZcQ4joCzpu8UuscLVZAprWGMmFiXpkaDVGCjWmkL8RIdcFStGY6m/D
0XjvEmOU8+gvgPcHEbmJ2zQdrYfGsypZFrBbnbOPsDM744Rwo7cG69tOav6UJ0PhGoXDEmRsw2ip
2VMKiIxXHlfDKtVPA4dnYNmmSg0Ry8GKPh9fhIWhnxtTyj6cuCJAbqsHu5xtnLB00ffWztXyFCKs
i/J5i7rQXqd5TIIO5OQOMtO/uhdHxnTG1TlencreeG/+SZr74Ge6CMmJbvFgWZAGsqE8kwR4ohEP
amrRHRyhvPAK6aw3jo4JK9J4D4R2aMQq+9QWBk9B3WHlC5zIX33v8+h1TBY2hY211iY17b+L5Akj
Q/ddHlGTG6N98nQJtx39ZVRDKSFQdptKwJ0OuPUq4XtNpP1Rw2CC6jGZO/OA0nqGuiV+hitlx88G
SyTjN3+N06l8FQt0dSn55Vv4PxHXA+oTUTvszZoxslDSJaG2kbepyaIn41W4Oq5rCkcPPeRWhFv5
9MfsW0Ljy6JPkV7LlqkzKiFhbgBKCZQKkT60NH3nlDqC9l+XK9yy2ovgcCbvODQ0B0F2SYdeqy5L
0l8Mj7ssVIv+RHNRvnc8jMD7ddl++XpN8sZq3CFq+Q6Tol2tfl1freIWeSeYzFYoeU+AZrQKOg0Z
6qqZOp8icAtKYbu/EXjrarS0jSkLR5MdRDNVLfE12YaJbPVsiB9voleWUf/jNwf1ze1EN4v5KVb6
n6Hg7leYS/0WB4K4/Of2EH7EobPCqAUf89Ig0eNbJN2zJvoyRfcV318BAXlkd/Kdlbrn6SjKzMaS
mxYhC6IDZfKvUxJKr+JCBAqkk3lAhw8gjqTdxPTQVJG9zo0vOu3Zt+ZEJ81IcvYgkADrkb7gu9jR
jVbPBuvmRTEnRPj6kBdEXQimj01Uce1XzJRob2cUkQFrH8oFUc1WUkTbfKiqvFFli/4VBox4a9KD
EJPL2KsKgUXCRLPMagWqeB/pgP1Nay89LAQIKCaq+/clbmK8hhh+wB5lh4M7J31pNTImQA3eQBpg
VjXvDFz6bNU+VblVCGiOcY4wGA88ga6qAzyzK6718aUy+KrBjCkWC8GRvV7DXu2koKHvTuTXW1gP
FNx1JlhzU9BV+CLqoQyifMH4Yt7GSIqwNcRFntHPRjOoKQRUGbygWmESuwoClB1C4x3D8qRhrQke
+xUpvzyMVgrLSM+OMY0QArXZmsYq9ynGiNrWnxN+/XQMysLW/lPuqSuKeVNUA/cy5ryvmfjF3OUV
zjt7+NvOMohhQSvLQdBLEm95SSc4qOqi4HZq++cW58j1zkjDYLUQ9V7KZyRAq1jDnCVp30gwLUqp
cNtQAhSYoWm6Nu09DpR5L/3m3Gw/vheDtN8GK5Gmv/bMCTSH8yO4JxClHbiBdVqJbc+wuoqEFrwo
Ay73viXKskQ4tKFD15APEHj42hdvMn4OgA8kw12gFDlg75tWdOs6JOM9fVToKw9svHB2x+aJK6tI
SNAFwR9xXwPKVWPHTU/ZY1oNnPNbv7udTxwNPyaT9zzcR7+qKljDn5gtDHZKIms6rSCW2Ix5TKf3
1UO6QHendFNeRKAiukTmnvW0Gk/wPyu4MfRx6qeNEaJp+uL4NWiPe/Z5msvfGUGiH/OKGSB6bl4r
hqPYZFZmyDiqhilyY1TkTViZ6UQ9KSVpcx6wvOZoo6PNU+446GDXkLTUSLSNWP4LSth6oZsdNCJ4
yl8i4+1efv1y87UJLIEXNLEqXUOlG2RBawU1fT44vIidSe/cfZtY6hpsRRRdQow04m12TnTmEfK8
aiAB8d6To9jZGOadDYn1neU56sIpmaYkhkBhsHcbv4uyFTU5EmdWJHs0dDZVn1ZI1ZYYz/GqObxY
/8MFUhhAPZ7c6vqGUGGIl12KRHlK3wWAYalxknY8HIcfycdSnP3sdYtOq6MiNtpN3ToNLDFuVJN9
dy5NXazndUHleJJpKUqIiL5RH34ykTDKLkD9MQTHacomQGB7oF3V3iFQLZ7CX8YiAhJ8japk19sx
omXNgBkOv9v+KRARsQt0jaxMg3bJLHZ3OpI4zIS/RPOhkmlVOREdi/fPzWEI6YiluQiIGDU4lUnb
3QSPYA8vhu/LysWXF/uvwc6LN8JzixC9rrgZPvlK8MVq8BONAWy5sYsmgc/+AiTf/ToPkZMHXIRX
P/RmmaXD2zBrOlpreCWt+9Fs5wR2dqT/Q+8s6R7PLp8DVkyuo2Ufgam+tQsA/S7F/5mNzAhop6Ku
Im63/MPKJ/oUv0j1oNOxXQwYPcEfp1mkX9l5+w+9RDiDteEux8jy4pRpPpWlAEsW5y644bLHdqAn
rU2ZhMiDQqLyiWmiQ8BLNkFxxbQPFDlvlSlwNXOqvAil8vhodSFehfsfmTRu4P9WWTJSx97upVTr
lXVxmcd/gcD42S6D3LJF1dzWooJhIjCjsqJG8fPIGhkZ/DNE6gsZigIM4VmzbI+WmfXoM9hIkzD+
PJd5O2A5aT5UKwtfth9Gfx6N2HvmWiomILsr3uoPpk3PETBtMd+tuYDOXr+ac7+IBq0rdkHAFo+b
Nyfe5KWU9uiDLpombuDKgunItmXxrZHXbBJxaCACDVmePnefzfyLvcdpdt1V9MCUiuSpz3YJDQXH
wqif0piJ78W8p4HfM3LFQv75ISHl8+5F5/AID1RVqU8X9r5DByWyJQgdIwpQzurxBSmqLSdmxYdt
RCUv/n8MWP3fWHZm86bk7WrF97HfTmo3nVxzDt6lTKAnhjpD2QTHLUzUlH6ApgyX8sQe8B2XPbE/
KAcmkyND8MMpbl0tPlBz8HLkdIxuCHDevNUbr65S4ICMN8yZvo36eqjQiXydn/nZ5Z6sx7wa+c/h
mHS56xG11Pw+pDCfdGtLISVCl/tcyyK2CaUu//74W/b9XCDRVuS9Y/vfYow4luRrV82m9Wl+vtip
bcv337531nhYhZ7OCuMjnBFxtLlHGBs6FZ/9aOYOnxINm1j4Z46Rjx0CK9PFE2L17CdQ0xqN5246
kQynxqL2zhg6T/mAKbsjAG1pT/FbplT8bEBKoTE2IwG0LU+yjMHGrgQ4YUIeXHTE6528R1gkdYYP
pXBucXpfGnq2ACy40zMaS5t90mBhUAKW26DQc5bXuPWMKdJReVSsgiuNvbigTs6O+asULBXMvldH
oZvEfVLZV5p8MdkYJUL4sQM9ZsTseluf1rKzHVn1R2CAJrBEbf3NaiSyKGqurcG6bnVFW8v4qXuT
uTsekeMMeJY6G+AU6Elj+WFwvqeuNVDcKJBA14UKh4xo2/cBkQbkd3hn7VKjitNf28RoPY2KBZcn
DdjD6SkBMk3JRhtCGzmD4cGYjuhJnyW3C4S+7e8pRDyS/WP/0/Qew1rTJj0DUa1uro9Qhe3+FLHI
wdkspEkVVOwKn62vpr5bFX/EklWIdosadN9mjweBey6U+wr1FrUR+NbPvu7nrYkaPFhqCfUIG6th
HRHsf2f3UwxKeETwqmqMR2PCHb1rqVeVJB3NhX78UANjjO9DH3sCVbJyd7gQRm7Oo0ilAAKN757v
9YsRnJ1z0HZlem4SLBy76advjmgq1o/8qzQGy3JnJDsijjm83pVo61ob/7nWKG0pqYHyt9AHgCvQ
YFKZ7CiU0ySUcDbqePK68tukQ+Zfx1bb7nn8m7dJhzalvP1RV+yXBiQtYAo99w/UVNdJEs9F5Iry
Ub0PEhMyq2QU30q/WLBXn0GU9Wy00yQgDL9nkBZNmfgfY7y9fQ2j1c1DfaWSzehcn+7pEufEUF+1
G8wfzy5/hdKlXy6Wou0hXq8wr0K+yuBGj2C0kgQpEcHU+V3BPZpBg2Ykw6NDcRy0y0lHljhCts76
mNgOeT5/c92/z0VDIlWn75J7p0FsVz3bAahO4OAcfneI1wUvFFyi66vVa5mP3ZsEusUYwQykETeJ
UajBbiUphIc2pZKgEQ0cY1V0k7LQyCT8RVQPakBKTiRpbfKHQSfIfnWvA0CJdIFRRfeeCaoIBzHb
zvPwnjS3RLqu22BKbkqOTGF6RchtXBKNYXeEO0JT4gTFyi53cUP5FGyrs0hsgyDBzCCGPZKMcSTB
WS/qLTuwZdapok3PIK0Ga/Fmn0RKoAK282h55DsI96cK0oIOs82jlKd/atoUhx2H+tfs0KEHGMjq
hqVFJvfQ7VGacEpPKU6Vj5L5aFFSMRG95GmS5DrYTNjwPBSmh2lSzWt75xoWV0YY+/hdilpkqW5P
S0NdR+UyN0iNRymVj3vsqfAbLMA6LVqZrM7+roo2jSSNA0dEKXVmZ2jJTrIn52KhyqJaawQkpzg/
GwcD6a13z5th0MimT+S+Jhio44z/QxP5uRlvLNNJKH7dfDLUbTliofWR8t7JvHg2wluYc9SWJlz3
k+hFQ+IebM1pnB9E3mI8N2iVjzhu1rC7Qf5jsOxHS7jS4UStlZvQjHXkjykxgCQbT33I5IJxu23G
IFrKryPeyM4Zel9FPlnVEIJDjoMgvzAR5m8T55pXQ+rLttId6+gg3ktFPvFjKFy1bHFj4JzgUNFx
0/ZvgXG94i/WBMzg44dZ/Q970hjM0PiCeEIpaanhvy6yj53Z2NtqknvoInx7Dc9suwSfGF9r4R//
fBDKsrKsmwG+3U3sjWrIXWDIs9Uo9Gk8y/LtltqW+6IkE10beViCjaYq9U0a2lfgeKm427iLq7PA
Pnxu7a0KALbIqYO8LERh9u1RvZHIneVnePNStLqAarvJlJi9eNJMi3CE7ive1s9n+3n3ed5FqyfO
lzRGUhPs1q3eMYL/D3E784O0iCnGTrw9BrgvOBXnzMScFKCRtNlq1GF9A9FDXt+h5d6BLzJHX+YJ
/aNvSNG8NgYQUoQLpPBspSC+C2HUWp2Yperq39Cz0HI17ht3s+WTJLfdGXS592Nh1INwTm4S0ZQz
+/lJ4dqYqCytAqRJO/hOKnWxxYabquWeIzVmDX2jPNjaZOsa4PMhoSssSjt86DvRJfyXq4wAzgoN
hIkA9bdsdhzGPFKMy9QqAhDP6HXGmHLqXTgJhuEVGCamhmHhS3H2zOEgnL5cBlozY5y/Obx14cb2
7vBKJwCGu0GlMxzesNoLMuntp+Orze5xY2JOOrUAE3Cahf3jQHXfZTKfsiFsqVF2RT18dw6B9o3t
c1ikcSF8NwEs7aeous4HD6eWCzDkRMh1V9oEtbienNVUD69Fo9SZuus9Y73Ic9bXW4EfMWL5oEVx
aXq+DZzptX9fBqUAS4tosPLtfkPXvNSo4pSf+CMp3QcdqfIkgeHremoTchltdrQmsNrtH03ckBEk
M8zQmuMhmVv7OgHd1t9zhH4xafs9JuoL7SklNlA/zoOOqfTqeFBrhOxUqXn9G8/fCkDlLhXQ2xO3
iaWW0j9l7cuVFyrwjzMgwk+F6bQMcD7L31arwYFEUN7MXSP6xvrw0HGBIFTfY8VZ7685c4tFNjRf
j2frMWZbR2r4RM5PplmIfLoAVpcFa1cpi1QHPddqokk/Tpr8O3+vZlJZtoB6AA2GqIk2ixxA/bxq
ka7rDtduqvVvPVOeI//V4/oJWhfut8k9drPuoODC+xnOVTlqjWa76zPzOoGl59Erotq/By6JYHNP
A5BW7qcipJw7BjAvSO9N6Wyftb0ZL/Wo7qQZyQvQYpyykjpfqBMLluS27QoKN37ocWgLi0oQaykO
SSRJQ5Y8B5b+TrnBSN03VEgXJejOBmTQpaUESnJk7uRpiYUtATT9jvl86kRoMOgvNnoHRcsING+6
Q7pFEsWBNGkqwTg2GblAEw/5TmFEIM2+731/uW1r80Dq4+xal5ovRVTLv+8kRZDuOL3MMlff0Tnj
dNulfNeDULIW2LJy06LI/IDraRdRQ47k1pvXfo7fMrzVzEJNW+fcZURcARldbTyNc0ilpzSa5ZoS
Zr1tqPezITE6y9XPx6YqbY2wR4s23CykAQbxDFYEjasduu6Aj+WNoyXeCpczsogX2mBTsIkjpm5i
145ZZfF2PRfIJ1H6zOGEaGzvqqvkERpic7EdxP3vt852TF0DEdFLssxzT8QzxeQVXGySQt7NO9p5
Grt2GlAhOdhvprcy2wAVcxKYE/zHZ86SN1uVPH4CXC9c6F5QQjXhylAdBdTpf8q4ixHcq0RyXULy
p65p4hFnQeL11ZL4F3wfd8HtJ3/t9j3ChLqYkzpVUnKverVf/5ocD39aETAoVd9QZ9nNT0pDs+aA
70xRXJ+XcDt1xHNgZaYadqs/7N1bkxdg9jvwPnHlyXLFHdKJTgcp1X1E2PaX+2qYLszz+qx7751d
+rP2uDrZPkdeBlkrH+BzxLC8Ncm4KTs+YvotlT2gcKSJ6KDxx5d68oV6NIc+3CtsKiGS92MLuhnI
yMv/HKkmpzLEH+rBXbeuFmN65pobVs0IRodguF+6P+wQpWq1/W0O8h6lYw56kAa4ydFpf9gZlxRR
tDKk+w5GYh496tizIpoUu5TiUj/ABxId5Jx0E3UNxNzwS0QlkJr9v2konmQFEMsltNIniP8NNz2P
i50fBp6T6gVLkQodGEC8okR6OGFX/LC3zOPgXL0cos7xGp6Yfzf6PlA9PHRJyL0NroUAgzZ8acxn
+n2MuT1bKRlfN41hOdAuztNQhwrnKWW5cniCCPxDlo51juljoHUuAn0Wh46EB9E0zUjA5YtdaDuM
nJeaTqHKkADfRV+V5djGBaOWyQamu480k9vvM39wdWwyc9kj3G3xYfRGh4Zk6k5Gf6jbvXzlwD2E
Ow/fN1KBNGUauQ5mcMm2GEcuRGg8dCndGmSv04J2BrVm6jxngDM2Q/+Lpq6MMIbAWdugVE2DAd6f
TbQupUoDgmsRVV2UkPE8nMnkYqOxU1lxI1rBaLjVuSlqeCgDfB8QIFMExrtdLb16jXFJ2Ja5RWwM
f/FlRozRQpfMhBGglnu8wiTUKad3nU1TOAbJO4FA8TejR/LXHEKFr/FL11Ny+RhVwru81blSMy0V
R6JwM8Umf06corioUf7x7pGUV98hossdGmZdB5M5wEdy978ers3+fh68qQFuSa7tu0cPvWh0amlK
P66+vCNFENLhUpjQAJn42LCr/+zI3xnZ5NFxlOuC68DEbTDtzVgA8Of3ASjcwDtzPpMZZTjzd94Q
PovB1Ft2+ZtTZwBYlktYpb0ZSKWX3/b4W1Xw0xIRJhwbMQQ36+GfLsj5eCh5Z6XIknRpiQ3yDizS
aOlguiIkeBm4vf7qkTrNloltqZyM/7/jiRTY1k6V9jzloPe5mL4PXcpj7AHE1wdXlz5aU2IS33eJ
sOTElODsbjP7dP9nza7sQ41Sd0Y/DlidlqWFpK1pYZ4m3EJtiS5cFaU5I2hxw0j2R6KYTLM4hDSd
9UeIKqof+DvuXR5NtJDWWcoBGf2wdijXxWFmeiII4oEs4gG9qu346UkfZlmp/0d08u2F674dRjKc
+FEpMPDy7we0zsEn0xzQEzpmrf34JChUhok9gmAyQfNCbHvBSfSjKovIgw3qlyYipyq4X22jCBhG
c7gh2o9yOhAFdT/q1qzSNsZRNbXy1BMoQI1HJ+X2Bu8VJ7YdNseklD2AKr1kB+/24QQ81CiAKZor
51DGuciM+9rbKOWuuUMmgrBuWKkOufMx4gqeSUlq/2xcIgGxCQ9YX8adaucNo7GnYFzHF7oqnKFV
Ga7izkRtcDR/c3pTHs5mO0PuyIvUk+ul3gXfoUL/1o98M0NcniKPeCrvy1D7qSV6wLGR2ttWOHh1
nltAMF8k0loeyUepg+xkTaCZhY1FfB1UoTEORguwzNTu4VUCz5Enx6KA2u76GHrlTIy0BodPzG5T
GwFKD0BtN9GIUoGgUe/AJ1BtVmsxPxrpRHfAnG6+p0CEUtvSKKVLbQWLKfqJBT1HlapKUXaNYucl
YsRsAKdHdgNgoy6V5HO17TgNagjg7K0OVWxDUv7frctq06Osfr4xNgq3DyyWKpbxfDBsyT4z9lfv
Px5IIHc2THyJ161vl6CUhKvEdMkxw60mHN/yH7tQCKQqbtgwWbaPGXztvHa77gtCSiHPulxUXaBI
hkUTeB7EE4TGxVELZqLWJZUqU9Y1iPIdjkRUH274C09X7slSbGrhs7m25H7Fy4fi/ig5UVtsJBIe
LQmLrgDq1E9sGkIxgo32Y4ZyjhyEKcyqMaBDpvX47huu990Fd/JBOE0T/MzWIGWk7maV4TfFS4Mp
Nf+JEYOCrSiGOSYzBnkbspIzOS8S+KVUkNayHjKWJhHSRlmOpYgxHsiPwRNGmKTvobS+1qtNMZ24
USWb6jBhfy68RjfprYNP8fkO6OcnS7g2dDfcv5fGfW00qz+5cJaAT+zAiiojOduhccwhVZ5BPSBE
6ZmmrmUkAuScUJWzEbxlsrpDpvRsNcTghkHAmH5XLry9v5SpoKC2/WzzbB6h47927Pxzgw6nC/xN
6q0fYswhAHL9Z10gD0Wb4w2r4iHXvzR6Cx5BPbtfSdh7XpdvUAYL4yXKYY8NAPZcu0kDlYD/V6aP
wVdu9F3S3QWwkEjZkCmckDo44taiykAyBK+VnDSpAnCgq1mxyRZ95opUFK9FRe2uaRgtqPV0MklM
1ysH4HPO21KAEkDeb0mtiIJaVUFIzow4y78f/h65fXWuLazxsYaZVkbucrRE8A2g+Jt1DAWhFllF
Fank0il81tNDHqPSYJvEeIixMWAhRh8vDkw8W/IKd/WJZv9d42N5kCw3fu4QU8SO9Gu3LvAUWBZS
Eey6QYBthJUvYBlyEoGLcvtBihY0aVk4eAQFVZoeJmWiRwe0brsg4YhUYrnVR0LGcOBnFO4cWECl
xesjxD25lLZCY6m7VoS30egYdrNNhmwzJnE1f8w3IKV9K0gGzb1mOXKqIJK3OPhyE+yUxRgptnZr
uL7rU1fbll+joG/xQf5ZwlipjsCTgR+EoF71I+bXShNJ6DcJUf/RxkDA/MdMllEErTF135Sfq3TA
RA6oFNLa6jsM8zIZTg/izbK0CmRTkauifj3csunpdQxZ/mKVelCnBoo1UEXyl2uscrcMQQvTJbxv
7wFZ8SWwan50tAFyUnCIJ6FEOT3CPLEe1PCgRBaCuwWGNu0o4wyNO5r3oACDdzC6GUH8tqOOXsp0
dP9qLE2recWXZ97U1aTJ1zgAgCFjxE3m/R0lrphnxKt6IKffug2qrIYNucRdsgTRlYvXzFJxjxJv
K5sG6sk27TpukZTA5nk5/3Kr0pRdshn5pVreVFPaOESZz/rphWgXfKhBaWIlFXXTV4weFSHqu3rD
AkfLD/quAJSfKjfrYlqMq57XEENDK0x/8/D3ir3i/0YpkGJPCPsPi6qCQL+VTFK0zI/ZF59L6gpT
GcyvTj/iwAoG1g2MexcL0u+rxcez8qXPglQB+kkprI4ofyun6+amLfoyxc+/StDf+aSwpuAGJsuQ
g9diBMmpaQP/5YbEv6i6Tw6YLQDsuuxisl34kYkB+wJmZ4bxl5TKQVLP6N5CQpFIUDyt2xE6Ijta
VwdUirqg4mtzAfC8G+J0+WMdXpf4YjYI/sUj1x5klSETQubG/HcgOqYrrG92VVCtZ/4u1AuhvGqc
4Xc4qeNLSs9juMa3CVET/s4T/5v3e95LVvSrVwU3yT9LR6Vby/3OD3l67Fan4+fcskK9+YgDRsh9
Up+9u3uKm/DPJ41HUcv2ZC/MmCdlak/6CUl13lJaNMQgyrOJa3VuvmHkd7EGREKsrS87TC26Nqln
XD3ZI6Mx8FFBRuaaeaitOeKVPwI7flx43YHaAKcmWrhUdmgDUJE8thGFXDzFE+puUMKn8338UV3J
mfMtPxVBxu8QmtcWeFropOxWXbdcl9fYLg6xf37lgigUeFABIkHUSUOaGtwrE02lZy2xnrEJckbL
bUyPNC6LjbFMOJ9fuk60Xw74TVPFv8AGIN5h/6oLSmvtvmQ8OxhJqMnCfCyBp97LQsH4TcpgmReI
mo24TwKHaWnY0cnvmW5PF05GCDE1MV//A4UtHuW3/gB5ucw99qWfp0GzhPAGDJQZoUQVWmRU5hBG
VJ6qAfQmw2EjXXv5ookjkh58sA4oDwNustQXFXiWkqn6l1Qa+FkxjWSU1tMqHUo1owilAAsQryQA
d0FRDjJNQ3ZigZJNvmsQIERnXG1j3RYx0ZO6Et11BBwiiMWLXWD0V/pY522p7kubD0qMrRCGl8LQ
B8+LCZKQm0aS3QPJ6MD7hU3SZDS2Hc/y0ascZmHsRQ7rRd3gTn/48SDX9QdzA28JNJHXGt55Vm7q
UKFgLcuU5cxpi1xDZIAKxclv9R4r6dzb9rVJtLrc0iH2b/YcPWCjxzcA3u/ZW6g6Q50Y8lTCaKzG
gWsqcYbn3+q04vzqZT6SpPzJI0JxTK6QPARCDhyJJtfRb56aEtGUT/WApHrQozLhK4bujbd3j0A0
lZD+tVl7Q9AJN/Y2NF+oUfRi96eMIN4RS60ZEihjYsUCcFgw3YCmB/PA8MrxpDNbMlekHNgROMtg
pMAo0uy6Lu6N+TKgHCE8J3aej6mJaerCYunoIsxyjY+xnc0VL1T+Npn57XuDBoM+GyLBSgTnxNnu
eq6Od7hT0SedIkDqfsZlH2zRZHPTfA+agjMeKhbEOVIUJ29ocTg47ce/BI7/RLuyF7/1YPbGCBdt
qODnGujzc9wel8fTXJ9qt6Zx/Zu/+6N65XE9pEbYAcBwywkgiUIHBxNopwfHmUXQeZ+se7tqN+0i
9iznv9qLAopXukcKsFRDqHe9yNQOXjGJnIzLUduQMckkzDMAcDmjl12/QMcZF73S5LaEbrhMSZ9B
QQcN7XhGwtQESxKnqKKulqy50FC3D9KognkKAdVZlry3lqJXxz3rW/0//6d8FOBep/Q2GcHhGoPb
fVTIqJP1ZrQ9D93EqeQYXQORtxHAZGdT97da7NOosac+QPaMM/HcIJRuZNIu7EolnyHHIjOWIe88
xNp1krYXVc6or58kNLwFZQM9kDccoTKvXmSmicFMA19DI3jyu01jvwFdr8BZT2zwhPbMqslBXBtu
aty55RDUswlGCgsRmWWPc9eBqVLcoUYJUlW/uBZOZ55T3F8eqMBniqP7NBwkuitlzl3296JRuqYx
/ZOBfhH5pu708BHD1PB8Hf/wC5qRKYnnQncQxWWWd8AR6cpunWZNqbqHgNZIrnEK0MuBGXhR9lp7
7Ab2oV7IZkLovKFEcaac/J8lt/udhsiq2JwAyX+g68ZkVjl75xKfGn399zPvJg1crWbHuqrApY0Q
wBGXWjfV+35CWS396IlzMbR2+jtIllv6bhKthRDLy++/FGUdahjEmSBnRRv3C8yrkNzm9FoNZgNU
HNe09XoLZc97KC55ZIsfb8rOqRFTLHaAfARNXDVNlgXHK8nPuz5DJDMLc2VUcpDjIFLx+hThJmax
A9EiDaK4lS7RSWa+J5ZRMBOiIY+r0G5U6FsnNaMptOm4MBvI+9vnRDd3Mvz8o8W5JhUYag5WjqVW
bPubjKUw/2ftpozClJGvJyRU5l7HcwB8ZmQsy/bobqozTqbKLhMbswJAS+6GV+jhtFVqQaUWOE31
EbbjTcHQlU/ZOP5QtmNZ4hVT22B0mL3rkKsyDCum2fvlMYLg0dF4NwankcNckH34571oJ5R1Zjqe
KdvqXHtgODN/GQQLseCEXibTRI21dbGO9AawG+CnYq6uxj4qcO+K9m/t1g+/AQ1JkmPM7u4uhljF
XzTzFcWigogMjPU4XFiPX9txUvyK7L5maAFJjhv8gDMkyLAuLdhWdMXQXEjbfOCtcgyqc1HmZABV
WcHFglcGAQXgh1UZs6BEvWJRDT4yf2nVsbUQb2OnZlAlZ9/zUooU+x3s881ggmMAnHs1Ze3K403J
x72VGvYgwF6pb4vLl9QzOMgKs7b4rnP3WN4IgyAb1AYK+DPdUFSuSifHmLD81MQAUrufv9jw97TZ
4V2y68qu3xcvU6VIvjwuXsZoOyUsyaKGSKj9yZuVXmAbo+k6E6KnS3wgm4G1Bd/SM9dS4WGKd88O
4+IwjVBzsgj/8SdR99hCVgEDKOCQ2gyUpijnJKMnBwL5bWgBMLcXbCmh2170/iqRaQG/m0adNcVo
5P76eaVSU6elgIQORmWqTurtDbkywLRVJkquH7nxfllFS/3wDb7LeGMgICvUD8tJckd6v45xeW9k
dgZLeiIVVVekQn0NTumlLzYQkgPAsm6meaNGAmAFvTZ0wuJso8n+RXbBfd0J+92EEjGhgAxutOTM
1YBYvfoOlR2/4zt3YdtoBdgyiP8N4uJOYkAhA6PNuea1lVXd52MlYRj1JcWaNAB1mTt9hXIj23+m
hhBqe/PHzzgzNqsI9D3j6sCevrlLgKAohb63T5NOOex6Ec8MemyxKi7Mb/ACnVDory3sYof6OEZe
xQwjl1xzYJF2fOB1BBoQGxmI0DQaX9bBWg4wfyWdKPXiEBzKBjZpaAI7gUfpv3JCVnpEE3+05Dxq
sLe2dPJFdXq/elw83U6oDC2qltLiwC4JNmUdSRVfkfjDtBYy4BADDaDnCHg8Vp2eG9hyoq01rRqS
FM9T8oB6e8vhN0Jn3iYSdZ5+RDiU4zv+ywdsch3qaCSJb/4X7/6QaEww0dUH89vYuO5raocKOotb
Xw3QACqsh4iEKZ8SE6WSeLgmozXXA3lIjPmZkcb+V+iuPJmxN8tz4si5G7/vbqQ1cI5Iuj3FG50O
jxzq34152gjC1BX+Ko8Rh7Y5mQyoOJk+VLRg0ghYWQbZnYrkE2VeDv5XGZZ5HG+fmKrHZge+0AU+
E2+pCO2D9ANgHHih3+9BtXwCmx+8At6NWrOs+Rc2+CAN4BYIk9+BxpDvUcDoSqhyeW9Gpu1PIATv
3TqI7fA3LQITYbuh7Sf5lqyzPFgWpSC6h80U+bgapwcP6CFhsFm+Ep1ERIchMlYv2icdkQmaOK0T
OzfGf9XpwLpv+LuOymmEbpFY6hsLiIt/2NKk+P2YAJO4ouHhLEWxBTJs1Knk0FylC9j8UDe6i0FH
wdFTf1f7gyIdG3ZydriS/QxJDiyFw2KZQLcn1C2KWuJaXhppvjanyTEhwOAt5n7kaNyWkj7Y0Zmg
Rnecefe8FWfAhsjzjcvaCu37qaHvLoG7D18kkDIN2shuIfCoI3bekaZ6/zi090Fy2CpAgib0IXiC
bRbO0Qb/2c336NAkRVzP0rTQbkCe6FNFTorSnPpGT8g4tIxOHZ+gKMUIx95zloM8eDWA0Iew2r5B
9XUpZs2z+b1+fcFENh5EE5++YfuZgXNyxsaYSrl8emezGuiZ8I3+fMU5yH3cUR8ufCDoRswxzwOW
hayHIb3g/zPGdHu7u3dionpZvuQjhQnvxvF4JfLt2bEOnTr3+TpNCkol/Aqxkj003fM+Ho8LMSls
fyNDoUyYP+VA9qWGOfUBZyi18vEFiaTarnFnvje6v2fnGrNdlR81DXckDAwMaecWvoGHSM2Nomd9
SefvCyi+2BJJMOqvwQMbOy8DmVuaAUpLsj5Tqlt61eembx47ZxI+oNiZQtZ6zJC3mk2b+X/Z5yWG
53mHyke4fO9Rahv/g5+orvbfyWJJEocw00ZFtHA44SJn1PzO8orDBacu+/uLM2fWK4QKZEjcqxCN
A9Jq9KJEwqTjkMinYiwtXGJLTDp88Nm/IeCvlebf8DV9A0vT+TsgtufoeMknJoVXBWa8+5YtGrmO
udDZn0vfL9ipOzFaVnBs43WIVjs7GnTOqzwVfw0fg+UMuRNWdlffl5eJairUmYWu2kqF7AGkrwid
AqWulzIL/4mQL18ySO0jXUuYwSg2qtPOC390Il2ASAfJv3Xl3xLKcXzDI/drY8hC0zcAXahn0Q8i
uKNCrrK8O+PrdSoMmytbbYoQJ3yFDKNH7s9bW0gU6dEaBMXb0mTtrpSwSpvl0BbknXnHw6tcsr8G
FD8h//Zipz+Afkzv90mMPVUIZjWrfJK0vUmHAKsi8Z2uYX+CSUvkFY8PRI7cpLfP1OMwL4zY27BD
wGYF1co4+UqnIFALpkE2Sg7XUiHUt7vXyAsxpZDMJrVnzBVCadoaUfRDhYkfnKWCeyi8fOfjlnQR
EmOSpl65kL1QkTg+Ix1YGsX1hAvNJ6wucrjvSVkeaUwKVN7WlNz/EqUEcVZcyLZvf4lHPw7kwQx+
5+5rzxczTRMB9T+ovFIbPzloP+Pdr9ffAI7bGrG1CUvFa5WmWv34KRAjzq92dDvsdxRbogHRSf/i
ydIcsfQKMXA5ba656cVQTtNnAna1pqSc5jYW+uTp2sqZjOhpEtLYeuheXgw4iezTGE3lNxF3aFwR
qIj9PmkNrXMOYstiAgQH31a83rPw2YrxM1uNEuuaDnEZrNYsSTXdjy7iWY9sc83XOG6nOWjivIZA
2KDohRxb/DOxRNhzwO2MZZUcZNqDp7SmmJ5dgEiyh1NgR/5U3HLWrb7+0e9n/ICnE8iscvxY2DvF
wMiJRbeXm6oLYP+VAQSzxwpYK9N3QkFymqQs/6uA3MrBjxZ66zOzjbQLrGy2SMKNuDfXMOsMZ6wm
Cto4hIbAFdvgK/hBaCi81rK65jD6n83n45bwPJZwRYxx7TKDk3pqCFHu3sWQZWfkvczF07wI9Nc+
fSroCOG3a/iO2Fx604hXfCeNx1M7NIVEH5eIFBKoANcFKPKaVfwLqyVy4RkrQ+AVMOoBeIcFr9BC
XTOjBUHu2RlNKQ14JKIlCrSKWiCK3X7zHGKv5+gizGOmtfbxmgIeAZ9eTY8wIa4KDmLzQiI6J6HV
K9DGKNezAjtGnM7rc6t7sxZpNUc70mi4y5smlKnzdc21XuMVyKzt40c9w0zgsUgmZ3YCjyO9fTOW
JF3QpXMtoUvQf9hKZUQM/4Wp5w7U9FVLLFTIquYFnNS4M0bqytzU+I2KhlS/pXZUg+FU1an6BdhI
j9WMIzG8BETNVG1nnLtVhpYQMaG5eoorL0LOeBwB3TQx9yXo6WMqGjoFQT0dCPeQI9tmKaoVhBBB
2mtLx/ulLMCtwbb+RltRp9Fdf14ppU9td+lSxqtvCx7xl4d80OfC0JR1ulncLskyCqga6EzzULxw
oI5G+0aMwGAyGyusPILJUUX5KwyPXDa2C+1mQlp/t5/gDAIAmmxSXUzpe85V5mKtDRU2YJceXMoz
rRgoxXpwUBXOSrwejbmhC0y+bFcU0vn4g3aEWBUlGHESolQx7QG/4188a6gJDx5N2TaK4bbIy9ed
OWlVNB4QXyU8GbwkXPeEeHIvea41Dhw6RIJWW+1c6bq+KwITmBEAvg+jkNaP8WKWlOjIDzINfgMz
k4C3XW0nIbSjS9O/Lm9tOgGhs0gmcW9gtHB62I2xR2g83Rt79uWtmntuKyEwoi/P7zfkrQO6WlYj
85HnKpVPvnnVmZaxeiPcVk9fqkK0RhNhyQC6sMB7Ye067BNRd53zNtMmZrtOJUuiOXU+uGP55Rxv
q8ZSwlQncCvGQ1dBQhqOjJTga5JzKALNEAc2AMV34iLZsZIkxL0fZtvWrHMsNNcb45FuoZLZKrLb
ZvqjYLB9SOpbaXEU34FNeWijX8LWwUT1xk62DZC7jHsLWR+bzeMhzD57th0NwXbe4+qvmNgZZijQ
Jd3nleXgtozePJfAFtESUMsVc7q1jAVcR/uRIGABPPVrkDO5wWMORPhbPDYyFEtB1DeBtcN8Xrn3
S3TfYn52B0uV0Bhg1ifz2iKZsUCL0oJyU/DZuMFCtS87kdSYdGlwM6UY/0o0bfEbauvvotpYqnOc
49KMGuc3aNhHA5++8ZR8BdiIfnagv2Xj7vEc6O2mu/APQ0DfXIhIqPUOmkBAHJIFOk6TfJfeSpDh
beeiUv+Vb4Oq3TfQHdvZIqfQ8qKpoi8o5I0gD2uZu3mzREHHNumI1J9g/b9MOrC/P07C2ITbJrOp
p9Kh57VbmrP7Vv1a+aNHSxYFgkqkNw0NDOHix+jqvT6VAS/TTPEvA3tGGPtej2Wu0m82Mm7ElNbN
DD7QrxNK9t9Fe/YGxMcdNEafnt53mVG/8qtBGueB9knsgA2sVlnxbRmAf34iX1C+rd1YVOtrp9lq
bEugEhMGoQ78wq6Q7RDG/q0XLeYL/H6O7uOS1m/ii+trVHO7G5EG06kPb2odIZXOLqTDiEFewPFj
smc6TIRgmWx8+6rOgzS6nqtEGLgFvq6V9aHTnpfgSpbbuUzLzmM4ypEmaUx1tuiVp+x6+JeHsdX6
mmDZYfepjOnUjfLMB+VD6MUf6N9yv+9cu7cZ1ZcflgQyl7fzAli9LtsIn4exrEbiVMRNNN5SEVx1
br3Q2pdK93E+znGsa3u/66Hb4haYKmGu4QCoqmwdAjzDW6erggV9dZDmslDw1f002SSCXX15rK9B
NghmqK+9JPfWtpHssvv2AyAuS/fzHZR7LbBKBsLAnVDzNVvwl88J8FL9QVVvR/qJsAeO87PpCXhp
o8a2AY+qT4ES/JuOwlNyLiFtIu1wQeQQL3pk4ewhd37IGfMkHFmV4ouhgfdTGHwLnSdxmS1+sw1b
zatnymepionGV4Zmu1MC9E08LPj/tizPHK+L6yS1W3zrWEcF8JGn4bR6dfuM8GPntUaCTfVh8H8H
uQBRuFzVT0xHtqIQHiRPs1GSjkNt2PeJEcuKVCbxqGVFiWde8jTNckwTXbR3+Bj9d8XlZlqfeGQK
bVbNRSK5rw1gPL6Y01dtX2cUZny8aKBRdJOB3zJHifpLG0RWgtDX/1XfbL8WGvtFj5JcREqPab4z
WWuQAPgjotDH6O7GLplCoxEKbtdWngUvw0nuzbQojq2x/Tc9LVRYlwJiiIBcILVYt/2ccz+Dd9Kw
+gWUpqtbuPJLU+nyf7G1KnlCDHcpScgP0uyU/4dh5iJbfe15kBWQSiQbIhMP+aau04yS1x332ZIA
pzOfd2L3UP+PdCtq6AXlawSX1XAlK1rqC57pXwiHWWetlSb5Y96Hzs1OOJYenrZN4N65d5CQebfH
o5kMkK7evQcLvzDi49yWfAPMXR9M4BqW74wkG24qhV5iYfJ4Arn156HuthUJ2LWfNv5r8/JmxfbB
mehrY/eO/t/UXSYGnQis9EMyzt3lC9FNI1majgSTC18taKC3vSfo7Yt+XwOpy6k8VWOaZhsA9zy/
VooFln1U1wTry0yasXwsrQHwIIwva5gxA/Ta5NeaZdSLkeqTrfJHKbk8n/u/F6Zz6sz5+2h2ahF0
Bm8nAQK56ysr5YqJrTggi27RlJbCpIQJBAl6XuJ0BaZBIUc7SF6F207hzlVUchuG6KfzlqeLZJCn
jIzoxw3u6d3QHMAZHkMI2qCui4SC4PruYwKm7LLI1cxSZrloz3Lqt87GyUd+xzD+ZksDDzQy2GfZ
qv3ZiJGXrVcnlEs+1Zs56nftoa/J9lLObk5bwcr5uP/h74EsemJZjrYccJ6GBBZ0RSOxNLxpIFhA
66zHO1JCPWpdUU3/K+FS+euROv1DkmWSroYMi6T4MTOtlYn/ms/ExtDC9Ew9DdyplqTQqIgYvb2f
gaN4TR4JxRdZTRVcwrXksFCzTyYbsCE7Gn0caC/YwLk2nHv4kma4vdYKMGD+1FEcoB6jO2ub7cES
MsOOiBvJ2TfDpe97rucnaFz2k4OlX/01dNlbDAnTwCxm0tGwt3nMATpmWPo8LAxHyDIX8hfKEnkg
vYlsGO5tSlbmh0X+9o7PYjs32NzF8i7SRa0HFZwlv+2pR0GMiA5YvJO28GM9G0ytkr7NOFvdi8lF
fv+2bjwqq7lAcORgpjnmVv3WuXmJrG7R2YRCfnJkdPkhFinKZZFJ4bY+f/z0/rUOYGPf1MRkUgzt
ODFhNh/i1+VJKKA9ThBklTyE0izDFxpGSoTp+ag9MvMjdpak7+ij5Q61PtOly7JAXD/qgxZpn3ZS
gKtqZjpo4Zh0t/ysjum9sokQYEV++2pMcyBTz+n1aF/X+sIbP7y6ALrqPFy/3ovS+n9cEmqVKPva
hUVwlnXkMLhF3r0lCc6Gocwy5dVr43F06m6GqFWOoi2/YMF1i/l3d2KCr3fxjzAIPqXdDavoH+X7
qdUTna6UzjqVZnLRKZEgfH7gVFD4NyKpKGbUoTt9Hbj45B9mvGvYaPGZHPKeOc3UL6EOzEaYyA3H
gw/shIts+MCESAuR/zmKqLWIhEefmTPReYv7FSCExb4ELcb3HJr0NGpi9ytv6l539TM5dmrhEQfM
I3hSuWmGzWyyK7rPIyirjKBaJh+ObuejX5xZg1NwCAs8KdVUj1Bjp6F4JEp6Dc2PaCFvPy1nvMsZ
BMfT1xIwCJgSfjZ2dPTH1jK2tHSqOV88JsnJIwyEdWlaqzdn7sqBR+Gs6r2+PLG5B2APMmhta/Gm
fY0cMyi0bGWJ2SYmRosSAYEEfJRDoiGac3jgvZcDle5vtxEyN4beaSuPM7eHaUPH6XkD5jcuXgt4
dRCxfbWBGE/bsWe4WHnrId4KZTrCCRTb/rFPWGkpvAk9rxzqmh0nTIqvfzSwzaoTJe2czoC4Qbbh
nO2Bv+DEHhFcdJCZcdzg4yVbmfFD1JU1C8GVNO9ILiPPyOa8Ar3AApfdjtDXAZDbsdKrIz92dehD
Kn8YNOuYVbyrZtbGjLvxeXlP4KnCyzeB0AGbOaDY4MYiYiQGDHCmMjejuNJv9jY3YTFWvWBv65AZ
vUhLFdeEtH0dPeLhH1mWDH/qve2XxcbWe8cAZSk+3PHB6Uiuy/scx5y3vXeLrtDm9RJCE1kMDjuv
arm7qjzXrv0p0ngKTejhmTlzs5Ozpai2oGjfx639/nRApCQ95jwTL4UFeZbbbvPWMmlE5OqUedUr
q9fYYV2XzxCTcxA073emZlCeSJctGQg+tIzZtcTI9O1655qzSsdjVsQf7O9Xb7J46LORjuY+EkaC
t2ulK/UsBa61+XahOkirJyVV4DYNNjSjhtKK52YCvs5I4mbz1paLyW0CPzUBRUkZAolEI68kwzFV
iy3C0OCuaES9X45ib2/0Laf+Y2qYbHSVn0+VfhMXX2SZwd884TfVc0zGFQKx971WaNCvA37IKMKz
IQdFZeZFGw7ngLXPD6UFEYk35CKqfxARdpeAfBZ/1qquNPLfwEuFphjA+VDHu9P6bYf3lDbllGzr
8rXVCS/33oMgFsy38DOm3H5B6iocjuIj1PWZY87DIn/dKl24Dd1B6/uZPwDzYTvDclVlQYFgwUcD
U1hm2tSbPYt4qV7L/fuLIk03R/W4BE2Utv76l/nVt/9PYPOZlaT6POrx7YwxJgUPR1TxasTm8Ibk
A321ZLxZY+4RzxzgCOyoGV4RjBFgXNrqUSzt2R1IH3PSUMqG4XXCVSby3kWGJJtBLM95t6CZ8QAX
XdYwY9xMz3bhqnpyk7HySwo04jA45/mKXPl8dDBROq8eHDFElt94ILbEkB54QNEQBu2vOSPQqYoB
7D4UoRKM4DYutmAD3Bx2QtPpP/OY9uMLklqszOX9KjHw1SDHidO/PqtFl0lcCM5sll5rjjb/pJPl
4U9s0G4VVnVzvh3Y7U23TKekPA83mcZK33ndvN+g84tzKti+7xPcPQmANNuJsmNJZu49UXXsCD1y
WsLopwkhcl7xBCoax8WRApWFO0L3ky4j0hJbWWuK7vjHF7+vOYS6tTPnnWmSalXoZfaaspUGJLEY
m5eabPOSyUdzwLObfHwKZrZBfectIB6ZGoZqQxrTUZjldJOoN+uU17ltewn9JWosFovdK25yQBpX
sJMUn0RikA8ZpjtB3OeIDi70P/Nctbv8ym6m/Aqdg2Ub+mGSLQNHDy5MOXROerXtpTqFnd74x6I1
vPjMbo1OhGpAeNY5fr86tII57BXEhpTrsej28vySK5E3RFxmSbzFFPzAaPz292bAq4ZA1EwglatK
xLj0aCISudS5x8VvZUpsif6lKYQ7MTjeOSOHKH1HsEa6wWBv4PRmzCxYJKMr1TSrJLg34Yg6CCk2
SsyI00ZtUt6zW+FQnX4FBVRsPchfCySicT0QGqBpLeVMhlXJcrjjm6L1Bk6p6v4cabJl11nGBY7F
WJulJUnrMYF4JMlxuo32/n/85E/co9TgyYYm8/TI2lUHLnPZj3HCYdFNeoKzessoN4uJx6zyJggx
1bq5NIS35Al2VHQaB4+Zh3lCwaLTwgQ+xIadMiRJeToOnc7+IouVHxpck4RcLgongid/3+at7zKC
jYUCk7gm8VFYNWF89yYzHfm92pntoFqguGnFRulyHxthsEI5vvT7LeT47RaZzali3Saopl75uayQ
WbCEW10AC68r8jRv5BmYQ7SPuvLII4w6PVKnCvg3EXxiOlsyMEj3bbHy4UHI8AT64pdSnMXKfsJL
6pOIUys0ZXmelcnxpcQ4sVF/XVVIZI5G3TokGOug76ttlHnkb7Mxswnx8T6Q/knXmGP74xwboMDy
bu+ctFdG1Xuta7cJpfVrEGoTkHeJY/10TDrh+er/6RtJTl0i73uL7ANt/8iP/2LIxJtAvCAIu5q9
j/A0wVkc9Njj2tSdw3+yrMhoOBJ7e2kA0pMWtqO+cXYkhUofxc5DFbbYrl214j+ZLBu21oaMMplF
U2cdR+4SRvQJtFMz5Kbj7TU9V9/2CiNcTuvse0Dak+HSGk3/n57BpvijMXUrqd+xj0gVE0XYkIMq
agvZ4wUb7qNCVBK/OEdSkgV1OjgzkPtP4HmRMsjS8n+rzRwMVogYhw8G+0QB+P3ASGG78F9XEIUq
Z9Y8kBqTeJ2XzAUan7lC9tsLHYsd2hprTkgy+75SxjgIKvqHSU4PtgU1+iw4SMkYzZgAcicIBg3F
7ttW1wd74Um+b80G57JKrZvSt9Lq/kKWAPYKFH9Xhvd2lI4mcuo8hIdcvSmtqC6VGg9riPfKoQtz
iLWKZnFzVYNurRACiErmKhkKv1x5NrsnSItTsXbtOshv1kZaUlq7IHyY8ie0kVTSCn8wjt91bBmY
jW8X6vNOBUg2z2stBFiMk1embYiYBudrnQynqVpGxcnsm0kW//nv/ZbUHsTxiOMr3UwMF0dKKvmz
CwsWd7zqhIDmPPufO4hZjG6iluz6vrGmI3Q8KwgFBab2x7uDfzpTx7be4nulNXwNZP51LbIiQqNL
k0lTYmtFD7ThveuE3QNvcGY+cd8UNNQY+J5VRjr1+HRzznCQAlAuqpduaCwmx7M8m95V/9Yhh9Gq
0dztqSevNL7db/akHehKZytTp01Bs1B/3I7Y2gfsmljMbH9P/+8qKoZ+eZozK4nSSOrzI2LhIF5O
sD2g7kcLqfSPAjrHmGfU5J12kAAw8bFZSNZpseh1caOoK5p1EcXCpme7zGEZMQBZfYyogSZzIAiW
gQV5ZqX6/LPDepI9NDJ8PSPAT/YddzNpfPX04fadSQ4fs3jOqq1mDQy58kkPXWUR7LuB6xSqSpnJ
MpLZEQyLs86D3zIZTEsXzBwOQH1eVO7UloTNhIe72MvOdwymBKgLlLlZ9mqxKFDBqx8BQ42c81H+
C2p+WC3SgBUGdBrB9Qg7HDVHfMPT7KibeV00MlDznxLpaXU7YdPabqTui9tKvwaVy3nXdxbHETfq
xQU4a7V5n+ttfuOWDqlFjzuZ46NYYvNZxUnPvaq7SeuZJ3RjD/GnFrIKgwuUMb9GBsTwWEoRo/C0
z7fe83I1dHOwqCSodEdOUbR+d92mcwIMu91+5TkVVbO4+/iKGbI9ZXLGb5NLAEdPv8qfsMlhM1Tv
BVQFfGfErGubV1cEbR2Ovquf83SmU/oBNTejdHJeAnhfeWrbSTqIg2ueKKx7O/uzi+ji/ohY19n0
DoObSj/+6FQxfg10QdlKOVytWJ+y52WJTW2cKogj6X7kfxGS64fxLPshm8jE+NVq2hxE4F5I1O7e
KmNRfe+7kK/FTo1A8LQLd1IyRyBaJyGQAONRsevA7DPGI9r7I/f7+21V4yRf00cJwdfkTmOdAXGI
1zF4Elo775tbP1XcnWK7vEnTtOUYq+iCdGRR/GZcnchsxXvjXhu7zeWzkLTDdZ8pXfrKsSybKBOK
6D8IpXYooNcaW1mRSWckmX4XT4ioEbi177xNkXeReAkiD52pXRsiS/ChdxufUv0DFmJQP13s0obK
+KoSFuQeEYYtx/lEQ7FndlX9KSNZA+krmneRVDHq7HABais9i8UOt7rvmNKBn7QkL0KB5Ky9ps9P
Rec1tFbF+2qf5DTSq2UrhSvN5vS91WX07d+dFYUAFuLfHxpg2WBN+mlROOdtN62LkKbyulsMz+yC
GBQ3YNxCpUu/UhizHVtQmTx2At6uDP9q/P6/548L6ms/Xxx65enkxbdTnc+1YB4Zx4skvVaLi+IW
ivFvNgdwMf7v1pbGR+Rq8Lpas29Xnqz2X+6L5X2en/9Ellp+YTix61Fs7KEPDKQK0TogPl4nLFgW
x4ylLJLMLiLqLImwZ7JLRnH47Q3y7CiW9Wyf4Y/1gASPta80ujaet3xge/YsTqThirP+4p0mnSPc
G4yAxcaePQm5U8JqcV+YYNo+ZfyC7w/pFYVrU68A/BJozteVMan2fM/7NlWLReAO42es9Rf5jXK1
u3Ek7oD53IIJHlaTetThgKtFBP4Hpg/62f1w/w1I5IXA4iLm1iYf3PaxOeBK3gpHM21kLIfgbcq4
dnBqdW9fcW8i8CBvQdnFi7gQammf2Nh8dtDzytnU+ki5IttfGEwLP4bq9u0WPBFhH3ukBlRMujXm
JGu3sFVpbHs/oH8CgYdAvg5GsLnzYlWVK+xTDA+m173E+JQUtCdgjquHnM4PdbdQGbkRcVS+w6Ic
HsXjkPhrcmmLnet4YDP6cHiWcHEUv3tXIQqN1Vq7K6aCdtwbv/zyvTI2V2CsS9U80p3rbMJDh++G
URJCW7Zj69HLkQw9Cc37jcRuLtB9f1aNKKxHEJfsSVyvkESrI3Ls5CFTgfhExDOefMyPUnWGNvpu
YYC+l+tJWuhRfxlWqeuMdpEr5DJRoNH8RbuF2I5wptFAk74LbkputbNZ2lPKCTbB7je9YldJK5c6
7hxqIvsCdTAFuniB0aRWKbCMDjOG+tJpGTBSpnBf3kMqpA2K+aaCQ8n/hHrWSPN8tnfTDWR4XdXe
ilBO/J7VX3Ql7Xf+5f7u0jYWK/iUrsSTWlkJKmcU5flyYWgfcaU8hyK4m+9lcOyW4G4oid90wHrQ
XQcXfqVuH/QYdMy+i3j2Ad/kneRXVG1GE5w1cHxv7Fp0yh2Bwm4E6pN47jr+3peEKKBkJnY4u01q
tU8/63V5iEqaRNlOgN9W1A2r3AOAoN2vmfcF7x2TeHQlMrLqLzVjZevCgGotiB2nMyj9J+fDsqw1
a1xoK/KDcvcrw/uwKm3fnjE9Ocl52J5AjHorjb+swrzhmsKLhUfuVyxylnw5fYVzHWHFrYepJceV
rkL7E3IM/48TQpK9QT5q+KOzs91odHyHza2Gbz4Xfmv7K1PvhcNPZT4QOykdkyywLxuB8xRKpl8Y
vPPJp32R3Kx4oyl+zAZh4K2vHqVLWwmxtCsOgD0NdayWGTlO0k/7rBC0rym8aZL+fxp0R7gsjZpZ
9f+4sV4G1WTzfCxjTZ58fSYug61wTwEk3jq/DJ34Tfyn9RTNDeeoy1hbOTHDzq20yLqfIkbnRDDs
x5hd/hCsOecqgH2ULP1n84k+seO3D3XoPVA6w3/zAWAklkfX1wp7ZqKdWhbJpgXSNcyQ5mjd2nzj
6apGftF6aeAv/gNtRwPeE5YvkBn0Z3vSwXCl5Ln34o63QM9oJm5vAZcknqEGk2+01a5P524jzViC
NnXa0joDk3S0IWg+A2k7rkZq+1wqxWGI9mhlIUDj+Z+PrDYMeH6lJCWbCaviXcXfHXw5yd8jyc5n
Cv2wLdjlyxifnlTGx13mNpA8YdMUhlmWhwT94Hach8XEnHeVDIZeGFHx1xtSEv+vphwJBI94TiVi
IUvwzYfjGY7B+7oDXyFQH68rAfxYpOFvyFHAffOoQG3/fTnKHH3CF03vD6w540ReUdvtJ7jFAyvl
hSzg6ToIjmZFhqXypU7yzbtAKZDXjLNB7RAdEikJNUolmREGqs8UTlgOiu+L9OlEpFgDz2Szy5eb
g816CyRofGjDWWaIiVjmuG9f8fuImmKcH6iRvyIN3i2JbzHc34hGGXrkWwF3+IWEqaoe+nu601fe
ZPt8oxMtYcqByi1qfQftWMZIyjQQC3xVKj1Nzi0iE+rSmdnr9w8xr/P2n0YcbbVWKV62mjT3UAFI
dydxqeA7+LRwL229ztENSxfs/NKif+OPqJobr5JTlCd1jbGhwk39CuhSb2mrsGVaUIWP0XUnhRQG
+IsXlAkZM8/6EjBa87YcKvGE3/0CSbKmqAATF8u2saJucCGvY9EhmrWXRbxEoPIrLcywTC6G605x
8ktLJber0ZslnQkuxCtQ+IHx1oYqIi0fviNMkr0pamtb9A+SjEPHfXJ5PiM6D73NQ0dIyFB+fzlt
gMytBIdaprsYwq3EN/zWXDNwLs2wAfvzVQxsNtCjZHsCuxfbCpv8FGUgJFxMg06N1YwZBZWwa0jT
GuM2fag6umnvzuIgBTdIC+oZa/YQH4Ao0VHx1AAQ4KQwbyzMsq4p6gMUUESSEfKRCKAIFlhJ9Q1g
A8J0ViSjFnGThAKvFLtwI5hrKT3iCrdqOszbxGq5h5XRzAj+Q4ZJA+hWBawKib5yUolprNq0ZV0d
Y8LIIfBurZxp9Tms4FNweACBayZNh3YOsx615pVm8HZDlv4Q32Y/rHhW3/2054QTJ2xVY2Znn4x6
IhPhFnTGvXalWF3vz6ilik3daSbmy1NfzsARVI9LVGTIC3MAjEbGJPcwom1xhfxvmfg055WTefd4
NjLGMKTOEG62seSj64pXL9bg2G0UGsKg9OAacI7WiytadMZccQdLgYSvdZpe6okB16M7GXmQC8G6
OTzPPSoQ5ruAjTmCqrL8sG8rpDLqIpJryH9EPgwmhFVRoxfdyk37O8pcHOessptqefW8/RIM1Jpa
gamW+2/iSdVRL9i36qG/lkCJlNfxyyGWbXo/+hz9ruJYTPBLatn35f9iH9eDTRXlzQ88lgT0l7s9
5biL1QBmwHkRFKH89gF4o2hoKWYVOljKRyg8O7mHIpgp25E2r8a3wV6mrmdU9cCVM3mlowhnxwQF
Y+HBGeT63euwdp3GJ8jZ/ZDYXUUPV9riSNS8DJqW7g5spW0deEZ+As7kJkK5wyB5PRCvjSLKaiEL
Gxvjj+RCW0yYmIZoUtTeBYFHuWBTAHiXPU872nNI8wUjmnoN6W2NjQnW2hL0DdsEvRFpGhPj5AMU
fZVeuRgPMSYhTX76ili7/4BW+c7dBp+M2cpqD32fc3O3uAY8innr/GJT9+YC6Jj1jIxgvhaHTjBx
72GFQTPZCxAL3gIwJSkiAd1eJM0w9BdMdRStmJ9ZlxW7KyZHsKtDeCo8mR6bFkpcpVLj+bAOztnm
v9Y29UjLpCBzptp8LcGywkHESMw6MWZDNe0A4VTaNjRpUVatTjcW0IqsmhxvQiPmWuiksm9LHG8E
bRnHRcDPCG+SMA69JWkvxR7v4X0t4sJGTaHKnzxFOLFGfT2bCYsxiRhj4ixD+erNUj93MrVtbwVE
0mofi56nrvbDNph6CgEQF5LoMih7A2FCXbsgCNzeUFtasKsb/sgsZ0jbf80kkh/2pLDhXu0Ur8Mr
XZr4iYTATGzVl7uh3f1gxr5nCFOIK9pQvHm9omj3YNAzlSyyJGGlpibAXToMN4idU1+VMbUq5U6l
QLsxIYBkaZhD97oVeWI8i9vdQedvYjkNP2oKynkK30QSZ0aw3iO53o6urODni7HjG+wZZfrbALQP
BlT5N4n1VkSVqDwdigA6+JcQ1GxD3wilHcjCzk/idQRVbKbZa7dZ2uQ2Cd1EMSYeMpQxNtibaJJ2
qYhJ147q1arQTeAt6ekb1quPT7t4KFmyeCk5PKcDLrs05PCmwdAIYbRu0B/Gj/pGYKfe9Vsm6t/f
VfgAkyUdR+X3Zdyv8bKBPkxno6B/qgJtIFM85nmY8fvmVbK/l1NbFA6nbyzg0RenAGPm5ikD6n00
k1nCS9dCV2iIf2hjgqlp9F1XMbMt0dTV+DpttkMQmQOyP9Ez/pdg3PciNdMVlyPHSuFC7q+zF7WC
82XojKUvYE7yCdz5gnDRIwYlHB7g95FIt3XADgL33Q3y6mlI9eKnxIVcemn++GkQcrBCgOfzePm8
qs5G8rDyzXSZsKu/Yfar4k8+4sVQoaq1QWjUpB0iPbzaCiNlPg13q8IGAJfjOoKZQcU2mSNac7f2
Tq8wklhT3rI9R7BD/5LFemTweOimYOCUARJWxk2R+rWHAZEIL/Q3PkwrdPExUPXQvTlRycWhAtQX
sYYR6fNk6IO6cQAIx6LnhIhroK0vI0pr6pH0oDPPelhR7KIdLDnwbfygCbIC1/ejymyERoq/InMb
Jnw//AKow79MLb5iNlfAuschsQd3HJvYcKWAljE+aZj1mrzK2VF/JA2XjCSaLv6VyUjMbUBDGdMf
EW8o0mBi/VkKfqbM9gYSsIeyEfGi7l7SaKOD+eypFSIco5iB8h3K/LXjfSfLDD3V93ipl113I5NK
5ZypW1FWBpn+QjydinbWaweJOopDQdHHHRG5Xo613qaC62ayHfUcU6jyiglfcbSfdliBeA76XGdV
caRRifToQWJDO/Gktbv6j7RFTKal4RwntxrVtWwoFAhM0ehbRbG/iFEfjhsf1/I6nleAdYkB3Hgd
PUvhqToqzNPN+ZuPe/V1jK6BY5b4uQ9bIi2gFmBgLcSPrJn9nlgDJbxy8T5ck56a2GIkJ4Y5DmA4
pmvE0Ax+WuQ8RvW1y4gqj+VPnPO3hz8dWVGvPGiCqjnaqQkjkW6kq/c2luHOvesKO3g0iNCHqpqb
YdM1pxrOlokmyUZqdzk0Zbhk63W27Iql+3TpE2ddYn0Ld4aAsxPMa7h2+5uFLhsL3YopG8skvB3+
KDMJUXUtdUEV36EGv0CZ+1YYnxi1EfpgCU2Be3EhnSPm+o3Jpzqqmn3nRV0GMkZoMOGjHAmQQ4AF
ESTmdu1LsVNJ996YvhfqVGVQFxF5LMvoOAjU/0pb/5b7jJHzkE1abFkk8UyrjtNPjW6mlxuQapvY
T0yQ8ldLxbApfA2ho92OEN0f+gNAGOKUz6XyBSRDMERTAYqwYKn4YzO3i4sQlq2vZfBUheXAKDm5
fC4FCWTQMIJ3olhg8Ws1WpooXgx3o9LretetxOJ1bFGkJaT2+y/gAA3jUDYRUsCDL5r36PZfq1Xt
LKOarJzrOotMm91eCY2DkKEPm6/nZW6+RDT2gZZb4AKv14A0KAiC6iNGHLAooooLP8SEEUclpJQY
3bUasLZkrGE7kJgA22QQvNwN9J2G2H6hhnc+QyYy+NysAGdRphc2EFfnhNyJ2LKy2XzGLTXJzW5e
kXQ4HhJdHDPREAgky5BRK/3XpQQoXTk08M+MvcvH781vxWtJW26MkX0W1ZJ/N4txxKo0PfnaXwI6
cbiaJTODRdKrTb2zbcaqyJ71kzccrPWEFiIbUvHhOQTajS+UnKVmu4m9aZpAa7IupYUzvMBNbOxG
rUUidd8h9dCr6gHvnHBPqbqmezhCUaz4rjhtfRORAbOtVxMz2i2lwpXa/Br9IlymFQLfKi0P2qb0
nYbcPgVgoMGvdDtoZhFNcpvJDy0h/hS6rFIIHdgMVLtqtcC6QATESLe9QdrpDv4ROdQXhL7U0yn9
IOSbtASEMGRnYOfQqK2YeRA2/gDBcPvAdo+tst0OuaFE4R0eGWmtsOjqPJutVYVU40dR3/ZtV5ZT
N6YGyEG0MCJc6k+W/DH9pqv5E3JiYfPrOGTXzdGLyi6NKCuyN2P7BomPANuU0eJCsKaaPK4EAcQA
iI683JD6ADchxt1LsRoiGeRkQIqPDwZjTYQJHdRJGXV3LO5vVdx1PiOUF5eNgulMD1s7dqy609kf
0Pui1Q5wYZbYtiWyha9b9jsiF/ztUJVBveAYDpoS72NCrdJAUHXYsXO7XxukplRq5aVLoJRAvVP+
gu/OR1y/URlNv4lfwIf52pBysSCGOgeXY1blqVw7fxCIQSC+bRK6W1TL3D7wEacU/W9m6pNslJd4
9tczupJapvA7dapWiZBdJDLEnHco5gyftuqW3ELFKXIH+BcLQys25+/9BnoLaNrOnpCvHjCQXC7k
yHeuokzhvhr1kd60SGLNJM3CRW5qRbOD/ZrTfDKHwtsuFt7qMzPL1dd1s73wDVdLMeDu/zHz3Iqo
Z3G1udbOTj6ZfX+YuiW0wAbOpGILhh6hLDjuUqmpWJGxRX2EdeSWP2GOz9UYONJLdCD0U9A72z9D
E5MM1Q/wUOjrXuNEFGLmwHgGJRtdZftUnks3XBazTzXvXJ7ysuSi2CofuL0uOCBwiImK2pRnkeao
DZgvtjjcG9P/4UbqsviYdRPjrsZRNpjQzQx8lciySfoYnZkYmZnRKZzAw819jQIWj+cy5QvIjCzU
KgfqM7SKSZ/PJyKWbcc56FgVlOwiBSMyMwkf20DdnI0prRVumRLLo8RjtGtQYkD/2GgGwKLiXOcN
3Eu7ZTMMQu7db+S3lkVPvVF9M4nQPM3XPVhfQ6hWdepB8uPlgzjhLvsVWosz69VYvevA7aBkKyrG
SX4Sh5CiBdhaSxZg0NONkbAC2h3IzSJpVhNiX4itpIDAdhuMdzscNoqKllXGqAlfbLHOPxxzzZll
t/ZAdhc4ENtDh/2tuKruw69O86r8VpUQXDOTXDI98VemRQlHekFxLkRzqmZ1aJwqk0taqQp8anqU
mg/PtP+1J+rHNwUf2jYdT6J9wYQg85M+Zf4r9VhVnJdv6CNX2pQkklLq5YSWtyHweK80wej3LDDl
7uKJXsbsRG8aRcakBA8j1Fr8C9MRbedVrToTZc27+IZsvNqYUhzRASMI8rgpCSTuCsBtK2A9jbOA
iLhXuXnm9AHJBRpnDuT4QehQ/M1hGzmoNznUR0robm0fXdfdSvnzqBIefzMf52w9SWvvzCWy8EHA
KboJTxzJm2gFe29B/ETHKRaIfm7T6ifTUfPB5auy4vlF7/4FzVdLX2SIvFZv4qe29Y9/TfgQ0h3B
dCsXPl5auJXgs2JeutUVF7TGD3h9H4SAaEnkVg3PHPvLMXteuqhEUTzz9e//ThziwGv0GA+Qsxdd
yFNf8I9lwyX9EK32fjrSlniByQmXhefAxsvcR6N8lJq8ern8UOZ6gULf/psdWkALklg3gfM4XznS
G+8zbx1l5Jg/WFVBjF4V+lgd/1RjWyj4mHLUd8M52SygFBUAQ0rL6IpcNpbZ0xz533Cd8olIU7CQ
xOvlZgrL26qPPXirsxrqrfejPLpIe2j6XPfeXjp5ZTvZKcpaaEMYg6ap8sb7tuctlYR7BzSH1puD
vgSqEfubcTk3d2MwTj9vX0OxDXcDcQOOG/jbDsUi9EIN6RLZrzT1930H041+L94hC5mddg+XUxGn
3JsleiwUsnzuVVTg7Oqw1v36HybDmZdejTzuAyTZhNju5v7BOXkQR2St9RYolxY0HYG7jP3LSd90
CgATvFJU+mVzv/aG3SPWpiu3bfKhlNBmA1yDfPp2dKd9cz35uCc0xN/L5GP0v/4RTD56tQsHjwP8
A9Iu5NtQL4eNxHXnFtPFD8K49JRVzBNJS1e8rYIDSwWnRkI7kyFWvfFUTchAbD/B9FYH4cGZ6Atc
O8nIgQp2I5eJxBt6GO6+pAI64aZzK8bsVJsXSZMFzfCJDU1Xw7HsF7WuXgP4YwTUH/Srv9GC+nv8
tKUxVtWH69HYQ8+xIHLumbz/RHryscJoP68EEq16sAiDNUSRgMzE4e7VdrPf+l1qXGv4FFb7qq5z
QVZryJLF3Hc8HNMlGUJw8ae37E9oSG3CUqtMNE4cFkhYq4VyQE5NXS0uSQOSr0IFW8N0/PxvMXeB
ZogAqqXzk73BpLh1sCAwKXWbS7dkGhdlwDaWeY1vgcEut2YlahMc7L+3EUh4qaglvalYBK+564OI
ZE/goEMm4IJXur7nj3Yj81Gjtjbyv1rC92UP+1nV+XHPfaph8hX5zGOoYqM+cb5xR9vkoUI50YKP
08CIzjUqekbE2afKdsnZSiDs28gkRO5Zb14jXqfpi71HEIdxtntXhb2hKJw60rpcHwOW/7cUemjo
nxysIeYYEbkNXQNmNN+UzJZTjO0SJGuKy73klYiIXklr7oG+mJD6FgBPgwAgbr02k0zexYE3Wwzr
ypT2YwMemgwQPULzA8Y+8/FPz8OgbO9LzR2HEty93appzRxdxURrYsipAeDYkXZFZmOU9CotOywm
rckWXc/xhE9dRIKhVQh4r+3HysSAP6vm1OFwQQpmjx7+VTvh5fsux8Beik/10B35wZN2bQArokTd
E+cfxa8B1nfgxT4b4hLZGPC2E9HMfUHpM30MTi5oNGLjv2e1bCkoErbfNYY8tLQXdyNNsreREsAx
Ehss3HrXVq/UjQUFxWBYv6Ooc1l47ofdhDLXFb9mIE0hqZ4EuuiFmIsBrIyPDEmDIZGUlIskUMQ7
AFZuy3iVWtQIPhVioW5ZIpAmy2dlpgbf3bdptGJonKwyP57Ad7+GTtu0m3SGIi1iSdOZIk4jA7eA
Z989B8jUM3ewCW6N5E73Azq2YX8iR20XBRVvtFewVe7JOZNu5z+84ifvWg6jz8CBBYQReLBJW8hD
aQikttnLHasqDZEpuqXaxghGFN/ErcG2bEAA8c7RsbCkGv2nLsrhg4m5y/a6OioV9lnuKayLMLw9
vMMv6tgFgR3LAvb3SjvA0jZPsmKLDcJje4z9n/L4bgnFEfR7OoBQyAsaQCAHqBdczv9B3GRR6rdO
T/QkYpYcaivfydeI9dnhCEgkwv8jg8Qoh93LH24Ch9jsPGrdGUMtUYvi8IjDvj0N6BrCZEGgoyBb
lSAvmP1pwpV4JwFsEdcpaaYI0K1qoxIaQ2wRrKMU/G3F5iVZ7DQeasrrMNvj6wLsIzZf0ygbKkgN
P9euohLa6PKhvqitFv9ytq/5Gv5vXHqIomLQxoR4HTT9EKE/juRJBLdhvJ8uez59jsFqusv69nE+
DBg9DmN+f7BuheOtHADZEbzxFPEuB3onsVguSjLQ4YJgugS7RV4Kc4s6pKuXfc6kiHfcrUOQSYpE
WTD0VKbuLSLmJEuvVE47MM28D10C2lztrdRhy+jYvA3+Qz9mLco7Q50NZbFU2zPErpfMvB6kDEOO
ZPKMDNlVkjJ79vWTje/yZvf+PKlMCYvgfeNzHhN5u8GWFR3CfJN+70vLAtCynjwVC+cTYAATKpLE
+AYU2Ee5fokEbm+Nz+HsZDkQC6dREFkANSUKQ3oOB1GdMycSpj/TzhKzYipGtGOMWK02EVuB0d7W
ywv6nn0ECSBzq/M+DRdGbbO0OVePt222x0R595jHcemMT8xHrwlsT93JAexV3YFo8TbkpwLYZ7WH
SKY3KkTpziIsGzzNgyh7p68XpbTV1r7dhai5nDAwrwZGb/vw+blnZJJ68IgDU0ypdG9NsvwU/PBF
6aFcBI+iA8V7+HkKKk7Z0ULQXcqmXgVeXBqDZH/SDBSk4t4icMb7oqpupcnXgV8KWZcNT2yVCW3C
s3JnPJnlWhjCuUQLjDK8MecXhbdeVhAh9ieSgYtGv4gC4HPNIVHVr7aZtVmXt29mBt1CSfW1VCMm
9mMR+/pYQoJhzsS6KEZFVBdYbxwcl1LgCzo3OXDzMl3oiwclNTI6F2400DMvKvV7ROHzv2BKePIi
JwWyapN/P0c4Agk/hGyfJfKvRHVpJFZgY4xdBF1S8GCEfWFSueCK1xq4BAMUtqOPytdVXmKL1Dgi
4s//YvaIfitaBt4E/EPYS6KNhP8iCM9ypLX9Q45h6PcBwquiZvn/Y3cCfwfKs0/tfvZBnGs5UK6z
SqTrYlHQYKYrJSED/dnJKhnv8xgZ7DK7MD6eo1+CgmhnfLCsBDBsl3OnlKTYz183B7gac7vEdNK+
37FzxSIkUiHiA7cE9TtRXk/Ddut+K3/NMB5SqYhVW+zCtkUVOjGZNqUNccO2kMJ+f6Y4C3mUEeaA
/gZTL+4kEi0gLEBK4+EzSGkTK4XW0OzCNHBN7WgLdGSPyZiRk1K5nCOEM9qjEiQSqJZR53avgWdR
ij9mXzv3aRSD874jAI86MGmMa4yRBi8CQj5RecnVI9jW6cwi9uHJvcBkgvhdvugd9Gy8Lk0hYvUn
o80s1Yc10eex3pneHayq2NQ5kmPCjKnWtuQbhTZfs01VMnLCu2DAJUrzy119wpJRRUM79LeSwXrl
o1ahjpkctnG1UunlEi/E/wk/avB+SZ9KWC0GjeN93CpyMytYutfVEqTTrqLyQZpFIBNWhWS/kRwd
mjddNfDdjw3Jt7b1npn8rL+80ffF0i+N5oFNBsKmZcUk8hdLBc3kgPORaQ90p9AhY5Tz3YXpGgI4
QsjtekwHBJgMVHA4IXD6dIZiDkRdBiV02TkROCHUcROgsQwf3kB75YNg2yswhBozOcfh1VGs56KY
unrKkIaz6HXyulB5tesezr781LV0UQ8sDHEmqdZOtrzuuf03QI01dyfe8RrlK6BYCp9mVs8Ixwu+
pYGsdDIkv2k1EobGKbkURgkPBSrcN6R6YbxIPYM43KUhEsdfcwLzEc0KrQLH6L2rwB8eiA2cQ+NL
iea/zn1riPcRPwTGQ8JHJpZ7qzE9usztHqQMrObTWjzxk2Le3miLLvJ6pRQgog0MU6ccPSuqB3nP
c0wQQP5ZUO1lpWchHglW+l1tfy88RGBbkvEPYSST5zSClhsZu+DslUzSj3AeWDlW6cig3OoGrQvN
TLDsTt+IGTOOqoZ3UqDchp2BkVbksjJdrXerp9CdWfXLYLDAOAQJqksJY+RQNjynk9bx4U3a0rm7
hIdP+uzPB0kvbHryJVmpIVoUQP5Mqzj7Wx3BlSwj6glOHzPoIMaoX5lM7Xh9v4zu5d+jqj5QbxCr
34Df6ItdA3MvoaxDHd6T0cC1QysdNfFa7XervNYAESe8JtNE7bBEQP0C26cjbRVDCT/aXeKft6UC
bmVM2MxY9oT5yfhkszDlbU53MiJsT+ji04XSLZw/9x/LLZBUGavDjTHTXnlONXJRZd+TkDIYKnGK
RBYAQXEWjVMAEY96brzKVhepWzUnfI0+KAhd2BbL9Y9vsRdAbzignaLZlTyVCy+QWku1Fx5qD0Co
j+/kw4UZb57GNXSBnwiEjU3DajFBaUASd8QOn1tp2Kf0eE88AGmPeMJ9nPZI0PyZqCT3ocxu7P41
H8MbhEcdlp2VwkFqv5T4xZaEkTi3Z+7tfkVkTI0YCDM2zHzaEg1EKSGAtz6jvew2fK2EFDb1Q0NN
Rs95rA5UusLxUlXLEdFkz7izWXsuaTRwiDbfGfywgxQjm5/DyAWYT0k52LG4fUeyVEQSK8+SSO0Z
u0oK6kvrthr7TNFHWQn5JSzcx9P/gtCFs89o3CtuyNAmMu6dxTOzsOPOYSNIcTsgwRp6jD/pqRmJ
MYdRxCRVw+A77+PrTFdFa+eWcvtFitoP1WDPWSCp+1JHpek+lmPOI4USOlhCM7aX4s57yxB9GmL+
tYPjqOXhf8M4513uZnP1YxY8sKP3Dtt7VLZQfFyJuwzg+UAgLRpmmIsdCzx+5xhYidrlhhseZNRZ
1JUymxmHPSNFBuH50SkODub5ozM8R/IkE5H5cOz9Q+Bk4vIC4TghuWgCvrj8KZWtYMeHXtAkXDVi
JnHmWikOyUYC82RohFV71rBGQmKGVVQDHE7cXnKMXCZLn9lqt1fPJPFwn80HQXW8k2PEjVzqm2BH
TsWL6hvJNruAu3+GpF1zj0t21QPlv1o4aNzaY8VnLu7YzAM5qA/XSyiXA9fStfETqVkqqb+/GFTC
VgSysuSsmcEn8A5sLWGcJiCBDaaSZKVfWLoh+1tZsMI1sumcJdjSQ0RQMALmsUjP/ZaFOvkbF/79
QNjJAJCLfL1aOdyRC0Cpl39Q7VnHnrkAsZayDbkuCceVzvH++lrPhHfR5vPNb+caRmg7Yhouay7N
1pmvqUuCgJMQ6VbxPH9dlpaP0L55mcuJnxcmpjlS5biPXxF5PRT3JgIiHuBPWqKHrxIDfqV9lVVx
nMj7q+TOiki7FUNsvFBUg5L1g4johxUQzl8X3whui54sryCfRPwdicYuQUs+vBMDkzK+EMWdPlFV
lChN8Uei1A3EW3GUjiqyDhsGRmQGX5ieIQZhFTBzSwHsv1hkPZxV26AI941sCYxCF8cyXCcSjNnM
KNF43YsfssgjiWMx7MyiCCgtFOO9gyffCdo6j8jO7/03zE0IMkd6fBEMjSantrNEz8Kai1qLOA80
paI+RptsXXaC9wM4Y2p+wHPZWrpvzBsQqcxX+0rskZ9U60kNgDq/5ERMbjrJyGRO7fUjT156Fb+1
JdDOrWfBt/fKctQ2ARdET44+ECkX3Z6CbT8yy7i8rv/Gkw+/+xjyJdzsVn/kvtdyACFQjtgaS/5f
sD40KqOy310iDfxVhAvAFj+hcQEQU0KEDhjqPcGEPzTHJBcXinlLyTjRhJLe9BddUf9phKNRipyD
ZA40awMv8yJfIt4IxrL1LseKlfpj0FNf0F/bdpVSOEOeAssIO6Wg9Sjtkntpq7JUDbWGYUHSYw5p
BD+57xrfXScXDJOisp6zkKtr1joxm/ArTI4EbC3Tibe3Jiy/SV69W3EbQFZVEJAn0P8P+Gcezcix
C4B2jodw7uwI5v9VvNpnCzeLOdEX6LbI9G9MNt5xtPCa8Ztx6MxUfPIltdAJkx2fwSrrBv8w2hhS
yKLIoXtV026pbXRqp59nl/dBLUNfZt3AnJU5WHeOb23mPrZH19jSxrizOw20Ccx08xKt/atXFkxr
OJW2I3A5qt7xrhPUAyXxlAKBmIyRPFSJ3kFvLksxhnzhOke1DI8Sg8UbPY69Bc4PwP7ywJsH1q4M
Ydfw6D/8DMOAysmxbm1Tf3eu2AgCpgUvJXmdedxfPWVHuVTkYJWQXuEbBg8T9xycL+lpGWRgFFz4
/2E6PbGwoOjWe6IORrYPrEJko1HxFNtSFPVa8xSRbcTpUCdUDb5VTa9ltNaQvCFhpLhNX/cbqdk4
UXrojJf0RxtaQsRMrJmyJyg4beNsF5ooJ/q5SMxnf5LIjbk20KOjb67+CLjou0+6ynbsO4SolWit
UFr6Q+yp8h0r4bC1+ibRiP+0GbkiMxEJvpWAcyKVmy8ML4z0kpTBNdAIGdArIAAsDCkWB4PCGm6M
QQ2QMkRwvD+LIjeS2j89y2a9CneMPKN3yQFp8H5hZhgoee+uRUoppChn2gQTDjT/Wii/q5H/28xn
9F+uaJ4WdWCZXKmrZBjBNdQb+md/+dL1K12ofWhMSkk26vvjWabDHv6of1dSWh0A4CITtcNFkqOg
pbiT+ezAL6If5OIocugUsjBmy0Leu3LMuWm6ar3DbFoKpmNImTT0wjcD/Z8JUTV0mBxMJzwc3aWj
WVwpfFI9zMIc9RuwG2tLTZhiywcaTRRuT2qvFpp0NH7nUhfnrU6F5513rntRdhLLGmzSYXzzqpGT
xDMAzqB+G0izRkdWCFPz1SQ7H+AfGE3hYB2zt0ZCNryMzP0JZudXmbl4lXloAuYtvAtg1Y6NUhXR
DmOFxzquo8EnMQR5rRPmr1ixCQeeaInGCJLqD3OxDLNCmopvbJ587jcGKOwouLvhYwS+p7Z3wl99
oOOjzcZ0Pmc3OfOLNf7g03WB+4mlsfKZIAjwMZqteRRmrwSPOfjifDjrFYM+1NzaXCLngAyYl654
LZJxNCXbPOYwnfVqBsyNRQS/GUS82MBy9Znqgpiye0IMy3JLwdw26Bl0AH1OdQayqeftXRXkuvsm
CVYSo8X5ZnXnBAiV6FWrYIReZJFrjjQerEddpeZkp2XBW36fwUp3mwBnj0JFpfZoOU4f6M1VyjrO
U2H7MKRjPt21zlytlnV+P9xmUqVpRK83bxV/Sn3eKn9oLt60EkkiJMT4JUe9M37MFRZ2xZrNCO++
onJ/WYHsDI3k0KuqIYAr4u9PeXCb2nMnpq+yAOvmaxzOR7osG8DGbKQ811p6/rUFMgcqPFg9PSVN
EL0MsufbarSHD96+wv9lxzeSftySsE9p+vk2OssjJlb8mMHLSCZ6+zRTEg9SXBdsxfrBg4dFs/Sn
GILXw/WPmVHCnsywSHoIOxWR4gGpPbkUVaCHqwH86us99/QTpG7akSWrDVpPYM1Hxg6gMgdsWNXx
E+2/OTqhPT1jjZMLysObK4P+Q4i2gh9owfO4LFbqRTRm/4Tr/9aZn4Ic0OmaVBQATyWQhic7KlGb
nrQtXdk4F/uKLd+Acb9QB684hEvGhJEl5uJPXJLj1GYOaXAWC0342wNuBjLfCak1Ktz61fgxIIM7
h98844ZWmetRZwM5jGtIROvDyV+/TXsvQN4cysNu3hVp4TpkZayJCNVpwbjDO1nwuuAhfLzCEeom
SShIvQnA3btbEuec2MXa65axngilElN75ttpadxRqTXBWu+03DJAIb+/cm6qLrZ6rTombNoE8KMA
XilNp63w5cw8TcsWzesLyAyasAvzbMnhCemx3PVTWRVow1hR8clbaji3kJyw+eDjRPsHy42kA6sJ
HK9pxtCy3idByuU+BqdlNfctCSCye6tLZPROI7TxVWQoIL00D7+KMBnUXDQ3IKO+SXQ2jF9m+uke
dX5NQqJcWNwoMiS7fVaeTc2rrRZhS42IbFfE0PKw+cYXzSbepIPwJuGeIBv51yjbtY7Hl9+9Mi8j
4ON0JozHk6RAxmZUcGdFJcPlPVlcOZA4VKXnWP2c3vpSjoE1Rc29Xv0r7cWhidpMRYKi2uFIfDuH
asDlIt6SfX+Xhv43ygCFbQKLA1BNZjepcFCj0EIyWR4uSp9O5+SzvayiiotcjBpXj6x2U6RJUFcL
Nulm4k6o6yU8JXLpkF3dGcTfM2M9D+vdFCOgMd8hIc/I3hsgOurKiEM056X43Qu2/YHgLd99amTu
lplp37gRcW3GtUZWHIFk0aQTbPXc+Vw71GF9OgXtik6Epps4fIz907Sr9RHiSD7vPwx+ohxzGmZe
7E3bDjt27+iPjZr3pY0lYcEMEb5qzCoNX6WB9DNd4cob9WRsT/pdfgRuHQ+JGFKUxbRNhRUgKBOz
cGssLNYCIK93OHvAQJBhfJinXg2ZAVtUNypetBQvz9wjQp/Ll7A7wX5RtihKA1vAjWW5gI1sg2NZ
D2mvgyZWXTRo9BCUIIfYmd/BXv8Uytirs82IpOwFjkNAG7qaIfKS/ZSILSE2Eua5PVs0k+ndDSx5
ACSa5OgtXNGlWd1bQmMkopljTL6ML4OAXiLLsLRYISIkZmI9SnmysLRuLNPFW+0+5tafCYYKw9mu
7+nZY7PaCOqTmc6L09amNUXmz7E+aiL2XI/eRDMXF1OPWx9IHSHmw4qkOcUUEMbsWAJ6JmlLt1yD
puQfxyYiDPJnugHUtXqfUZDVZd+7trAeJDDBbRxV45SF9GNbEASlS2xhc+QgcFLp3ltltSE6iDaa
AoCEuCh2SmaqypZlllwV9bH3NtTMD6AnT7WnyM5NrIMsyVil9o59v5DwzB/okSndWbxGeFsevUVH
Jxvn5Xgx/6uLu+WDQA/IpWoA5WhdHvuHtFN6fvcyEF/gA3cXFsJZnPMhcXBIorRhzORXFmWiqs8l
ZRoZF9lvezEnURdpX814CQJZ4o3dt5me5mgk7f/3KtTYCfCjeGIJ+Eu3+Brf0hlmtcYVjexTWsHg
hFlf8j+JuXu9N21NyXwDHIuNpN3JU9y7AQ1w+sFltnMxcwdckfwP/Hdr9NZw9peWo6bjQaTwZeFd
zLia/CmvZ1ydyTgFA9CofEngDCuiszbZhf1iF5XizATmg7LWX8MzScCO+CzwAlb3S6qrUNJ0yme+
hJh2hDI37wan6Q2Ns7VvBXDoseh3gZ+BuuP2cNoaAqdpl/HkM1YhWCAgGJDE0U1u7Gaj641FI127
omOmK1RTu3M6G/R3LqEe5LxIIfMcw3k3EEpBH/aiQW2hNvwtxRW3e86cTdccHE65KIelvA7EQ7TM
bUgBdZLbntu9fFBHQsot1GmksyDZ9ZY+QZ/gwllHb+hU7fwx/1np9U13Ey3wtrdZYyQ9T7dRoynr
cGioCTvly76kqnEL++9IawXDChe9WBuoP746GvoWVTQ1+8nT3KHoBdszSI2x/DfAQNpHJsWpUIYG
h0wrqDR1bGtd3SGdLrhJPbQaFSE36xZaxlSkmilkEhRu4F5T9wQk4RsfvEPvnCHtUVZ/g4ZcMQnP
cT0fnt0nT1yM4cbzVc/Ph0kTmLYbl0k7IubC+qF8RIsEPFA5/HvDYNcQ27yvig1KOSIo8NhM+oPN
U6YKDmcYgFCmk0Uk42CsSaSqwCBXFvOAs9uxBevkNd4L78ihIwABl9yHn294BB5NNdlcxVrwNpt5
9KYZPlV3qLV6KuSzGot63P1e7Q+VJzRNArJwVHGVHy7Flm512gaANv7t8v8VIfyFCBAuYOqhso2N
bxQAw31YaoKkg2zroUl46r2fzz1ulfSqfnWs5BIwSdlw+PM1NULMMk6yEnENc8YWI1FgTL+k3jbD
6Wh1T1eekCqK18wWDTqGnT6DknG0JUXc6ZB0HWr5buPy4AOwqvcscw6YOgE65pW3hnR3RIksFRRu
KB7fZkCQPCSDlcAhipdqm26f+PBon/Rx7I6AMkoOTCzfgIhLh59EueZYcm2oBuLPYO8fN6AaErE5
SPybecVRaZbT2z/5sqO+UqCM1yCBMtmF7vfNQGd2pET1LFbUcURjGnctHckDJYl9TOld2BwZkq0p
CyAAyN2nm+IITDtd0nUVZwyEGHhbAS3kPHrNiDFzojTpFP8i4HF/xmOj28xzJkRa4oco+B/hs1M1
Y1j1wPCoGSAPODFW5sY7n0jA1FdZgpjlS8AVUSY3UIchKo3XZuUxZjzGCj/AG5/0gDIAn01y1yI8
K13BNfzLmBhQKZDe2tnr88OlNaDgGfO1yE/6va8b7kJIEQSV7YFt3O2rBNMsPe8krtIHb1ng7PSi
h/hx0EZJXYhdCzlFuf1SrH2aA2zZdlmtlauuEbiEAq+r759y9B7FXM0Vh8LsAWoFxRtiPTZCgbDz
8xeBcCmVKH+JQFJUwWoJ4Af0OihSZoQtOqB8nyJTQLEeKEiYRCpT0PXMMlb+hmCPB0GQeLpdRvfD
HowtmLvoLg11EfjjvnXbuFbCF4BKTnaZDn2p0UeuMzYbEiEQx8ABm4FY+SgwZ9xsZ1SzTLv4TnOj
cfgbMLCFAtyTL6duM0QoDm2mtkiWT82Da8tOyw2sznjuJ+ah00hBaLId8UBqBTUr1kMU5x3O6Xcj
6uKASZjcj4w5R/OeoihodDDICPX1PxxyfFiQKvdKfgzRykqFKefuIvzStBuTww/AUssC1x8AsIbD
PEBPrzkInlU5gab0KnmJoLBHzcCg7XA13NAC+wkgjdhAWuztlvy4LMhqm/UGD6oN0oTDOrcxLOmL
A6lNZKdTtSZLYjIA6U7YSbCI5DNVn0P7Mmzh1NDvzvVyOG36NvVUEOrQa7a+1QOHbRXdwKnBd/8l
NDXsNG4BhoKlEl7kjJ1jjGRqvdpoZT2sTB4qauL8cnpe3AoPmkQMLN2EChFhqH1Ln4XMAUsuZpoa
tYzoLm342jzrqwzc8b1MvRwSmKTganBQeBXaBoG6Kx+1/3p/b8qusI3t+Li6E16yFRQZuI54o1SE
cSk6OvG6ZYgiKJvIMDby0jRa2CxDMtZ7FbmxiztPElLEboaJ3Ehkjk4DILWgfPNaQ73dnjWy6CPC
Eqy1YTL4R/o1FekoSD8COpjhyHbxUcrwvxcf9SBTLWkmVSh5BR08MhIjJO6f61p7r+LEg9asjxuU
Ptdwcs1RMZbYBRpehmbwxyF/iIaQA+nd5G0ows0+QDKjcZrhlod00RN0iFBHj/2dIQZzTFfyQSKd
bLnDG98FDjDtqVApYLDtm1pS/s08WKaycKPk+giod3utVkRk/EsCHv2cCZelzLnfU+hugecd+y55
n1UmwNQD55NDojy2dLv3cvYISU/Y0JC2U/aHdUOfEVnSL3iEs76Rsf8KPv5/O5rzFBc4gNvSVDHt
WP8WW1kfyxvyarIpwpiKHsV6M8g1u1Ulfxl52wRmjsz1ZJ5xwyKuM9b5KPRxnLDAL221BggHP/8I
3zJ+DSXyJLOsn8SNXT76ltGwMi3JnHJMMv36Zqq/fA605Qs/GcNIEDAFjwRKkMGt7on3enm1U4/y
vJYfsm2tlcpB864KazX+3Y1ifd5+2m9P2S6mV99HGfar7aq1d675XM+GKZTbQrMqghTM76fRE9XO
LSAk41mQy9hxWxcj5YV3x0cfssooyhtBvpQIPLwzxm9AR/MSjbiGFDSCHCz4FxVszpvnjHNsRVw/
y2+UD+T/n1ELkxT8jZ7d9VqXQfywflfiKf9aWDPrdbq25rdA4ULGmjCKScvqQZkjLMtKSYS+p/6d
ORPv4EiDEM7cTRKlvO2VFToizDn9dHD0TrMc9tze/0WfEyCLyeAlmqjG3EY5TkblaEoZ3M2s266i
v/HJoS5mW26EGbXKPb+5LTh/cjb5ERFqaSFlntEdYWX/D9tcx/RNcefNKLq2T+Tk6XH2NgvPQfqq
2sRmeDLcEioZsLwUDdvSLdt0LK56vGP54By9HMMkFG8c3BYBuITWr+iJU17dA8gCYXhsudCYpEP2
E11xqja6BpQcV7KmVO7q1HpTV8IcAlG49m0FLiEZyY+5VebHPuY7pzee8cj4QMJLd8HVI5tMbOGY
6gZZGSAbRUsKkKfpshcPvijkn8yJHzfxCNj8Nial0kFa/SUKefTNf95jUJOi8IVspoMD9WkoIpdX
9s5KJXbFUM684MhRtp06b4ZPKH79k0UkCZNPOgS2d80pmxeob6haK6skI75vXz+h6wDSSuoqWDz9
+ZE1qOh415v8JCRqXxnLr/nlEINqOdtYy6EIInLHhLBc3ii/eX9klz4zTRYkEmi/s+PMj9Ljsc0D
EBDp7p84WYLrKmiquR1LVUsn0D3Mf4aOWIkp0Z+v1Vcj79HdCcjleAARBe4kOBslaFJjtqL1Asr1
nvfGofReAommEEhuzIfd9lfFZitm4XgQEGDNLVu/78YukL0h9838UF4iixYbyHlXfC7PHLnCNSWc
tjCTT5kJDW1mDZyacDaVGP6G4uNlyYg76jbhN3YUbyR8ECXcAXgCO1cNlCUB9wzA5RRtPjtyenD1
85y9Ix+W+iySRkpwjTQgXChC5q9DYqxNtVR7INnwpCMfOlyo4byzZs/tCiFQw2VT+R/kTofGf7+Z
SCZuqOJOW/oer72W8pH2oKBTe0mghvKGf94pLmeHhiwjusKtXsFbfeMC+m7pjR5/ge6hduv1y+Ft
VXpVgcMddg/eibg2dk78o9iw2zL0PcrfaoNnzr54t99IumVnvYef1WceUxnNipF6LYoXwwBOLceW
fOEFru0T5ELF1Ack+z2nT4BOBvhNMha/tUdTfaH9pgACAsrEWdLJDIHi6kpQCIeY3oW+vkJNJPXX
LJP5iZVn0VUzcyHF4gTUq80KnnlKFnXUzI4JeSQcnV2/QRUIAhsHANUZw/SbSBAEDORabAPBfWYd
uGH5y4EOCcHTB9AfDcHtaEQqS7XOf78Qx26zseKlVBI8+aDWLe9oWj7kxqcfxZDtlXdPbVd++pbk
TIBcmdi3bKtzmWWV1ZIAlGKSQX2agal9xDk+IrIL9izKbsZB2D5tYkaUx3iOtkS8fB3E9PMNnznW
idK/uRSGQ6dIJUCz/ClMX8yFQm+fUrMBZxyMogWl2F9YiJTM/bewgCqcVAyLgUZ3f7AOZrV7Mif0
fCUbdwHW5hXwzK1x2aRomAdPmVTzZG83hJ6bxznSVUuOOV1zLtZG+7tu3jzOVle1lxrBcZY/tuiR
G+SPC9OSMEgwpPwcNRvAd38tA97shC6FI/rqJ5NSeSNXkGww/2lVXvrrwhIu6vIkazXeciW7IHy7
EmCtIyP9XMWaCkqHAObw0crLmlx82nqeUboCrdaJysygW5YqnSVEDkJcRUkI8kvI75eEWxFSKLgr
aZUwKj7kL8qQObOXlXu9WR/cP/S4CS9ptQkBEZHlnFMPfHMQmcfoVO4y3s1SszeyjYk+vLxdHgeV
nXVZAsY+S/fiGIvr8lO7sBWMzdC1v1xSZd4UHk0z5pjSRY1s2uP5Cu3JAUeC4mvenG3x7xRlkk6w
A0ssQMkSOLBwvLUTuk6UPnMvK2VlzUmuqpvKapo9vpYVzRVLP25ZMOoYEOUWu6xKUQUf8jNRUcs8
8ecMJsfIxKm6J0HSIMW89MqdHAGXPdsMo50iqhgKGqirVWWV2pwkw9biIzRBDTPD0khcG8h2ZXHo
xKOUtbXbzuwO/e3UtqLhdK8GzP7cdxmnq1Gh7VZD8vCEtQC829yV0nNqWhin1mPGXwy20Y2vOBfu
o466m0GgvdsO2Uk7YS22VMxnATNr/1FffULYqXRKLK2pdblElEXAA5mCpWxViMwNe/Lg6/Xx4zxn
vcujIu+jErxonn+oZeIYvtLfyicMqKpl/aBLe/ZtYsOgxwB6KAvSBdgMIAD4wbzGkQloMfxZwU7k
VGxXW7bYjbaqZf0ktCEkv6+nKIbCJUs8ZYtm9rPbNPOgcZ0hP6AsJw/E06F9eRc08RFbWoaV5p7B
B1iGEgiOLCclxopXXUyDsgWXGoRbzeGW8FYWKiQfoCiS1GdvF9yivRIBt+igslhToetlpb4AC/b4
6vcPtdlgzdbqGC85woEZgueFNthUIvsxd/wT7bg4OfCOcGm3j1kNJzTdewl/tC95Ua6bBb2Vdt1a
+DsAG1RQ2Ue++J0XKfBrPKAJBQT2G4/x2XqQ886QuMquToVklX82afKel3Y48xRNwWrGe9fRnYib
k2ONZQuE9l2/8hkg8pCj8rVVzf+/nBPbKml3E81E2EwqdgYi58a9Efqbx42+su+7WDvPChLkUS3S
l8xPGLXRZUtn7NQOOhTHfDe1GJleN5kHm7R7Tpjiw72XtQvNwRG2QBZWPjKCtIPbfOUoYS5vK+RC
FfWLM3RSbiYKt3WCsnkSPVUsZCt/V1tK8/cAVzd8B9uI4soDOnZeahJ44I27xFZxmSHiFawGcJtW
voX4WuC+R9qAbFjU50unKkcwcX14UGB7WWcpFAPQ64rZjxh+nc2nGedRi9iNQRU5oEQ1G3ZCUadl
2+EAplg0U4Uqxu0Agp+w0H2lpCHlGJrYArYuKSchSDnv6/AYdQkIh3ryllf3p9mZccRZdtN8dfTp
IwJc1x30bVYNhSZkKUI3ZWGlN5wqCFZ1N8KEUYOau/TVz5v/iIbbjB/mwO4EBXvjTwKU1q/b2284
goDBkMY2DzulsTsUnVASjnolLMSic/iCXGnWG39sqEm0dbuYUkffariH1vV9GaTwLbE0L3FJnHgG
BB6nV4AMcKSQ2Gq1bg3yEizmdJuXS/cO/Uw5C9oHprLeLar+2taUrzdCc3V8nK308JiPr4fjQT+9
+uCkJL+vqsqhgn91eI4RB+pXkiw1mAj7O7bUlsKLsT77SX3Hx4uHwOR+DQOVogPQnNiJRKU2ap0d
2NmRJGr5lpBpt3xWly3WsAf1b/RvvkemQNBHJQ/IXVscZssmACtogtj0o69baFxqnPFYUq43Ho1N
/Zk+hEG10f6IL7a6bNJogqgmXHc4qjmg2qMcXl2XDkbdw5x2MKQO8LTmpQrXPCpRNwRCD34H9t+M
fDArfDlDrbND7sDKFAm3+V1DqWQaYi6d2yNLqBk3S5JBq4PalXWB3ztGDA+iQhA61iP+lPH8wuFx
GmX991UICxR9dLUFhfOnDRjVDS/5IX5piB8452FhTzut1r8bhe+R9c0UXx41mto80/QBQkLZ+Mio
CXKiXDxmI9j77Cbz9D68D8VwmAnZiMGCW3EANXSLtrb3XoBTast2Vv8eAyQx2YFChw4c3j4LSBAX
9Rylr/Ss46yt/u94/X9O/kt3dPt+0G7Cen0iyoYaOdPde8BaZppkMlk34+FxhZPoF8nzqG8wyJjU
uSlsvjqsRznqnmoHEdSQLlFZv0jrjmlFyDxGlPb0rJ5+4IxdWkmy8x33bC6wADkmpURYtydd2MPh
M+EX6R+k+G4pfWX0d9r5iqRWYipG7mn2eCtoqAGlK4GkzMmZUHEEs4ehYzedjB8GsmAtR2iByTuS
GSiP1eX3Lnd6URl8Q1SoCZIgHc4nfhIYO502IAnT7hKhp5NPFwfvZ46D8WLd/+kTmaGSX4nKJ64n
sBKqk0P8rdoG8MQOvihpH/m26yvTFWyvXtJ/8KzV0I1RYMrcGE4cKTrMCK/mdybKwKoisgdRV/1I
14vSToP+w5Tw5Oqr3Fk45f9BXKbpvRXipCQFr6wXPDowafIjPF+4L847h7GwmC/wV78BgnYhKdUT
ExFiqNjFiuWI8lgs3aCWtvCo4/slFOZIxgLCTdXBw5OM24QjOOmVveGriUtPI1dGHWzQQvwfADNt
d4ObpyhQJNgIyG58Yry3afNsLW6gtMkCljFx2qq5FXRihZ5xRf7L2QPwszb+mpe0hVGsiYstAiHL
WkoDu4J1DqmgbvYSN0jtBiiVErniLUEROOzABkrw6eqqHOSMw0skrubWa8P1YfzCyegZHjKI9XGk
HuHuKLYasF+sWIpNoLhGijkozjo6YYzuuDtt4Nv725Em14bHRmD/lFGP6CzIvjQff8CGi/MEpOVU
e4OVZmbNQkiS8zrs8RCZr8TMgcMQY7TEvnz30PMiPlXQ2jR+pg946ePZHrSq5Io/D71Z8lG5FkjR
5PaIaEXKYM43ZobhIyxJIIxo3rsSbTtmybZHFyP20Knf5OTAJDPycXNDpSGlvMsT0ebzalACaCpQ
Pb76ntjUNkiyJGlY9bgGoO8D1iXgIqxOEQKnQohiBXC/rUOKVk4Xt0G4YYVewEN7cRRubc5tlSs3
PAHPGVJRSB26Lu9V7tjWotCI1F1Xc5z99YPiHqRh41G1xJpPEoZomlTwnbYZVoMpkApk4pux0qit
rXYgMaSlZUXG4zsE8x7wG1m6TVQC7ePTXr7sKMQC/dJMH21RbIEk45lZrHAXaMli4HI4VeJpbbsG
oDAc1PZTuXJO7Q73vyC+Bc4dzSBLW4f419DqU8UdOx3RR63iD/AdddUhT+QQShUNZVwxLUcMDgBi
+YfZD023WdVYFlUDdopZz5+NtX6z95RACeCPBoYqUp8IEuLIzt31+qYDppAfDW+fpg526AFKLLus
Ad3RLNt/wb5QOMrWVM0teZ8HrdXaTxWzP56/ReXInxqzm0QHtR17/RjmX29zWOXya1lnos4m+Ib/
Qbwma1xq0SLA+fS88BdxjoncqCBdbLPPuH+hhLjCk09xlXKo6CCvyidNHm1+UZiAWWu4OmT2lOfF
g5VQhTPQmlqJboHkABgAUpMGA8QjYcVoGoG4jfF5nxRp3AwVQCYYyz1lxQr0oAy1RA4bFbtnLB7T
QUWnMJ1q4toLXaU7phslhPWo9zW/afnYZ1xUD6CfJU1KwUao6RMgFjb7n/mbMkvmXPVqiEZxnfK7
y3sRk5IdRSYbjE5V2t/6/I4A8Ayn4Lf9yUqndeIfBR/UCUGp0wt4AUWH4PN9WMF9MwUK0JI7WUHA
GfIn5Q9K/+F0SBSXnF8kwK97KCt148RSF1i3bvQtrCtPJJV7ayArEG3op3YamQ9FgQ1l1Wbtnghg
O2ft6MM6MBrTKkUAXepA4zLzhwX0JeXZqWWzUflGMr/HqTIsO2ZiJuQWhcFm+gd0M567/UxFjCEf
8epk5JZJh6Y7hGEW/ek6rDndLs+Ms9T+cBpslFUB1tRgxnhRLWvX0mE6W8mvCl63BlQnXuX2XH/Q
R82RmS3a/AoAe4X1YzQ0LfpeO9E19F+A/NlMSiTTkU4K86oJN/SiS8ISAsXMAYmWbFgsAJRs9pOn
b+8C/P0MTpU9fMaveghgNgz0SEwkjsRxzUC/7RKcop2E9Au0rfMxc4Pdfcl/dH75TGP61b81KPw5
o+Rz4rxPjIi+xo90Ls6d8B9H1v533xE8hVXHahU4tpvOnMYlK9vgzeSoyIbzn1C2TaiIrCqk+TTu
t6X67h2TJcLcx0A66+DRrqHusOxjFHCMGCeyert4BZyv3JcUzpZaFfa114ANQm/CMzA2s2I4WlLa
oAAUbS8Yo9/pqFYU25B4A6XNXYrJN46tfDmEDyufGMzYAU0UiimXV4bkhZ36b0E7StMtk9WEMtUq
WXSv0J0c2jpZ/xshyjh0GxEjB472WVb1whzp1viLxcMt+A2Yc1AIdTCsSf8eXWG0xHIVkUp47dE8
pYXVev4ldIMuSd8cl48Vdw3N+d9WJ4/BryRJ4BPzBFd8BKqgWux78kcJ7DUYSyHwvc5Xt7OZxmMm
uXgP73Il4ZgRH+vNqktAUk+qUfbd0EVx8fc0iVBQ4DxI3LpuvhIXrRpdPUBEMc5+R+IASMmjBWfJ
/Z+Seh/uTJW04jIDrw/v8xVtRoBw4QcVp9LMTlN/gXw0K/fuQ4CHpixCKloPj/9+W9Ysj2mCNzzN
TaQeS9783c8u81RgM/mspu7jAdvQbzq42H/r+F91UW5UxcRNeXRJG8hv6PbcXGo16TvCGiAy5yHd
Mewu0+CdqMENyep1quveVs6L9SXVtv72WDbcxhzImYxPLCA5WCTLF1LK8tB5b2HPHg/oMowo78uK
40RiDqejIfjo0SelT0rmexVeeI3joolJ2Zm5pHuraXAFOHbLwBwNdWVqqKUqvm4kHCDKvTi9jV5T
rv1c/sQqN22u+lVn6/VdX0+Fp5hI+g3uJqKtGu/Q2stZIfm0hn0NHk8+/S4d/YZiuXnsxvr0KRDC
xE3V2hTl1v8tyv4bfhJVm19xXmw8D1q9D+URU27CqAIUy4TyWxs4/9HbNR1HgC3zU0Pt/vZy2JTV
KyQJXClsk/xNhoZe2xRDu75YkXLe0HQCiE/VrZwwIfbGV9tPtHZOebuxHx9gx/axrGurnw5Qh0Vh
4YkzKv36Fq+MO7N9eLrsCMi0SrABqwlhurHWVYhvhAVZz+X5giAr/ONi15fp8ICdovtIH3fowhP6
BlAaNDYcCyaN3D7voM96TLaAWRGc0zwyjzMQXYYQAy6vzd97Pdl/uEAkOFPmxAipTGlstVKrzhDC
EFroE6zCx9NwRyXqy383fukq1clqVdtYVEQoKm4Mbf/TJaPUdtwYJGBfPeSF0F9So+S5+/iJTzp0
zQrnwtG2ZCKs0EJvbWVCNIkTFaPsYuSWjlVyHfO0eG1CVTLbynlNym9M1J0TFtmK1Vq07/fJzDp/
RXe9ZMN0Df7CYLeWzLH26nGjc6CEztdTWsD6i6zSrInJEG9X9pKvZsovgkZNmiymAKuMuukPZIVs
4d+2qngPquYD6Czyszy8krEYVHmkLIksVL3F08uLcnKi26mosM4W4vANa8PHpX/A50M4EUXmYTBg
3gFcPz6PVFZbWm/kmXlD32YNsrjkp/8dZaiGVD8gsgHX0RQsNLfv35Lgmm8Rj+rTnGsfYLWqG38G
f+2pBgZ3JkFecLqK9HYGtQQ6d+5a/ikaconPS6re0SpMUQXN4beiChN2nAS8pD8TZRbig7IKf27Z
qWHpb4rWfhHSiTGn+yV8WTYiOel2AYmGWOx0e6vrGsJELr8+DajKLLoD7ocVzSDCMtZEReMsNF+n
xNh9zAm0PT60FWbcO9uV93PRtM0pC9ZEthU32s7Uwlv+AIfta5ln8cBsJfkcg1rZ6Emb+rxDoPJR
pPzBTuoTjFP62cp4w10qg77kLgZXSMBtL7hJoHEt5tkdMSw0znWG5z5N3MBg7W9v9d2FRNavs+gE
c7ihNqzafx7UfqYrwXnZ2wkLc8K7YrcWotnSuyq+fgEU8YI0ON/daTj1lsJlUZ6hiuyXeIJFybfQ
az26fulmPnAhBVm8Sd1AlE+s9nVySoMpXwA77bNjOVbNIqMLAwYjnNCcPah8fIJE5+KeEYptWbkY
wvqi9eEMbWIdtFlYlz7FuY61kMe0n2BzpooQcCNsTdF+cmNItjMjhUisC7IzmxhjNVJdE9NJObV+
wihXSQ7bqBvvtZw6Nsyn5Gd6rgbb9ZuGQtmOoyXclXuS3ECffElfjMgIM66C4vh/ZTfF+ETur63W
r9j/T7SOTh/KbwRIihv0OJ0Su+vjl8803BHDCQ8+0fnR9bhl67juGB8uZtbcLyXCS2V34ugH5L8X
HHn9EdJFV3lzcn4dhl3wtEJcn7WCMmdnjaA9KblQOGKtYSfl8GcqpAFBg1WZ0/tFZql/bAhTY2U6
MRnxojGpvCqTXU6vPKK8GUmWYsMFoj4EcDzfz9IFfTO+ZxgbDH9HIPdiFmO+uk/Ox3yMjdax3GA3
fypv4uohxo6wlH1F9lvM2j5+pRbz77p53eOubsoOdxTKanhjd2Nt4ysMwRiKfe07LfXUBPFLgylG
XyJpSgrY8AwLth5WCIbeNzVMAPQjA5+Fw9Yf01nIqBRTRS2721YLiVl0ITIIPGKIfmc1l5yeyKU4
0wdaGZwIVoHzf5rQ/YKSTBOO84wd1+OeGyhXDIdXIHy8xZR5GVe8LgeiWdLZK2SmWNOY7Uc1ANmp
y4VyP6DBtsGntQeMQvbKGSFZeXb/NYnMIDpX505GPveBBIaFU6Mboo3qc9s7zJLMPMyf6H/+FWnG
/Zh1n6xUCSK/BppUDjmi72Z+9Twkeb+zZNxMGJ0VJvOVOxnym7lmrO/c8qbIP3fbOhYazZOxrS3x
OAZDXNFOriY+YugGqlh70HfyLanhtr45vN5ecU5VeGUNtJPx5q3gwxWiC9xN5oPchCY9jcTDEXyl
e9jPl+jWQ8zdoBCb+6kF8pyDYvacNUH/6f3J1908UjIRznWxktcWBrvt95W0BdKmReK/dpMVoBbf
PxFcRob6Cea8FlV2uH4gxykIPsb67tY4ZklWVKsqWu657xiA5hA++FgfyrTv/JII+W9Ozfiym/eE
rMTM9njlyz21RuQbv/XIT7tu1J9bCTdS+9onFlawyKT9J7KTMpE7C6kKYdQlHryLhfcRbBj4DxVD
tjw/5poGJF7jPaPSMv/TnkKnLFwTf8Fly4Lpf/pXB/TfKGa+bgCY250LplJjRtrQq0Klmnn3Q3WV
LoUTh/Vrzbr3EbGIidHyxM94n5nePQ6QZIwKacU0f7DGZgr6zLlHMxsD0DG8he6Or0M+mIRNnmDV
q1dizyMAGc6KcOZf9dCxND7WWQHqfT2g0blb1eD6/uqRjHJzoKnqqHzCFMn5cecLIhgohtpiVfts
otSPYRBJBUSMsUg16kU7gVmbF1PRHPmt/Mq6kc4saIqPYQr03eN6PksEyo62PAJPrAYTv2z11hci
qW+IcnjJX7a+GJAKWS/1IqQA+qOzb/jxd0Nd3kWn0ZHnC0KNUAwD0qx9sqQt0AlE+kZ7KOOYRxma
AoJTnOLNGlyabdhSnbj7KGrk6A4Nx65KS8LuPJFHZrvl9OTl+UkhoEhW0R/DExvBMMpbL6uQOhhx
KYJG9YH6twxZZaV4Bj0daTXNPOGgtHPmkjXE/IY+45zD0TUMe4HWG0F4TnhuJ+Zw7V2+3lbtbp+x
csoTBXJFcu3hFi5IEziltaoD+Krzti/o8wIvl/ObJoyAY69eXPP9vv+gRhb/RjeEgTaWm6NALrpi
Ns2BybHmKQfiU1XxBPUfaSUd8g3nozx20l44N3WPCwUx1VjL42oUIvlEivprddgMC38Q8gZrOsob
wS3CnBs99yUacBvOooTLsRed3kbcgt+rtxuAOFyr5ZkbJi8QMYEU2qMo+bj5hhQWQ49Dvi/7y2G9
s1UD3vCVBp5a7en8qUyr+9t2XEwPFCVLnWxODTiJjtinowlgTp6YpWKM+XdG4l2v9/IZfrj7bB0D
BKX+VSRZUOSBdWYTsYYZe4pUnewZhE6XH5qb3Bl1Is65SfAbXaj/3klPjlL+0NmGFRaFhWHqhB/G
yQbMLs5CgRP7KpkRXQ/4CC1y4M2be+m4/h5IN2FlYFNmWm6sbwismnIJaYlw0nkQWv0Gquj/sfA6
bzlTYHcExLJrRaXH0EEr2QbgJkecyZH9QclYyy1J/PqSjoB0LnPyp8NLXdX8fq3CjWhIOLIE75wf
msjbwpAIsPVyAfHCgatOWcIchq4zSEYE6aS14xm8+iu2O8TyMGFG6W3p5PRhBasses8yWEJ3y0zI
yWL/fH+0WOEJ9NYqX2tehJRETpJIAepomBRyzgrdQvPgm4JYg7X4EBHaXB3hZ+77meII0qfIPppg
fNuZTFntsyi0BgldSbzYixuwtgl8+yhqxLUEnOnd0aSZitRALonesEDYZqK9WD1SN541ppT8AIVA
sHk8TmQewHcqh5ZAYGQMHyjXRd6l+kpMnKQXrFzrY3mRMReK/7OV3Kz2tgrBPa0+D9/XlI1UneUG
oS53OSThY6hNqaNI+zCLH+23od1q9zTJ1JOlJXrlSLc03ua5B+jLaMXvyxm3yZaR3imcu0T2nKp3
RJqgEHeNCNu2dEBunCyfpg+Xju6dMc/fqujEHgivGXwPmfAoGTFuQYx5KVBNCCnJT0y3fi2VLcEA
d11q5hTV0Hwmwpw7ABeQnAKVFdU6xwPVh1W5lWXC+5fh6pkLs2TRm8v+Y/O/eWH4DFcrYZZb2vBg
IkvcB0lqEpIbQ2S3mGXQGXjIrV9YghvR7k/ARVYnGRiPcyAbeezY0ocFhFT81VKSQvF146CmZVi+
LkKHPgWlOisOjHre8mtjwbAtGQAwBtY7oMmXODYUQj+gocEVXw27Qid8yPwU1j3J9IlWAwfYovqi
v+oZu8cEukPNwlrzI57SRX4cY1lhPvdWRZk3BKg6YCnNJMX+89oMXBERbW6WtA/xZ6VM4xvhkKur
sr3zDJFv5VstJsTuWx+czLHtfY+rzvsv93A0japQqfSfGxcUncIwr283EmXqQ7bKh2c0fcXz8nxO
VVVW8yiYirs6atBd81aI6b8GPCIZLlAiOC6nnHiYTmSNXJMfo3WKglaTUqKqlCnXo2fN1ClVNSTg
/AwgUA4NAk+pf4kb/gvxqytysfNLafdCP38ZHATXhYC/j8XTNNxnrvBxN6zhl/MmsbRlm0wv+FhP
/R2lZ7ptBuZMiXqfk3HHSuEWCK5BRniiijEkpp9JcrN7OSsAUYKWo0rZpApE429Yf8LiBxwaJg2s
/V3j6wN1RBEwd0UOV4O1ZVXF7/qIeS+cRLyYkiQtLJ8wFT07JfxqcN7fbsYOgfS3rNP0smIkke/H
HJOlITPKHnAboL2v0dOOoclAuMDm9RuVzjqOWcoyrXGhuGqgLb1mXf9K6BhzNtM7u/VnohXHUSio
0njcJ9k/7D2gzpnZpZgWr10zOcsP/XOSkUg9cFQ7m01zoVf7a/gAN2eXt4DmfNKAfHfsV+kGe5Z3
mouxW0myJtlN6JCVq4gLXJFPWHHwh7O3+vNGhF/3TogYz6g/2eE6NsCc9aOSwE+JW2rQ2XlmS8hg
mtWSm3fzRGE1OBS4dRWtsirKsK6kANj5go4UiQ6q6eQqOAzQ8PZNCHtHziCYDzPgOo2H0iNuL4mR
PBuY4avwpHBdY+cI3WZ5eLj+6It2ci87Kj0PbCr4v2w/h8A82YVcLpwwOUXarigWj/o23nKnutgS
sB+kU7iPMbGz19NCHVertqyA2Q9bT7NTRZCuiz0wkMcIrhwfyJuA/5QnRAhMnyUgNWv6A2ceBcXK
z3GnsPC+bWonP2UXpm0heiR3ubuFmjJLqvAPNn7MPYyXmPdkFLuAStP5TXWmNA7TD/WajgQ1sYuF
UoWViqyG4tJWzPFOBug45JnOf0VISgs/B9aSyX1MxbmY8hr+z1MEbMdbpWScA3OB3/NiWMJpHZIz
VL3zu/afHFC0POjzH+YT+1/7VkscUXi5M00zDVdSv/z4hQPD4OdWGh697+iBWBJrqvMJFIyGH9Yi
Ett/GZHJEolOnAJD9SMhhqiD/eC9PeunI0UFPXeCBCsSrkfLLSB+6EzhXHhaNoa4CAq37rKD6jij
5BPXjaRcMoaGHArMx1hnZwPrl/sLx3tBS+TZKt2AU9+su5uY04FagdC+hfgQcZ0REvy7R7oxebQ8
evfwBx4PYkdQ4q7bnovIt8NcG1qb+dKh6pgsnelgRo+w0E9qSD7x6O5PFdZB6CatUi/MlGvgyEcX
ITl87rOn9WGSeCNOy7eEqRv6VEQZn+icb+gl6oRrsWXGcF3XOWFou5Ld4ohvhWF+jzdlME9ujm9F
ecqvm6CE5f8SIpTVjrVR5n6fdkd3Qrk3+/SFJlQh2aA4vCpXSpS48GnvdLRnvX+Eohuu/0YfMwWE
G6Sqjt/K42575a1qXbQPQnZf3ItDdk5exgnkZUU2Km5T/b4pZnywGGPvpa9/M1XvVW9PP4g3GIBe
mSd9QTaLZubpCRSjkEwAn+NqwZf/IxWy7mouyOlJ4o3U/csWCFshlLVPcYZlolBKe26GBNT/hNTY
c5VNhHRDpKGJs6+xm/iSFSyTy6sQnazya/p6F7CG0HPXgS1GUp7FX5wE84E0s+m3884aJJbOYaYu
R82asfTt8B1cl3UPeHXnACtCF5AAmZTwuJyYt2c1JChAh6kFzNodC7H1MaPgvDkIgusHTpXM9xe+
3ZZ1c/kEw760SPfA7dc/D7vhu0RqbQzlOL9oPbnBpFtInJUYpNxqo7k/3n5PAFbebI05wtY2cV5c
hSsQJ9gj2xVr6O7AgMxCUwm+ygojuTRbS6Cc0VEWqFmA0M/prKxSFBgKzuMLOTdb+/CTS0E5cRwz
SU+gMgUubJm1P3rOlYNQzH0J7F6XeiLPR76IKQBH4DlaVwQnOi1orKPWTYLp2vXrMMVrWrq4E+gO
gjo/twb+WeBbRhH56v39/KCDlKdXeWqGwnci+X3O1aDBffymm/WVXMcY8fjnEXqtdebxMyf4HNzU
cibvyForTlV1/44Le716e27qNDGNWKBQH1JK+g6E4tPY0a2AB4C91goGXFowYti1OYfXR7DHOpAD
fv76pDncxvUiREo62lIhouVKGiruECMHf3vSJA8kHKxifAPotgHH9EwOJFPzkNnIul9NDBwAwo+Y
qSBUBl9B8avnm6alvn6N7zwWBVwHwaTEjlcS1uEknCwLvDZrpKVO9spSyBytOttKneke7iPJYvhF
vavifox4RMXChUX6N/LjI0M7Qmee1hrefJDxgo9K5vpVbNyeQutWbXuzj8pWjxdRVF+Hx6LbvQ7J
3xwvQQcXLz/8iZ2js/XPO40eVsHlcGuFKM8FebRGn90oCs08D80G2TjT7Ny0xdWFbRX7n7oybIch
z5rcSoRGB9/Bu7H2Y8DuXWS1KsJS+LkBzx7ZxzPYb3Y4PvyD9V/nzDWDE+xcekm5Yzg5AA4/b1BN
PGAIoYXUvMWy0RD3PAB/3Ke/+CGuMlNDOKeRVSWC33uyR9TYZSLvivmCwXViDqUl2iMSWobfU6Ix
IvxJD+GVHMnRUgVgdJB6KNTc8dQO8kvKaVv3ET5wwinLDYrxmzTKA8YLaKEsYYTOCTc64wOfRaK8
iEVhsIwnoH43DeRfaSSbhF1tYZh7PaeHRXDi2EPqSc6BUnOY5O8P66fvtFwv+2wucW26UgSyg6N0
EOcemx8LibyGfnvA9XnFZoRFBlcNB7VxfhKz87IJGgZ7P3scGJBxQLWYqJBEikJoGTl1+ey7hpeF
oR/ot+1DDDKAXgkdgc+K5CsKSt+4BxVkVWxB8wH3NAWlx9z+ynnBmL4jlBetMyc7ZZtYOwVza8k6
hXBa6CqRblrukj2tVq+DKPj/1uaPvhgebVglABn6V9PLkeMFnYlNvAClJad7wDQjMoNnnTECxRNN
tBv1KYYtgY5b1MGJokImikKPrqB2892WsfqYR20lZtldsUm5T15vyq0av/3JvG0qv7P8QMquiEar
Jl7GKv8qlhOLLvS0neKsK7jiFmB42CIpBeMLq4cZpYLPHKWD996GpJWsMvkYU+yYJJ2erl7SokRo
8gQ4IJ/Fwyl0IFal/VUj3nL68pbg0HxUmhtkgEbgRgWXy2gtd/wTKp0wAZ0oeevnJ5Gbaqj6cCrz
9zbsW4tHCdAjPKbuY/eYHOJxXrjaNNp8/um0ImHLKXvraAEkL1zPtDGBVKoMeivY5AauGDvQ7Eum
lEbK4y8VlxKYHTh/0I4PzBoLwUlT8jplhamTbxc0QKTPjNbMtzrA+f3IyY3h6r6GwOGS/mvsvJOB
60X7KeNcMGrNbkI9+c7j2ihwdQcj/N0IPE40RwNmmrbsG3JrMG/uvBqxZCpeL7IORzHLk+0a2unM
HLk/NDXADAxT+4Tqr0DO4Y9sQvWKw9x+Bp3WiJBMLIGHeiUFBmhYNw7N+cYcsgm+3HDsIqcBt8lM
K7UMt1RgmQKtR1W1UfEyvjb+WcE55L0sofCb2AVmVHQg00ECRXq+mn7nOR39w9M3NWpU8hNY1Ik1
qwhc6wg/yVvGYP/a8qv41QlKuoIM9CCRPpxQLYTX5GB6RRTVzJ4Q5PG31DK3+ZcwoRgKf5311uLs
7DwgTO2pLNU27xuWgPQ+CM8YZlQiA3lFwoTJY7isYT0M9fnuzx3fpTH1BGxfg1bxjOGRNL3kCXwh
UR+L1NhBLlgFOZ3ZVl5j56Jqs7wpymMViw1L9VPfgo52V+DPgrJMIBqTQRYHmYOkvYc0UVuXatnZ
FVh99ripWrtBetJAB1vxjrYXC0bmJQksSqj30/OR9UysexJnvSs8cywxR08e66oaWcrNfH8L71HM
Ya+Wx7Wu/uWbjZ33Vcy5eU7lDJ0zy2G5wu3PL5AN6Qcx6ChJH0kNRBdXLfuC5dFXm3YFyl1YXzmV
d8HzJ92Riewz0egOcflsGH/gLKX39rvYTl0nvtY6R43BWrmQQYOVqXdlY4lBE37jJ6cCOBkH0b7n
qpIZGlzJXyjVcz9n7/qpcBlOnnO18qn66EBnEoFs01my2vWHybFpUakEPXd68akpitziUoAsNihK
isRjXSNQSRSYXXqWYTCEDLhymjf/c0ZlUbjjWGuv7gDx4VWwiYNZgJYb6Fp3U5RpgxS70doS6TMI
8VYrrbbSOz9CWuf9Vy7p6zpSJDnannIm3LYZ7tINgBMbdg0nIJ5kBG02TpVcCfsp9RV7J1I5Ug0U
mB7tcM84rF5t3s9zx3E4i7AnUyoKo+uahwDAw+/liip+fzzOkZm0QGowlcEEzwn65belWB6SVAPj
RyGSSbxyhMDag4tXSb1riZgmzhju9kEKF0XEfgHnrhjFHuKDCfXkNAiVsdCWDkgEpddMoEiICc8C
6qV7bdaTd1wK8ODsqjKYgI5Kt/FADdIIBo9+BnBgVKUqPSU5wQFbKSb5Bw6k1mWidX4sJP9jQ//O
xdCivIKuNh8pZ6nvzVqakZ/t9yNfhk0ST1QFLoxbTf4+139T2GgLTREm3v/kY2Ej6it9NWB1ZhtD
slZkPN5MdSw+8v1xPm6GvU2yyzfAELCOvwXwizMTwfnxyDnp89gh0KzYsFmeY6jLYNZpSzwdvSju
s0DKON4CCnS4HZ2njzEHhNpNv5EqWJCsS4d/UrJf0JyjIcFThVt+qy07vRhLDw/FFXCECf6Vt4IH
qNNO32VFzdwM4cPbuz+bOPBO0pjNc4a0JAmeRnr2COX+aKHehLeas0GhFl7RIlOI+hG6gPLa0JCj
1XV0JA8j7jLKOudT1XN17fKfqxN91SW4LOLKIocZwdgwNmbEXKU/CkB8pUvDiFbmcYuKxM0fzdnz
zne0UQvR1VCc87hF9eOztcTDoDfUI5CVss8Io/g4rwNjUzuzF8sEGsox9DCvhnNaBpAfl5/N5dOF
zlvaa5XqiRkKLYMFUXdgloEkwZCkxMC2Wbi8es1LTpSfguzTv0Es8Mch7xe35RZ71/aBdcmiJ+o+
FJrOiyimpdEKAL5h+mimTf1dRczVlHaMFqfkNP49k59izQ60X7o6anoUJsaJ/KYX7gSUCpruZIR9
iSGPwPTs1nvWaZj9TTw9GY3GToeif05rRTeHkBENebNLSsNyB5CDQvjhCW9QKcf68HsZZonyIIrt
MuZxYPKTJRY0pK7D6V34q/WjnwgpAA4c7UWFJ5rZW8789wWhIdvmOxhfDF4cmWYSVGX6z3b323ST
ohgG7+mAAjBHo/FJpU1JHcDHtT3yfCz/KjADd0nCKA0aSsVuA/WOMdFKlMAvYHOD1h26a08BwesW
kLIBcl2cpha/7z9ouamVnluasOA5rAsY/wCf8g9rjgEyDxK5aSiAsFDbB6c1PnkHJW1gJSRniXbB
E33DQsNSiUmB2PJaEQimABaNuTUoO5SaFTcuNG2UgacblISyNHHL6AbJ3kiLw610bry1kD2V+qwP
hEGzKOTAKRsdVTe+/7iYXEfLtMIZbjmCh2XM+ezshoSGovnVpIVJhdA0+RyFj7TUj3y/dsSLvq0V
ILYOlSdhuUQ25WCpMXitH36uYxa8Q73D/+2XNrVdXh1lctVhy/1YpLp7IXxdh627oHum5EfjatYK
7arvLt00SzdSQg7JhrACRRGc+t9vnwtzjxeHuakugptyrIQYvzoNyb/tI8WFkMvb897bZeFBvw3h
0b8GcgKnxdidlD+pQGROSGJwME3eEquNh0W5F1ol7Oju6RewIRJslakV2KD7umUY4aPUcniEFIbl
jZIOFLyx4/YzxNDoluWNqUWT0ZJFxlM5jEFMbMzkVNu3RroAT9epllT86Bw/eB3IiTWhamQQ9LVS
/KLn/wXvSrNAXpTmPFc3N/xG/qESs9jIg75Qa1ixlEkZx1xLKjemuQasK5498nSQtiK5cSu6wrua
MM3Zg9fTpkwKvxaX99zprETwyIFgk4i/7Rlj81KdWmx4VjU6ZKm0SCBb8aoBcju3cbyTLkRsxIDE
mw/GgZi2NbSChxAtgubvKvZGcvUVxPTRMt9Wt8jyDIAIDcLfkRzxt3jKvk4xMCk8dumF/rQCbKSf
kFgTR/8ELeTGa4pnB7m3G5VBtAHz8Zz35Z8fricXHFv5IoGfddEehBfbeIpEMmIVltlM6/QzKesP
8mlwpxtOHFfgtxv/f7IoY/A5jSjdoMamoAzpIAy2FzJdeBoDiTN2T812hY7NV0oEy4gs3+BGvyDK
BLw38c45L8nELb9fNjhj44tszIhRLYyIOcSX/CaRI/x+iN4FNTetJlWkclDgl/qVSgkyDKBAswuY
xu2boKf/Ngt/qU2V2ki3nYl+IsyYFbCtf8gH+42ibSL6X6iyR1nvrsQQRpCWd6IHNs93Z6PUxhSl
uHxq2gXC4dFtymz+ZY62ktiQQ+ujG1j+mYuhXH6x4i3yAxtcsA40eaXPeGFSdzXCGSPo+wKVuFeC
DNc32acQ6s27J8LdUTojDUv3eAEidvmrpIfzv7Jg6MsazyQ7a8tQhNh6Fg2XhM2R1j+uLkoPUQDC
jdii+xJmzEZzP7L60PBCtOs2ABpr1+effGwnw7+ldK3X+IB8nx2dtAbsHSV3G8ICOpXSz75fADqy
5ZB7tv731H0eq1Fp2DGb3dyX6NaTjWqQQzn1wmrknRsQCPY4zCYKg459JCyjimYk9DhH1TFu5ttW
h1G98PjKxBBUYemMqWYmJygXT/BfZv94p86AHqfOJdr06MWHFjH2Rr3qUhtX5T6+2ZLUqTI/lrmy
ylxnuxsLYypjTx9CpQouxAbshuPW9VcPH9s0mrcX+UeKGjGFSaLUuChoCT+Fpfqrpp5BiXnUFzwM
06I0CC9Ib56WFR66KJJQp3aAzM5MkBpFwrHmIAMmmw8SOh2HxLVXT6CZuPR6CAw26lth022uNMSL
uUv8lxtzyey+53CAyAvt3wBvfFwu3iZoTxDTufx8GHfPaC9BxtK3STJ71ZhxURSkTm/ASmF5jkgJ
fJd+h1xOXFfoPyi6anQKz0rXdTsKUKZ0juyYcgdhERBpyCcW913cTZv6sGppYX/UUOvZrHLNL5Bw
QCOdKtWo0uNW9VayDt34ihmuzjJtZ23YINTUrWCmK/ENp+nnVNQ3WblJkMmRNYzwa+rEBedaZ/br
kAR7Y0e1kfeB080L1Z19Uvxw2jg08mfl+7t6YvOLhaA1W0/ct2oRPdT2jkrOTYr4UoYH3FY4Y6QV
yizI+W4gU4J9FQ1+vwV5SaJ6qMHcxS4pI3/pzEdJ8WMABVytT/TtlSPd1NTPapCYWA6YDN8iSGjD
wbCWEBsfWZKB52SLZy4HaHQDnk1q/6UfoRwjzShr7pi0dVkuvi9gQsdYj71r1gtPjAQ0/Hr9vOVc
ahbHWFFPVLRpbqzLo+rkoO+wvqEW7HMmxXOusYw/HZYgf0p0pLc2mvyLECNvjVZwNRQtzOEIiPZb
dW63fJYBV8XzVvZ29Rz7hHH0ipSfmJDjJy6w02W8QCIhDjouGU2tulG0xl8hjrm4kK6GLC+CI1xr
A48AkfrB840YF/nZhptd8X+3pU1BaLGVeIA3y70pQhoC8S2d1HVtiZbCW40VQKgrRbQdhZhk7WTx
XJl4WPCyQBLcCBme9j3ZzH+aGoTsiqvr6DjCQRlJjPbAMiXZNjlBSYW9s6q2Rmrppvw/XyRPi0Ta
AsFY19dNGuOaCCq/yZAFs3HtRoWv1djOJqY2TuowMRg6a2vRcTHQb6RxLZUWnpPMQTmwU+ndvFue
Zq6guPVz09vvRggpQt0gJwmMaZGUkcBw8QFORSt8ScEd4CpZfXz/4knp9iEDVphM5iK8FKFDxYen
eZKYVk3dJgKKPzImz0ilVuepfUPRqzydvmgD1l9zkb9YrydTRs/muOG9fNQYeB1fZbnRD5mZn2Hj
AZh9rNACDUv8S+AoE9Q5mr5YKfdQDcrl7vq2vlzggXjX6oI+74vWn4WFURIfsGUHjxnQaTFlD1TE
PSsje+x+6wBT6xji94Nt8vNTRJ7d8bzgdVasB5U4rPW2p8Fi4LwgQj9QOCejPuHKXB5XlKASprZa
ntWnWOSV70jtv1AQ1ffw6dCAyrGjrFl8EX78TuU/XTqYm6nJBYL0tsngxhHLdbJegjTZBClMMhA/
1OgXMRKHrKI5qurJglOqeZHe941hNsjW5bSwcp4gL2piEVK2xPXcc73WQfOUH1JoM5YEXyzHDASn
9e44lXHepUaDDbiwzb7w5hRN2CrbXMJ6oc1vB8c715UvYHQ/eaDWysYbhvEIrT57Mn/o8tBxBtFj
j9Pw+aBOeyqRFQrVxQleUlcDqnBu2S558epuvmiTduKF3T332+RBAiMNzQ+S4MNcYAbPJGtIFZ45
OGE+HqBYiy3K3bbJgxgvAz5AdFjWhDb9ubzRAX/dCG4oeL2Cux1mDKfhffnb+l3WJ8m8rDEJ/AON
vIsQUe53vMTetvm6QbgVycY0yLz5+tRlycmCb8nFM/o+8o923oFMy56CtKcZaNjim0tGVdn/+YKb
11wnOdtxxoguMwRPjyv9oZWaroLvu+D9F20TB6SD6mAZu4yRvB5wp34qPsggUYLZUf2v4I3dbvDy
J0gFoG4FMp1jUkxQuHRAv978K8vf7Rx2iy6b6pciYE8WAwGKeUMVJxmnVfab88ZKnyzY3eA8/QyE
9j2dfMfax4fBqX7WIX6HjL4X3kYdansEegwDw3QepOWc2n3iexBTx4SHzEzD+ivwYbtRL0Phwj0Y
sHXsF5NWRU0Wm5klmDSrAgFd9VGQxNhbIGBKlrS0R1Wir3fc0VWwwJozJMUxNMyE1XhM43ICIDnL
Qt3N3KmVyxQvaQZgbH0iHdv3CwClOsWg1nbN5PMQRLgDZJ26vSyDjyODOYDQlPw5yHQY5CGXPTpc
OlyYjOIDeW+7lFWSZInLNlEgC1x04GoVxKJjgRCItY6IdT0zF9DACnY+0XSURI7H9mRrGMponqYp
0Efpjg2fiE2hDnFrAYVGxRfVs/diZcG3bfDFfl6tp/d+2zNqdsBYnyHIr23Qqp9nmxhbjAIHIVFT
1INXUy9Yd787Op6JMrj/j9qsmhzhDn0gPNdcKte7I122Td7Xw1Cr0rI5Gtoo4KS+VPo1uf7SQnc7
K1IQoDSfWiE7Wy/RiLS8yURkZWiVn+5awK6N4h1P0+zakX0+mTx4icTsdNLQXp8sCBAvN3UkO/VM
vOSeeKSIvQzRyo3djlUngVF/AZA9lIAJU3eMKyHZIPW8rMjcQ0MrQb077sAnJb/14IR+xwoiB6q3
npyEtT63lGFPYoWQ3SLIzB5s4mlGmDvIFQqAoUEZtTO5C0lstaT3yXbRcKH4DUYC2hpVffSC0viv
U5IoAnxGfXBW9vwz7o873dxrVPYQsutjkT/xgK5AegKUTdyIhubRYqhltzDn0X/K7WrZPgCKQQYe
ShFt0OTO2R0ISc0T+254hAExCVGDtsn1tJ5znn9Y2Szn6G+cUPT54wiGLDjtFYEVJoV1KDAybEj7
1e6aDbOA2t4d9mXflQ/0VOsw7jKgSch4BUPFEBLK+eLwgraDhPt1j7/L3GoFZr0Tard/l4H6H6sf
d41CYMhzM0z1uenDU0TXmWGHsXLEEZt/flPb4EgCEbiJzid0kam3qMFr8p51bkmFo0sK7IVsDBj1
mnpYsjNApw/lBssrIA3c0DJvoV1KkU1zHYD7uJyJmQ5Og5UA6l9g2nD+zDYFNXHRpXTZCdH0yXqS
FY80EexsgpACUBD8vqNb/mslhhYWvIt7EaWAC/TRX4aM0hx7fPinV84sMX1OBIYB8I73XcdBWCak
FZZYrkzeUVcBvkAcwezXGifUZWFoJI8p9frZ07sxRzp4KV6if036oY7Yv29VLpcjYKMTQPnPx02F
BFEXqF3QIcm4ACUloZK8yNm3kgt+jGZX/2X3ryqA0+EcJnuGUYU1kSQZD8yDLwifB4GMAtbQNx+s
51zrGEGRZVJXfvHAuIZqHX9vmozWkojUrmqF++i3LvBj1cM6woVtrStMV8sXYCSMs4mYICWJa5LM
GX56o2jjlXQxYMEqU3IQO4nmhBTjJupJfgQjdN+wCK6+FqZNem2AQlOd+cUdqLslFze95E10g8DU
13TLOQK/2xaOyZzJpO8pCpIewGQL3ki5Tjdc9N51iCsLWsmXqgTEbtckvmY29eiF1SRnetVW3Phz
BEGD2t9YM4lI1V0yRM42Nc/6RDxqua/M8HRSxf81U7u53zmaQo8L1Wkx9+VINMPqDDMWyzAv9DBW
Dv+JP3lPd5YHv7p2B8/5zpDrT5i3+/BS6ctplU6SOr1AJQfeAqxKokglxae0wqjduDsKAH7yasfi
yHVqS3bUIXNFITePy6LxGkFFpyceGfLEHQw1Z1Vt6jjVWrdP/kZoM5djbK+DuU51FugYHERFQ7ER
UvLAtnyIWcuSCeY6jvy5OXU1Z4I83RbCn4u1EG/KjF0NnNouxMK62o5NXyyHc7pY08a3RIFbdqFJ
EZH6C3Owabg8xJtEYV/eK93IhUCYvclxCX2N7RZCMYL6t+wFVp8agsZl6sYqUDrmixlE9aN7nz7H
scxumTrqaIzCXin4ubrvL+RXOTK+0GAeolscD5wTodhSSsf/+BU305CeCMPWUk7uzwxaU/dcm29S
699lGZ4FCA29Oqzh9GurkS4cmmJdeEgQfbfdrWo1VtpPif1PkThfZi3D24vFEd6/+zdiFUFcy2WD
oIWw4GZr6skcTj4n12qE1cEIMQqcmAqPIiMJGP6Jb6TWhLZ8uc22Oh2irw9INKxayqrmv/M5DxEe
1reRebNbeBtgTTf9Kqgtov0CZE9ChnsBmaaNZ2quGRoDicTRxGudij8Ec6pX68CWk870zCuhAU2l
P7gc8TAedDCpLLNe8td/rPODpHf5ZY2hV/wUqNEIuTq7uv/v/2e1i8VAikEv591Y/vOTwuLmGu2l
dtUb37zGGkMpnFKCVYvk8msSzvQyqeCgOJ8P27gsbp0MtIKGKcJHjPeqhKxlDZtVOvlhwbdNwpWg
lbQ3GiTm2ZiWScqELJU/m4ICX1AsJWOjNCt8TcFuLuhh+byda7DzEwoW900Z3fOnuidO+uI53EZV
OhUqrckhm+1Ix3PA6S0zCZ1DWTyBx2YRsy6aj/ynqd3kWsUkYtLHNr4KPKSSadyY2ST7qipwhwXp
aJBoqwnCa6JXYk+1h7iZz+KwGewZIg8piz0mlSUCPpIZtGHhDayUnkDCh9hyI/Lyz/hIaI0d86Ny
yw8VJAL3Ft9P9O1yRuRvgRJ997VMLKSkZTGrl+dhwRXc4Ip9lj13yF8uzz/Z8XotJLrWPNxk35xe
xXjKcrRcBLJ7AhfdrpNJauyIZ1wW9vD4N1JFuKMG/vXw2ruojLScqnEjkh681ERJASR2jJxIL+iJ
fE3mdRakR22uqtcM0TgCI/V28WwLlEB9HOpijPXiSbYY0WiMWP8avgM9X3YZUn6ODm1ETZmyf/5+
FJ3wod1fDXTko0GriMDSeM1ggtWWeBrsaDo/20kb8XoUhq/OJp41e9BnjYpYJe8uCxuVbEtHqEZb
RxzywDu5v+9vtRpbst/3GVO0mgQ345C86eVkqjy2NCiJbpAfOks3g4Uh41xm/DpTr3uIliIN4msK
UNcbstSoXnKOZs8Z24KzFmHJmiSdeu86EHgEie1/8RpQ+KkGuVpx93xCDjvS5HhTINPkemgYnY/h
7hjwjP/KQTKmHLmeWoYjuq4aKvKw8CiM0cDkPVwnPru1cnhHUsreC/rs2lRQd6lZZVHgVDkXc3Tg
IhhcoS9g64YvooEoA+EITeR2baw5ggHYGqFFfrFoFAsyBUomkfBPrjFZCpNMTSrbdvFOaw0RUs9r
hShBPlGxH64198AjU+dXtwu1WrTrehQOKpWGMuhHJZ3vfhxSuoexV28Fn5Wl5uO8AKHb9GaUqtqY
TGvp4vLZGpsa8N3qHOakjpg5skgmdGyC7cFTpl2ZfGYdQSWbuAAOdO1OFAmp+UEiZwokZRfmhSJK
FSMAPEuBLYPhFjmIQVAZkBmOr1M9Q5/U5P9zhHOx7BW1INRHJi77RIAsyHLXV1vupk/DKQDeIe5X
0WFEnQ0xPJx3+PyXEY/+qL/VHpnubpv1Hpf7EGtCT0t3RQRZ4krCKJjNQYmnuDXgFyD58Z5rUmZa
bpeV5iytOhWwz3KU1IeN/dzYw8ONm9Y5O/6D6m/9LKWI5ltfNIbIgUIVEvUYf57y2MUVfMSfL9uK
URS5NSR7/8rNDGxn5nw+iIYrz7pphl9w85SbZMgsUf6cxLrimsc/BbWK3OklPHlsbvut9KDIIaj6
78EGyJ6YQ/rY5xtx+foBAJz6NQC25l1/DYrT7TI4iCQLhld+U+GPYgn4IXdXN8ZuEnv0UEnE0tq1
UPvhCrcK6tCUh5TwKvZg+oofetY9DZFBfSiy4/Z8Ad1OrA4HLUYScHzsC43LgI3VIcFss+DnWOfN
BQB6Bm/ryLuWi7PKkSYXCD4Eei1HVGXgRDRV+NULk8B6Uxuphfq4mYN0D5/xQzaRVklAr2H/IuzV
ajTI69YP9Ked3ZqLyan1tNjEfRzTcAbbfy8lg3cL63Tk8ZxsY3Yoim+jPiIV88y82tFMYamvtgDh
cgQ76cICeyC+I6DmBoWcDwjzlz3z7C0aY1aMPoGyZ3Gm4jt+d/PnTzxwPC/C1eX7q9amLVUE2RLo
R96QuqwrHTU7g+pi6ccxqiatb/NDm9RwhZnQTKvN+PdQVVYc4JSle515KcM2pnxLhNwZgutpI3OM
SaFA9V+RULwKs0cTLFgjG7+5p5A0SYNZ3TcgNX0OgG93l3o1g0A7cWrNFD8aWh8IBa3T0vKwVWyU
0J+LGD5SwvSpiUmdXcfQkFsP92BNKlebrzZdfXNKMMDSeScfXt9LafVjKZfe0eZ3PDGLoiLaqdID
+YS6oOW7gLLLG8hebkXXeJ4oS78HKjD0dPNhTteC1sePmC5XoSImLZ+1D32uKT5KTYFlx5dWXTTY
gqLMkrDBYt0cRGsGfr3oyLvfJyxrZ5yc+PAVbHx4G50h2eeMZvcKflo3av357Lg/P4MUd2TeFh/x
ldzAMCoI3miEV7sgpUgZBukRnf7L42/vf3B1XSG3VE7cYqWbtj6OtaMtbxEvwLGHVpX7v2F+vb5I
gfR368okIpAU0ijQ8h7/GaETEgGfcWnoJtwqctBjkqfsg44DytTkqdDZBL/iBMNLloPedST7pPyY
3NBlKZFQg4VJ1MntARpX6wk/hsN6ts8V8CE69EAtZSLrmdFan2ICnIP+cH/tHvm4FBQVkThoylJs
iGROdf0Cavibi9FEERtPzXn91nkX53oNyXmpM7bNl2a+j5Q61enTkvTG2FlO6DkcIHA40DPZo2UB
AgoZLv3NFOnUqyWLxAvhkLNte2eStXw9qNsNSxjgRK4Rpj52EJGTaJyLu8AwN9ZfxBlLs61xudrc
9JdAz3hciNkzjvDJzfcpEEI9qDU4MvnnSeqKM4rPED9gkC+XRjQcjeKww1lGULq1yMeef+A+fxg3
qeUWQYlBeFKaa+fJArawItDw6X76rtpos/EgY6XLKGBtYPCpZZYbAFwCvbj3hbtv2XluM8593JOz
TqrNdVlwKspzopIsnPbArejHNP0UXZYI90Ac7Klen/PZoF5CL9PakpS+42MFxvvOOBokxT1LCivj
xl+k+nUl+17fuChO24pgMTdRj13tWiORloOhL90FOzKdaR2ihEBlPoLEPES/TS3I2NGk595qZgmc
gGq/TTdMt51Vt8cTuf6msFKIyssS1rPkTqw7vjxq84YBOZmPvRQpmws9k+lv51qFt7yvRudDMJe3
1zc3PVL3N+S6n3P0SC1U2w/QsvL6+XlIqalfdPTbFzkZ0AHaNlqHKIKbntBePpdY2dOJf+qOoSWp
BS+VDEFbH0Nf/lkRZbMqRn1lfwZvqigyVCk/cIeaNBEtJVs2cNOknAGk5UuMXJL5UwophGHuqnS+
ONGgDxDb4Jw3DvhS2vvKj+BL4p5pJP/suF1vfqwTm01z2f/fN5h0Sd+KaXUy3lRaK2+F26FLyroD
yGqWYh41puz8b4V9GKF2kWwRrGOf+KnFzaXp7TAADKreWQOvprjN4BGjqHyQro74Qp9WJSkcsRln
zo2CIhHq741gg84WAYvHdFg2y7xz1kwQ37W7O//7j7wsT7cQlqczpEnFHLSPAnYFQmGson5HgjmD
AKT3QHa65bxxDApTOxrcX66WWEbJ44QYW/llSEBwpMPWEPZ4yrMQN3uwtwdM6EUqZniQxarBxTxb
2YHCnWXI9SCwl3hEZMlsHRhU9DTLYlv6LRnpkUdRUTNg0mrlPz2iLtbU7p+rwBY7urIaKj+sNaD/
6IS7EFRtoNt2eOCk+6qc+iIDl7kA0yJtfX8+RcJwpVNCswPeCFFxujWqZBiXUH30mey6LZeFMhry
h7/ebsGTmzyVrDMfxf377sVo4j9K7IaAOJpREgMxcVm+2jbCcf6PRRFEY6dmEmkJ77mJwGNp5OGj
yYWZ6pCrFRmKcho6VR6xyYqdcNXDBuLSze4Xe3YMkBENK5DEynfCFgLkcTP5YJonVh7V83wB1TKR
y1JnTOEDl8NU0p7nU1GOjt++j4qpaB5yBJb3ug36cRF1B5C+DfHUQxgOtqlRKuMQSKx8uPotDoKl
1jznP7U8iMdbUnIwF+I9k3/300ngtgQL+ZCNvFfpt2F+65LM6HSYm5LkaSB+LjoJxmasl8F5JfbX
lMf5MRWXluuw7YU8rqWpeicKIyxkPLVJUn6eT8WQFEDag4qsvy1aCp1NCB5SYPyh7uHQ5H8bpogr
g43LHuq+HQ8e/b+NylEPoYOe8LbDBrDzNivzj6Khf4Bnu9GJKGA0rJreBZJbDfJEzjiyfSffmeZp
e3jq3Bri4ofKy2yVOqOOm0e2gbsskbIvCskQtMnbn4kQX21wTAYCrKM+MLUAFv9xPi+VDAxIMpCB
gOei+fEKGNhxEw2rII8nTf7xTi56pI65ywrfJ4b/HBL/MLuzivlw/gzbAbnbTItF3GD2Je5huczz
amp+/HD6E1S1TXhVaa+sFKIDfVhpvlh4C5i8FJSHWo0+MPbEMeYE5OL5TrA4Fj4BqIaz1UpQYPVo
QMQVYk9JMfp4CsYs5YRSp2eRHV0/ct4uHSUVfPlPkkaI5QWPzHpXJVwLWh4rp2Wr9OMeLa8UZAIH
wd+T+M0bKk815uiYaXWCd/RZkdq856wms6zSBc02CV0iVwiso9auvqRzwFa/LtcESfBg/vh2oAu+
AeoeylORW1gM++YqdvD/nZFPiD+xqd3HYcJRRJNoN/mdarc9R/Eb9j+OmkCAUQbuIjyBYxyS7iJs
gHjD/q5o7tDZ0RvrF1pdDj9Tw5aGJvVViS+caKD1wKaq6QuqaR6CTFm6kKUWJJs0OZkoMfLstvXm
c1lznJg0L/31veY12tgnaQT7gO5NOvDj0K1gtISRmeUKyFXuFdbXfSfhWEPxiorCwSA4D7UZN6Ju
3omjYkWKPtGr8PGFDBczdXysgtKv9ZgiDcGdMn6p655VW0NyG0D2mXNI+mUnv+H+FqVJnoQb2hF5
2tXn8oYa86n/5aoUhsb7Z8cINa0R8CPfe/w1DLzuVb2Fsm6HszYU7BgxjqVXDBBeHYYHJtn7kWV0
RTaHf529LDj4+u+rqtgU8ZqG7wz8YFXZJcEds1wY8B66AAgIotADaZRPY8741zW5cbfR4YqpsyKN
fPUV3B2zq2XiByE0ZbWR/eqfoQOGUqvjhNc+kzaEPsRsDqZmaIQe6xN487zFxX7PzZK1nU+Utitf
kqcfxFmaLA+CPSmB93pN45Sg2AGqiNAhNIj4bX6TGpQyQLuO/Y1syZH3K16vXi4pQdeAVLt4Tt2W
edeW5hYCYJ+wNiabyUDoW90+Stai5iAhmeLVCVgx48ENxl5pYhYSwsXooBEgOohBoDaPiEACg3A/
c5YnWJPL2+heZVpzdsO3Bai4UVfdHnNDxE4cgt/pANU93Q3/FNdC96q/SVI7qTejdv0rE7ycxKHB
NZghpoY+GOHlOShijenc8f7veupcnPdR6IfUpP8K8+/yrlzG2+aL+2Zf9KleC2ZikNZXUMu0TmWZ
Qus7wc9/JnXwjfR0WiMDm8uuG/GLZhWQ4ur8snlSD9Z4qr6wxRJu++OrxfyGl9nwfY+hqWZwp78E
qj5G5wY9dzx510ix1rm81iJfwuGHi+Pvgn5zvIL/oMXENevQco7JHky2TOnPWCCKjhMP5/nTRLLm
svkSUxi41PfAUXQ/cDRXrfzauEuzh1LHJZNhonAM/P16qe4sAwhl4ehEalibPLVe8wuthJVaJN9F
kN0jRMegGmyHTBE8k2+KGk/bM0EGsJ+xnnMuBRIr5DQE0/Z64ZWRE/Lk/ntPppXwXzUjQy92+XYZ
4wy+Yh/nhmyeCGemHyfirHXMsPuuWyyxyX/nfoCtVm/l7DJlf1IyALsTNe1FXvOwPMPSPlJRUrmJ
2csJ5B10UQDWb0Xt2s5nsF/JO8Y7yoX6PEU5HqNGIDWiX5Dfqh+MuVcDYBIv+IcmrEukmdy5ZkKV
c5gO4Tpp1CDwWKFadF7mcSHL2UcvtwkekeeCLsG6a6zQDWeuqJz1PyesJHM1Fh2V1cnjtsG70nyF
tksFFBzB8mwYuobRj+t8I29363Phaq1RbASWuL5miQNGG8Mho0R8ul9o63Bpsn7EBXAkLTe1cwIq
LNa3A8rZYfxRBCUshYypFDeKDdecNEBNUlbMnIeXio9YNurz1oqB+2YFkSh8tgF3r1tmNufipHZd
FdAi5Zxy9BNg2UMu3glbTTS5MKrmn8waIOq4TyWsRx0yuOmwuEbK792q9oIoOjloM8axxczI+SsC
reDaPvWoQSZsEQdjQbuYuZMRk/QUM7t32HCjI8t1AB+axyAGDcfLQmVr9K2e/Z1PrTVd2AoN8Mgu
A78YGVrDIRV6hseJ9EMT1GKkfdLmkTMwwjcpI9y+kqPv8j/ssUGriHjTDEPlXkOgyI1/1vYkX+JD
FvUBKJFpVBTg45VbQpFPXeLaGN7KRqMaHdt8PLMxPfQqZm796Ewy6qrE3iZoXgGYUg0EPE0TACy9
abTuZeUT7hK4VxQyGwWmoJ66j8kHI8XWpb+1l3abV7RuqAWmyklmLNm4wEmgeGTWmndHI+8/btQy
OR5XGHIRd+9BqCW8OfhObBHG24Yc3/PD59LR56JWSvOAdnmXZRSoB0xmCn8R1s9QAn3Umz1XlrNy
oOcfSRZpwRZ2fJOf5AdZEG8utUsZCkU1dnhHAEtqtozKYoL/xGwpL1bCgrMRAGTW0003DHqec1I/
tMO5Pm07OU78ByQXuebwMFHn4GhGI+QrDqh5i96qKnpa7mqQ1rQBquQihPJmzXfXjNBbXxJwlj2i
L1Yc+fxsZI5HDI0yJeDlMJB2ZHOCz4E7vFOr3SBeoTH8ckKQjJ9y7ugYq1j51zD6cGCyi9gmispJ
RRpLwnqmByZXS16Hce7HlGK21Wv2P4ZsdTDWOAd5bGG+LNF5jW2CKRD1Gdnpx9MXTHGv9+YGXGMe
dA6+9mFsrQzA/n4oeQ552AlQzz9wITUIH6s6N7PPf3NgI/GztFQoLs4cEZFhXJvdGtB/901MlGuv
+x14gC+iJbV3oDZwWbA+pmR5wAUjX7mnOScKBBOrw9TWCdmtujpHOuzLyYHZNkkTYbsy/pTPkez6
yBR0cbFYARk5Y5PtrJEj2V/kNJadABRjEEohgfg1HybOJXd5UAe4uSkmcSPuuEf6fe9DhBSOsSCB
vh3KYBnqyG07W4w38pigaUlXQBsmSDcOKAgiV089Jw7j3y1wBrnjcfmUtCnsHOifFkuXG44HKhfn
aMR9BEOhSwKv88SSviixwH4aX8I2DZaEYVryYoYU5hWqc/mFLIrCO+jY6/M/zyhcxMHAaI1rFI+6
phu00z2XlpykhRhSMZFtsyEPbe0Ub85TLTlYnZ67t9WoTgsRj3GH0uyZ6jl6M2suwSAJ8KRBxFo4
pqvHiv+R3k6IkYGOSWUMTrSShrTiM3k5bWMetfQTiLx8fhpUQf/nWm7vOEOHfg2/7W+G74TPuKYz
gipuTVaL/ZCnwL4tVszPXz2lZGCwiKspclPPBpBq5SUFXfEasA4YW/1kOUHzTc7sZBJZrF/RMXFe
nDnjv31Ik5VcasXZrCXPr2lciGvwj/5cpzFcVlL2hdn0YYg38orvgaJ9UwAHDqEdYHMrjQul7sKk
wZKUJBiq7ry1jyF7Q5RJKSkiD5PRy6wpk5DbThTjGhsEgK9fSuk+I3/ap/oOJ2XLXGV5YKMchXSU
pKQ+KUQW7ri2uttNt8P8DovGwclwfCL8TnM7GDrTAYTukZztU7LK/NnuUG0OIaaTSxYW+Pgle9ex
UIxEO+paPcwlCVAzFprdAPJS7zXNz6psQb1fU5mCNPRb3v2xEe65uCb1GjKmLG25kVUkEjK7dXGW
gbHBo2/+f0Kwv2Dg+lDXkGaResl9lBFEviZixNNIlY3GKTOd/3SJyPFW8bHoO9yTqFo6oYkjwwgT
MZEFlEKvKdIadS6MNu6dAdxoKjLNNqXQ5/1HpRZAgfEK+xYRTAC57qxq/jWGEDMVxTWCu3zRSo3l
RUFG3fm8bVt9PrfLqj/T4Nt/X7ap4ZyIqzKQky4s14QF/vxEiTvwIjdqmfvtkPKjdOHM+URX4SB9
NXdBuxSHl2phQ/1Wb8y186AT/CJeyjiPLcONMc7xcOue2FGsgLxMsEvGBmSsCjdEbk2RZH8nLK6t
XyLOBUu9kosbqXx/gVHy/BfKev5HsugQ0z45WbqtdhSNu9YP8e8jiD+CuHsPSLBYB62evfmfBLJq
zzBmp0lGYVcsPhD4jpd7BkNIQU/p4V5L+CV/wLsoNBlTC0Nq8YdAHHcQ0EGE638OG9ebZhRxazHk
9KebwysO4g1/MCgw7vfaB61K/pcvOhfORftjQ+y9WDD+fi37GnLr9BBUqytR2q/N54S5XzK+tMAW
J8QOGN009eP0knxDkj/ZX6KE1Yw2Sk+3LBcWIhhpSq4wkFBC6l71PLKeMj5rA3JkzAozxt7BpBUS
Z8Yt+IO4d7mRDjczuq3LxF5kXV9JBUGaxYjVY5bQjrBZwx8m7bFJoPFNX6JhBhkVkwZ1/AjxjZ+4
BwKDoGV4yA1xBNSKpuNjUvSxiXuT/RfaSdue0FqnejDZdTnzEglYQ81rtki+F8p6I3djSC5UDjDY
ZdHcPSU3TKbzRvuN7Bzs5aONFj34KahezywjwQwgpLvp7YDcuJwWn6aDSZHiaUUqDLpFkb9kJ9bK
y3lK1bDncDQz7rFwy0nqFN/uCQnjyKCU0kIbjjw47iq6yXbhCm6X94meZmLUaOAdCTYeFwVuVPTb
RKwCOdnKF9qk3D7yriYGuuGXmFVwPdiy5SMPmXSnoJ0N6lAllwWQ64pTx1BxdehbogSH1wEXgYUC
Fmt+tv9oj04fSGOcGjpHeFTcKfFLuz7K2gVRKBXzTIGiOpJBDMgS3r94ay9KOAshIh/wS2yVZzMm
KWMipXXcOQ4p6S4/uBJ/akqunKv+v8qPpXE2G77GBFJ3DFk+5Rh6RmqV8h6jFwm9Y9+KP0hCZtZI
gHvcfBZ3Tf2PfvJwyi3kq/M+7gXdK3aI1rigj3XXIqaQCKeSIpDVZdFf9pz6q02ceqmbFmcG82EE
nQYos3bNj8FTbPWEduUH/DYbDjMBv2RcIw+zLqUhIFTHEmHeTEDXn+/Fceb3rycY5adH0L57PC3C
aeBfk6EJBcRgYjD8JGqjDX2DdGl0ia9l9X8nh1OEQJ8XSeVWTlAuca4rsnAvn4DNFd77aML8s8LL
2RpjjXRpPN6jTLQpH7tvBmXkd5eJ4wqNImvKMJtad/W4WLl9XfAHB9ASFck4OJrTfTLXbZUBo//f
ISWT63d0jv4xAQ+H5zg8tZ003EOSlhl+duV8HD8eYqAsRD+6ioCB+K0uIJXQ+aSBhEFY2d3w7O9G
4C9fJI1IpK8ddXlxWh6EvfguDo4sX3q7+HUqhQVIuI7xQjuwtQOAZkRTuTTE8mDrq8yYhbS0ZwZz
7W9bVoZAeagedeBUBwYdnHtOITv+4/LlSYfDBIrmQvyPp2b2oO4sRlN5aU2FOAu1O4SCF0pYrTIq
Qj5GkXekoVa5IPjsLsjD6q+WHqE/cxAuF5af0mTDhIv4TPI9ndfSKEScxIK/A9ubKJcj0LoBrI/3
gzO6JfhBdpSBn1ZLh0rApdAtsbRNfd71iJWylGyCYIcdZNyecPTQMeGwPA6VsWA/deXhmz3S5F8U
qTbEroVOehduSTGsXXuJMX9cJazHoQGlR6MCJdyg6u9XMnIzOaWdaxhdBzQQro0BeSp5xN8+JC+u
+5+G0qMHQtIb7473RLDSBMYdKccADXOTJAurxoUIeCUA9/314q3asuV395esXyT6ERT7Lg3Nz0ct
rnFuSaYTeENu1C/q1tcaxQ6It4YfvixWSjC5cliw+x8sAbxlNnoyiQGzH87TP+5oAIuHdnNXn2rL
DD3kiSM+9LY5VgU1eVxduGxTr2N1nzx7+xMJEotktCLZTfMhwhgp6s2zQlKQFDyMw6gJ/d/Nl6OF
zJfgr1h7lDN6ACTKWGrQpa8hz/uFEvPLdXFQ2ZzEVJBRiLmW1ICORwozyqRzWNPTrGQoL2sPtF7c
XyuMECaYh1v12j6ErAjrKp3l8uEqn5XcPR42XlVs6gMAQNBkSD7fvnHGPOX9WASW/zF7qWMfOzIz
JBS2xYzthN9GG8gSB3jcRDsfarbYWLYyMHS7gFrtz8CUIO+JgutfKogixR37R6yINqO9Lyer0uww
pFKM96p7BYbU4CknjbyUOzhYz+taM59edl86eDj8tVPFkKi+NyD82FiT4WCfTKPMNXo4JNEbBEof
E7/GUccIhrQNeUHIFZdShetGSUPXNs6l/sg8wx+JfDy2WTyefu0BlMXj/8U6juhS/kgWwPqw4pw8
bXizNLtw8vKTu1RhaLdRDpwfU/1s/w0c+fek9/8jc3Juta4cLVd9YcmY+HvN0fByEkyUoSshrvmJ
r9DztUJCJgl5daKmCDY4+t8gkoQU4ePpyTXaWrixsc+iLfMIuglt5OR2VCu87MAi5+DVC3g1P2QD
x7wfzm+7NQTzYTXLjtoXX2y4fw1zmF5mNjVqLMB+fsU1/ZY8rz2bIYi5NSYTx5pUtM8s8kdMrgeq
btEEmJLyPyghJ/6f7uvrFqNerdTWpLLdKCS2bQVpfCMTCepSWyhKIC336QW/0a5wg3YHRURYexrq
JWFn5xx0V16uvRX/Sl0bpMDADJEs8or2Nr63wZPyeknEEZT2PR3eTPjB5gfOoQW06auVHjMwlSbk
jmvqskL0DbFiOhYRJYp7K/tC/u46OakJ1/xh9SnQuI1Nr0Y5L01sOIRSv0pLflscusY8AKd8t2Sq
8lTpv4zjKl6HmNtYy30xjUKYHsujELSnxVtmXgHRGoxlyWZ9IwP/01D4mOdb2IkC5erLuhprmWGn
D/BL2eKFSpQGkXaKiaAMfZCXJp/9VxbcHaEq4pdUAfeAVopmwqKsuVjyOFMD/g3BIsEO7jyxiVz1
E+DAKf8yeQ8Gmu/wad626JbySN0T2cgrAcXrNPVGPKzfluwU5vrlzm7cDMjaKvAiwR4vcZf7RmyP
MaJaUtvLgc3BbiqlBJQlsOUY+WFS13TdFUJrSrX7sg9auQyUyq8StYCteBdnE7m/Vgm19qe4fFr5
4wAsxGvxuEDizcdtqd7hxpBh+1eNH1ogXTNZYhX5fvtOsiAPR1Ri+uR3lKpLCTkbwvafOdUMrYy4
8i3XjNT5EjZ1pjukFh4wt7ht8iPtPGW22lTMzhjus7G1/0tiMrs0K5jw4ejymvJ6gWPTzAwv7d9f
v4DGEKlPt4SJ/VY5gZXwbakQjdTTXgGb278XKANEbBwVSivtTHg57jLZ571JMPpcm+EzoyDXL232
74S3X1+5gdHWaJUN3xi956nyEUmucJbzbSo2YtG2EZlWlgs5+PLx6uSae3l8bg4J3Mg6DDGJa9xg
lfVJhbk8ClAXLfk6OTdDrQGOXTkcXAD6UVN5oVNxMaCWUM7OguCLqBZYCa9C9mB9HnIcYA1JosFq
drUvHuLYDDPygnNOXSX+yQxDr41m6egqJgtETZSZUqywdp3xi5IDhwQ/ii5WX/9hs7eey3dbHJ8P
Kznq73LwdZj1XHfKmai2O0sxpLwhRgOpZELjxXKydxtriQr3KsVhxqsvZuF2wF452gNFy3Bn4DXj
AH8Dl1HpV0dQiIBEHY3hgJstutPVbp0yD6KOa+at7jo4hfJ3zvBMIqUhfqBz5z6+Z4nUW92jLX36
kqom/VYTwCbVnqaXrtPXtVG78Wvrc+tQllbi3uHKRoZ4oHaF0FHEIrVjQqhM4wHEKc2f411FnFjD
FrevAURYpXGAmbOP9DiEgtQdw9PxZ3gvPD9rAaMQW3Pa6fEoFFTi0uWq+M+YSJsA5/Jx7ymKWZxS
y9s6rbbSKyC4hDY3SlNm0RSaZgWPe6ez+AEUIBo8ZQs56o9mRydyxgsLNhWFO+xSxYgdwpPBN0P8
bcsyh2UgQVbrNA2dxgrA/4jusP0MuM1Z1XYl9y2ra4gvout+FQvDVLjZwPyTwqfEtgcYcz2mTRJ1
olGa/chiOpZLsgBJuvQqDkdzFBvjPSNoJMkPRco8OxPSg69l7KoHKyvdwgZx57j/wc0tIn4R/N9e
dK4QatYu3DJryl1jKf9msLaA4d9nhn2DQxcZBIUeaHsQJLKk2SQBhiiljNh1mHmREKEPOG44J/TY
qXHRkZCZCmd/0Z6v39olrlMZvf/k2JGS/Sk3pxvlHL8dS9ImlhYuW+5jzGwMSTioQ2RySOjw9d/I
j9HQfxVdftAdbG/s0OdRaGQqqK64ZNyQYmcj1Q/YQokB94LVsO44dIJrPyNTo7ZaeEfw9m7Up5aO
Mq3WfWX2VdWV4Gn4qWH5Ng4hkkPAQUr1Dloe87B9Cu6wqexcPr2z4mAo8+5Y/vM9ZeNpwt9ZG/xa
+0ZtbsfrBZ9FAXWrrnsOVss6d2fgtVpWK23zQfcYFUyoXjZZeyO0RPRhlfBsKQdhxBxC//oejtmH
AT9jt48uSgZgZz44+BxDcCOzXMA2bCG5vM8G0r9vaTq/Tv6Io+saDBCfkagcL3aL9lO/d7QDL7ja
OkABW45sUpWzkzAQyngaq44oo3GgpqaERiNSL3WOZzCiYZ5fZtQrG3ML2WS/k4a/JLlPRTU0YVIc
uozV+oTgPqvQAXRxk5Zsn8Lyhti3NcEpoVrp3sHgdI9QaV5HvoQrivFvzBN32ow/I0iuGRI0t2EW
ADtpS6xlp7k7X6rzT6cE0yNAYjWV5ItNRZaubb07EFgRVmH+pbLDel7c45dcm1VaWbxugnjOyhZv
om0fqn/U9SlND8rbLY9MeYDzPOcOUiVBbYbaebFOxAKNrKEqZPOdqUMehSmBSqrnsrAHODuTlaEV
5i4o7A7hg699ZRa4LFqg9sVLS5ZXn2dWOg7YEPb+2NCrf2HRKPCGGdNtRhKoEQYdLehOEb6C2Mx4
TPabUfqTeRqg+dCmsVEgIdy0vmHtmYhHFfCjCx81TExO1MfLTYAG9uNQd3Ca31Le4ik6gmAQgYkV
vVLvzKrZwwaXkFkaaRpxzUrHnZfw1NeeIE1TLKee83NvIet8pP2caWLuseIm/GGkL6SkLwkb1NGr
cAwklI37ncreJ5APLSH4ppMn2b2QQ5dWgLeJm/xeIcMSw3xgmTTOqEODpAmkdc1rqEj6YK8EWJqC
K8fq6t1iYs7hmVCdJmiKJdUcaWxuzzmn83MALGDUo3BBTOJaVQ30BphSFMvtCJjwb6AgXQCycSRX
LJzZSZAoCnd7q6Si1ovt+DUAq3+WKfLOo2r6P8OphtQEKIJo39B4S0mEL61Pu3hywD7M1PGTPoaC
R3SA7DiqesFTqxWwOio4E24JAttbO3QPcpnPxRVxSyWdbNBZWoSEm9DrYQb6XEIUunu9WZXfHJLp
6NgXgMx80EkA3ZT5roorcGKegdod6U9Jm7etqFqkI+eK8CDJMFpYH674Hj3qOTj5eyi457sAdQBo
KZ1MiHEUKcn6q/SU2DsvXQnsAhDQa4BI1leuc5GhiXN52ZfBr4tAr3Gn30RWuvwQJuhppuN3WGWF
p2gj9CuZ0gB3Ajr88W/ftfpyt9wcKsebOrAlJ/FU8V3UF2xHoYK44Yf8XK15PrVvjswovylBWSXc
bEXhYK4Iv0uSJKBSbCZpyyXPESZdbLWCSAQ308/XvFmAbquT7EJ31JFfaXkpcz2/5lT6QCkToZ34
9CGSjMA5bG5KQQ1LlnBniHW1fC7i2QJoHY1hKMrYPeh03tEb3AOwgGzSezQRoT9zrbmJz3BSm+on
JTsysfadm3d6IwpIOmX2AmbdJ0SFQcshbkAtHs36V847k1HVyR8GHfXslRGWzNM0gsI/m+xa6xjH
zam5Qpia2imOeFF3ovqoub1iiu2hl6SCUAKLGBxYSzUv9TUMAoysEUJSjloLKUmkCgL7tpk7WOwp
cDBuBtQUFSNtg6KkTRMGGDYH25ZMbTzH7hXDlsLdO4FvNHYuDPBHN5WVD5r+ugEEQl0sJMf5tsiz
mm6riM+GxPq2/61tfP5IDxnNrUaR+snGCbMY/mh9LOk/wJ2bLW2ZnH2UdDj+ViQIl07V6NSqcx4t
COj5xFx/Ha+7I9oQogH2Tu0HgHL5ECm44IAX42YoSBlyg4HPtpHCaAiyI1FAYpNWoaWEHPT+3CzA
oKQ/fEXRCurmv3j69TcnnWxPJIb017XpXzfNDvP5DcyyGrYyu5mdxqVCbzp6dHN4kvJb6CcHAn1o
Jx6KSet3F8aOxYxNO/ktBg1PsvUZpAZUSNeKEfwAfppHSkpkMqLDPrGijP8JUdnR6knyId7DGSTs
TH+ipP6PnW/y6R40wAjqkn4fPLD5jtOBJrwsaS1e1y2wuJpjW7EAYlLASTusM/PemtadircNzJ8T
FGiswtM90SJgo3wNJtvH/Q4UhloUhNlnDBQnSw+KuVv+H3DYdUioJQ2+kUClCZ1tt1m+BkCYQcQC
MLVm9jOks8w/wqo8aqpadq+CVgsJXDdmM5Ekgl700JHWnLiAVZR+bp/8dyMiwj+9jwg6v/TgvVMY
eU/CTLe0aXIRrLFEaHD1cSK2mfXydmmRqjFRTTGs15wTwa0ibMUxgq847tZfsscpfK5o1MCR3ZyB
q5yZ1y/PR7PRbCEdV2jEjJLnMHixFnx9bSgqXnES+EVuM04DlIYlKUIZdvOuCv+XrUW5hvnoRtBs
NbzBQGQrek7odZsQaL6FqrSNCnghJsHeyenGjG/RKq8kB7u2NWvF7oHjjslcTJSyXIVf33GUO5QA
o+5SpAHdzCGQnMTV5RRqL27cvvxCeooCyiqSCqRrDoosUhx1lzkZRRxPd6t7r7EQn28HJdUVPvcg
3jm/EGOp8/e8fw30xA39A2ic5LFmcpXt2iuiSIMBhrdvyppLGMFhmUcZooNg6MAwh5qCmQf4uF94
vm1kr1o0xoWhdOTDrJ0/LOm5tNkmORMwO1r8BgO5MEhW6d8pzCbSlq1eZC+Pg3/RmoaqnlQB1e/P
DGRH4LcWbaj7ouZk3tDAJt9bUIke8jIUYINW8P97tbWzUA7g04Dyr5I+XWAc70oEFzKAQQbG6eyK
YxJC7BrAuUJfloQp5sDCWgf6dn+rdWd5mnZLl5Sacm8njeOa0E1JRiRfLrwSDkmF5X3DiGCUSGki
xxo5/yEcajL8DkOmJnpDNlWfta/CH1dZWju0pkHfoFfuvHwTLrUb2J1SfJ4eziiGTBLCAZyCRONW
/oYbd2TktWsknnLwSRfJVxiHjC3VRh/Wf5EnbWf8DK6SddD6jRcTjUKZ2w0TGn+U2pydGXip6dXx
LFEKmaGRa3O0oNqKV3idSNknl7uTFb7G6T3UoYmdw6Yui0HFgJ5DkYbt5kAHrhNKHKe+h3Ox2FhX
2NFjUWkFGZiewAlxoYGRtX45HdpCuwQEgyHkLt47/bQeTJIdY/r2e60b+INCsiYvMjTO79KBCiTz
bHP0fTvdST22O6MiI+maouHHhtzEzLyrDGNmlDDJUbVluvspJ5Td/CwJPTXWyNvgh+XAZ+FYN6dM
RFgdJHjELaH7d8SPN72IykD+OpdejnWc1yBXJACOo4fQVo+v6x3C+ilNE4NdLnIOW78OEjHcEntQ
HZ/ehtRpYX9nkMNyWOmvLxw5eedTey/b0WiDgyn3lMb8tH+gCM77L2OMVgR2twzNXe3G8comFyOY
RS+17bEo9sPY+9R9n+PgZ9yjxmBYq+aRvIhqG9M7GblRFJv/pYDX1HLn6J1s0S+TIAtYELtgEsT/
3H1SRxWvffn4ECrjPW35I2MDPpzGqNKC/TuRIUTtzt/L7SIMs1cWVZNvsr0UtV2wwuXquc3fTuSM
8GieVXX/+brHbxyCPdZfB5tExmqWXxrWoFLui2vIU+5aSVbV4xakc1cFDkVHk1QmEQP3zxXegfxg
PxUAsKTTYjl7mtNeyamf2NGW/u0RbVww9IAQqcdv+0IDi7bzHuaef69D3CkGoYm+KOy5k2zCFRSZ
d+1wSfov/MDUk+Fj3lR2QGK1d7SqreDwD/6kImbM3+RbibZmWp38UiKq6rRGMFseJ3Zo4//CoF+k
P7dS/5DlBNTk4bdVinyGJATmhL1FwyYDETMncSh1XYgS63pqbAS7adMnvAKe3UjaZNkg0ndhYSG9
efoYkfnfaqhEOKSKkVrbHxas6ZW79UIgtn/xHjggSlHlZ36JZCDNnu3EYNNOMye6lqj3KD5smEj6
+5skQl3LLGFsGg/HzZgef3FPLP685owKkAzdfKzR2BUmISs+HB15BWc8olyylNS+lJwv5nbJFB5Q
yDFmaqg1UkWbUIZtw+2PvZvtF9kYnvJQqWEgTDTHQhYUfGDklY4MAlb6a3NSaHx88U7eYcAlQy4C
KixtkOOEeuHLl3SnUf/dBn+tQzyuCWFWh0clIeosSQ0cwit+QANwoTLLGNtpPH4pYML6MDBDrE3z
dtRESrFlmZSGsyZaE9u2KSFMfNyg0QVjgnWcvU1Fm3orb/XPkMyx4IWwOUAHGVGnGLz81cHoHkZL
ztyLplZP+4JPeFkgxSGS3W6MKNK/zolWAq8aLE6w7+BhV9T6LjHDiGFWlNxPpBIQgzfXT7sECl69
QaiUXbVYZcOiSp7WOYvbRwyAdkUE7NAL9WnQ5Kpbuh7sMPujnzjJfvH4Nor8NqfoVck3/jTrZbWn
hOO9gROTYYucDeQd8jkueq7ELekCTXJtKBQYbKHyNtAcVfYohKdEyq4dsW0z9z6UDFcZrl5X82Lj
FLG8bPZOZ8QW79+pxNa3/I+5zBSYdUcxKROOwPmBvgVKIvv/IQpmgglEXBLhK6qgiiJghpobQuM6
QgqEB+dIcw+ZNlWs4XgIABU/nYu6dGqg9RD2T8ZPoWE4oODAK94iYNyMEFBknGNW6rseQrf3l/E+
w6qqzCdmN6WwE9mmO0OJ9Uiepc9X5dVC1n36ufGXsgngD2YQp/uJLcUAdNCaJ3bT7px5S/uYmRd0
AO+oAQ2qtQtgNtx9k40ACnlN3tVRhorvvZ81WYxf0PblQGjKqjJs+FMaMIQ7Hzw4fFco9Uk8CdaC
SOpaA01sSmF+jEgHAW/YQiMHJCiZBsTa3FoVzJpvO/Wqq3B3ZlYTCBMEbcfmiB+k0eV6C727lGE2
9K3188G10zkTFGyztK2cG40c4O2eeKpeIk6FZFaOwfaYp8IfRt3cITDunwo4wXipiCfpFQmJVUx7
zhHk4AVATdh7hWhq5bAuaeZz9faE4p/ymkhewSJ8n2ZUDgPUdnzWVnaoyWNayGQgyoRioYKCY5Ly
cUnUpTn+sZNeGjR8ORCBaEpt3b5XeMsXw/JxByhSglnIEe6rY2Rgz2YCvPf6sNyNzA274p/c4Q4J
gt27jHifGKOJ+5GOJEk4FFRNF7gacDHHQxLjR+fgCbN9es84m7zmj7CBiNQUPDksqWxi45pMcZKZ
n4tcI2fLUXyUG7VT4KftkLFew5kvVoCcSiq4qXM/+DS3svexESadwZlmrYXd5l2QhY7im0151tXE
6lsOFuEw3MHW6RylSUqqDrFeXobY3d9lAz3Z7muWNTGuzW3e9XdxZYFTdMUycUmO64ud8LAVTbJS
raNi8uSg7cOP4K9SjGosJOxiJ9IgAwdsJ8nbtHfDiScN2H75gaUkN2VNKLsTezWlVT6Y9uc9VgIj
etbaFnDZZB5iHIT57dpXmYYxZ885VcDoVwzKM3ECfqMZaINO3zcl/FCkhguGXJ+90jRT/XI3iGPs
YOwv0G/0FAIOkqnXl0ygWRikKiuQaaJhFv9rc2e6J8c+xZA2vyBwaCUjOfRnNi7MTVfeypQvvlQO
mKi4ycFjRV2lLTX3nso3b6C1v4LB7pDf9eMCnkWqC3QOJu9Cc7QChYZWnDGUGL75gqoNMFD63OH/
fx+hfWuYHbOUBZO120cTEHG2tiETLko9G3hgXZMuabWngiQlBR5HxU26rOF0leFfZnMW8ob6gOnF
ZUooS21n4HSx3SLjW6NPIGemv/xPAdsWLsTheEPKohEooP4ZGKQPUCxt8vRWGemdB74YbihTxov1
ZCtT+jtt9pAVfKdpbAVT+Pgx5oKsGMIQVThM5EOirMbUWqk4lDWPYbKWHonTnYwUw0XFmDtHMGgT
33xJjd+2VsUtfCEcyq1pfFw1+ihAHOG41tigga2+QHWyh4dgG2lmx7EroMQ9Qrb/Jv9KJhsn96Kv
uMpZMuobiAu8pl2se72GuYEQBNOwQLuB6iMt/2IHl79i8pF5StFeblFl6TxX0sFxOO0QuD4tlCBJ
VOe1kkFbM6iAjwWLhFq6X6ND+F1l6b2r1xakuS2MVrET3k6Zq9lZh7mAUl9fa9lHGSLjShYIMQHw
kyHP8lcpDZd6mNg0YS9D7s0nslaIm6KwOp6UugfNEgCABod4SlvyLQrw+HH1C7ozLCY9s06Jg+H4
C9H3t1ZeS/Fp3gsEDQIYiaesulN7qXJKhHBM7wo+u/VzHSqOo2Hvj/9RtkDzWrGjO1L4Py5OYz9A
BcISnB/+Sedu5rkYvnTRwXm4q3rZLuzg5YMhL6hBLk+ns9PSHowqa4ftL+ak+S1Dt1qzIjX0jMy9
J50KZ/XzoN1M4JTQkvX1msXigXFIKlH9bHeFILyW3+lXxGHWQu/f5jr88dirCbYacRRj9JnVQ8rf
IuI/VxHMQLE2iowFtt2uKoSSsBwKSWbl0s2HJO6AIlGoQMgDyqsDjVkHloVgM7hhHyb5caySYxJv
2GudfIssSnpgTTgsMvGsu5cr+RNv5V5QCN40OD+/xVyjXtLeqFF1tElEiHd71snVMazbbWW4cA+n
kkFcwu4cRFYTubbx6cwmSToSBFF0WfbwWmYOGWbZO0dvjnsetFjtkGnksdsl565ATxvbN8+DBiXN
Xaa0xsiRNnvt4IlCqhIEHXFQinwVfENZHTjc1F9xgdVOk8NuQkJdBymIHofGL5XV3mRIsHLSgAmB
Q6OZ5rogIcjgnT51lUhm8/kribwE+ZWxv2xq3yUuVVlSZ/jrdxknwEfo13Ud6ng4BzQ9w6nyBbJW
FRolpo1ailrwR/V2/aQa34skbuH5XrWiqHWXHiNUsRqxPp1FA/xIj0BEIO3LviUWldjWr+llwxXa
UfuFNjvDCEOXsOXrBHwAy1v8Zu8IOFEhX3nm+G1u0tTExl+63ZhaDoQ9DTVGT0TkRstXsLP+auvv
ecg0XUE3hiqAR9vt4ZsmhI0gaIvqgX7ZoL+E2KdwmojcWXbaLKII798NW2exfGkDM/XqNskRr7+u
pwFlKM21QDJVBK+JzGkZsSMc+YmQsqOIGdYWJAo2zg0vFAqSfHmz+/qnsIfdKJ//byaEExF3k2Tn
QBu7JTc3FPdwp/404h0YFkSKI8Ps9Wx+JwyeS95RSR3QOM5TICYZtTgINlBdckIohDjtMV6uAJyQ
PYvkVSCFN2lO4Tz9O5dKBm0Q0uIX9ptRGYdV5L/6UbeHacAQUPvpEUdldwZ372lQ8z1oq599Aftf
VZtBtLCbufluupKfx8yWmY/LxAo3QxckEAOZlZF/RDZTrNqcwisN20C2QpfCgqr+DUyYf3tOaBaK
8iLXfhK4WMqJM0jepkHgpcFA+hb/cZA89zoufSoq4qWCC+qlxaaIW6AsLw2fL26WXg0wOamW51aT
kig1C7bV5cxR/F9fJCkUHU3ss4dJ5bxtnxQCZh1JOFxFfuSh8xT4QGWcivyDmmoWQliTOtB/thBr
vNxxDd2ZswpPMER4X8PdqpR6kP7vjfLPAO8fcsFh87OV+qnIINoNSS40uc3T54yjELQtjigvIZBK
8UEhJVVLaKXkjiXdzrRMpUspSJ1Ne+G4KQRPhXZpVKEcZR6cBqk8JFOjDWei3KSkil3wxs9PBJ5e
EBBdwkohHYXr2EvyuCp+HDJ5TlnTUe8nmDF1SBEuagKng9JqZJ+w2D9CcP6dcY2EbHY36dhiMN+K
KCZCL8uc3F5xgtSxPWNmeQq3r2yL/e6RE5HH3f5igur3BCfnDbpiEePZWsOsYaqEBeEdSHWFEd8Y
fnV6kdC+A6Hayd/KrSqzPZjG1igL6iTl9K14ullyl/J6Z3VrvB+C4fPmXWC+orBjiWRK5qhRUGX/
2HCoN4gA218bU6U2Foo55caMUV4JS32eRvC7Lctoc5g0c0mKmaj+WEY/WXqr1c5IM08+Ysqv2l17
gLRhTMIJfHFR9fx/n/7l07+Yf1amWdlU7xdQUjZR9QZwrwQeXx/iMOsFE6Y+3IWW9bKghA5TNvzV
ov8Bn82u0qgykgIHxMDHUzyUekegcG/T/93d+HfyRJ5HHm2a0susMV10G+dztod2suQc3goK+WEJ
8SDGNs5pz5VwZt15gVQxgb+D5wmSnHrKnttLrzOJ6i4xcuazhg2ahyNVXfuIIOugBQOf2mebR8NT
VeJdECJ8XC8ouVDi1X+gpoZJWMeLN8eo5zRV0UJPrxFok1x6NVoERB2mPwb5TezfE2/9/os9ZEec
RnbgGYYFuEez0U5cNxbyCANQezScJ1dOdQJebhvyFwiH3tEDbfGiGD7j6BiCLXNyDS3S8e7GcV7s
kOeixCOG789aTI36lVXg6W8V+NJfoiyr92a9JM3p25o0ml4RPrknu6nZ77TgJdSraYDyXD+0eTIC
m6lSZJk79ofyWiF6l1TSdhxs5/A0YyOBe7NFxdIt1E5wNUHipHdKn733FDmECWSkSe5nn6Q0DN91
0nRxknnArb75KvB8NIQbAogBgWE+0XpVr/nWp1JsmdJi+ri4uRs44WEuszR7Gul6rRMbGp6Hwrwx
/T6oSDPTEL4BnWfIbYrng8wz1tgXiC+x1/Dmntg4fuSu7O7wvya6tp6lrL+HZjWyAuekhDJMON2D
JbHHypYE5FtOR2kg5sJYdEo8PH5jpB+qkmCHpSZfdYHryAU3eT2GS3MIbthza0y5kZF0iyG42Saz
VqPXtWU227nAQt+pVt7QHLaw2i8k07+ESmRolGmhfnScg4sNKy2OFkC9lgB+EB5IFm+2gHDjF107
FhKJTb0j//QFVPkw/t3dsZW1M7+rAVPu2kqweoQ4ojqmIV7TLLQYZdJ1oomeB8TipTK4Xp6VEA+q
JqFIfTHSDYUvbLgHV1JC2PpHgGZVzxw140WZJqG+yL32YiyK9A06LzJLdkqQj+iB+pUD8uq1fPhp
kct4S2dryJnYDBAZlc4F/Yokl8XM6IKqXxw2Ccjv4fkBmdUIXv7BXu/AFaLBHpSXOA9sUqrOcL4Z
UhZ5vIYvxEP8y+M1rj2sllgzXpgtArHMJUehLSQMskUHtZB8Gwsmqzy8EiCbYk57vaY2Gl5OAb8i
f6CHwMYiAFpmUbCDT/Os7Syp8JqfRhxh6jKjNeGUN1lK7jjvQrwzvVThcS7NvnS4/bTtoH3Nx3lz
esebJ5O4siZ1hPWHBpD7K9JyNoBJWc4Ym6pDIyKPiAeEKrDY+3VGJ2BMtPkV53cSyAREExC2X6/h
hlHSB88H+nl5Lq2Xzgc4DQB+8Z+ZX4GwTQlRku5tw2yRmSTRfjqUp1DxlS0wXZTvZPq/vxZWIBmm
9zjsQeBHdCtgeL1TZZUf01xyYJembSjgNv4WZIchCEgIqdgkz3HhU3QdvIk3Taku3LX4Ybn2u4TA
nWvcy1zRy+nxSGibKr+VVhvzlBpNI7uiyXzVwItkMuczuzGDMBLFy4w/7FXazdt45bnxEEYvmPUJ
C2oSOSR309VnqMNyDyYepPrpXMhwWM4XsHoN0Ep1r0KhCq8Kfe0baHLFUk8qO5VMt1puMBmEAcKr
8KtHwLPncQaTbpO+yX5dUmuiQr9l7ldn8fA2MkDDwX0Dd3Dgodw16IJI2D1SF+Kah4Q1Sqr3DokZ
plxMAVhqtq0c8Ddst7MJDQgB81AzPi0iEl9uR7Bf/Nk3HmHPlis0iG7ZJ2RCrVqqucSn5jAV/Fzw
rlEVZyLx0kN0Va/ElZzIouW2jxjQCHoX/tY2aiC7IeI7YgbqzjSyBfEQx7sF5DW9YhyUxfvFyx4U
rf2U69rY615htQHLxqfh5ILsOTiA0ErFmtyoH/of0nAq7Q8LV3KGSA7ixW76CpvqCXCS43BgPT25
/JNPo34uxe8TZ5uiQrr6YQaBiM+rQxQFInQpMeFCSPf+uaZBlnJOR/UN7ldkuyJxIOoBp89Yjaab
3aJO92/6hfs/duqJbpu73QKBqVeYztHTWke61JYgtK8cNgPxeN6A5uYncT7ZCyFWWSh63dXPzFTu
nLeQZmCHHoGF/nAny9x3GEDUeNsW0tZgqqEtcqwm1dWRFkNZ6dW0wiVTKwXv6cW63h9WirGcU7lC
nltSxYwTQdazq2sUxsp10Xaz6LBqVOV22CKCb6O/4gEefTv96J0bOD4NP7NLQQ64gCFgWTB3xTPS
e0iimA/lo/CZ5BLDfAaEzDbi+9kZtVD9J9yLPrq6Hnmz8OcSwyJyYXDi+5N1+jR6+zO60Vjsjk69
Ta7htT5Xz+6wJdVpMenMi5NvnrCe9lmsNHzwi/dZnbFtJSjfbBwNRGEuUL5JgZaNBEY66D4p0O5h
eq4IXdJyRuyz8Xs+nIjHQBpHJHDw2IggYqbFYVE9eYGZi2ebwBVILdxr4NmoJdYV3hvyN6wegaIQ
Ek/cpdMHfP0Lf3fsD9w5WNQ/YcEvPjJoggrqxdM+p7PNj8bXA/p5vfqufGzwGzQIqCjfh2LKzGtK
1iSnxpnfcIJr40lc1FeDf30Zkh2qBpHTI55nRfI7jlF6qifVqgDOrL4U8xIwarfE/LHLbx/834gW
/AvvIdNnGoXFpMBms68Yqe1utq6CUEaYA+xqmejb8cvy0P9yipSEIieqM4fAo6dPFFdy8Ry4QOiK
1g+guwgMuHc/btbX+jTNxrQC77rJegQm67UAuOaYQNOOI53X4oTqfbgvwj8oAG24xxXysmErwESc
7yGi0zK5wsRBT1q1YWtKEXebCkb3MeGNdfmBnM2bkfq8LAV80L2aE7969j3cwBmVYL19VE00Ivek
3CftcjoJWoZ8ghIzYOS0zvsn0yPGaZNe+gHlZbYeuX+0KQsYocc7b1+cERLHlDyLk9YVqagyDZmk
Bmi5/6J3M6c7EyJsQtEBkyJI41LbfHzmKvLsLYkZFLUTjUjQeocHiNzx6CZ91O1sxsjnmsa4O2cm
4e1jlu8DMhvGNFJRKuJHCKgvycKr9ZPg6yLrZCVfVEhRZMrJGMk78zW2PrqzRS8vjKPYovpz+t7d
flQu3JHg1/PRM0x/Cwb6r4FWPqsr8r/gmtkCvbuY5U9TgS6ZjO1kQAzeRxgochwrcwO4VWXH4Puf
oOQkwxw+Co0R2sdxnG+4sJyNmXvUolTCO+mUtplnlcNzYyPyH6kmdozxe/EW97ftUqOk8OqrwPKM
SDdYskA9MHL9d1Ot6lWHwtelmN2ueIM92qTXgOXialtqmohPC/3+Iy2C6OHjEk3j+rP0b5X1c0fM
gNA5eTpFqocOt+3J/IiEK4Jp0z/glga4qmhMKVHD/6KPnJcJuRl74I3h/CaQFWOrrXkE2c2ckrYW
M+4rCeyOTUs2uhruTno4vFJG+ewOpZIcTMb6xKxqTNMTpY8rQVFGL+G5BKR+94brI3pBgZORBSoc
ZYWtTi1I6oTejB0Yn6t1HvRt0I4yDvFdXOxxl8pvlXLc8G040z5Jh1c2kSaVu/cnEJ5RDEZc8aDV
ssElX+jLPgNxT7aZ68RHcK3hgdgpsF+h7c5bLdz9KQImnSYg5di6/iXZP1TofsIAJxyBP9OB1htp
4y8WMeT4D+FhQVzr5Lz60eWM9uR8ORI5Cdm6iSYawTmufNzZOYd1Ip7Hn4DJrCtST3tz6GOg4S0M
umkbtsmLBFNxDGHkkbwiMEXioMboGiDscNXQ6UeNzn+tMouiqTaUpErj11whKdqGnP+kcCTn7zM7
NcibilNNodtscXN5VHdbJHuqJ4xSiYE6HXOUHmINd1z9DcspTYxuXH7zSdvlk7q3blTVWXLkOGg7
tXjw7InkGeyFr8folWmRhrA0Q7kkFjSDrk50QuefCOBsjGzwMO4dDaPT88NsiCzutgQBcgTaSvl2
xcXUX9g93+ncN5XvG4RIvXZTo+aH6akGM/xDpFzhT6Wpa2YIWmlHinQZlEOLml/MiSTQjQe1kEnz
Dlm25aIjh1yFeRW/AsOfacFqptoSose6bSHkcNoqErz1aGQ0piTXTgdPtjOR4RDIYLzJ6R7BJO1P
mRWUnCGDj6Y+RJPe7Lk1ttz7mphl9wbMgM2xuIzOXzEOxh69kKNRoyyiN16jW+k5663zQSNQ63Dj
QboEMGPPlvp7a0u4LgrKx9DQLobDWpK/jnEBJieUgpPLYhdbiRtC8Q7OhI1+bfJ6EJBzuc8ukrK8
I/nZVUSMl7D9v0iigorEOWfsxQ8y2WtQueddD/4xK1ItRDGU7BUnoseaeB/DD4EwdAW5xpk9ReRj
s0ZjjmtE12nY/FJco1jZL3ndyzE9dXDxgVckPBD0d2w3fEtruL6aEjNkZLoaCMoI6N2Vdn8seeLV
u42cusMBtzOhn1pjVb9cRlT9xnhp90EvUMyg7w+/shapsNhLxRcwcryjPm65HXkba5JGNd/T2NYe
YyVDAmVW1MmmE9fcNp5/AEm8/fKawlNX3JbMidpfRJ/IdqB0pPKG2udU5fN1USRF+w6U66pszCPy
z07jIXlde6rDNznZqH9SBkmP77MI4xY9HY1RKkc+IGZsNOSqhiQgkDbtIbLeU11IhJGJCGZwPGSs
kDBh3bHkBmAaHOXWdvMxrZ4or9M8NqS6fKWIwLOWc5WpcKYp7evCPsplamVEHMCU47PT/Ib1sCBQ
O/BXk56xLyK60WVqlOhf1N27ORiQ+sCBMyyufZ8GEe/QnhNWhAk6RPgAlXDYkQyKK/hGV/MOKjpk
VRQc0dG3FkIlH03cBVjBHQV39ANpICNs62RJE3krHPu+rWL/GQoKvECwI58okKyaJ3Qlz09i3M3o
CJ+8+c6IT9Nm2BSH1Loj1r3F8LZFwCaW1DMEwJdvElmmpWgvCbqa45nPpsyJXhypqZrbx3ydvo2M
84HoYR7Iwwhahio7BxvAbisG9mBuwt16yohEfRurGXcgbB3Htf5zKTHhDVZ++qEWOQ7b4jxoNBME
eDrSNWcnC3BccF8nptpqt6Nv1uFHO+Gb+kBf4dySwwiEzpy/Mf+zHqp6i8eS1jXMsg2mjyNwCN0N
o/LZgDOB4uWIQq5PukXFPbDMZQ63ezJ8iftzuVhTd1k0YBlBRfOQchyFNzK2MArr2FhJd5XCITSV
1STzHRKO+M8x5UTfgUelGvWbBaAcTeQZQmf5EIentvduaPAqkdPSw7792n1IakwlYYt8O6jXV0hq
vwxbsyL9+GimU5AnO9Z4Un2kDbxt/JWb/nPCSSAt9xL5nlx3OKVvdTR4V4pev6YCD3WBqGL9KBmp
/4s0uPDcfK5vPoXCYlM+C5SlkKNbE0hrpr8IMjXyojqo3/v+S5+nATsgK0sm6XzY0S3FB8VnPQ8p
E53PpjYsHV19PAzryc+Jbt2+nKBoZbbbMfOW+1szKtKH0yhDd8x1OKs0yv8270kvCqForxxaj4jx
nFmaE31TeNMWPNhAwTyb4B6+nsgbLtbiY9bBn3ZoZ5bV1sR09qqkj5sJia361DxDi2TMs5366i01
8h0kLsOh97ycEZJsz+BT7fY2vaiXjxyx0SS5rXmBhXK7QZycGQVxZiBRaND5/ZZ1REhSOOnJZm44
RAqATOGEPDW/3E3XJ7GJDrCkQaAlesrtDSISiiMINDP1StpaRaJFqBe/j9tfawudEMObkAXvkj8z
qM38fLo0UKATm9C8Lo3xKWxh5ZCBkV2su6pSqO24ShkqN8UGQqaRTkzdahmxAxFvH6Nnmi93V1rb
PnVdWj1gp1ZNdbymwVAecFiYG4nbTesoEq9qiXDFsnDHvtqRXwP9qIJ2yiT6Rhymcijx97f4c1S+
FGuPj/UNDlEwxtYRAM4LOQQCr1+42CHtqraPw8oyli+4f7n4AKk49wPvVANk7IelgbTlVaFp8mWP
LwmrPOvQnp+5A+D+txIwW3yXTfwsCoD2UkDrZoLqhO3psepmjQN5OvgvMqeIzBNzxLnwK7I+pwqs
q0syr53TRNLUEo80ElRQwW1Dd87wsgd5RoX5VNHHH3RsZduUSxH/i8au9nSyulnUmNCYygm1h7fQ
sFOST06XVNbdauuqGSOcDHOu8IIz+7ZJHn1gQhWLDmAdEIxKUqCKodK9Swv8n1Xi/DZvenlgqR54
RIfl737Z4pLmE4Lk21DJGXrprFkcMXAp/OaEIqNHH0eHigV89oC8kJu3pq94hstMV6cZjBB3rG+9
kVQ1T/+Vtyx7x7pi6eehXk3yn6In0auCluCqhMVCD8x6TjF842/2nGObUZ4xhx+LQTXWqObRSd7z
/NudRbTmGhVjsH8AhmhfqsjZQTHr76gP8KMyNFoyEAozgap5X+az/4xn+kIzrd+QRP6vnZrX/XdQ
F5qSzLxRBL26ufiPYqVPAcdQCAXGVChsWF9KxAx/hsDRsRqzztfASqzPXHtenDcAq+s7Lcj2GZ1E
GeL0mgE4L4Wgry3dkpzDaCmVSbO8KdfCz6uv3IlVXPx150S/JEBRqSSJMm3mmk0sXFgL1Z+v4Klm
i+kB0qGuE7oS0PkQ+Vhyl//qHshQr8jubVQl84eXvWNSyGYhvlRkx9yYidgTCCICHgPi8cTroGIp
Aq9hV8dciUc6LwuD4rRsj8Kxf4r4VhZ6VZxZUGS9lZ6AaIKKML6jIZpip9vLY52jUPgA/Ge+W60X
GbhIKdkWH7TkcWHdSsjUvExCa/thx7a9BCkwjj52MLTMRDxgNfnpmyGwC9CQk3JC+k35x2rEhWJl
FtuIoyWaOjnQZW6JcRUQnoABn7yf+OKGMPlSzLjrvBytbt7/3DUiZrrOQZJn6BRrumxGjuyxSGrx
l2WLFF7KRT7s60q1pif2NAGRKTFgvWyLGnYn7POXbHVDHjFGJ809CsxOz8VMj9B2DGe+kfYgjuD+
3eXhbji+f2zmD5IND/Gyxtu7ZG0VBDh0wpaEV/zjsdRXJ//AQSiQVFwvIc2a/2RObvZ9zxjAZij/
JHHmhgBwnY+AP6zqXy9BJ7QwX7yTx1Ni0w+6n8AcWlbYhjOUNcux/bpbsiuV+HgvMHw16krDp7qj
SXA849HMxh8PuU9q/5lCmxjIQpjEI2gmPgBdxxyAP4sNSJ7bOr8cm1SQ5f3fs8ii33eDpgPYbf0c
vnBY9rPAixSDxiRNq93i9U3SD3CODBFrIPYOriU3XLpPMyXg/1r7WRkcyZuvOvHzCn7dkJcmzbT/
Kuh+g6q6fOLZRpyfJXV1vV/8AK8ovEn0mlMCbigBwn4NLrrbqeHN18JgwH9rVFB3rwbIb8N+wNKq
MRyrZnBlwamwPUYdGkQqC6XeQIz2BLye2uk96JR/71rRdUOS58bweuSox3zxEvF+Pcz5RK3Hz/Xa
XrWZT+XVR55LaPwcprSZNSKRK7Y5ZMMRVLcpgiKazPdzm1f72/dnJRsJVyregjEZt4m3KyK3HYDQ
sD9MPg7pEGy8IZ3EpaPRh2OWt/qyORx4eJ5nktxpw3iQepWkLuvJtH+9bIO5qtsoUksB/vNC9ak8
gXXxIcHDz5v1jZqo8yq2fCqAneCQMoX/57l64Dylow4yVcB7YHzm+86hGilI3eWqsPyKUc+AZEyP
aLAgg+FEY8yxAu120HuCw9BMrPKY90cJVNgnHJP5fg5IlhvyRxM9jR3yg4U8azZHeGZyngz3s4zg
smJtnL5hDPS96z9jUmm0UwbHC6MicCy92gGmAJZ2C8xXbXs6ZVwSvouPu7bENhaGXo1eCSJsg2mv
YwXPqO0XC3HMdvs+pW1uBjfYHZ8NlT3iJ1EW/+wl5bNV9Rnt2reKjHbVSJHyzMm0sWwujhrisblB
KL0acZsQ+dD0X8KIkMADcJFt+0RfjCDswIgBXtaHaLyT9SWrAaOyh73yiAg2T0yVLVKGArVM3uX8
JQxtcjI/uXzF4tkIbYH56u4B6QWT4ALsQun1j8uc1u7WWwsuR/6Tennif5SYtlKC6C7BTaCwXTE4
m8popK40g+MK6iFRExs15CO+fxcMnB7m7oqewM2hdm3VW9otNn7CtsF+6dH1ck7oxmmODyB9cAI/
P3aoDe8Hn0xuaBKoksKxJEvFUk34vrx+/Wp336zdNF/b9tcGNx3ooWhFmt7oyZCLJYG1TNZUYzNC
3Exa5TpDjMXmf4q7OCW2l3/iaG7KSByhrZpILZsxNkcjs0sCd8zAVnvhwrM1D5uCa2va4aMUXLwO
Tr3RlFU976OKvtRv+OhHdBL5ufy8Ya78cnoB7V/jUqpxN+yZRFnca8ftiZq2F/ByNmftfTv1YSgZ
4y5+wV6Wv7TJnjV4JKmPwaqjPMSiOTXLP2ceW+3Bs+ID32w3dFB9lmFCvYC1ObP9B7jklXhwCF8T
P+W8CmtXH/s+Ymd+3FOhjy0UnBt2FnbHVPnW7nfTTHTQcxF096z0/wlwQ1+8HjOuIkoVjodmGX2P
AaoffxsTJQEGMwrhkkD4Ii3YorYOWLXj0bBE3sdUbOAlXXjdIOvWYNiBb0/QbRWJ7/REUmrCmi3M
25JldotRkUZn1/sjboMY33epX3XXgcnz4BF6JEiAwPUcYF+1yZKkBnlG+4iXPpFJHzF7YaBQKA2b
6jk1bKwHaF5hIvVGZcaaRZjLpL3OcdpcnBc3rTzWRqJQuhxUmvLdlFa0U0iFmcd9m2kYNVd8+rx+
B1jSEkMytV3ME7B+57T0oOAbOsx1A06r9nO3xRyJECdCGrQXDN3RDl38S4knw2+rBYG2vXJDu93i
jc5dWs5ODX/4zIeCc1Z3lPe89IvWZRbpsC/gvsvjhGI2HYvg5lQxc7QeDI/FklqBdUcIA+OxaaNQ
A7OB77gfllFC+3KT7Tg4OXdzgvGEg0Z9eKWJ3SN0F45SLqIEP4qtDFO4LSaB2xd+3owHmJryYBUF
VWIFp2FQlunS/bTn5oRg8Nt2rvbTx7++6pmQ5fb4TKKbssLS9Z1Lxxgc5FA7AZtphWJ2zBTonitc
vB5EanhnCJy//Z0aTiRIxOANlkAT1HnwEac+bal6BPY2xX61x7lQpYJhebmZm5QfDodRk+Bq/ZKX
VKhj4F4eWZ53tRWoenmHd4HhTawbkaTm55I14IEdinEjNflPgMnuqsy46aT+8HgtpX3lsAjJIC7O
BnqCgHEV4C+z3b3dUiOM2ONCY/5ML4iP3IiWwO2sotz2NwpPvv23Y5ta82NR1nd1TZIL0J9u5we2
qVaHa0lSv/abwK8a6betPor5ie5C/8jCHYqFp2kXlShb9jxQ7ACbgzBcUnWb2Jp45NFD0/86t6WR
vNtWLp+6nHBBo7AJi6jbSQMUkE30mRIFx7KKxpl0Ksr1PMPrzfhu3cHNwG7jsPPQ7K+wltegi0IO
rfuVs9WQPoO8w9dO0H6RApejskgmIVIQJ0+B44xPIuSkikvpgqVGgjIwsm+tdPJOpX+daH83dRWN
AvWs5fll7W/xd6VLO+PnyoEEO2xCnsbF44GfzZF3lvRVqTSOOFsyM6cnl8bxHUvAn+4Zy9YeOolC
zuddZdlewqnHz3B9/bxeH+AUSX1Y/h0ZWZcEVuR+PyNy0teVa0sdYLSJ+LFGjAgE2OqB6lBkGdkX
RqOEkeb4T1BmtchtrP42Q9NJp8GtX/hABE16+bZgbSvYeJ/7uMe3FD3gcc0yJOhAmbLaZxF9VwUw
1JvVa4DDKKz00y7lnt4peP9ZV7rB2Y9NmtO7T+HaxppJrt5p0v3WCUqbNziBr7OFhmcErg0PJLP6
aWt6LtpX7M60cbT71cYWPZ60v1eMeG1MGqLtGSn6uluKAfTncXukp35XLtmOyxFrErH6ccZ4h215
vCjj6CmSZdUMqsQQJXA21+wJ897YyA+tgoZR7UHHya7/0WEODkRe5Vi+/mgjmLRypR6bZgn2//kb
bWrzc6/6A/kPOIo+rYTCEnEnsUjWZWuPP1pl3Iiwole6PTj/3JqNSvaKwnaDEo3XbxEX8CGkacSh
I4EYrj1ig+jT8Xqizjn45vY8IIubjQ9YhoN5WEX+YNgkB8R3NceuxXuprMj9rVZzw1tW/G/y3plS
o0Y9cvI3uGHdmnI1KRQOFGtGidOHUdo31DV1SW66XldVNwmIYZ0+sbarxBt04JKrItX33qALSbLn
t5z1j4jalyfzJLrKtaJtB4iNAeos7pkBGeloIpH0BHIcxPpDq6ALrDkVRieOr055kwaBWSKpbLZp
UsnD6Jc+rbzFEFbZmssbPUn4SdJPIZY/y9nP7VXevytLz8r1JZqjqySpYccEcBj5KtJEVLXS4WJm
nvZk7OtYy6on0aB8KOY2ogygew8W7SMs33ChilUL4dJAJc10tDELDhaqhvUC2SamdOc0yxuw2XT7
Is3M+pD2VVghECC6mGRhmaGxeogIREolcBYvRBuVzpk39zymeRI9tSpNVz8cWEFsVUjeDPYbSb65
u0bTIZy5r2n9WOwErW9/OyEBd+xpfLIpouOCDlU3kKYuIK/2+eF/aWGJ3kNjbAiBeQC5j7ROF/tq
vVhLGowdqGmAGZXRBTIr+RFcOdu1fIrrJONteYC0anGwzQ6u/WdjMO/Vl2E/S/JSX5B75MT3a/oi
No5V440o+CxBYR6eI8TwCSOrK0QaXuK1sYQazbLUozZR9o8sCmG641OyuARmbhGBMIDDmEvwsDCr
rIDsh0k29NHX7U48P0U8CReDHOQH/HlFYFz77JvpWHIrKasQWuYboSzn4nSTLLmjOPMohPdhha+e
xLWSCcLNLDVRFU/3m/5ZBuXFOu8q1fQ4RTZeQt82CgT3Mbn7Lqb6XEXrNZ3ZKK/L8s6Ll5b1Pyph
djiCPXU4SCGBIWAY8YwQSlrQwUWBZFuUMTvDvvD7MjI6rnGjm+HcHrffgK+K+At3LLUmXOHIMapr
RHK/dlHKyOTQtOWpikL3AZGi+rnVfcpqiNTMoEIPZTIIxMAHco2+dzzEVve2wPc94Kfcpi0qNJGC
+WyuZzwoPfEmAmve9TVinfeWy4Qxj9rvKmyhnytqYat7QBlYTS5e3hQJ5Ab9Gq5WGxE8Fo7BboQH
WJ5+fjN7EBXbBI5FJNIBQPx721LIYLjMvrt47nmUzJpy3qwvtbkKw8WlLssW78eYzHN3i8Cu5dS/
roaTLcmkyPq/f4yZpoIqBKg3AKU8fDCaQsnt6eveUZyhy5uhhUoA59L4K9vJDLjBk1EykBvjjJyD
nVy6X2QGkRY9Vocvqj0h/ySe3GFgUZqS57zZYH8zBdljO2wNXF0fOXYAJEQjFZNhfY+VOVgbw4bb
0TR/JDS0YGUMTyXLLurfs+esltLObHgI7asuzrDfNLphZ77qaSfI5Nx2KrFc5mfUk3LlZ5EgnqCk
DAiBeYTP1x+irap1fM3gndX8DaDzYMf1PWCJ0ViYzhZ8Pg4nhWKaC+I0pqnIfWZMSkxciROpMxrr
1qEzgn5K1o24ddGhQkzBzdQXcShPi/izm9X7ibJmLRln1248vdFjeo6i8viSOAM7qoi3leGGUC7M
QrKhYlqrTG1eKNgvlTtpg98Amw7aXip/AAtQ0bgSM5pKF7dQGLLawdfBzOwkOA5AYEBXCERVhKUR
AjoyaW1hnnW1yYyEPH/lq42ShZ6Dqp8Mm5TEM4ItnwJ8ffV2X8Z+1ax92FiV0pnAum0zA6iUq6ir
/jrI7yIiw8IK8GTzzLlaCkaWXpA6Inwmy7LJuS9Xp+IfOBc0S68q9zSYyyiB8snbw8untQKLx7lN
X/gL9Ndes41PIh79nRRd3myPVqNMGNyrMxHM9qqiumsdQ2xwkt1T00c1EhT1YXMkBaKR1aB3/WaC
QM9fJe2LhO88n2g2jBf9F1Vl8fe3Qnd5dzdW9DK+BhGLmtc15qNIl8VmRI/r9yNalAPS/2qZhRgt
u3gMJYBty/vrzVKFYnNMz2yRarErvpvERmgzrIBvfue/KyUsxTUO+pRoGRYgzoj6g/1WFoD8TbLJ
YjYVljysF4xUflydZPtkqZKsgFHOfKIdjuI+BF0V/zp8wKvFOZhyD8mP8S9s5gcWqbMVGygleMRn
6c7AH0dLwfjw/I4AQwPN3vGOMRXhQUSn+K3fNr3zWcuzK5VacjK86e5vbSDnoStyn1G0xmJtsbaS
IfcO5LY8ok9vZD72pZpdc7aw8A80dDaHqb+1Hv9msOSgyZzHuOjflVcE72S/8KPgbm9l/VWqPagU
AbJsw1JgRv4MxsxMc5t4TUWvA4+Cbz5z8NqnG9rYw6447hSLeD0TuTbwjytNCWfQFpQo6dYbVi0O
kYh2a6WcA/ld5p66Xs4WYfuYL5t42e4nCx8kpezDOYX2aujYrDXBQe6e/DaVmi2F5Ncox/LtMRcC
rgg3Qvhgc22STjdGDI707anRhm2NTJGGn3Wb2TR9XE29Gq9i+Gcc6xMmVS1HhePb6mfubdFPuilO
Kd01b4GkczKq4aJzcQFaFREvtLR24Qcs0kKVXDA5Gxt6l3sSYB39xmgK2eak7Rde3AAe5io3euQS
/EynLTY4Tj0QNQ60P+ymkawzpSOfGz7kbJImn2MMrqMUmvTyuk6ACwgdllXub0YA6rezK+fAvNMo
mSiEwzWdzcvCzCm+J7NyaT1bbiyvu2QLOnygaw9gYrvJpso3ICa6Q+Kt54p0wc2/ov5+rFIxLoNW
3hhs4sjx4i5ITaRdmTUZCyU4aHy9YIXN2ILsdokZice354umWhCoMjLdCQHucxbn8ZTF+6dX7nrf
aNaKIiksV4wjf77HgESLzUUnGLRnKdpLnbHDduEAO9Yc18TcHETzESeLK1v/fDOfGDsLaxtsry7e
3w8VoIpvjpztU4aqW+euDWJFQt64jRmZ4CqdcJ6Us4mz4zoBXJ1+qiaxaz2UZZMvGRFmrE3jV7fP
WJyBMpxKJoBvo3tK/qiUWMsN81B4YoLhzUsdftupzGBJGsAheja/CWQ+xaw7+fwDxeDewt1KJNVq
/BynS2RoUDWJ4OJq6ZQc4//yQJohqJWe2H78zGsvqlzU4TcV6qF7t6eRNoOVXCZXsts4X/Muto6P
H3A+YqT/k+L7fhPHEy/cO5xqtNG5DSL9eFSFFOe3LKI6u+Xqm4VQrzrE8Fi6VjPA/YMM/VbglC9Y
e5HEqvowb93apJQvV4+VX+gQ7WqjzBUxI4/cdgC9OPuMc3RtKPtTccHp3A+/NuZfGYwL63YTq8un
6WAuuvRaBL7aL+tz6gc80zh78pF3mAA+O/11gtKL9aQvgKtb0H2riRYI4oS/GnQ7p4p9fsgKnI3T
XQVQDCKvKWcXR3NWH8gcwQRaevdWNnxsecrGVfkJlNK2hWCHYDCbWXkw4dBotdHhQlX6+Sq+feqF
Y/rzk8aKfzBHE5fIifbITW/cY/li0IGuYPCgiibgizBlnXW+j7z8ulwRoDNOitHXZ+QIAtrOv0zV
k2r0uRePS/BLa1EE6kHz7fD7/4e6aGYcglJWqrwl6f+cFvi9qG//iOQjHjYDtctpMYP8DiUk2qCV
IB4V2yYFO/KZWvVQXXY2yU20yjJtOaee4F8z8mvyHtUrJfW9TXB+cRdjusqHsTJUH+PAyailkEuJ
+JYWvxnBGEdJtSBzuE8bwt9fIuqMc8n3mwIzlXruo8PqzmTFnDJGYHjhWEOvvMgfB9tR6IClBT8l
t3gVBmUtaRZSaU+XJTVlR8oid7kc6LFTf3dE+TS/4TwlZaQsBfX+akjHGWcWV3n1KidY8r0uwZ5n
SYnHW/u8LQvb0HkbQ9oWQSuKBz3+zvbLlihAZMSVLPqeWrYhitmj+eDYyVimVxWfb17+js/Ha9i9
9PUKfNNVMvJwzx4JSJ0NZbAl6bmT00Qxl1pLz6Z/JGsX8AjGoNnsGLXgJsSMDu0qbsVuy060pfhp
NUG4yVC4Atw87KMsQZwNWdzW11HQ3KdJmsrBuPHLSd8Ojk5X5jf1phcT4gMRt0mSIUAhT0NyhXlb
b3Y7j+kCsVAApzq6WCbvXPvWUOV88C3rLcbNYvWdY2sIGVcv8Ot1NTjLhI3gB1jS5Zr4357Opi+d
0SrAfLYMAubfNu4NvVoeyINgJznTSTniGnsqpSX0ZYViZJUWISlHqbf44fiyNohluXwfB3HH0Raz
b80T8XnhrF/LfOtEcql21fL5K76Epb3TleyBZhqYEF6wFBJgXF/6+5u9oZOYksQlxBOjrC8hCCjf
f98a9g3rAeDAUFOv6/6YB5ShAbejhcxcp8FDXALhFPgvyevykZJQ9tOLUvVfyowFRuxj2yYaO1IL
OU4VlLDQpmTXGRDcTd+DsHpvZON7OgD9NeI43OLVqRrW6eEzZj+Rg5niGmJyRnWCi6dIMjgDEhmi
FknR3jimJJrzRAN5PIKnLe3VxoqurwvXbOyVhnLjar1YusqfDSbyfyCCMsISUo7+8VMnSDOzOSKf
6N+tKedt0PRVQWhaDGrNJIm9U6EzZt7Mqnc+ix8kn2BSztUGO3yFlSa/oNdt+wj94tyORTAYxVH3
pLwwxZl7dKNih29G0cYywocFhO33QH+kZE8pXE+Z0SXYnjB4WJP7XBjwgggj/IkLxPpgaWI9j/kS
chUbB7T3NopRv70P+Q3Jid5Qa/JwIxd9Ne8Md+bC9Xc7fiW2/X20DufSUc2RZaryCX9wyg1yYwyW
DOtS3tMaRr8lXkjC9GR5l0M0c+emtaB5fP4HeHM9ndL9XehpaA2XA0ckD1xynXTZmWyKy4aeo3z2
k1WGxqfAUnaHlSxdxgNbFMeNRYBL3Xi0osf1fkVcmlEAQiuCQNyyJO1Airs7BUpF+yOAFdPZjRUO
XAIxRYf7epZwr8rKXvz3IOPWGeAEuP2oLIekm5c5DtU81Xkm2DFzr8c0cF9jsihXUfKMNS8ljFnN
wqa0vTZPIOOszvTvcFOiwMTU2dq4dK/ZcDpKHo7hTsOL8x/zG5h6KOsBk2iw+KVgf17wRyZnuGJ/
JvE2QutOuyjTnCNy3ZtYsc6s+4dC2uhDjU9XMlESHjTmuNemQ+JhAXP5KLfPs/byeLrnmbXUUdQb
3eX1VpXIENRoVlPu7hG1lPjZPYzBHS6YuKFN3wIeAE7m6WdPWHQlNwpOLGH/3Ibs89ybKl9jAmxF
I1eowCsboWp58HFJsJe5/VdjNQLOqS+AaoqTnrF85nZZGcy0lwc/nWTelWfCbEeIUR42RduUstLS
WszVVK87e66mNmATaj21S0Srkg1qE0OvftFn3kTuGuHSz8zOLzq46YoLnU1609/Ybs0qnYOOUHs9
b3n1SKV2bKayGNnVjONIEgkh1tOkJTg9FJUR9RnJgdy31aR/fmGqjKfP43wclmOd5AuFbjfn3Fnu
wkuVVd4YDSlyoWLXLq5kZ6XbK6efSnWKrpKZXM8gHS+BRulaw5u61+32QuT+m3wdu1PYsoN1whhA
RHjrTYdGohAeEf7htQBSUmQSa7f65YeKKCLPbXc3PPGsiURp5zgKRNsPGER7WQzGEybToJmk1JrJ
RVsbagvm0f+XPeTlJKQrzBT7Cbk5g2MmOmirFnWMJZrmekx/JXIPd9GRX7shgOSFm+jhLByOA6iF
HQgtSfhU2m/Hi24AG+jwfzW/DnxwUmkLgLyI7Xcib1xUHjPoezIdVjt/gV/z15A0OJdYrvs81SZh
lzwKZ58YuOnNQXlxiYEbqhVgoTC9TNrREOvVwxBupnky0whmAmfFwLFNyUsUxLvTYwxU8Ya/aseB
l4tQgaEhJUTBL6aoPlW0ioZMOsCZThG+9ym5REQAfQMgJw9TgQ/RIvJ8cROWGgtaHN1nwcbgU9+x
37601ORdFBnkXfhX46x1hERwIyc2AGPgZ7BetazGAiUX9X6DI9BoxzIfp2bY9vLRtN5c24nGTdRb
lS9bnPBqUtK30LuGAxqdapGhqbtKvPQbEJEUq2NbrtTg0yBqZ3BSwbFWZAWiiiH7r4qZMV6P8KAO
N/+7Nz3QPXrqsvtNxnFZ2MNCj+HJ6BhSLI+cukMxuloTHAbPW2yWE8nJJCLUw5822rUXBFEewVno
/ZHGWmJR/YD6+nU4bwNMbWJVE2/M8MhlWIYfCWNSo4zLRTG+fX5SBRFd3s0ynPDwnvz890ltqkkf
8m9G5OTwEpZqmby2T3H5FtQcAMZHDcokSrky06SUH/cnAZ3FnHAnD2QEVJ8SSYFTVVXS0ZP9A4Oy
lO8+voNvo3Vkw8FX4NKGL5iOWH3tf2mnTjj67IUHzQ4rR7bM4ZjEfiq4c/CK2iZJIW8m/SVi7Klh
qOx2ToAqA2/cFr4XlUa1+oNOcKiGpb2VdyqAssln6GPQaogdUshRNH/HD4GuifS19hDxuIQp5WVg
n6NWn+UlR+kwnsJKYBG5Nd7kTaSYvF2deqc+Y26egfZ24mK1eqidqxKLRquFh3CyIzjJXgcOHiDB
PsAwlGBlsPAwnFWcio2squ7Y9TIbhyDIji97M4BW8hPwwLN3iLRADV9YnYepbjDiJXmHHNSwVVO8
AJKw2SqxEHTYlEScRuITN36oqJIHrvvS0a1cQJP2u0YscYkDOV/jGxpJ7QjcoKU8OwwffYzZpXln
9G9EjlwUwo7zD7+LEqp8tog4rmgUM/bO6F2kbEryOoa1XzYRUEqCyHtbO9rIPCJsI78+8XMGSY7c
3K1GCBJ4m9ERwu1fq8TWGRr2z2SduqZPMI0iT++IONuTrQ28yMvUBgbuNnaurMF6qDLLc7ErJaTX
K6ra/tlufqzNPnkqo1LxWqhz7LCWCCUwibplhpcOzRCZZ2OgvW/cjXqmVdJRImxkaHZHaB9fUua8
BQcDLifp00crBJypTay6Q7AI2FpdJOC//RYRPBAZHkDYBk0R5J0mFLz3+B22q43Cz/VUM2BMqsnU
ykRAGqYFehAwFe9mjbCHFejVSJy17bVn3BV1w2dou4oCq538m2y/LAn6chBqlD7o3WALv4lf4Odc
x3gLd20HCUBHeXbAGZ5Pv7IiEWaQXqfu08FVOzrC7gpQ3r50mOFzlBlqy9Zg6Hom3n14NXRANsqE
AWWKtR1Ghn15iT+Sg8e3D3nUG7VOLnRDwaz2GB3q6OTZEt7Xga8rYhEUSEAygNZp4kddDrrnfMxL
b0e1QalW8bzDJQgrnf8/NUEWPV23HN3K7n7AJ4O89WC9A6C1+d+rdc22Ev62hc7xAbcWTSkoE9Nb
n+Wim/DV3Gf6skpPZP2hUxxB4T5OzZhmG3Nag9jlmwZWPbJDgYyMCZCxepHyj/Xll6/9a4JRgrzC
jgtCY8Y7jQrC1K9xVH7Tm+m4+bKT61/mvb5R861mBETduA17nK1Hja5OIv8osCyLiGywKOEK2Cx6
n2qsFyaknJ1j3LRKkZsxCyzhtQQacVt+x+pTicVa35Z/IomFFRUuKJjpC9YpzsPTMXsxoaW6EuF9
2wWh4fNXYTLXIIyInzkRmIicRgHINVEi5H6RY2q+Bs7fF0WjXvLaPEsHte3BFHZtw4g7afxd4Tyt
grYgATkqUEnZIiMwq80WNjNrFcSEzJSm5EQlSa6XvprzizgNZI0QJfrOTMJx1T94TUrSuxItwHwM
PDrqMsHPEiko3Y9nn9nWJijn25JaWLJyqhYlvNVgcQdSO8A2Y6Pkw4tX0GrXgbTxwqUX/ziqC8WL
NpFXEakq0ViX0wWnSiTYNFyw/Cq9+Eb8gkC3mpAdIJrYaGIx0wWraU0h9BteaGkr10t+MZ95ntEx
pRwyGGKkIPpNATks+dX1kXuDTjOWVWhxsQVYwXkuMnAJizvtoNyRVjGqwQ4Yiqe3lsgnvM6swiBS
5wS3+P1UM1hL3cQ3XUvnbU8kqsPEOOpqohExUnWz4JwWWNPcbPAvCuzJy9uZcTj80hZZ6dTcmWLf
vfTObIrbefsNRs1N1FDpexJdbgCChTOlckYaF8H3q79jX+8cAYXz5Vvv7CHBXp2moLd4FjgiR9KC
A2TqCIOXu8v5bKetnNa6gvCkZ0ZatxuLM8yY4Fnu60jO2yps2XoOE0qWo7JL+Qi7ZWWr+vSr3nM7
22XhwqWR6SSVVAmNBJJpXGpjj2WRFkUqQKog6L1JrjdO6fk9c0I8/rq7vgJlsUeC1bI20NO8YygK
yaK0mQc/d8ZniJ3Jv1nZpFiSOu2wVpUX2oQEXA3byj0LihwzcOLhe7E6uRtUJYp2HzW+i8R+NUWM
riMdlm1MR8Xwjcz19FAsH3IDYO8Xd6oegrtNsDSImkqRxNQJDHINtg14Re45KLROSoGLoYgx7IQt
Vm7aJyHm6JxsRvUBlscfls1hIjv0e93imNPCYiOPQ+OktxPq+hdylLJYf/sqpxPK48K3mVU5VsMj
CEm455Fknl5Q77I4oi1hjSH2r6Ye0vzh+OqhLVaxagM7omOu7oGJhLhhpZFG6hXEwIbABr2LyVxZ
o0X0db6pU+6tFL8KZE/CY0Q5tU4KJu9y0H3lfZJ90EXt62Ik7TAV5TSn0mmcGIkgL7eluJwPB2rR
VqE39nvsdJ7c5eI04XRQfcKwOzxluRX2m22zDBjugzj1iFd232hc6IHYnM8uBCBIRPt31Saxv4QI
O+zfQnLi/NinPKG5K6oY0U9p7wOw61/fQ/7CFeP5fMz1ZfS9FzE8MOXEIQha0tBh8cxv+mAj4P2o
2u+1v92qHeMi+70QXdxeu0M0/kQMaG4leunK1bf8vW0Sh6gQ+P/EQBkUsx//9eDIQeFuaL3opmNd
ScUjNptLzbcr/Z935VzISy69R+TiFrOX1ZwiqZ5wlRJOVDvuE5bCuyUe011arVfAlyN0KDQPlK+S
SHKzinxJw1gSi+g10+PBxoPFFO1lqqEaKBhUkCAXxJf/Z92kxQzTpIQ9TPFr+ES26z59n1liRiMQ
fdjETUtTe7TNYrXqDGkykV79zpZ7ibsP6YQoocldClxKTzWf40sf+0rHd/4ITLQy+/A6mkCU3ZZG
c9s+eIFf27xXKdlxApLeuuZAMsvlgRCgQLSDSKunlZdR9SGJ1LjgvAP6S/ueGCCqrica7Sap5Zwe
B2oVd3tU7NB/QUaydqnvg17hgspDXcgktx9a3aJvG2pRInoESZHKhOKWZarEeTcTKBKwayUJGwCC
pH/cOii/OfBj//9m7AFGXEGxEjolU5dEvDnF+b78mhCK+P7aoIVedSZhtgDrWs31imQ90h81543M
YIpjN8zFTYnGDWSxXHuZqWDGFWJfzcjSGON0D1F+bH/ZUdtUJdYC161NWr983ut2UmsvTeIOTksY
o+/Dl2DopxrLTxCMs4pgLoOiq4zbXg1dCpetvz0GrzRV36mlz/b522Ht/1A+q7X5AH1tWuQrQKYQ
0L8zobZgsDSJQKdY4RTxnjSRRPfn6+dey7xqpHxlHHAhH31QuZiYl+0sIn/G4BHc0GSdX08w4Uw6
m2SiCXskQBSEX9gaZsq9nF6nn5OBcX3jjiEnzfcMlCzTP+hW/DKh1gxxhvXfV3FAC+6YuE6CYmzx
G8dOazDe8RurV6X3ein0C83odHFVuY2inPCxLJfQ8v3K1h8lGv0L8ttT3QTctQGbPuzLrhQIjof4
+AoMAEhn4E4VPnVUhSgLnpotapH8TzNfGZwJTkHwRv5iGdiwEE0s9N9MYjSqIjzM9Ne2n3nva1xl
AeNi/ZdsE6RLmNgU38hyxTF/ct2qm6uddQeTQvdzayVipJnf7bwgDZ83+52M9Le5s9V3/RLk8Orr
DXp6V8zCMTv5kSuvH3/n29E+k5F4PNyKSBLmoMcz5S56RcseCS4aKRlnEDr/KkI+W+qk4nMFsSvp
k6Qqj9SrwnfzKcVsrfJzq1K9cF8QoxwoVzti0PhqadDH6UAayuqAfxUenrUeWxCegw+tA+tQDKtP
6RPnr+e8EyC94/0RgAijxkTXGr2SiBam57l/ybHVbztDmmteijQEKDUWdjaJAhaLkwIUg1tIUN4g
uzyn4Zphi1ZOHB9kgKFihjqCmYbSqJ2bdQycL3xy3MYmBScLItx1ENcN/67itsAyWVwfHcAdj4/+
MBEjMiFXuV1m6omnpvlK4Ea5ySYhuni/r7v2pB8TVL0LbIZ21LE7F1eVg/LG3svMHFsuoPDBS2Lt
ufi443z6agAQ2mZ5AmysGgFXyE0sL86E5R6rSBXKuAU2IEEEcYF1dqwgT38aN0Kbo8B0RMB6rtdK
mIT5xYN9ItL0hvDmH5BWQbCMWCZNN0FBipjmX8RU+jhkzp7SgCoAGPPxoXPyU6bHfYxAc3VKWYXF
zw7zAgtys4o1BtSvCGv7SiEUWN5Lwi5qPBA4BUAVww4xkpFcxBVWt/ka1owKQgBUi/Zuj97RWHFA
ryzMM6Km09wrGxrX+0eeegv3uDjh3v50ZstuC+rvxcx4JQPv/AkqzHxVqBLKbS3jUk1mr6RYjbC8
Lxum4Nh/6zB7X35tc1gNhYoxTjBkNB4wv98lqYUPrnpaE1H8s9UOCqVw90HEtINtFJ1rS0QyTz2S
TI7K7rOMfyhCqaSjSCZRbN5c0qzeC9+dMtYobbu458lCW3yJ9ZwIvD+aA9zUa7SDjtJQ2cUrx9Vy
MPx/ht+6FP277MFyghkkVh/zWssEDMzdet/XYuCHzZPiRMytYng+paeWm3TvKXjzxKXZOL+rhSkC
fu21Xjz7ZMx+X30omrU2U4Gjh1uwzANxo1PFHu28mRszHYktPolp3Phw5ElSKP9INgu4Fza4NG7D
WbEmw1ZAjE4330w4yElqzRBpiRhKubzClotwjcfzIATBGqxFPKjn4k+ppYfGqNa7xbuXPCT+t1DL
rTPmbL/3JR7WwnCDHL0pWqWBtzcsgngA9tdsJJne0uACw5mzbpv4ir0zzAWQFdQJeMkTjPK2a7Hn
TH3FBEGykAJeLNd13f8C4J0YwShpF0nxs6gmeSYDzjibbk+8+xBFsbx63x4mxTEKL3jxMqMW7ryl
nFgFkIh7Q8gXsYk9opqDBfDte5TsNM6xkiw6rU+W0nZVPLqSVA4LuBSCok/bSrE0aAW+CqDZ73lW
1O3Yn0ua8JHN+KYJTxd8WbCP6OnBJ1I+QKf7pDVBiG4UPlI2t87cLd+ahQFnvmT3EPl/NPDqbAmU
uN219D60M8xzrRf3qMES8lI/HBKkV0TQFlT1xSfXKrw3JWZkqlsnR7kCKdQg/IgW1IWT3ZnpFsKj
7gRYoWZWMsIehXTzvmfavKnr3qtcLyt1z/Dr/aqsseweWnUjjLRZCWhvsxHsXlfsbeXMX/F0LcHI
sQMD+L/+Mdo3YMRh+WI62u50d05JbTrCWD5b+6Mj9Phi3ec+oQxaIL/ivTRE3XZj+qDNb4mnJQjq
S2YV6uW0qfl+3Vv7sFAAktlfrr4uO8XZ9Fn/6oVTEa+vjTQyMEZ0vmA4Ky/jrjDvnCw4XHIaLTMK
sBfAyJbHkyjMxEMj0g7NnNUbNaWzrYRIVV8DzOPsTmbsvU90Kb7lQyCGjm1TMs3QftIbhvV3NPVK
9MaA3L9KdLbo+kuGZEEi1QdW+7wfNW+oaGEWN/6tyW8Gd+utXDwED17jCDhuDZgu9rCw2bUMomKS
5P1C1J4ucJG4BYEdzXtt86hki62TxYgMEtipNLJlGFh0pIpbQECTDVgWakDG5EbQkcJ7nzTaTO9d
ygGXU75UCiGSVEJJDjlOZUsXaOzpYFFQ9hSvCjA5f6+L/2u3S2fmiVV6ImTPlWxcq8T4uDcxs4yB
D1dgWNrWBhYA1ITnzfYbb0ejcuQPFx6yrF7xG9lmGNnoriBiYHz6Kv2m1A7Kp5oZQo1dD0thloOj
ivqvmEVm3qGEdiL/ZkDzXb63OsxLamKfzX7IgCP2HT/1wyc9dkAkXNY001YZ3RZQ3ONlWonI8Rw9
NOJX9Vvvvlw3mw2PDujs5wSzWFd+avaR46BqPvtbdwZAZOKF2syHbkIfKYtEhiBOapq2rs3xNsLH
anj8E0S54NadiAXRA4c7ddTf4pYmQcnVrz31f/nD/iM4KO3x3O+i/2u5/kSa9szP1z6hbYo2yD+h
spTcSqFGYBsj4mlXqqyMB3XQXhnXdrSD0+3k5Nb3pw93tdhLGa8BRSkZYG1sHXvKdXkoFZegNbI9
4D3kgBUNAotYCSlWQtuuCIq9oOdVQsSFpYoVVUQT38kPxR4V9EpLnB288pVD3pgiyqAvBAfJP+1t
ujJfDduixEnGDg5MbiD1RlUWw66Wmhc4NxIly3TQfpRBxTU251IFS5A15qHVWG/KCo/bEv03AKln
aDYPMuYJ+vujvgu3T5NVLhORoQWF+4GqAxcjX5XFBy2qqajuZMWsddXYo5FQXo9UrJW5s+BSf8+m
m8C27Gbjsj4NBuIn5ziJ4BQgq8hCNjkpw+jF59d+LkTekZLW5ZG4EnuRi0g9F9T8hJ+nVogAVPNv
2zvEIwQVnIpPE6Q2SB1+kZZH17OnPGfZkfdjHu4UYEvw14UYgIxxwvMiiVQknF8Ag3eSMt3JyOL/
9dVJv/pPBIoPTgH1M1FnBz6LADEP2i4M6N7yNt30VXzNWqKYJ/XMG5QhVjqAlQFiUw3g8pGRUPvd
sAB+3HIFNvbr/rmHuC9vqpQP7p3/893ZrRfFr51/tU5qTMjqxR7FM/Py/DSVvV27dARnZ41SUJFP
085/KN64Ag+eBIrwWQc9g8PC6R5sgvgP7wffVSys/lviujtNgdTrp3lGbAD8pvCeUDyAmCQKd7VI
k9DQL7ty1sHdNFlddgFEwglWG0F31q7WGB2eqvk4jrGnHvgnMJVMQutQZJ5T79eRk5ODw/tIB3Mq
2nDr/ASr/OvtkIoDeZHA1od8DEvm2k43aHPg7mFMJDAOj+gUGe/Sn7iUmQOnK0KsyW4wpekZ1W2n
UJMpar4+s7IH02PQzVpRSwt+RwsHIyA/bh5CcWYf36cJU4vaJBA9BBmsBGf8Cti4za4M2KzttU2E
qPm4HpM3AENShBt3dOtdjjkdMkq/k/MIpgNwa3Rsc/UwRlnvFA/8kgNFtXHczWkEIhMU0SCI6Sep
b/BWIEOZ3cH7ky3hU3nS2QecVUXzJXXgpg/UStFM31zEc6RE2Z5xdk1S3UXWMw+rscu4kmbidTWt
VRZ1P9sLvKFAHQqFJIL0rw8rwBZN8CFDyld/k/5eFWshXryzA0SwJK5DvHb9tjALaPDf/MeQE24H
AGSqO+I4JCCFBY0I1YWLfGtVxE1tXpFMvm/dfQ/gqboXt7UVoq8jCBrhkr8RHoS1RXPwcEcwSoRK
ejy+MXpXwu2pzO0pYmSjWjwDfDpjtPUcGAaL2eSi8DvcYcYAVcC+z0MIp2h9pFArhF8/cJ2CFTpU
X7pQN2a9Zo9tfkRBRUpjP6qOWy5g/CsVggpJPN1R1Xx+AQ34aVLtesiLvHksxnTOyAUwf4h91jjz
hTnOKVuF+1EvDdoOEfRjT8tmC+VsMVzFsTsA49LTeupcULU1Bej7xhyUuMYPG9PjkQX4QOL5bxN9
OxcoN9qb1Ge0Jyo3V1HT9x7OaLfaf5XzmlOzIUTizWffgXd8nK0FARbQ2Sj//Py3GFhCon/3tA7O
RTKLSDy1gHHcT6jxanq2qWycIL5SAfY4tR7XyGz821nvFlT29eSZoGd4ksqA5aa+mj6jiMQHKIEa
qGhwNeXuFiUjtzMaEIaDphjxJZEW6bZGR/cSKiUKqi8vPoXkIYzWR8sC1XL6O7xQ5sI5xRX0w237
bVkf3yGIMqs4cGv/bXUbN5wArSVCJLNlgKaaoSgq/eicQrV1U6/8ZKVwf75gxKf0t+FY27COgNpL
XtrZ5xD7y0MC4uFICHqQnVTRzgEYHRqWsY+W8DvEjtxi6dwZqcPmvHqzb0mHAuNQkJBVAnXWYhR+
BlPZ8pYyszFnCsQ9x2CAwDNNJRg7PmvnNDrqZePzFG8J8qMZMF2aasHkaja9IkL/KWJFJiFfLGJE
O3/GmvVbia9oN0vi4jEPDzBUAI8DhISaWozw68R0G6kRKOFPtnDksgLP20rvvZRiZaaZ4n4KxWlI
ZIMH9a76b9EtC7BYauyYy/6vmXif/FisW5FyxKq4jKTo8pcKBJI1ZPFw0agZdSs03eyl2QbUrKaS
6qLUWvDdWrJmNyI6rKvJs/CDDMG7auvfRhDh3SbIFtndYVjw32Aphxq8C3IoA+y3l05FP6h5PuUX
rPOH2V9xb8lPwr6Yui3qFcUln1gCb8cmqGrFwPZiZwd+KNsUSPJU1XtnRdZNnqdyYF2eBmBC4u0V
S7H9q0zk/P7wtgfrQgrgsnQnyuDVmQd3z1JhjP0wB2M9NlZOeLApsC1TW7VVkxg6w26FYB/HUPKJ
x0eLsLpVT1P5bCFrLNQW/ejFrRHAGFyGqwEss9PZbEoXVSwb9h53pB+yvrgsrvGeDb036IAikuX0
6IzPOyrQdJSHCNNojJ0GbA04I0M2nz2xE3j4hI8MM+0C6hZuk1HkiiFqLmaI5K8wm2x+dUG24XCl
p/iUKxNvk784VAgEGdVygcciRU2+wdzk3g0n/QyY5hsq3xPpGCX13rWMlfTWFI5evnilkhy2uCmk
bZaHQs4s8TxeNW05U64WqzmDgwM92vzjaVI0uMoa4x44Rruyyqb2WN5T2ky35abSng1HrgRsfUpM
y+pqJFiZ6rYYxN5QfKPcsOTyIYwjFAdnt+W9nWtrAVAiJ12ajKp9HtED8EYsckLKUbBe1l8B/34e
qj1g+hlo3Ej5rSqujNvo8pVcpjt2SZAB2JMGpnzna8jxSdWql2Ui/67aCLKCcs7uPyMJkqS79pvV
neNFSRNh2hywRA4PhxnLbGJx9jX9CbZJtwqVDKd2Kbed1sriovDEQVilKDrya33IEiBOCis+1z/+
e4Z5grP5wqMDqTWEr5IFd1+r4rH7l1kfgJkEPyDeec6IpU9zPGoOk7bdwyAKPA4R61hVXOvXoD5N
ffDrVwc7C6hL60mHdjFBoE1R9eRKNiUmQFdDFl+JWSg8EHsu+RvmqnainuIQ1vMEMvXTB+zblUj6
SNu0NZq2/CfZllEHEHChKn+KijsGsLtMiOJEaTa48SF/7X+/5oCl/Ma1hTsK6NUogI3xqfYap4c9
bE3blYtUrP08vYTNNh+fS7klo7QiUo13SngMSGQ3kcmhaQwWMc/g9ucnu+3pm/PH2EW9yHchIvUP
VIsnZETBM5pbpIXnJJEIdFRfBnahKJyqXk59WCvrN1aOx2pr/cPbYHI36aWn8MpJouPLdM1kHlNS
+7GnXFJHIL/BBqVbVcu5+Tp8T/tvNu4GQwijmwNmm7KCRy0H6imRc3BuP7Z8XfvrptdFMqkfSRiQ
3TqD511+d6Gq3WMvuAKSH2l1By6nn8+DaY/tgGYDrlwd+RiHUZfmlCwjDid/nyNbg5P1G9dMTwJ2
Qps8HB8BvaDQ5e3JZxCwsvhs2uKX1P27qp+VEvPOBMTLwuK/Q2SZ51i/T9/mAxeqkcObCFE0a1O5
cnci+qvI/3ToXOBQdXd+CDWE4GOD+AvBVzykl+rJFe43iUFDY8sFCkymC81hvP6plv8xVnYm9MW+
x1qn0sSckeHPFKVLGL6p3ouztTcg4pWAkk5LzydmUoCEtonZvQ62NmBz7Pu2HvenFj2XXEbyLDZc
DzIDactGrf/LmxDaJldAtGExfgJS9taopG/xy8M/Bb/zAsb1uyEBvUgCp/FsoIxcrnJb/IQeII8o
/otwMqeHwhjOtowzzLFm2zJAt8YKZ76iAkIgECs7ktBd55L+i+s0Uflq1s4PXV9j7e7C1+7X/g9x
n+kK594+gLp7Awr8JKqMEketSA1bOwTyyfRT8l56KAIGsba7ek9NMDGGqRXFQYeGPByR1N+LP6ly
OkQwKJVGLb/HWTsA5aGU9u+ZUSCeDM7IOkk44m0A0Y3nmfCxEnLjsuFs6oiLwyt5S61pag3bHxXW
kaCNVcEh66YUnms2nVdPQeUeArTEuQQH5aJdnhjqhtexhu3UoZs1yU3k7Xq8S/CWBTtfzyiwSPEk
aQVcLHFd50GTe3cQAn4lhSbyI6sA2ObiPypeAOH0icblAr91W4cYw3p6cQFZ53ba8UNERx+5RUe6
6HvaR5CKy2r7QwHwYUqSzKiZjVnOEs3WY2w1BgMmhIqlWyHjElt+2Hij/Pc4XYv5XKAnm96lztvM
y+wBCwuGpRAn7tgKMT6F5nyyBt+T/AyvN1abWFNGrB2755svu75q4upBVA8mhdzHZyNm8Y22WnlM
S7e/EgkLyu5kjpk/rBQo3qOYv/TFAyMixjvvN9fee/06OE4o+g/oVFjoDuEKe+kd/DRaUyYrQH/i
Y35w0LTcyffwSMAZDJy4YjOU1DWZUNFvrELkeO4TrjwIVwjwIDQ2ikRz05w29eiJYZmqw4g4WnBk
Cttdnl82wjxXU/9uF69/qWZxG5C3KlbtiN77Dwz0LtizuVhEUW0DZzEx477cbD1QboFO58xPw1IJ
PEPzHjrKHgFzzLIPqwu1CktKYIzrqfFwutwN6Dkc0pXUMjFJ3NRXvE1CF/kn4M1QtLmG0GrO8C7I
GDsJH097hgAChYTraZqMXSizQeUfjHU/OnP7AXvtsSY97tdaGeE6P9QsFbMkguoodcA1AHWK3Qpx
YXAyl3uCHCwr5qxouF4tHTcbbT16TaIvhgBmzYliN4jraaGR6PCiXTybfz35L1LrIYyv0zmYvgto
BWFoshUCn1nBkrVEpSLaANFKvtxYDL+F1cQ28d5/bU6yW8zgoGKxjGLqSUnl08Xk39OqFxGYGJ+3
k40m+FXEXoCy8dXQp/tGB7SMmhL17ORv3TXi3dfI67nNPqcynPeYto0nuwPnCVbJfDHgADvAmCbN
Tkw6RhqM3Idrf3ExRgwLD7DD3qSenY4zfbYyQIRJ/TX0K2bYbKE2dSi6R9E/ZTCJEMp88xS3im4G
VchphTK1IW7Rs1ETQ2xWYAd9h1q/A/TXsFJIjNN6KhUxzRs18jVUgGxVFJ1aTtr2KyIXEeHBNwth
Ti8Q5+cunIafpEPMjUvUMkoArSnKTe+3C0qdrBTLGp01++aKwSLUau5YJ8QAS2huRlCs23Vkd/tO
FkPnIMw5kCJ1e2+9x6Vb4Szo6tGPyRD8WRkjIzS/FipBTcMkAgOjNK9E/SCTmGtIPRkiSIDz55Zg
2BbBr9j7muP6w1WggT7HbMl3V1IS4XrFfjxa7I1UL0QEmVVPbjqgQllQs8FNSBJzX8vnJNGf6M09
SrA2hpJBHOytERTWQCz5AInOuZYUX55mca4T5EvB3NiNN2YuQeLmnDR+mqKrMDBbRp9Nuhdfurzh
A48hK7R5wieBDXdfWHGaOX6wm/jLdvd0qLmwos+8lgRVjDTlsVKj6FH18AF93vzTp34+yzso/MSQ
9Aicky5K/FnbaYezVNbBFhgwLz3QzV2M40TzXjZb8sR4xx9SNaT4U7pOcdNpioNACTiwCC5C44oS
OjHx8xkwMOZ6Gn/sYS9GYOQcb1nyVTiQh9g2cA81hEmlPOxDuIYo3CyhYpaWvJpb0yX6H7tGHZkr
wIPW7n3gFKLcHIIrEt64dzqqcIwyi9FxnuYHNHUQWBd3VWogg4e/sSIk2UI/Z7yJVFcnNszx0r90
KrDn09rvfbf9UUXMe50OB1NtTk9D9uw7PDW93NI5dr1B9qNFDteYt8tlsbeD2bOtBR6ns87cqAu3
kJ9pKd1TeBb9bhyZqjGKOVp470HcPuQPvETLCE1dOebd8oa2Wb7gylA90wuNvrNMghfhuScFnkCo
exM2giKRygEDzvZ1MqlkOL0AvGM5erEGpN9+r6mthddtjk1nZwiogHG0Vhkv4RU//m0yj7NNqikN
6u+ckpv3VCWjkAf4wwnEbF6C6/riZ96qTUFSoLyo5bKquwb3b6KSvN4co00pIZOSv4FbsoQr8rYQ
EDkeSBwyqhjbqN7E1FeaSHI2jfPx5lPOw1vKJk5iatgIN1//DJOFiV1/CEQbO35dYx+BhQgXXuNn
7iRTw8CK/qlzcjPSpnRdUj1mleQV9yByTCIKJRgUUfgVy2CpfgtN79mC/7ewY5hT1PromsEYzls8
te1GNH610K76cDKJK90jbNtwbhxNzwQbnwnAE64McHHXpQ+5sjWi6bBOSaq+N8zCc8eybBGAv1To
wbxce76Oms3qjUDMrh+0ia82FpxWlmcwpNdf52jxlR+mK6JpTUATCN7fmt3EIum4z1YjGdkh23iu
e0Gac1bfagpzcC16g7+QYM/uScHx1N7gJ96SaI0rOWFhs5eKZT0ReNcg+lcXdt2A6TZrQkrvoFQg
8F7esEWsNaELlMNTqs1v1Udpk7QpIUEoaXtBPdqmGaf4R4Lv9CJTLDRHY5vqQR6gz2gc+tBnoG9K
vzRwPdM63pVD6GSmLtcxR/1WZfGYVwD1xziohSxjiXZ3dtxczjfxlEWYakP38jrCTOQVPEMJ2FCW
oQaGFlX2MCFD9Q0DKTVr+edWsLESnbsnWW44qefN4eF1t8yjVVvjDb4xoUWcz7ULzTT7Qt/Q2UxD
Q7ydaDr05VVr0YxQmKx82kkk64kpAFwOfnpbWNjfwdTqNutnJDMms79oZJ9/ZtlnV2f32xctWEbn
vM4tGHbZPvR01Npi5AMfXb1fIpBIbCrBUAkn+xgIcxd906h0W0h+kb1GD/FvU9DojtJFHrT8e0n5
uVuqsWZNFT5dSF8mvuiaqlB+nT67y6tGsSAsSa2xx16mGyIIzVfFaGrgdZ0pPpMrKZHVHiPWHpjE
Owj1rBCtdEmOBHjFowBEo4FrwtaDRQewdFSCbEvIRBuCXEJwlpX/BAb86L3L1s3VhSX1KrOLVm1y
pPRalxLlpVmtq/5r/HC7HOQLFXu6qdipn0KxsgI7E1T/pUf2/8oqe6bXhTl0p1YE8CjcsEOEQO+/
qOCM9zkub7GsQm2iAJll2IYoiWpNaKyrkLpFSgObt6vhcjIfD+ZI8zXkD39xVLRzEAUSP0QTW0n9
mq445cS7OhbPf4rN1UGIsTC2oDk/vhTLycCu4MyKNoxpZMnFbY9w8AiZc63vS9H+1wiRy0X4UF1U
vn94iukCxxdNxzsUEiRvGc+BAYwXCQ9R/4yYkLsGuOUlkMNxoBMaKdfQd0YJolgRDAVXWKDI5JxC
uk8Aig3bWgOdm145U6Kc7Nq84iV5DGHwDERSfp2fyOsJWibkXrw9+QzC5t058bh2C/1ssldyzUnO
a+IbloOtPE3Yw0lSSIMuRAhzQl8til1O1gNLnA4exYZzWQ0SzhkSgeXgp5sSplwH91n9Qprn0Yzs
QhW1H4ASuMqldGgpFgUqV7fYOcIEbo2r+mmC+kB/4x0Mh9giOwOsiGcPDGfhzJGH+DXq+lip8qPP
6DOCuYegeTXXMEC6miTlYaltrM+EA1hCcaGVhMeD2RbwgvjjRamEGjimBlOfWZsopWoz72Qzb+72
zYVCKPDrHkEifQFc4BwXD750hjdXp6rEb+3QJ6Wf9aDfchbg69s6BCohNBf+PLtlOVKMRwvtI+bA
I7RymNfRBQEcM2NW/PKXpHBKiyl86SQToN5K5ojTIJkOWHRuMZWu7n583QCLdwH+EZdYJcvjkl9S
ezD0zPj9RRvNcCET6RUSFPSsUc4/aEeYX6V1Hft07eKMW5lHmrztJyhnUmfloEmcSiMUE5ioArw7
Ngn6oYr9K9kHand1+NOUXol9ia50I0Qu3hWZRtyYX+3FIFK5jAYnL5YJIqTO+EUjnNQwq9IZeyse
LRwoNuQlUlTzpdaJF4tfU8IQ/gwD7Ot1SZdM9kQs1MOAqt81dPlHhsbkMqLNz5nsdy/MfobQM8vo
Jhizvj73wP9aVBfyydtym0OVayLvclN77gKRKIR/A6oegVJds3uQTzAvoziYqQmENVGp6tfgSBQP
COvIO2ajVIWCamW+lyk5jtRChwpzwb5oKA1CQoKyJvwffewJsRc67I1686ogqMSZyRZeSYW5acoQ
pq89SoLy1GlOle+dBRggSH2ZxQhYq2FCFgdr8oIDvdcFP4xqoxrV/VRArfpO1/zMEHv+2wSAhYNt
55b+mbtqPiJP2OkonYzFENcaq8qP9sYR0mi91KWoXiQrOCnIKFf4D+QNwePLX1VGSONuCvGtfV+v
rCXpc/sVLC+CcWcpfJRVcwIvOwkksm6+XXTg4fWNzwsdBRABW9xr/KM6JGnlIMinAz4wEkio9HGE
MX0yXUwYEEYzj9mu99VhKxPbqDkhfgx/s+gAr8WeBIWiYgvGfJRu5zsWKAceGsvaOTTtZb0Nac+B
NLnnkNKd6VHFJ/FYBxv/XuzXvvUalnJoAQ5lDXoBPvBlzxY6ZHjQD6soALzTXfKUmEZAF5sm8EvA
RS2WU4D0//mGrXZkYusaWuRUOIH4eoB4g60wMHryUIoa2QtNmFYa19m4oIOfnOkAjPydEJX2ZChG
s7uCEbchMULVuzghDkC6gzKmOF0cYqgTdTQ3hE81d4jsiEzlcZNUze87NYkvD4ZZtUtdIXBcvLAP
zr9mwNWESqLJnlTBdDFVidPHP0A5OTfNSSfAa9RW2YpLys35a6k193zQ4EAPmVApFWoo5MSXs6gV
M9DyBQAxMAgXrkA+bYpWjZmnmbD4GVsHN5O02tRV4G8d3Cn8PWJhbf6Su8X3TZWiGPCej0Phzeqn
v8Cw3/UZkDw1vlKBaBG3ADEyyQqBKjKcaX2qA235IJZZ4xHjZtGPNmfCTIKBiMqcwljCzOnv3V0a
dfIiQ9rnNZLLQyCqIIyFSprzjEBj7+3bCFWzL2sxhllWEjL56A/PoPrdSYjbRYI361CXFCmnxhVn
xTqHGU6IfGmOeP7saH4vWyVPOi6PepSUEQuRBAvH+ORp9nbaKY1alVwNDTyqe/SbclRgDHewJGwB
Hfqd2TseP/KzdmhPPY6p4PG4+SNGkRCMGjzLMvFP5XblPpGRZYc4oaD0QTRdZ0rbOl2Eceo8FBGN
yYYTSMM0OBTq9CpzdzqzVaQyJJyzZUz4R6q4uxJtPKTquP/8icnAb4F1f4DEW4R3+PU65FTbVv/Z
0AWKlkVpFj2E5mhezjuGMvzfHTWQrttcxu1PcnaIJ64Dc+d626r5XNYys5+PG6tI4uL/Gr2dD8Pn
m2fNRui0FdiVwP34IojS0ZdUGK/gIdN9FxJK51JupBBrs+lY3Ge9rlnyMZySDPdm1F+kF+gAYZnO
PgsLW4IJjhMjH+bGXxL3ClcVdKFgtZG/d7TLuxTDxg79rPsz8wdtuLT9rcnssUWKvcD6KTPlQO1u
0VLebrlN3GRdn5dG9z7ngyYW1+AtdCmUoM8Jd61rjBMU2ppnj9XS7DtDzj9b/yTffnR4EiUQGA67
ETfMQuGsfgirukDxj6XfSx5p+Jj2jzmm0gafu6w5vzlUiarDHVOU07vDal8F70l3IIY6RUBYhTJf
Qo8t3H+LYLsDuYXmbD0qOaTdK4Xaj+KhM7kJrIy39o0aJiuhQCN5FtcblDjgD1oMIPiIqWeEmS+s
3ZYyijVshphvF/4J2xUJAyaGkcsBz9g79jzyWWROcESSuQ9LLfOFhbNCJLErWIb1+vyuuDBUkUA5
R9R4aFIo/tj4Tlyygq7LWByczElRQN9N4+QYDKXLUKdDYEzCAptNrOMJkIKyNdlaSC0oBvAXjeyd
AyNkiEIw8FB9Z6fg+oLED1DdWYCC3gn3Zm7F2nuV+AZfLPU4yXVFSWwJasixBCPQQReww6VNLS+B
JjuOQj7t9KR1miD4gT6aEFhQ270+3SFAL2yalEfwRJVxM7+4txiYcmtn2s3lDqKsDYIQcbr20NKZ
JnV/j57S30K0N5bxsVzG6l8PblWm9DJupjQqaksgpXkr+KqjHnJ6oZf+SsXNC3pVx8Pq5BxcKHFQ
Pnbx48ZwAageXRVLyPLdKqEvEsUHVdIOalwFtLhWrtlRqwi6vi9RyPm86fGcpnIJAXAL/KV5DUHk
am0D4bIAO95i/ph3ghhXuR1bLWXdZFRgTxka/RN5BDWqIBcz/vmpTK6/iACwke50pK8heVHh5cgf
LFdy10afYw1pMgEx01c5PI9QoBNjtHfiP+4E11yfjouex9hChhZ/pVM3l0j7/OIPaBgQWQ52lShQ
El7emHBtenwRgct7vb+R8mKxPTPskcxGVzHiX5bXTWwCb8ln4Hr/0sooQOAIzBk4RgHtOIp/IrwD
veAw62gEI5VNYo8j0pxTl263IrHIEeQ/NCoEez26NstggqOmRFqf7rZESft4yt2jyWAswMH/veeJ
yRO29+FAz9Y+uDsLs5EwG2YaSshg8zboNRaHxzllcmkxjuCvabT360a05njv56DeHhtIA/tw0yxI
rV6Wf0o3+63IePBPx8QaN6WJR2vFZmHaoqjcITkH53AJFIqgS4Z0qJYUbH3CivOSO3DyK7v0HbMA
MTuFG7WYqYDi6oy9fYp7zjCnqrtqKJ10KZatrIqzXEM36QcfbSdqc+i0Nt330h9e9nhh17S5WZl8
d3tDv4V19xoYtDXDIgvpXYIdyJJrI4iATUjI2cmoXEXXpn6gwgHkMOgk22/ucaBPABrI2kl6mNw4
8YDwzJRst8kgTriMNIZATzAjEww89VxEP+R5rM8qWK+yhMlxxiHRlx/vDtosUa5l1e29QHFylYde
vdlIZDTAKwl64JT+aURinoeHOMljwqwU2vyNA7FRPyoITKWkkPCZrL24WXuuZdy8B8gZss00Raa7
UAIa6sVBB9XezchWrCILX//rZg198n8BjSQiLhCixl61U4CR5omMj/YsZ+eFpBKYfqtYPqSy2OoG
BdVmdVnWZKXNptnewMR1LCr7rvOf26qhHOZIqYkzgqXiAaUBziiuMJ2HWdpORH5H9MT4JxH4rtsz
Xt6/VoKK1vD+ApJe+vKHtr4/SrrLqfljK7r5SXDB2/V35pZ4V1hwLNZKT+AEDxFYxMXyLW9k6tPl
jD88dVNpO0pe9Sj49bi7Mx/OKWv4EJDpLq18mWYJy4GQDQ+FkTYY78qHanH8Hg+HjgDkHgulLHgn
UTAwa6cRqJ4tt24/H2+lJpS6Iw18pJHJTXOlJDXsIdYLg+L95UpWQlIMssLtAsscrvAraTXbJI2i
ZXbnC9mJvzgQUMzaDsyJzZOlAMQP4mGJqDDM4pnS78idYKXi+7iI6jZWzybTPMFCmNy6hk8zN1pJ
XvbXDW3S3IXxaTZ3z+trSNQjcZdQCO7R7JTHymytNKX6Qb3hrn2N3IgYRkCKZJlPWMUoTjexSGI2
P3CgFDyrTtgJeGaN1WfZNEdmEmDSl9B2HtkPUj4iE3tp/E6ovNAgfZKt2W4/OmXNSI2cc5zJR6S8
/AwYMDf3BaemaZDeOKbjcOXC3Xj48XICkTt+qA+6Np4ujcF59XEdArMsU414saUXkD7QtDkeyu4y
jdi8NXsQvrKCf7ONDLSYOWWzKP3hXbSfayHCY71KF0lwiE2BQPcGfqoy1sYXS9RFzYv7nA1tNLZ1
VEitsqLBMtnAcF/Kd+zLnXgV0/cVutKMRQA8jB03HtnKKdT+BH7P5LuF0X3xCnEJ47bDP68apJFX
+FNLPgFIuLKcRWLx071C079MG1wpQAYCOi/IpF/KlY+XvEvbnZGJ8mMauSSbF3qKsSUKZx/pVz73
U/DsyfA4rG9aIRdFC/qj2lvQqbYPqpvTMmYAk359tinPZHeT4V1JQNnwrruMoF5PA2/KVEBVimZF
lDY4xj2vx82yaZsGQ9kM1kT/8u42kh+f0jnX4IfdYk0uX0/uIOMXjw4JuJwf3jwBVe2/7R8dmJVX
D+W8Weqt5/vbzXWSpb2sXo6JSwmamo5ByweJfWe3eGV3dKtDxoZpETOjY/evGrl+DUexRQt4XkOy
nA+ABGFIZNBXOl5pmfArNvi38MUwb7YJMZIf2x66B2BZis0Wbki0AT2C4m9dGxkz7HYulG0U9TF7
TN9wexg3toIUAS3BV11LVuNLaxF/5MvryU/70awotdNo7Ws6yNu6kpa8tTwNEx7IG7BP0k1Q6Fmp
/0WnRQ7D6NTYyJ9/7vcM9fB+ZuaE+CPzKalQlS4s/2JuUF4c73ofshtFCpgHavY2Jtq3rp0l+eem
zokAXAa7B56k8wNha0JxlDkaIAcpgud7JAKqfQmd8gy62ByO+Hs/MHsD8As5VrZnf19QRn3vGwXl
hkHRwPGeasFCxzTqFMa6JFR/aoDoLTiDHhW1WLeItt1ZdiEd8uHVCBUrlCfeeaHJvoTnZYIEmmWw
KZJnPR3I3XL5mW6gZjUixeIPWHkqvyJ2QR2Qu56xXUtg70oZvuKCQ/5ZDZfCI8OuwYbonspNJWm0
5abqd7G7wg0kKRpPptDoodsVhGh9NcqapnadCK1QQ/IJqivd46MuK4UNsUH2QYq+VW1UqRCIoODa
xtu9tn2DvEgMToRAK8Uw+bQKf3E+q3gDxVuH2/+nxi4yRpRBwKxXYVSDyx0D/ojAAFpaaE5AwWco
Vb47L/BOSM9gAEcqogGthknCGT2O07HjXTB8dSXqjsCeaT48Ica/Ny+5/MrSRtAiXUYaJlV3qEKM
xBonz9LCFNH+x1wfcWW/s4cMWkzfcv0J3eqw/MNNDciLnZhKUFddjSIXiGFcd2Y574rAQf9bwZzI
+rCIT4oHqfRo5NomjZsNK0v4hSGi9uNuZGf/Yo974piRSSDZhK5U1KEdO0cj2mcre3erGZhjZIMB
gurhnlMuvRt3mhvcal7E9nlACdkzu1lymVnDMkzwyQ8vC0yScsncBiko5m+Tgwg5KGXrmR+wttgR
GxD7DC1s6M6zn8cYdui8UHUXeSUu1Ar46zI1BSQkeiF4NY2KurbLx3uFiHmlZyoHn65PgHuT27xG
9ExeC5Pc/S4e5zmSFWlU41quFW3fL9+SKCiH1TXaymS4+7IhM9Z3VDE853vu0SSpFzZt/gXnZvMM
mKvNSaxOdiA8z3UPtzTnEDVqVOY5yemcvBqY7CmFlBvNXm076BFZ8ZLUHxGKDlq4LkoIcobWrq9X
DL2rJRzTZm/bt7BQk9e+/ZeC+vQ1tHl9a5UPrCu8i6BPo1rFpWCIOxeDfu109tbrl+EFDzVthGxr
Yy2Zd17o07BneUcTlpzx0K146ehFJede1h+m4UAOy7sMQM0WG74GQ7IgPQinduFCjDu48Q08SMSD
IEXXf51Q2Jzp0vCmmpA2ftTTB8gl1Uy9d/3X9QpUlbQvv3KEZRYXJNmSjwJn673vH+jZlDGrPFPh
jRQmBD2RXrltBwb3fOzunPUQ4CMCUzBYe/jUxkF6cvX4Y7X7PrtdzzyOQ6epJR9bv08c/oLPDKfP
IrEe/q9uUDMaCduwTlz97NUWOdICoJ4QrffKGlF+9+FIR5k5YrdKYSUoneZS/s1eiVmIWElEQdtS
CiWU4sU2rgvugQCQEwC43vpp15N/MocmCvk+hPCfWHHBEiT3Y1nFk/oMfgqDxgsgD56hWfdKIeew
DL4FIqz/PUzQJEdAa7f92IVhCGfjCLv5xQ0unelaHGJv5lAXYIAvNgZSvuD89YnCM9S9KiyB2/n8
1JNne0DIyktWxW3fF0kZ/1W3ucyzW8YvOGM2FZikMEYtREeMNzG+BtO2WpD0IvuQx0pi2pdv4hoU
ni3OXjoEocKrgcbljFZ7I7II9pOi6V+HcFmqVly8ZQ8xduFSd93Q9y2sWdi4yOflqV9r/4hQ2/8j
PMk3AanN9P9i5CQWv4Ax4LW3uNDFg0dV5pRHiHdOhhd5uaBsFVRsNieFpwN0sGWeTKfd987e2PUx
UEc12PufjgXtAW8Z/cKvnYGcJ07oD9eP7w56TjeyxzGZVUIQ1ZS/fA6KfeUfY8OCRI3kiKihBzTE
81srBvUhRmi1gtOQqRpP6dntcBF8VL7JoyNn+IsZ9AZYPa5ng3qpiNj401pQzP7XQE1lbrwc57/8
Uin0obAz+KpmScP2ubs0zTv7Z/J/BZX955zTFwnvlfCGqG4co4ixoh1Bb7lRfE+7DSULKWaqH1xf
YkwjxGiIxNafk3PW4tEo0mftZtrso0Yw7k9OIAeSMoM/GryPTUNqIrucL533jVHnSoXNr43lVgeY
ea3/KrcwNJFkezXRCfwdhyLOgR+551eM6O7liHAv4zh2CTWmjQmmpmmoQCs1pC3z0fpKmgcglFCw
8Tl97It//tELH3O/FZzT7Svv6q9hFDdT6uGRzbBqeo5gKKBrETGYGZ1L1YXi9gqCzEdiwyXNHpAS
j4WDDB/PJQxMNWTTUNhfnwBBRaSvFQe1XRcN2IaLu4x1nF83MelE1EFng2NxLuWW82HQMSSFdEuq
MSrySMpsOwiLM1JvU8o55A9i4l7qLO1IqrfDnBfn0kNv7z+1DQPZYSds+mDEr1uHQ2yqs2Qkc7W3
x1rK1R5si0Zg/E+ecsqpdYtLja7cbcFCqbGG3knSBkVg7WkeOmhRYg6CB/c37JA79A9+sDbeWiiG
Bw9Xt57tt3LWQHLzAgKjrNsEGliQ5zqiuixS8p/rdvekDICaJsU+FuX2EQQqY3bA8V3tjdRa3fYv
5+oXFEQwFq2jlKV6Q7UwCleswD6QdhCZ0i0HyNo1aeBH86RAcDi5nmcCp1HFyKyiC9p5ec/+xwNC
Hklr5JgCBqtrWlHVM24DdfbkW0bZYdpwnkaZ7DMg6SAMDX1sczRxZLrFK8cD47P6XkkNCK/iwXw4
+8txbo+JH07NMudwudWkYucw7isOKTtumtmJtWV6aRHPAYpaIzD+m+/MBNBg7qvSmg0H1Y8PctY+
0IJuce/YJJ2lxg0x6Tl45D5VRkOP2ZTfGbm+AcCWFcIx3s3it0OPDBfcz00QVY4VBYsaE/otZARE
SIR6sBFHyLyztTLx5WzRzj5ic7T9pJme5xnw/IaA08/8vZ11CHoc+pkPSnRMSZyeDsxG4ltWslam
oBD0sdiO9ZnKLHGmvJePHmq9CDpV21Sg/fCmp7YWkT+qu+SpOLurv1KZ+YRx9JmyMsRLOaDvtNKN
wy/Ea7HSfGSY97IbfR/HNqDdGf8/2Z//pxuSa/0r4if7ueLNQQ67RrqFXTVBa1ThsOdYWhGaBeaD
qng9CtwiRAMjrq+HT2NHIuChpAS9zONNlHkdhdPMQpx0OzLLJOP1QWXprqNrE5gaB43+fsvQ0iKR
Ufsnqg6OKP4w8W/AxS2yCp/qoDEifZK0T9+XSvUc+/xW6a/CtyLo4JryPxnJ0uEJ+NC94OguZY5F
qC3MCGfgWcB9su695OITSCZtCQgLTAr/br+meBMTJOYCMBdYnqAg04ByuBZsZUSaPUgxMrjL0EVw
ayMleuyGuVkS7HQD+/TLRkRSuT5YHSjGXloKBASfNQwkRdRI+aWKGzu1UxnEUOmnMDxDt05NCChl
ub93bAyGUfi1bF7rHBbhqInnNYj2lydoQUUPAypwZ6uXVq8XjkgOfx83AypIL+Bwi63gCJ6wQeF9
dxIhC08aSuXxqy6lxj8D12SR1yH/U+8K1B4qhIa1TxIp8LCitvoLKvaFFeZ+gg1ysFYNyPN+e5IP
JnbnBH40tnbbIa2qKCvhw03iP5MNNN0DxKJ5DiuYfXhKvdxDnfp1riOaHZ/tGr31IOEr5Z7oHVUI
L5F/LCc3YRCLeZwVwWgaew9DgKksdcuu69pPwxQPbpA4RO2gAQyRts8p+/C2Crf0uUtSzUv4bjDR
jO153ew0xHeH8z/BHYvVhswjhUz0JGHPSOUO5w97tLY+X+npk6OG3H0P99slmbo8IbHlo8wUmfvy
MpVifKNyWN8jEuQi4bvbjThsDN2iFb4ZITd4gULv3gtCMA5J2BMWZuh3Z1ulJLjWDnIDFSOS59Wa
4gVFNRrYM9PJvyINiPDxSYWcMZ07jyWNMULvwERzc8Az9ufObMd5ozvuxk2QxxUMlmYrejdff6Nh
Z7sbYOAoNGZUnKkTiGJV4ZlSpGFM6vDGKTIKJddcOdlUR/s56rpXHSzQ6RQCJcI7yWiPuRiRGjud
Y6eq519rkEPnnUr5PyQTn/rSobMCHUfC1X77WZ9LeRiRHtbyHus4RXwOZQU1apqEnMBGttkFZDzp
j3SnMCpaRaf5VVZ84++RtA4pBjeaMdstVpjQK0Ovsdz2SqEEM5zYdTsKG4/7/48S79nTbwnSux7y
AavtIXH7260HI5oJh9pAZhkN2YDVHTqDAB0hn8RwJPSGP6sc/17OSF1xHxaCEqEpUleWLyuyHwUO
Ws5I4Hekyk29Mg/6w8h2Xkp+almkZlhRQkCHq/UKWBlKEPq3jiJWlBhm1NGQGHKs8dSbjhrmkx7n
mhskqaMy6DPZPoiIwjdIFpC+hhXF4kAusv2jjMEv3cHxfKIHW+pwEXSJ4CsZt/NNnUfVf8SIBKsi
DmAG+g7mGrDOeYiqjKhdcy1yFDIPs8TSIYTp7CLnyWbqA1aXri6ghxJnzXa9Q8jWuNbgEJ3mxk5B
SizrfZmb3wNVcUaLteSuGPjpbPeqHc+4Kh5oJoZ4B4r4x9TAdusHxgK55Xy/4Iv64MyUHigwPPN5
drsuIrFqQoK2+ggxt1+FVAuMqvI1qENMWIF7QUWEijZuSCPfnrpghhMuF6Jdz+esry7/Qcsc2e1O
+PoIs6XN2fCJAWlg6ik/BkhYk+bGgUlH6vdP3ZARIfRavuYjchB57QOzI1xwVV0kGi4NFxWH9buE
nOnucibhUbUZjwPtxpkLhXl7OkwHGkqJA0nGNVCxvj9wwMdAaUxdYN2urXvts9FKLP98+jI1t0qW
VzR319rxhmh8EmPk4x+NieOtFDqB7sQI12zgp4/LhXmnFi6MvlvAKfzfWdGg0rXigcLmaq+QCYQX
SHQTs3UzyYpy6tMqZ2Pql6PBgfZCY5DVC8HzXgbsbkDSX5RkwH0o2MZ3Duk8e/0g+Zxt/LIcox0q
T1dGeHMt/hD4bOpCgUWjEZZuOqORG7TXGU7sr9KXooTIWqOs9cmHW01eHcHlizGZVgs/AUh3/Z36
SQutZAJ2noXsdkUzY6z3OKGLEVvC433Dn+USN+gtSu+LtOwMB9KEsM3RyAF2SH0UtLlfyZRpfmRl
8UFfQ8jTi6y1KGQ9qLhGEweheR/XdS3gsQK2z6V+9AyUnqzFmvfCipqbCd4Gs4/MVXxPGvZowqPN
17NGLB9htC6e90PmikwNnAYq/rESQRl76exYx5C4EBjD1GTjowKl4SnyxY27hyC0u/pxWJ2sf1Y6
QPaspTl0FT4rIdYyO3fB6UBMqKK7a5BW/z+CSS6yu3uO4X5xQmNywVfg1ZN/UD0C9eUE4XM/GA11
m94fzwohSRUSxceO3zL12XdkC+V7M49ekB+1XEtaQO8un3Z+Jl0b4a4/GAq03dWHDQ1guprPvlQs
Gf3Nj9uZkm70YlrA72eXtpfzYLzD+tE8i/vCBzYOCMpTZHSGqwU2in0/zxKVU0Cnyt8dyXFiKuGM
cbXl/67j5mNda5MvfVosR+QsH4qnMcQeM1AlEo8Ijfsm9Ew+eHDXnkyLAPwoxvTXr9vtjmIgvIuP
EkxgIK67O04zcCIuRxp8pHH8qLE9HaOlvnGV/FzAiWsyW78B4DczXLdlGAbXZrxY2nrDmAhpOhsj
yenL7r5RBY1SM2vyL14CGaF0foHdsXONSFV6ksRTTFOySvbtVivNWkUI4LKW9wzHdTVStCxrbZvm
uJ6dIZVLlLbJNjOl487Tv7KZhjCrb3Thn0ZMMuybsCGgvydHXaplDe2SDHEtp04ie/i7h8OaXomA
r2vAJk9qbHfGEa01KvEgL77JxJ8rYR42ZdWZW3aRCZr/3dmrrbzeBtHOrX3pSokTMprqiEmf9S5t
y+iHdX9tg73HpvD1bS5N1EMO9+fhM1TOVIykRyW3zN1Si55wf3ei9GuamcdFDjYPW+RGqPIrS7Yh
ol+yV7r0HLEHS2zbcTjjHYTEptbGfQZMiKicwX84OTqqJcuQ06qiFITYT+TkfcCvBMEpoMbga2pU
qAfF3ihnHbZGLEsTWKS6p0KKrelxFJPcYJ/wdBa0SZ+UABluI2kna8faqZem93It6uy2HQA8GhIY
UV+2Bjmb9PPTkX/fiQm0VVSXc+aTsumWMtkS9Kd5sszBnYA0B7ck2Zl3BctCu9ZxpU3CHvDG78e7
wsk1oAWfkIOcSnmlhqKDj+4n6GRk16pM6T0hVWNRo3st8J2fDTVH9f3Depd4Ix3mbJTgrZgwBkzx
kzCiXQ1PrNcvXemEz4Cl4TbNu8N23AFPs0z1VPLbnvzHiec/444Sq+3EWmb09wDlX7Rxi/5oxGvX
u7b0JrBl7ILEErb7pGAkiQr+yF1LwPk80JMDPRpSS8Y/xrAhWgKv+zXVB4fWM+3MAp1RWbQFRlyu
9bKqSTSZeU9jd5kKZn/E/xJNSlYawi+X99PRjYUJl+m/KK7RLRapwUz4IhICcGkf28A9EIqjDEw0
qmwmFuBbVZyW03gWBumtauICKF7jzNbPeISnlpkFLOA3z6pPLYOIeM74HP4GSXrEi8E2STHDYzR5
8Jz95Nr6N0ulLQuZRoc/RSmJsIwXDI0hXPqKwmi3ppp/bbY5Ui9YYdux7FEdhVaHbh9XMX9dqBW3
qANbcg3RqJ9IA/mviDWBHCsuB7z8UkPrgFz/gs1NnTlzr2qByTmnIlNmzmtJkamY36xE10o1UYmD
boYxROmWb3nm4oIvmvM6JT1OknCrHz4UFI6w4Jjk0UB4IBcH2VWan/1WlVUPL2ZOmLmGjqxIIAd1
KSc1xS2sio8+i/mVEqWEQjwtqMld+JPfmP6LBBvIycALmpS2dHhamv/WISGfMKNwnrLtqtMXmwwV
5eb5K2Tu0dZGdYN1q38/LfYZPnAf7u9T7g2WbB/JUjUH/HjG7MA6vagdqSk2A5Z1phIVl65uhGsP
91RUmF0NB7oSJwmd71zPXFwrQl6LCpay+CKVXgr4ybtNozdqLIyQ3mtIPJ9eLvGOLPy3rsBtNam7
r9BTVeMrZ1dpC3M6CLK6Ly0pVfNJ5yJCula6c7wNWm8O57a/TPJlAm93qv7oeaLP+7Mu9223h+BM
YOxnSmjz5cJCCakGbb6CsvJBJBZYCN0bkoJPSR2GsF3f3xIFWeoGCJBMMelKVf4Gm6ZdCZRk0iWa
f5KlVanFskERzxwoJQQnOO5jrPLrOacMRHGfY1wcKVTOBJtJflri4b35ch+QnZVVD4yFAELi4DIe
r+rn+nwPuJTStkakEqVNOukQsFnNsMs5I02btWtcXfCSUC9iYAj7YpYEgu/jpvuQaKZkXSFAGT83
vT4xlZUuSQ069NLOeOmVaovA8AwJ4V3NKoJJm3lEgfzKpiT3UUGInClX04J66ot1H2ZbbfcW2jMj
f51HDecbYZjmUOoFiXycAGeDMND3kS2h6wySXP0nicBYn2aRERrJLC1qtcW4cJuarSxKNqAqZNVR
vXPBzCVsD4OMZYLkO8MAR5q/mDmUepRuQb0GfLdg/qdrNX+YVyc8CJKvDS5l96MKNbLVjYp8/kvx
fZtxBZLgw8caY7QRESej6Jhg5tRWoZkxE5q/Xa20TqwOvL7gbUGxH/QEFeMDjOO21HAHewNkF4FO
TJ3N4HYSfFK24iWronC7jwlPs32YZ1v9TI2vIwM1+PzydqrY6fpX4QW2kQP2zsyT5JKZdMCWxAXs
k9GOUCTQzbIchIEYjiyPTyl7UBtzIzxF+I76CcrLz23yjMUl4UiIEJz/AygLqREgeZ5Q1KxgsrRE
GnaWn+zt867pe/C1tz8VAZF/qgbMuj2PefTJsvCVtlM4UHE6bKlR2m7mu2V5vcE4pT9hx1Y6SLoz
o4+VVaipX5WdN/JCso6VXTlFnOrn1np6RqW6CuswqgqR8eBZIxWOrFDv2UoH1elgZTIlQ0KJQzpb
BuMhclr/Obs6q4rbbQyKCnYhq/80gavgT8kmnCelmc8EyDhEGbO+Hyoyw5rkcOXb+wJve2vHoUhd
/D5nKi4VSFePpobEtl1ro0FSAErBVzHx2ddOom3Qh4swZA8dBNEgSd6TwgvL2UHAJw6nu6ACCI+q
wsT9jC+NRVro0dV/7fy6P0mZDyLvhbUnRTnS9vtRZtT/g1Q4RT501J22dgjaRH4vpL6kJC2HXtqx
oLMjahBKnCv1j8br3afuSOQ025gqSh492Rij7loS+l58qKDGFkd/lQ5riddLYHUbH5tSM416Xu9B
7sP/OV22oj1TKUIi3AKnyD7M0/Ic9Gb1hW1GENYQcEKW/IwDKT6kECvfEyHbXyh4ouYMUmo+8Gh2
Aiqd5OliAc7QRzRzgn1o9GgE48BbxU0gUxzomNt40DjlWF8RU4bHjPkaV3fRvcjY8eP3Xq/m925m
8IVHzxWCtmpsN/VJ80tBXhQ8AugDv6hgb0ic5EVk1rd4Mwbv+323NMwi8zyJP+fz09Jxnuz1HTSh
KvOpad2covIRvmt5BbM2H7xW5DINnGWjB91EdQktVBRnp1gF5DB6xSpIt95eR+8OMb/zlfazxPzZ
pQY159+ndSFnlxIi+/TfGb/qGbCWoLIty6SHIHmUS6edD2qzv75l2Askt9KczMIkBAM/Iy/4QWGS
jHFMk3heHvJZ7ABwl2eIHjA8kzpgCDIPK/AzYJu06k3XkSHUZ5cQoJyp+Eyr6k/9euIkbphYlHIw
Tpf5WcKiVqso+sB+H31k6yN3mDpVzlIe4YPfyy/ebFIwq4TI+/RePdkIRvxiBgdFlKumAKd2UV7Z
h62j7NDEHKwnTUku7FRNT4tbVS2KoRw6mHGeE47hm0pT9hbAm5AH7IBDlRRyOrqMcA1SH2Dh0Mx8
b1bhk+k0mQHwJrjz4duAey6K80BCBMFmnHURJASp5pur/nlfGjZnGdgkHwpxpRxjG/8USKau7uGD
+/OxbqamZhwogijLnxQI/Jdepbt4paTm6/Ek8f5eB9v+btMcfcGbu/IGj7qtlc87E4QdUviwXHlc
Ysc7KZLrkNuWqn8OOca/4MPu4jgo9AqQnnqIpEczn9kMBSTA6zEqNA9kQAKTi0wHkIjLr4wWT9no
UmP7AzUvN6fCaZ4awbLjFMov7b0sQMaB13etCaB6V8cTt8jBHtYBNCelvgxo2qWqlpjzdS9O35iE
IZjlKu4kFeMQYQlsHhl6iZTWwk7IwZDnPaKcxw6vAEO+ZkNhVPgjjaClSylb0rtnYP3GatCJS9ue
73KjsiNGlU9CTLpAfQGQftFo5sbffodashD6XBR3GWZuYPdoC7svljwJTA6fiSB7oaqwZH5JAli/
kgXldDDkekfV/OIe2EFzU3O2wcmMI3zhODIWSt4uJsxEq/rmELhC6dhjA9p7RRkIc4wyHtgzFWI0
vx8HAO/0Q78KpdUQaRDh9wqce1viPFFGUV6/oLEddj5r1enuyLNuWUuUngR4hJIsvw0ry9PlY+ks
1s1d4uze7cDwXhmX916yXozE9ssOjL/8pvhWXV/wunGsaUD9BkH9VKB3kCT25vXq0Tl7zW1wUgcw
YuJi/ByjlBNPmEHUmQBTIHaqeSxwqnGk7lL9y54PWKmITJdmIqArEh9hFJ+u0jW/H4tWxmkY1IwZ
vpHAN3xXxcyM65aZJ3DyGX8IOleTso72iJJX0OxzNHQexMRJouwd3kKD6pThZsoIV8bjj/ur1oMs
Fokj5pNk8SVaTjGAjYa+RUaD6+yvW5JKtf7NeRWwdbo+lV29TZJOIwgqI84LFcp46ITXMBPwTqc4
2pfvAzxqTiRIQtZuBafQgPmPxSrDfw75jD2GWs0jZ5PKPj0aVI6Z9ngixlYRRHRSv+1wgpSeiIZv
E++sLqPPE/ud+HWlAFKgU4xxb1pua+BaMwFkX9O5NMYwsbcZ7uOFsk5Qte/DrnyGHAFcTUNG4H1w
pFrlKQ3XyqI74fhIeyisBPCiHgNLI878kco01WnRJQRRtqHfwf/aMOlAq/4NkgwiIB7xKznK+F4F
cuNqiZy9PZit1u95vZ9AtHEkAKN3Ls3CIbdg+Mnmth8/EbKzZZG+C62sKa/xDCy7pY7V+bC0d282
l6ZxRswZQOvRgfFFQTI5a4WaBHdYj5HzJx2I2LBCOfM44Yw1I/FdNzQLGyJejGjps13DT5TwABZs
uzd7BCIBVZb3AV1uErgCpmbX4YMF2ir11lw8Fekg0JGLkMLvGBsVnw2dFhRFZXtR99NynnaZx447
/zOslinREOI422b7yUw+VTT80qD8IGQ5+Ri4yX9gSQleZkgnHz0LhGz+zMocawIA3GGKB0rcG/6w
Qwh9aKwq0T2QRejCe9SzTTVb6SLtS4nDMqIHu7cMNSIHx376tFeI7IaHlOEkTcmVhqKhKnIJ/nqG
0V4Ji1yqYAz7Vstuzi4/dDOCvXLSP5fVTcTKtBum/SCC5cZCrQw6fEfgHPUDFCD0Sk7YXPaLgoRK
sEEqB+EhfPf+nMSgP+F8Ru+yz6SYxjGs1KtMoSWUJD0P0D37tPSEuzUS+IPk42bR24Lr6gkMLBk5
1AygLbixQTMpQzgdLAvr3DxfWD+QaO3N0vmsM69vaRwstzlqx36xRrFwcmEYDO8zgWiWiTHHJR01
aDJWVdkjrb9JEpx8u3mnipezkDro/n2NU7oQE6QBvbyRIphC/oZN9yrIyCEV5yH3wbRwtScKPFUq
S9JUDmWaocs6K5b/O7Dpo/VSAoSGki7y44GTawtC+kM2RjPpU+OfMXE/alpw6N/t1vmeBSx4Ox4h
8qpgNltduFJy3Ib+crheI/QzhK8IN3aggPK+0fzshc3fqAye/XxlB8VTcIJ7gYrtDr+Rdc0vTVmx
gEAt4qEqA+uSg8ElILyncMAQX7Y03ylCJwQvnyoNHi1D3zqfdNp+z9ot28niyVaRyh2bVHbTaOOW
WWUHadfzuEkGEl0K4ouePldZ9G19W9CroDKFewWrO8tuhcjYrPEQ2EGmMre/hjuAmmc6k2Uk5Gxj
A6BYAdrL3nxLmQw0uxgIAi8l1io8Des1yWkH0a6IBlnVVvtLJcsFluyyw2ZlRlfak9+ldSUE7E3F
+47x0RcLDSAT2LBG3tWlC86spqNMaVZ+/Q8n4R6bQXBHpZNDtb13aX0t2ZMoHjL5XHrNhEX0muoL
4WwuVTKNRXPSNGAJZJM/iIrMbgUiB3/8jjawW9ZVpyVVnqbYmmzqs2yf8GmS98AMkJ8FEyeOQMtc
aR5XItAqPVc8bK34YZWkTJNUhcgRJTB13fKsEPU5r24l7zJsdeT8Hk+aQVdn5qcNLSjL/n5Vq7z4
Q3gclgOC7yIWvOjLVwvb5wblJzlKSI+mJrjXV1yFKsv9OBbpVA3h7CniyDoyflA217Bkdb0KKJ0y
FnJBbOvbcbvGnmZg4vgsQuoBmAX56iDZuMr+gZYkH6qRCO3luFvTHF+xheVP7PKspkH/twwOSEy2
acQRO6E1z2Yk3kLr1puwMzmMB3Dpu9AW6vkxUZsr92qq3lKNBSNf8leDKGVk+Oa1B8Vo/mwLerGK
0jSIa7CfLdcWlHRf5nwRgcSoEdNSgytiB0QTHk08JXIuBXXFXZeg3UMf+QHWsS1eCJkB4sSbQgFg
T2YpWX8gdIwqbrdgUW9ZQ159MFmHxMwHQzes28Nq6P2IShqXtCyOnr7cypZ3xZi3DjqrBXJuS+A3
jpFqXRsJI9Q/VYUa6gNAERWBgkjc46r9rpYxnfPUWTplA8BmUWJrwgORAPHN7Ax9ExBaUFfjJwLe
Ib/zCJ/5npUhPAWu/ceyurowTg3dXIA9H0aKNpg3pFu7+bkiL7/pJATLASmUUhHb6wVPm1a8XSLO
5v5sdZ3hwn2P5+VApZICocYug81HWhJBkVbo/DGPrem8MyhAU8FNS+oJWzoS94rxkWKmo6gNdEn4
PRS/ikQqqCVRJJNLE4c5ylFEAmALBUztuHZ3CEdaoEGMlMW6GKjmwLmcbvOWe+w6bKqU7wehwwx7
5QjwWEYG+pOxgta6IDmPfg8V4MEDcj7uOgoVWJBMCcWrPjAZoLPt+mr9LE66DWDgoWu/+ZFAIpSm
2hBTQgt7bXTwqdiq/xljiHEgLfSJop8b6Gq5cCylGHKmG9exJxOQhLRaJHc/S0IWG98YUkc2uBsb
I83SOlMwOqMG3yawW6HPuaAEpdJef69SopdrS5/qSBt5CY2nJcyihlOxEFyH3A5zxPdbhIbVHAWf
o2MBayQ9CSk3r7/EgPRLbU+DXuX79ryz7raHlgtxRJ6KDumhhkgzg+4vkCCc4jxy0BSHYDYD6d/P
0L2XU/Kp41YLs0hxM43QLHDfMsBnAAC85bHo16+LMFG7vUrYt5pU3BY6HpCb0vCXdH3RBPj8dfKE
6+9RSGOlvmaF5U1fqKTkoaaoOXIDN8CROwpnae1mzC9N8xvUdpCn5bc5uAWsiF75/83WoOY1k90h
Zd1bqGLet/HBz6FGipkJZnKcdQUW6MC3MXwY09JynTK7C1bT4U5A4oX8KhFlr1LUduGd/0sLQhHs
YfzeSDYrPR59qZj5sfbl/GhCe4lNzu6faI3NIwGA6LxfiucuG1wfJmTZcOluMBiVYJXjhtRBmvzH
DVU3W3DiMeqH+Sgx9QIvIP1JzH8wdtfj2kx2OuFDSKR2vEEW5wXgn42H5dXF7/JweF8i3XFpKTt3
1ljZd90lyddsZ+EL7r2wZikd9GgPEHf3TYkj0KZWeyD+UNsbejIeXr0qFhr/xorFfuwNKrXBirip
LnUPFq7Huu0FkhjYO7i2qlqLdE/xjgLMwHNyDm/gbiYAJLCweGoOjo9ozgHVa0J4J2jJwH/sOkeR
eYcVBOX9ZmKL90QI2ycc83jrNfupFVS7sHBEbIf28aZAnXP9PQ/YBrDHjL/87vDNroHNsW/BNZ/o
mLvtAYpWRCypdrrMoFs5j2a9HbXt/onKrT65V8rII8tU6T0esAJwg0hLQTSNK8kRO2ipT+5Zp9/a
/bAwoA5ljrR4kr13F0l+EglXX5uRCAchpI/Ztjw4OWddna+EURmRRKXLs3GMaK8xtQf2IHJ6oKOn
usK//ahmHMRQXu53tlpbyFvXdWK8ZKGS8NPydtMAeV5QkQL29Yec6ggwc+NXLr7ZXQo/rQcIXkdO
uvRXbSB+EVnRysbP98Q7CkNUx4Nt0te+xGqzretCfHFKy3U0V45K4wDWZhRqQa3mT1yNVX6y4evV
kTZ2L22MqBtPXDS++pCakERWeFAcpi2vWT6Sm8/s0XJjA/1UoXzBA7s6djsyT9rCw5oriG0y5CCf
g4GTpySP2muoqR6Kc85FmzxwHhIWdbw999IzB+kjE6GveBY0xMcm7NT2XVnJNLbLk5Z21tmm/b3/
TLUNcr/gOwyXHwoA8dW4hZbIP/h2pXW0l1GeMoEdkPIvfFBfimqcSZjSHGz0GCqloMjAUMVfG/Ng
Oszaspz+37IpWt5dxI8VX9rDsJmbD8kr9epC5xVgvdP7HDf8TcP82uZdTxGcnx7SlrC2ibqme83T
dnZFe4ArHRz5eb+haNDJnH4CCrF8IhvrmK76F7gXFUmxjEOhVJiLANHqKgvJp5TWECXYHTAOBoTl
+RwIe3ApIN/yUMIYCGwxb8+Xjsf2xs6OmNv+MwiJOk37h4upxL4L6cY+JGZNEeW1XOYHrmw+f3vf
R02uutP+/+OIKSXN3zO3fssLUuapyLKYlpupr+WChg2JMLjgIIAuV6lZOnPrXGEmeN2F+Kcw6VMj
fLTC0VyBi35bR1K5m8v8lq4MS/CHrdAi2Eoh2GdvP9Q6v0GggKZ1b07PwvKmwiZZPexKYY+65R/i
s0tlIvPXvtcqRZER7mcZHTuLn7/FwV4GNzhmDmE1LGdb95DHnRteLagaUnD252vShmGcMhdeEaAd
9UR9r5GDqsiK4T/OrFqEpbVmSpIzziY4pVsygkmRvXcSuiCQrbLQubnea/MzHGUFJgJ4kPspiaqB
GB5nDQ62xMxVQ98SdXKu+ziymIf47xQymtoiOLG4F0V1okFbGIb6fZcU9DpeXfbbS8oOeTeAGSUu
u/7Ii8opir6bzV1bSsPDJcaWNWVsK8Vf4eu9De7QtLF42/gMNSM72EAnld7potQDEPJ2nAItXzm3
9vG0pNSfG3mnZefGsO4vrcUWu2pKDLFCkhKE+ARnXmCqa6A4WWvw9fAyGej69nzXorU2T4OTptOk
mleAtSztjw92Q4YudsJL2CrAY6eWPHA0s2NYavM2VoE8zC4g2Se7CMhXEkCcLpD/V/PXYbpkRdwK
ALqwz958MWqqIfN3FohB+UrHwDH2/AJm8R24Jk/xSLK1mvW8kqrtPgdxuCEXFrYD5LulZOzjdGwz
cCATcVhHmRLB9QUwunTl5VGUTNF3eQ+avtXG/SVquICTWZXH07p/yjZSzxns+pJ8/cFQGfn4dOPq
Akh4kFdukGUQ8PvAHx9rVz7RSQtLnHv3ycguV2rvHWqOs4eEUpRV7kmBe73hFFIHqQmYb+Bk95mj
rcx3HlmB+XoZ88G40J9cu5wO9liCBxNYnalFHV8EG79hWomihqLmMOS+JYq9lU+RmtJP5QYuHVOU
GjFVBTzGDWCzDDOrPK3qaz9wUxxzm84jJC23mYnS4K5YxYGirYayPlXVF2b7O1tbCNjLr95TV3tN
ES8omnvLUeOMF0BKYbxfp6FgDcTBWkDtTZFzSvLJXpyIOVzISIng+hc24Ay6jB+8M+H/UMHRZiTW
B2MwmgS4hfbrDdyfK+u6b+VY0FGLuaFeRfXZUh5U0ViB4Y9b6aZieXITNeWBdsMwaAniNF4hDYbT
whUvD5C5zkauRF66hhIMXr9bkXVMl4p9pcQbC5BwkHIU3PhoUkV7A59y+zEAvBb8P6LRBNzZdcOO
1iFaQJoM9PcPD+0eJQhJ382WgbgDxTDvOGDw4nT3hfYFz5PDmD/0GApg9dxAiwMSqxkonqAoCcJM
JRfQ/uBqcsOif6JR776v3NN5q0WECdVgfAQ6Aya2RSSdFI3sowGyiD/CZStatMqc67tVw7ocQwHa
b8gT7U5z674NJ5/wiJRhDBJkPXzu/b3UCZTkFbmEIf427NLIB31FL996x9zqMPT2l329mnX7TjR6
aNU6tr4CQXoCs7uFy/7XfDW/Mjk1RkN2C6VfYd5PgdRTXpZSaFHxXBKT1OtdcgV1fwB53+oDXsmF
vF5Q11pWOIPJ1za0mLOTkK/gModrwQpAmBF+/R6YbySmBLZX/TKnlM/JWV9k4DxbnSi/Rp3e0oYY
6dTpTR3CxcywVuGnB+LACZUMNW2XMooXb3dpohIZzNT5P5BtqdYCQRX1kTBjvZax2LkOvnEC7uBE
SZVSuBo+8SDD8cc5SbkYOjjOGwSHEAyd1W1Sks3ePfSJ+R4Mz41minvf/e2OxIjZVgsEhNaID9aZ
KYh+wZ6VEqfxDFCcfdGX1YlWtMf8yvQfUj3Ux3cAPn2ztPtTLlg4st6grKSIhINMtKsR3XG6bKHR
rY6jodexqwuMQ9hHj+j9v5aMeQe8DgAqiRYV3LzPSOrusiZnITQ4Xa1D3/D4w+hdFaUxdEo7mCxY
xHlQN4gKQsGisDxQjD/wtDQDL0cbLPv6QY9EHSWCvExhzo4VQjYeHiVZMG1v3YeO4toim/bJcL9v
l9/y3QwQ9zwFMzz2JL6AS7AmVjkfIQaco9z9apQtqgAsjni7IO1WCeFg1Iv8Zq6tjp+l7UZU5Po9
4wLiJl60om/+SmImelkWHGGXn9CXMN3kPeMoJVqR5RbEwuPl+2/JGa6I7dINepRH40KObl/xO2d/
3N7kFUQzNtcVVvUO4LCc2Pm2fJYRl7YHfFe1rSGz08sXqfxOyXIEFFXwtsXzRbjaizGas/PSjh+M
CssrvIjLcZJkSXxdrEn7mU4m/4TO0W0XYFD8qfRlEJCPLM5liOdxuEUhlRd/M87/B/hP/9HoDcX2
w+R68qZkEuTn44VgfReGrl+3gT2K9HRyJelodmTZJiMMewR/lNHn/FAmiz9ApXlhbCgoVosv1H3R
MR0N6qOAgwL6IM33lesmoHvv4CTuyGnY3gbE+gZMXlGNh5e2EJFiRp/Gf7zjKwkRrEhk8qKa5zQC
K960cD5qvprgTD2rU09i36dhAURqJjNvZwEgYrUDoE2AQVlycLa7fCtoZxRswOsWVA2m6r+Hc776
rVY8slESOahEj4+D73s2yjnTdcWDHgVyKsPmJHF80GiIfvd8+uU6gmiTnKJTDmNjldretvWlhSjN
vFY6Gl4pBBkpRWSpC9koOzk7j614ZkZiIBLTSCyz8+4zSO54f9XffDN0WKggbDcVn5N7t0zppS09
e9s+OM39iii/YWrgezxeFuJt61DyXdSbBgGyNix+YiHRrzMmxT1GzLDZFsMwQRhDneTwMIPRmu4b
SluZGVaWIqgAtZardjIZugXEE0ACO8F15VwOkEs7+PIQ46bsKQ1acprU3hjLWk6fH7XlHeTueTqz
rIZ2PCQTn3QC951XIXi4aULH3U7ta5DLc7s8lm03frvkRaGZLNPX6qKzDr6mCw/oQQ7ISqmVGmwv
lfUGcXps87IXVzMd/gfjvHnRa388Droc8B40+Vs7G/ZZTXnrU1Vdhn60outGWX2whIugwdqZi5D1
IKTyspgHko1oV+G3YDAPjF4Sl/YYiTwHJrdoATkcwAqK/6yjfpAFofjhf2ju62QSwdOI3I1iHXBr
gyPJFUxXoG1hvKT2Ln5mmJ7JSNlIwA8USu2QqLMd4UH7sw/geSBV8og6oiWyV/7lqpK8kgg/HRuB
620NrAGxSSsyC1ZSgOTy8ke95c+viQVWNBZB7WY6z91WB85HDuBBnb6KIGrO8tI9ObQUJmrjWC1x
JEpWd0zwAkPTW8L/NJtKJkjGg1qJS5tyYfTzxUvs7pZ9hZWxSgAOz3KupSJOZzEiZmniNc0Ws0J4
0jBeZPYLHDWaPz+pSgUD2TtZ8FDQt59KCMK0dVLfRBjybMN2oYiLltidTmP+o1yb4yNSamLjWE7H
8CkiLWNSUkl91Q6VH8MWCxnxYjOchS2/3gL76uoJFzNyY3x0cg4JsCW9ZffO98WBKrpxN5HMUw2n
Z5U5rtlVP/CCwJzR4WaD8YuZNV2dgsA6a+i8IJPmcusnqZVLBXKVzLamZLCPZw1U1uNXm4ZuF7SO
70xDCnChl0yQy4pKEfXwD74C9e/Js6EsFj5odQwUuiGv3m7WMdhan2OUknwjafZrkqJEugwbecWx
0jRQ4Xfpqv+Pmw61+zssPGI++gngOvJyfa+X/PtJY3k3FEE4zBuupA2Wb65gpvRDnmhd7vNICImH
dyy3GnuPUIpNV8kgHvGKiwwX6zxYEPt1Sd7viy/wbratKQdgtHm5sXpn1Ph5e2zDYTYLHowE4j6M
yTZ7yfzgb38yDYvfXjUYPWcQWi8tUT/dzmDDIAbAJcguoXPw/v93RDsSKXTmv5qCf43KQBe68yel
W3Nla1v4pLb+a7guSAYl6Jt/ZIULnyMqu6SVLzD9x1FV/EoRvUsHEaqgVnq67CEa+HwZRIAsUOoP
n/+SaTK5BhykFb6DYh1HhR3YIkeyIo9r9qnPXQcYzGOOl/Ah37JTtd58HnaPsbu/HZMSYv9ilLcl
wES6PBJPr53q9n+8Ug/Y1fG6iUNpP0N9Ri93fnNjmEV5g+3ibzMeFKmZXSInykI9E5uX63HbE8YM
Hnm2Rx/YcoNEPUQQrZQQBbksqfMsqW06DaO4bxssWJuLIspGdhEPF+iTmnNkcT97hB956fFzO4PL
9faslv/sWZ0lrjLAaJ0WVDwS/QdcZmWQ4jw9NAwIzQUQ5vYf/KNFQ4PePjUjAJ6fZQyZgRGOClY1
EybexpLAf5e+mVVLke/hcJf8EdRnABDbD2ppXhvvQL1xEON5Vm6jyuApe6tZmw5ZGlom8EH+zREn
YJPpHWfCCAZvSTomcrbXUHGEVANJrAnIuObYG50+GF23e4MwUsnqrluBx1otLU3PD9vacHn+Veda
0qCxmiAd1vyOEJLH8mV5R/sYUO6te0/vzdFJRnqIPxMxbA8JCM0Fk1eY5/OAowJ6L1WVLEc2sIsw
gKzcEZc48gBgYjSj0iuNfhv+6qSiSJrvUh9O9oN9P3rD3l2rSmqQEQZSc6ewQ+JIT0PtD6i8NKOp
g8jPdfZOoa5YJOgr1LefT8WsEZB9R1VnYZv0luohuW68qG3Omg7OQsWs/NkK9p9MOgyXO2vFm151
YV+W9r5NOHTIkxqIP+LpwWCOuRyy6l67mq9ugdzxCZXKhjxzM9HSDa5lvhOgZh0zvqDiuKA7ey5y
DpKQYXYIHZcOP6fqzE9c2RMKiUAgXStvgKJOmyKcsoJmNaBs3lEJn1qIbK3CAGAWwIKqSlSXEtUh
t1IvZ0pHUd0muckNC2xB9P5FhqV/Sr+pvSDdOEFkq7ORJ9cBg4zYmqO+wMNCOYVbSgqC/NCZZhtz
FQ4PUQt+L1CCvO8AiQIduvZrr90rWMQUs0usqGgVDfw5y2NhnnOKAE80TkB+7HdLx76zo1mH/RGm
CLxJR5Y+qYXELSqQZ9MRI+p5KBblD1WDDsmrl+TMOn5hMDqzAXmuzRcgakF8jgRi7lqinheSh8/O
ZveDSnR2hfg6NqOcHPLjTe93YLAPSa6vaq6siE4EtXZLrtMBrQ5PdXMh2QZ9WEFewuGJwNpEOuwk
/xWAJhw7UP7pUjNT5vNr6dj9Ks2pzYCVBREpYtoux3rQaQMXw9HVzru5amyHlqzFp+nTtpH2FzVS
ZVi054QyQOIzomkakwc2tY5oXoGC9VOq5bj97wK1RaxkY7yMZScbmWv4pu1N/gQJVVRS1n/mfuPw
eWxblMk7VVrKYQ7axwwWlIEUyCAFdQWucZT1mfpwcNhmbw6hQKFq+XAdgIVYa+rVVjnrTfv3HymA
lFWjzIvZWFEvryb9Q5jUoKk8FbiASCZVsLTLGCwpFi58dpfkpP1owLINSHvQdMozWOB2RcHx4Tv3
R1i/jsKQERNKaM0Xb79rnyQKNanpkqN2Jz7RlZ/LZsfyxnHJLGqJzkjVjSygMtMMHzj+zeillruT
uOkHJWZaCG5MP9SWldZUJ1FfuaJ93CluS5FDnDQD8vCmmFG8oU9ktBvoYNAXTXYrx8iV6PjLE6oh
60+yda0PRa0QYMGHiIX5l9UwOpmcZAvwXublEUtsBYH5LvZYj8s/rsXMTrCsCV07WEZixw5pgatd
P/TcGoMR5j4QIF/I2eghWno/9gDaclew/ZZJoRjU/KCx5JqgpP1i0rTRKNgSlOqiATSiNHIqfb8J
hMOfzoN1N++gJck04E+mgHxb40fxrgba+uGC9xTccI7tgrX7nq4CSfhujRtFFWGIcB3V/9YsqpXu
pagdhc3G/5tKNm8hPn3kLP8f2T9VPLXSYEagJZwA155Ha+1BlDTb88yLUIuY0101tU83LV06pu5O
ryOJ3a+HT/uRok836dxUnHIpxZHRRwrox/vOSUaTY2ICLt6wppISW/MEz4XxfuMghtK0sM9vMgXE
0tVv+8VSmmkWtUqXkaIH6M5bKjJFTl+L9NdYtPo8wjcrJJc7mdB1N460TWI2nhEJcBBD4cZVO6oI
geFVxm5RmCqjnwAhrsdiIl8/l4flXsnpdIc0HXTW1CL44g1G3J1HVvZtpnI1ap2qkixkpaQrGMD5
8m0HsofnHT9n/Xd+psnQSotacY3UettvEJi1B/eWGgbZcqudjk3efEBpWbVQBTkn9vPRjqRCfdM1
OvMB+AH2AyElGrJn+U9cTsQbpRjtAe9cXU7bDj3xgRlpOhIOF/xAUTCoC0fNXi6YqXfZUajDrkEk
yFafDAI1v2XXdBknOyQmDbSuRyLrAowOsZe8N5Uln3ngSt3EzdVF4HtCcrhnDnREhmNDU011YGel
24EVlLq2eVffjNhfbnqBD+AYnrzmvELboMqLbyOAFGaUGc5wcrYaGksUY5+9E2PeE9uErh4ifWjX
JrQ88hZE9yidA7w65RmOMdkBPUn7fNI9i7PqthEWuytejEfo9jUcs9LuNbp1IeETyVhBrfKW51ZF
ydRHENyhZHV3dgdeTxwZMAO+Z7xLVF0yswAYPvyqsEXtpcR49dXz8LJeKNbalWbZx1cr3bCOdaFR
t3ztryCDUzONLa1WGydcSR/noWDcQ7Vu904U9ykHqT0HEWaYklVG9gZ6KWh5tPVJ1wnFiC+sx3MN
SOycUnScUATGVlSUX8x/HzBRG84vCptExxUgzgJq2Uq0I6o4bT9AoGTTjfJ8kHcqmFDGyfQulVjr
BnYj4/BmsuE/+1m2o4GRN3lrHUiJVm0qDUWjRpoFIYTuAG7kf8B6+J4PNUXGMl8/r5Ahm5BSVKLI
1wng49uIoFSCIThl4VN2S/7NnytVMU9WJdjFlPwyBC2jH/kPnHjOhDPio4V9IHTgKpGYAvJS1Xey
gJNKirw9pv1HILnxPstZhQepKZ2pnOUp9yL2Vk+sWbuCqgZPPC5ePDxG4NqG6YD0cTyz+nbpaO9Q
B/kKNa8zaIzuK8PTKD36+3QLcVOQBcMHdGdOB+6C5ObW2XN/hq5G137xxo4fGfxA5Qjs6QonvDIe
ibwKlslV3W0yBBN4iutpNEuWgYQ6iBRhNwN5sZd0FvAHKbbBvvVwfh9+NCg44Di6SQ/Ll5jS1tE8
bgDT2pvXY4e3S6OkRb/hgA+0pJ+NlN2FRCqBfJ5m5o0zjS+e+WeV5F5tJk8blwlkXoc9ogR8Di4Q
lZBlYPkPPOnYMPPJMTaKANLWUt0nSJ1jnX2MCqMgKv2ZH11R64AawqjA+uS8W7mTLLz9FlDxn4L8
sFVGqX7WDiKxifEFKVhLtiWGTO+XLESqMGKoi5ltmT1qxH4wpWBEOAv4272l556sWCAaI0dMk/P+
vuwTOGbVimmsWndFvCmy3qcoSmGBUHJDEtXSrn8XBOyVFIQn0eqlbxpCiAQhfOKzxp3qZDXRsQIc
JObX3BxGisMky5CESvEniyTP1DOlx5FGMuP0JNTNVp3hg8o8AycPGCGIhj7IG5MIaCqgCluV2sMW
ecVyXCKe/HricmCNipjhdIqx+P5IPFkEqE2tidcTBdGdg8HV7uRPFjFxd5EjRrC6pBu7O+HpEPqu
RZhAWaDn6Tu+REQKxq4bkOdbdOj/soSgrlb9SBDnmFuMihNtj+POFKJneZBVmxqr7AKc98PyzSv3
lmlQCiuzzsebL5NfLYaYaoesYvIRWpD1+ZfIj7xzkajTBVc5bMA75uW7BhFBIT/7RPRwSUHagxZR
qUTTH6kJ/O8GsCUs2tOMyIPng6aiGczBYikY+voO2G3VaaZLhwf9rNnpt+uAm5Yoo8ClzcTF/aZj
fSzekjlbXeVfCi81ycsWHmqZMPLvTZM334zIwacrgUrXMpbb5R0n1kdplU83pNjJ3MTDuGlUlSO5
u0VpYFrIOCHCJCreYh8h8wInGxHi2VrA+OHMK2m134kRjFYhOlKj2EPHZGtaTa4wkDByggC/WC2t
Sim/mDAfOZltetlRQpgtx4xKc3bjfR3PW7NfR3qZ+hUxwea5Gb5d9ZdvNOY3RgvSOHRpu9URU59E
Q8fNZh48k3ACWJFO5WKfKPVY+IrV8TpiTBjIMdMqPTrobe3mwen73QiT9g0O7++MXXgk6+Bqb0Qy
PLKDNdJxxOcLs4UM44O9Qg/c4w4yFwIyuFFnuGJzkWQuMaLiQNL9zLzAVKpha4bjO5Fb0s8GhXoH
WPZTcY9roupmn2mgaUgxzF/pBP11BMu2Oy6T4tRCaRUQqHj1SbNo6ZR8uGJX3qoi1Ktr+mcIKMRO
vcie3Hakut758krVMFHnAIV7WfQRajzr96ZRc09v5H11ahWSfHdwj6PQZgk/nfdfaF2NsbLHlpg1
vbHZKmzwmZuWt6nYP81WW/4cr+pH1rEDjIXxNNVkgMYKjQ4REehNYSaLd/bkn5FJoLdJ4riwoaQW
52gfBBFzTtvLEqcjm+SlwAnF3PY6FX+Aso3ipKjQuUqBTtWiUyoMbr6Edvlgix7Qz0zm398QnzzS
pZzNURoqLqqBJX7Uxrqd4A9vEQg1wXvRMx/FnK82P8FSGg/EuF/vgyWW5qY4/8Pc3LtrvFYhYpi2
8leV30LKnvlTpde4OxKjrORDvWcfi60+xLmsJv8VCAmdRI7YMT78Ix2grK9Cc6VsjebGEoRni9AQ
6i9qhDbX7hAzBSg2j5782b4UIJVjWTFxZgmYXklR2uuGiBa4NSSNkWOiytclG22fGP0euGTwZ7sy
CaD9bMPonxLpaKSp50Z4dc+yWCqywn9t2e/yfFf4BMt7i5N06RdDyi9il1eOfK3w8wHP1H92E7X/
MRdD03ue34VpfoyvM/Qfl+ZUs/DOR08z0evAsYxqNpuR3Rwf5K4rXHNRa+DgJxKbyYOdbD3soSU6
9mXAg6iDsiTfrhwm2J4qmTdj1TNopLe/ElyRt5hAVoEzRnUWvs/KrHSOx5hVJKKLoxkCkD9u6zn6
MYfh/DFb63upJ7mavnLoEgMrO3v+Rc8/VDUgJoTemxXjKA3sV6mCyAsy5Ah5wZ5+4CjpbZdgUq1a
mzk/hQVsR4vJtjrljVUVzb3ASg9epgaoeLbkVYShRz8/HivmoonTu9kpjPIrpKI3c3fjWaxFRwcL
ckGSrHXVE3IUossFta7gVzzppTdKNOmyGCNXZobsP0RpG66Bd/SAyVJQsPTdP5E+nNhbmzHmB14l
8v2zy77KgiVx86ntuSipYwFOYJtVsJSFpVfyB6eUyf+1yRpQiVM3ZAn8J/5t4w5PNoDkx5jyY0ZP
P/kC9HESDe8s7KUfju5ttQSZJGa7JWg2Bo0UvLoFlIokh6dCu61eGXXK8bR6Gt/PhtLllVwY6OhP
lgErMJ4HEwg4ZPKTsDbn/7gJaLugQpOnAXQ8m5Uo5psRtZzg4VAWMeI9YjL1wPVpP563AHjyfPcP
dhH84173s9+T2b5PbIfWNgFPEV3P353Qk+sRvTsX7mT5QPxw/DTC3XlbgVsj+shYwA26nGwJ+x/A
DIbv/AcQmHoouNHMlnjd47sdfAYXD0JFgo2vkQQLUP+b8JIFmvyeKMhLf3/WabAzPhIZoxehbjMf
AWP7wcfRQNlz4IQJY8WeB93nLpK+TekNTVDu8TqHAXPxRvK9XJKJ1OzRGP+EZNGeN7pjFMNmiB8s
Ox00Bysx/0NiNhdK9sLEL/ZCPBvVgPMHngzQStrDs1OIzo35pMC1R0zeySN2POQReBCrkdoYDFUG
SkzAys0Oc0xMB4rQPeL2p6fsF3IrIeQfUH4yOZagrXAPu55v69/+4Zm0Qa/RrwX7h70izNo5kgY+
8qkqySTBMviKe14BFO57fO2Bry9RH9yXYhC6WaywWAH/4yWdgkYsM9mZkzVvDINCxZLUdsDKabOG
BWt4xikft/r3ue8yQnVyFr2f4ElAKgb5TeFop53k2Y222w0WhOA3hEb2e5J8bWtLP3QUup/El4HB
0xtCAtGKsvVxXteuIezbyIDOB/N30ut+4AgzePgv11TW58DJCAI5QkZQDTnymZfXNoA/7vlpiwle
njSNb/h3IlKlAqUipEOdxgx5TjKWWbl1VuafbEnc9GmYSKZiC0E83f+e+JeUss1h4aQ3xX6KMJAM
bxQt6GKeBYkdMRmHoY+HlIOPIB3453KXCSNOJZuQM0zKDqbp0RI0XenbpkeGiEcTNTi1FLVLFGin
UFaJqbmrdKAPhkeZ8tW+hvj44CrSpFAstqW9ifibeLo9pk+5iK7zUYyqBf8Q/k/CD2HhNa6fRwnu
VE5HyWatW37yMVfoOntyYo1QAT9dU1NDSDKEbz9+k4HmIdYrPuUyKfEzXC9pgc++ZAX6YIhybN62
qM2wRLK9J1uLVCWBOjrGgzOELHgFWx4rQfpaXvbl2I4rkEYMEXnro2tgKNB7SyV00oxluvKXmuRH
47SmeL/2Wa0FCr1ZOE8gUW2dE81hyVlglRKmQYJFaWgAyCEnwov9a9vjahmg0u5aRF6n/KrXIwUp
hodu+c2lzBoIeeTxA+9iVfxrIoBMWYWIXqziX81rUGxnHLODEqRD0RBggkiqS9RMigLtt+8R2bXD
SU2d33jwAEhNjzeRYYHgrFWbn+D3ZpVYa4v1N1rkkt6ty6tmyxHOpnv3het0fJ+AzTF274uNkEOq
hQ6Gl62bkncYvoycHCn8uZCX8s21Z8XEt4sMikss8WGxOzaA1pRXdaaZfTeBWAcFE99rAYskMWSg
3+rRwNgPtstqzIvsLM9mVeC+maLwwHOcDXdHiAnXqLxF/nQ8Giq2l2DBw7krRYrBSuDKkAeovQaP
K7FLXfyl6Up2ukeu+3DnBQkBvf2+U7I5/zuvhKNqhko0f+AKHZHCT14nVIaKSlA4hsjXOgTCcsHv
EUfHIL92VaGbk7mRk54oq5yYmKhXvtvRUrdAY/SkLfPzRM+jmONREMbd91RLiWMHJn+8jSEQYI37
0pdqam5G0SIHifasZF9rum927dnR/cPz5kV8GZbJBOlZ9Ylus0HYlRC60jtrEfidGgHnfyVaN9P8
ZSFEC+A/BAFHKQ2CJDTnmBHRVu5DgmWpdtTD3uzeCpI7zS40iUtARfRcPIL7j0gLvMV9xSxo+NCb
ZqhIBvjBXdArvGOwJhb4lC0cH0Bi2YPgxIbS7D5Wdft9mcgvbIOgih6q4+blVn2uSeeDyKptZ21U
vZ6lhFiycfJ/Tu+jnrujN+B+16faG6jH+Oc5YcwGha1OurLapR+yZBC5tSpABpE/pJZAkyErmkFs
s1uUtpwkVFVq0JA1RWONzBetVsaayiNbpqx7YCWCEA5s6jTVI8wNae6aP3xDjSeQfum6QY51dC8m
DhVy2aINl5sscLSW0Xb9oAPAvw2qXiHwWf3jq48Jx31l47DSULreC6DEmM+l651TWLBAhqDzAzcr
zeg/9dsNlVmkUgKM1OFcPWuDH9lhgWhANfIs9THfeDHgyoOOb0EWi2QWQ9yw//QmhhoAQP8vocz7
qCXlYy7Sr1IBoPO3ECWz+E8972WvzdZ+jZd57FubbFQCO9P3UnreEAO5/FmsbRN+O+VfIk1b53oa
UfWjYXOUG4BdXeC63I4pJiXcoalXFv3F3CDDW15Tr55yBei15kAVWRPz8+57tQ6W5UByvuqqyJC8
9/YXHaK9syZaSLTbyjflSvfq7bRYb6Tzc/xi81bpXiEi2CzwknaUmijxtv7H+ePkYF03Nb2QIKyY
1ZDIUcmaGoUtYzuF59XtRYIAKwJriPBehJQ39TWrYIqKtdkf+/bgzZv7Bz1dtxjJH3sQ6wEerM0J
asVVumQ/zjTNydkDj8Id2ljxdpOQrWpef1PlYlXu6j0+SCPNdA2COZVpmw/5obxn416EYR1MULuT
QvmkXvG49BmOIOpqtYohjWfgM0z236AFGSQgAj2qFsqjeSk+l2IdjFQXwTcMk3FAlThiKecRL+8A
xkMeHCFN6/JLLeBaVYEBGYS0VAVzIDnYLz1MPRLxur+QEXl09JrjrozNt0p5x3jzSksNtfvG6abh
8OdUBm80RRzFrzSD8BU/y77ZuOrDvPn3npenh74aelqHB85K5OVr66dnwJ/mgt4oDL5IUtNbEwRD
76tJk5AsjsrPekSV7yFu9iIHLM+QDBuDgnWofQKJfdodiz+XhPgfdhxxGDyj/3x9nB2ApJAa0drz
/46DlN2v8meWz6gu91U8MKc4/jTuF69uf/KQjbgIpzd6A+gyMxAYwmkWlz8SbgXjIoXi09StNM6M
zfPNXfFxhahE0gVUuYyXEFuxoZgyNwrCxzDxqSklJ/xbgVS0aIQ6L8BUGEz0EZn50XTx2piAx7Ud
pwMrIpcrHQYXM8W3O/ug3989hzmJXE4Fs3jiq19cvA9xylV/sw3PkBsK/cl+ws5Gzpc7DD9ozprD
cBwzwSRDYhq7cIT1FucxJeN4Dhdb4mbJZ0jyKQ/T21YAkbSBzbdek9XnDHAsexNp3LizaL5/Rg3z
sbOeM4pXp/69fhdNmcyRUWi+q2/MpxIeHvCffqKD86jFfROU7R+qNLdbVMIV+WeXjntyAvY1+aLZ
Dy59CwNxMZ7jNQwnbhfbyzbEFz1YzXA9Br2kJ+jUEs25RuEL9nl4uHqKFdBO/lG0vMAWV5CxqtdG
xHr0ByLIZaw+P+ypAA/b7zO3Y3Bby2FnxpOaVYLVI8chry3qdpbK1p0oOXEsg1gKIqURT0WSun5V
queQInWBivvfiD57F0dC9VHFApyyW1/pWMVM+9i9vK8pys+3Ff0zppWJX66N1nXEx97663My7DmK
soOxFQHcQ+4WAhacSDP/B7JriAR/g6bdLuy50t5FcztmiOI80p5XTeo+GzV+qD9VpHMv/xmmYxLI
21J6lIdNuc+b34rbBPkkAe7ED1PeS0QXe4EXVTO9jEY1TNgaGGniBZs8ZZzB94rlnFSbu17uuTeQ
+/OmbwTJhTrI1Gee711D6vLhQQ3R/YUs1fth4qD4b5nk3PTzKxldxvL/a/IUGfMVz3EZT1p38on+
oo4VsgFdQLYZH/grGyeq3dP33DeCHB0B3YNYgo1DknijbvsrcfZKjq3Oh4c5Ovi2Nrkt7t/SbBV8
EilpehxsFIJSloxBViZ1V8Ja2CHKphz8VogmmAFsB2PiEPsANNxIWpKAq7/cHXDaKvaAEaW30uzH
vFwJilhrCNDUgCcQeoLGsBk0ERiemFgofqmenx1EVSYrrIwYfhZSnFWzJXT9iBA1gJ57z4xRywrM
wZ25S/3Kev7sHLHFmjGJFEsBpvI+JTnCZ/pVhG+v9kQZbxbI/JJ3YoIcJ4tuyk27TG6eiTrsa7Kd
TcKJJmBhjh8Ox981iQg8Kd2H3plIccnsLaaDEMOCOmlgDjhRGcmyz5xk8Uf84azdykQUHSzweN98
wQghr5cmW4G/3o9jAOzY5yBnKTPQZ5l2t3xpDXWvpXeHEHQI18ThiDA+688bKKYQyeG/XPoNT+Tk
vQReEM5jL39nrQ3BLcG3dn8+tVeWV7CRDCxgkjc7rRGW28zIIaQSSxtfudR4A/UE1pMVZ5jOkmLE
UkVnHCj6ZGbmGYIbyKAFir8xYGgpfY9hkSSe6+EfT0nZCwJakzptMErt41FZCjsk44Cd2EcgvTDH
Q9v0lqEIluoJ+a12ANXYlefc+2tKbg3JaN4eZAg3TF5T4dJNdH5oS1a/8/tt3cmi7y2gvxYBRdOI
pqwkeiOpO/6ASPl39oL2bolsqZRwpDXIeozyYshK7+BKx7o4d5hDZd3IeLolPNOEytmf9reft1lO
pxI0mjsK+5AnnusBZohlso+SKfO4b7bY3qrdj59YSTnQgR71nz9fxXMcK7OO8vd23yyKpzqqb/jh
vhbLPMgn+nnKfT+Yyc24ODU6LeR+qXkKYzu393usIs6QuMacm4p3+WbhiDzHhQJ9GerTQwlfPBWb
GWyY1vMPBAG1W8tJwWGh8W3pybO7So6LCOM3YtRgXW6M8qYB1dcDBur32uOyp+nf5pRjdPM8Iv/7
GJtUWI+mnMWmjoNLyv87JJxKNGteNTFecG0G/g5yElgaYjg1igQLasrw5kEAsDJkS50oUWtP6dl8
mZ51ivHcT3AQWE19AfWTupbal0Wfw+64rfkq3NbUDuryUfU0A8aePHyLd1B3uI0CqZQe1cRiMd1A
RuaAITBdRNjLhxJgsB9tQAnhUWrynORTwZx5L5vzxdxazczGlPC4wRrpa+1XCVwcIT2T1pVkhw+4
9hfjKQXJwLoZm864Q2sO63zSWMlPkv8XOc2vaTGop2gcZ8Y5N+GGXm3ccDb1k7eZ5MUTeop5S66P
pAFU6ZerF4544qrYLxAlOiphDehbBwQWFLYKoQDYLTveM7MxLy6LT34kPzFXRln4FxO2VbU9VaOG
SZGmFEcr9xwoj0+FkEC8J0INL/gsOPi756uhYk3wpDbQsBO4XYKTOqJnrDdWqmMrBCkXM+7zvNAw
2afXVmRMPd3EUDofkoIXKASAvZp7NcTk03PLNxNi0ZyWqkKIME3WVxzbtmxrF2Lsj+MKJlZpC5Ot
QnvJuCog1t4dWuqZUOvOhCDUKWMPm6UgWCdBKxQXmXu+jbA6bVd46fRH4QXKzTgClLoPXdl/Zfhu
xmLiWfoqXywxGLY/Velg7Z3PrvtXmycAekSFNrFWTUPmYO5P6RUgDFG8CWF3C1vneFYJo1J/YGNG
AVH42Dg5GS+ljGvzqd52g9JpKSn54MzxioLSmpZ0FbInnxt617mSx6wnSZfcp78YL60NjN3NgkQr
xI+bhHRr0Y4wMCqpIJmGl8onIvM9Q5AvSSq/JqwBPn7jJaq5yCz3Sm94KreIA3LtRd8omU88DLH1
mbIyAi+pUj8Jjvq18Fj+R7agc2eh/Hlzb5zim4ZgPGzlcTNnAIhdsPRJ6oFfXrXjLJNCRIKWwRtr
3Mu5Ijfq+9x7R+djWFyz1G1W0DkSGlU4d4YfkXlzFiSbVD7hOC24TYxvurHS5JdbaHv0oIXT86UJ
3enx3DYqNlgK37RgsKMlafCAHXtxpk+qhpjjGbv8eXvomsbplUPGJh7HFcSuYfxSCrmkG3OmeqBA
F/hWDeQc/ylw3mo6wiQhmbDc3ONDjbQtaUpH67GzGpr7IYGdVdDQM3j6fZAitX+68GkmCHbaqeE0
sxMb5aT4pt6c9buVL3ym4o3p+60l8zeva9yH6twLl2rnpDyLPaBLatXcmnUeck5MdxZ3onusnPMt
BY7WCtMmJ/hMRus0kM86JaopCBu7n7PU4sTuxT0PerfWJ+c5zmkz/YcDDYT9QyAVJtk6jhuh32rG
+Gkqwk8vqSEBc83j8S40y6FEPS3PCcU0jD0Ctn0xz+/yI7FGNbe5Eabph1lAslF6o3pqTVUfc13T
qxhuVlsGjAv0LJfpJS5zYDN9WX6maopOCq0gNKR6ltVr2F2HvWGlzmhdfThRq9xNE5iDgGWUzSqF
qVJuhShdm/idf10/Mn41AZFTadia9I7DiKml6h2OeAZXPXo3CC7kWctExk9r1UjBflGOx5BFgXBJ
fkLJpAwOa2k/sQCUH6JxDn6wsXoLUyPYdy4mHxpGvUWT0kMfqWgzM3jgA0eT1N+6YQDa8HO9S1DT
mI2aDlD+Tfm8FrLSGJqPVCYrDg+sJXJPnfnNHT1Y1wzAPFSeUi1KrWie0FMwyoXXiGnf796VXRmg
EThHd8R/yLWfl1xkMIjSwx3EaxPyAPOxJ0upQTcKD9sI18QDf/P6GPdUug6e7wCeJ7oVDhDXIOCd
SqOYmTOsgA67UXNx4qUyIu9dVeTuStPazWWiEnWIm2zxahJDOr6T01h4v+z60QPGNqVRUvFO51pM
wSuNXErvj8lUFv47rKAvnx6zhQ0dRNuw43fIf4NLAbf3JWZuYh+oY2bo4kaAhrwCmPR4HsmhAgK/
e3hE/RvyZTcvUm5droDFegswiyWY5XIvUDjH8TLMAbwGMC8oLOvKH87sBZYP4gCRtwjjZjcIjgjV
tg980U/mr1d5g1K2moQb8ifSTsGsrSgRkWV0vetwiy+/O6rtHYn+aMuLQpX7sZ2MKiwhIEDKGUWN
Rh8PsuH9ecT4j0fbIWbAuuRpyqRlz0ZlbVqAJpBHdNXdJJ8UT6rrhuiGedbV2hu4TGu9Js19H3+P
jcyhO0GF7xwyC+LPsSGA3ZSWxZ6mA8Xl+Euikf6hUC5ngt5wRP0cC9g9Q9EFyGtSfNVNSVAfqUSz
HgxcwRiOGxaEn/V/NLCchIO60x2JbQwRaNKXG0YVqd1VJIgkjCUadT/QU+w2mJAc07gkAu5Je9OD
igoJ8tPohfHPWyS84LW67PTMgSOy6lu6H1iJ/timgkCOLpPrJDeieWBNK8RXnwjDS9Y+spnB2pAu
wZS2w2qtMC2jqaFVggXohJCzSHqsd+SSA3Qgdiu9Pkem0Rs2CC7WdZzE9DhIVufEFu3ZsMG5xLF1
Fm/fMlRABwLvcF4hJw8RxL3L1UXSy1cFbJ34qunbdbudDATd1XL7+IrcYykE+39kt7cxVp6GKvbb
po4niGLSjr+w3cbXLK7mtezxbszEad+wGi1kp78CL+aDTV696UvD5tvVwHE+zS26RKZTJMBt00wi
t07tJIByffyMeODf+V5nC+Czw4NeJ9p4odAo2ekDtLSdRFu+5Q2i1Oz7XvK/5IABO7/8RUwOJw7X
/ACHWfFyK34OhF4waTw7K9e/ndpi9h5PseU6b+urS5hUO6YpAEfXh0hdfOIHwl8YCLvQzcT+Bh8r
fZGsNfyZ93t/wbbMzzzxTfNn+wdCHQWVUOfYzOkNCTViCVb210dNh5Iznl9KHYAayK2f455w9b+s
BEJRcNboyxxcwRLzs+DzU540ao9Jt296MFz00NpAyABH0worRwMVhb2VPNS6RATLtwR3+T8QSBM0
dP32EuVRCIQUPoI6UC/TPHEY7Q+Ue/9PRY2N+j0hvvDG7QrWz4p0WZfjZnvXky/JF7MwQiEQFFZK
ob1j4IF6VyJJWacffo9VQumA+1xEOGyAkJNPD2CiEjXe3B4+nzgMjJFqvvXydXDnZlFLNUmOWac6
Y3EIMRUc8LW8tzQqg/qaLPm0IFnawBk/vw5osAEp4PJKNZihXSCMXYqFwb0RMyRuMPg+pmq9Tt+H
lFGY8mzoVTrluwg47wzoItSKSFrTHNW3IEjI3KQdisH9nmJj4giWHIiDsQjq4mvjZPvIckwte4Cf
EcB++UyVtovKENaME6g+qq12TbHpVORXtY4QyxtLyMhM1xNbAlHrpufj8TpOc51LgXLNFZPlnMPr
vJYwXThhCVPn+HTr1g9q/ML/Jf9Ij302qkGl5Y0r47JTaaaLT1vMU9TccGQR+3ON1ijzYqjQypsn
g4edvHDm444fuUE0TIC7UJ9DkYL6tw51nDc8AgDE6sMED3Kwx1ExyixquUEoHHoa6FrmJBjJcNpB
NXRVkaqf/2ftQDbBhVW8qB2ukwG/+E2yOdgfiT28D7x2zM9VJbjfrcM6SUKuDwqjyPgrHT10FfIJ
c0onWL+p2Xa6ZbtONZk0WKrJxqrs8uAwnygfASyrYVzy4JW5FugS2Tqp7W+XP2TtGplSuIjd7Gx2
ASb9VuNoMtZn3mkv7KCKrqn818l8Sj7ltnp9ywrG6yATyxBdAyv+FSfL/BNecUoCBUs+iCTgoE4W
PEw/uDZhcnaK1sjhMCILOmcWpFPCzaB6K7qbzOs7Bp6rGYNGbtUD59RITdrb+wdpI/3PQMf8w8hJ
fqwcjegK4tggjAF53wS2VE5Z9yNTLc0nsm52QhvkFRouxOFxqpmEvawuULr/qIOpgcg4EUjdRLkt
Ma/CQzhPqAp3H/Z2e/uVMNCFHk1HtEL1NjxA0t6HjmIgfBFLsvYA+1f3a6UR/PICPORQMdf+567o
n5Q2zmv6k9CWl+JEGvxh3TpG47DA/tHklkek8/ZZKkRRSj2gyaioB8OtP9VBtku4QQr/n4kUZ/6e
ZlAUiORJatKyG+fb7mLoZhah1LOUOJ9p+kbeuhhOg9NP2M4IhbLUXbKeV3XlZ0m7kMkzeBRi40An
XggX3Bc/mXTQ/mM78TTH2Wo67vB3096TrE3KjUZCUEs7J1vFH18zmvdfraGEFS3sW65tkxcA92Tm
oc9ouVG7PkNF511WWn2f3YJM+hNh6UPms4tbT1maF8GVPBPHT7mGHDWsJfwDNHhKUUu2yQ3cJaNJ
DLLlNvTzAjcHir/1XB43AbEaMObYGju5+AA3Lu+h0+CitUg54Y0RFq2JebbkJItKrIpdapbGfs8C
ZY1nqXwINTMBaxWN65TcdoEMWAR7P9fcMst9OGuoFhM44llQ2SgG7WFbAOzNiiMbWTEOc/q84vv0
3ZRo1wXzDtMECBARnlGhVvdjSiBeR5SPxuZf++eNd+kxhM7E3UcgAs8wYb+5re21/+Fn3FZJVrva
EslvTCA/+8X8wOYnqtvhXASm5q8yKjeRC1+aeHUQJwKTSVLhCKo3uLuikAiOHqSGpzDBPcJiKaoJ
QbcSNzzbtVoYYMgQ3IEGGXXZwf769dUCKKe4AULLzFyCTkvsIlaLwbrr/lIwKOh4FjMw3vlxdYTD
589t1DtMutDr1Gc+7eRg6dfRrC5dbRYM6Rh2ee6dd0e3CDhPzXL5/E9c6bt5EFzm2JTN8sSkvhHJ
JT8blgtDjRMI0mN8W359zk06tbqCXORdQnyWlokrmQkVv1uUu5+PJsJQkdPbWwdkzFKK6Gp4boOs
GeF7n7HVKoSpNNUehaNU4M/zT+M/+Ipi5NdtS+kAVxhC0sanpxci0FYVTUSG98mV8lmlD2Qr4j5P
3gIEyCzBJL9yVUI+qAavUmGYmxYl9YTaFpO1FZK8Jq9Xn1Uip49wJRyFOA1deDvULc1Xje+qAjk/
pefAEdcR9ufioBC7MtEDZPtmAc1sivTcjlu/s7BzlaQt1smGnqBTCp+XvxhWSHCrvi0MDVQRDKAi
uxoam8wJ3Vcp2JXLOrIs5UXGxg0M2q2CDgp27+pkPpk2G0itqfjiBdnINRz0hficdldz+Ey9iwMr
BtLzFaDAgxJNov0cFiYDxSucqiDLC2lufOuMYThpJea4FxLHP7GDtkqsDyH3ka6FyFvtAmRtAOk8
XTNj4kAhc4/a2hpzfarP9EltDf4roCVSZ5ee9F1s7V/SY3+sDbGrb8qo+QbRQ0F6tIboDZ8UyIma
skeQp+3qyLp/uDk9roh+mmlU8U7trevwwRkpq4mJA4O0CARNZkE0uVeg7nW4gkFGvFmsMZkWFGji
OpyDT25Rd0vx9khETqHSwNithktmV9zWUzbtCArAF4UeQCc7XgPVY5LKveF0qYd0gn67Qt22R89r
WZyowt08S24uM7WCK3YJFbVXhvg7gM+QrjN1pOPFu0QJ11WyToG9rw7nWOjnZvSI6qAj5UScLmGO
J6v62tBeHeaVsVdGFMn86UEJwu1WftL3CogiMb+zPldjzDXFxQf7exIAgtNA2xsKBjtV43i4Eop9
vpTlVlWeLd1ZjW0JKNMA3IH/atRBL5p3Ovp7bziZ+972jEMkuUXwP1IJQSYeZqb4JChdOgCo7A2b
ex4IrrbgT6FvnUuvQSjGh9mdkD+RXSFPlIwL1/sC8ZjsxjhIKkUD8u5+RWxAu+bS295HsmjFQn0d
hmGY7ZR4EPeudEMhjnsZuqi+UIvU6Q8TkDqoJN8y4XkkYGN9WYOeU/frT66J9Bjsy2Fnnw9QmXpm
NEFhQaSbI3lZt7ohaogR83ipt7JUX1Y8bKjnzC1+ctpVGD0Pii/c+QCR0gm6V7x/6yscYAzqp0e/
wEyUinR1eoLNbSqkqMdJi+i+CA2nKJ4WrN4ghEP+cboddXge4CkUD6EMya6TsEh7rxTwrHl298zn
hZIpDg5g8ET7wLd0bIEM0+O5fqOk4W1y4LxrcCa+fyQpdXPx4FyIFXzOMCYEDDbMcTRvO11nDLU0
WHfdtDP8CwcwYVHPR+XxZKruqMU2crEKOJoiHjG/gG2sKjnozA9GM6hYDVgcS/5jdiiZPoWbH3Sp
R/nwiS38Lt0kw1MqxwjYaEav9WCmedzvGaHuZXzcZL106YSkVKNFHR/W7KLBdr6MGi8enIQ3LI0E
Kz8PTNYkwNWBnTwWvOM1MiHKil+LWLAFif/Z9JGOJGeCvVQiuV7FlXk4ItBDD9JQN327zbuoET/Y
Jn9e9hlNF+iaeBLM7BiHMJHjTmwaB52BaSOcyx4SFcZ8VNQQYY8bcpnUfeJcx5nBX/r7lcgO5xJA
keShEc9JMxd5t6U9uvE/nBMJrDRuU0h9kdNrLT/EqB41s0tSPFoXy/AYeVORKT9RKvNZS5exaI+K
L9Wmvc9ErRjTIsvyAkxyyDfIKDA8TGXEbhTY4yAEVptS78dndvkItRzU6KzLbNByQPdvmwO6XlyT
8+dHBMb6qNNLdlRJMkA/oqe1dk6Vn8gT8LUA3DGjUkqmcoWuS1+gXXi/tG/JQIrxryaiXN2SdUjx
ChcUorccbYSxu3FBiTKb3MDavWDO8mOVXWUwDaNwUpBEfCW7Pq0i3/yFEDIOYTOpTukkKUoZbgcK
px4uUJgeHf6/o4m6kWbpAToCnE8EvD0m4DcuyOiHPrarDM9ytn+Dt3Stj7P3HISfgSUuYt0H3bol
VuKsS0k5Q3mopuIqJ4ZAVkhyJsfb88/11KCr5dhZntxdZxoMpaFhCmzf2rYDZ7qr9vLiuAs/qO4F
3ug+X37hLzFZfxbnyTo7hY16hr15oz4w+4+4emcuJZocPr41PLe/PwoTsV+HhTOpLU3sWD+dZ3NA
LRb0zCIv/sIH/fO6nQGZkUnU+6QJGI2XstKTagjqUw78/o3fRuwgLwqRHZFAlZoU3ljtVPL4ESEC
2qoGU7bUObmOCSCLum5OTOh6vZ60Qh/YEDNDnXfGH6sn/T2/OBJiHeiKgFCR2PIw4YzRGWAPUz2p
Gx9JDbRJSXpNDAML7NQ9hPdb1iYaBydpOJ1mCrlxlbmuwKsPpITF+8bYBEb/SJXd3ABk7ldDkRiT
jQD2mehkKuf3RvLuv5+AEGqwxtI/1orF2tK9kNAt18Gq0Bv1KJ6sHRY4g89efBBt9AkUP0i9VaCR
MCbn5yzJSGHgTdtjig6IKtUBamQQW1Jisokru2KJVy+YHoOSoNEGoeUcyNej5sQYPrmKM2qSFVYr
Bj5T3PLtBGYIXnTslrYWNJEv0lm2dLaxRb0dqLc6WUecgfxm2yakQLBI+qqfvpdNVm2V8qTr6+Nq
Vm9mzyA7xNdEWopVxfiar/DQ4nmeLx70NftBFO69IMEikQ7B1YuySTIM2qO9aY+A9Oq/FKjPjOf1
wLMhAV2qkEzCgo4scteN3z8eIgLHh72kxHx+y0UQOsiuNFZuxeu1eZM8wA5flrS7MUTSw05C29wp
gdxJ1nKpzvmufl1/nF1KKVMDS1eQmkIFUUBquyf/623w/guk0qh1YWpxYYcJJUeTF9I+Oaq6L8lV
DrUNfe/6XnCjtM+8nzaNwcF+r17jXwumxnTIcqTfXAhEzzq24AqprUw6mzM2kcDph69NH/VhIyn3
VCC+RLH30Wehg472/+zq8YpAlaZ2JzI5Bqac4Rp4D/zjBHiZvgv16fXjsYrXHOcb0tfwVxgIQ5oo
6CgWGRdLZ8SKx1nGog4FETQa1XQID589G3E1Ru5VbeiMf151PR/PAQFy0Q2tAzl8Lb7xf6Ef2RIy
VPzjhShNeQYj73H1hm4hSeA+p4Jk+M+SuwA5XAqpbP9RsujEC6EqSLaW36U1YHpKdwYiE1HgCxk+
KDa2srIQhC+YQZfPa4GAblWtQT8TchwqVmRxjTlX6D8Vs+JQHMdBIjYJUhGl+SuABX71YRppF3PN
I++760pSV2GfGKsUd/nixXDJzygKsB8/6blPZOaNNf7QsKqOQPI2IvtgV9Cg1d+fA4d3Ncb1Zn26
a1ts6oqB3sYdZJz8byhCx/Q/VYE0+oyn+Q+lp10IUZ0TFp0iUtrv0bscyiGfgTz4JHmhsVdudaov
zD2O/phuAp0phLI0E9iqW8DPWbH5TxGj/isW4Jsrrhm/+fcXMEF9UKJHdQVFraaaxmAywkrwSSDk
w8TD7CXv6LvoMMl2kRCy35BcFS/gbrLqchT71CMj8FfPmu3qC+91EFKWmsWDm3M9gQidTnwQc57t
FlOfGR6loc4/KGaKgJSbImyJRwo85FCGRKkqkYQ/7gQxHv72UlyZKJ5zCLLgbv539Rge+uYdRLVR
lC88QV6QEHkvF1EeS/YQLkRbbzsWTYpAqHPekLEkASa+TOuNL3udoF/M1eERGEadIMs94K+ieHu2
cwYo+0fttZ7hqZYrPGSO9SeVwHliVMQSOqu8sPOCD2bP37ib46J9YmmNeaPRFOa9aIYjuDNkC5rw
qbrhv08RkpRNDRGiqOPJ25XAP7KTpUE57XoQ/Xqn9/CfgNBbEASnsJY3rTz2Lj0nmBT1V498+qoA
fmDHCaDLEmBUDMRmBun+8j1Hy/jQQyFL9bXknMWjB4TV6pNDEiYtITaWrF7FHJNfjPsUuNjEXJm+
zFDVNA9VhJZcT2cF0SPljXGT6eG6AdrILSnY2zo14lGPMR6JXiE9kycX+MlR6HmIj34JrwBfAkvI
Wq9fDxRY0zAYdwLBPJZkCXqLwHY3tyZVfJFdw1gewobVUvXP79OkX81mRIaPiU3/ADeVtQqz/vPs
WpIQvf5RbBEErb3aQVPb4uuhy+pD2HSRQOdd6Q8xs0xupvqWpZiffJVeA1L+1XkASUlehz72aB4q
k7SEhLTFRxKUAiKau/RwvxXGgTf/DZErvkyClCltIzg9Q8wDM63DTddXgUvN2IVTM0O0/k/CI2pf
AV06MJGTBUo6bD/tCAohcXRUcZKW/3nUvl0hm2+I5aIyiuqd7qdHIQUcG25NI5aILJGjSl36fIvX
HXtJXXEbE54OsvVvUz3Wg3QBZHm53B85+1xPSkUbk3kho4L0mpCef2FP87Scpvn2j4Ttlxr1qQNR
BhTwOpr2/cWhLgEvt+AkYj8eaGC6J+arTfH/huGBsjCeg8yJhizkhxUbcvzHArAOZBs1SXjRZ520
CN0bxSIig5DFq9TWbaH9drHqoQ+yc4jvrBAFb2vtH236yH+ZVQnZFNO5T32yeoJwWUZnYcYc5+Jp
LSjhhxTl3R8o8bz2Mz7lLjD8Ujo5B2VGl/Oqg8pN2ZVtwmoBDqLgUXW57Pvo7s1+rkv4Qju0SNV5
Q8fIjas1EqDuINQT8FtWVeywoDAmOA9W+awHWLl0or4r3ctnQSxa7Lq7tVxvfaJtkjgUfdfTnujx
BFiLUeJE1hfgnhiII7wMVJT1uK3AcrW9/7ctBldEH0GMVM+nfz1PM/Y/lkRtldGSxJTpbS/JKMx9
PuLyz8sm2EHNvHElVpUHL36lHRVhBVzxG9V5YiCo/uqMJwDsPl6b9Y25VGxjRua2/40UUBv2DodL
saQcpWOr98OZMQlFPlcJlgNr8QmoZj2T0OPbtfeIdHc5W4rj7zmXQY/ynjRRez0eeUH4BjquEOt9
wDeYx4O06bUvxXMyC/naBMkNnDI0Hww5xhLarSK0Z1Kb3VtVB6Jf5SntA2c+ECNDSMk0MILhatJ3
0BYzmfpix3JeiNq8m+KpBRM/p2hS1Xxm20DOnekuAqY53UmOJi2fx06PtiNsxUMTzRtGqOLzqs9u
dLXss8VVsCVrxj86c2oqug8kHPAGe80V0DqBGnUPcunUn6bLyKL45fkfNyZvadFR9+yEgw5Qlos2
sVENEXVi3mBLzvnmi/Vhs32q0zsbYO0ix/ThfMo1L8I7MnlFDg3j7pd3eqI0JVHJxZGCiNFnncAo
HxBrmziovU6AMYYcPzNcrXps9fofBWu6wx7HXpeiHm8g7iVZBUrnWMd8NtcQBtuJb+9JQuA6JYJF
tPcWKEpSQDBBkcsdNJ/HVMzZGwu5i7NkaIbuFpcU3gm3ILSxSm04LFhniVmYntFpNtZ8ojkqem1I
L/XUco0z3WhZrsnyxG6fkyWZ00RamnNTrM3p8taGcGzJYkiVkCNTsEsOfpt8j+FgP6ZOxQA+XuEM
Ft5DELfwFSAmuMUkPJG+baAb5kpJFmx4E+FgHmAHNJ0v3DkCuB2lwgPRgZnIO0GF8a+LkTEtXOdi
gYOy/sq4Y9UKhwLKii9MJ+pzJ4jmV7hff0HLr5uufZ9TiMjRpSDKavZxdFzm5BGFTHKee6ydHLHt
hrciAH5j94ewY9yHmMbKm+ig0gobI5iccK2aE/WGyPMcJeMsmjOe8uREIRqePAXORXx9rhHqylA9
OjZitYbsdPe0uOpA3NfbYfA5OMHENwkI4rAkZcMW4oMPtnb0Oqhyf2eKgQKgSNrj97fbiyHgkpIP
YNxKzhOXqDagIH04yqxew48RIt4oo5B//xwZ/wzLYOtK/4yioqFpH40oUssOTNJrA2vhRs41dEWX
t5wGnYJ9tQsDtwoSVHE21fJMXGLy+zBOn+xduQ2Vuk+3zpi4haRviQBJdZMOkw13bAwm9Jv1Ls9d
YkON8g9PMFWwDVTWM/gJAolxyWEcnVA3sWg9bSxS5duUnlhBJ4Ys5AiK5eafgqVZEc9D8yNbSs2r
G/Qr2jOlNlLY5KtGaVVty2zf+W5Hzt1qjLQw/UysInCFAPDEs0F5d2xZgIQ9mfRkWv5ni4MVStVg
vzNxUw94HdQ1azE60kyIHEvE0YH8bDnI9PPVP6iOPs8o35puO7Q13RigPOOfVav+ZbdvLDlaM16J
4587ekPbhfXM+0le3yVFl1vDPsoZrxs9CyJCAc4VKrdFq36taDwlKYliNbF+IEbs0mECH8z4EodI
raj4BJPARqAFIdxFzPZNBxoNfFMc7yNdn51S3FfrDLXjo2o3rtji8KIp3nfsjalHpCqDx0f8x59S
v9mdCrWfsViQ1jCf5CueCOcm+hcSZxgQBQTiX1jsVW7Qu7HOT3tzH2bOHERIpwb0UGmS0IX13gRp
FlqkAzxhJ+KO4h7VfvqrPfNlhixRuqbCjmPlaw4nF23p5JbHTcvscBTt1UXS3cxot5q5uVn4Etbf
1cj1iEGc8MWw1lkKGNBggX3wdAh+54Wg+101f2czbbDuCTFvZTJkxaoPWR0p+Pw5LgUMr6/nFN6h
dohq1vgHVlZ+LhJxHuH1uCALOWj5A9RFvil9xh1axd0eBDv3rA03pLk6DpDg/AybQf+abVPuWPd5
yqQwT2vbaWXZSrfS2RymYlae4L2K8Ly4om0vY6RHknsQ1tBdzoCA4U97UFdUl4c33d+DgoAz+LiJ
tYq2o1J0kvn6YcbOZcHHMORt+Mb28SFdWrefEXeNd+xRFp0yNIb6VoL5IY5PGNKm/ZfvzRO2pZ8i
ZRyeajSzF6cvTR3C+z9Lj+ZWxxq1dsaTct9jSloZyb+CG1cQQZ16wn458T0mYzOhyNZ6fpr14jn9
mg0pKC61+5YR6g+xvBKqO8Q4+x83YT9jxuxLZf7sLV9h3E47WUG5bIZgNQ4GdCtx4J97WbEmQQ/M
k5obbv600goKz2INA8aI1Kx/+qb3v8cp1q4q2KGy1ntmdyxdA9CQ5RVVGboMm3Zi1h3k6UBtk3Ud
w+OYk2rNwaSEZeTtD83keMYIxMoNCrO4Q4Ofq2ZglGPh7z9WlQs7un9jOhSm8Xcw9pWoc7+IZAhx
XiW9H6dpEJE9vrnUdQVRelRBLjf/lregzZ41bT4Ai7aOG4xrqrtwAI8O6jmIFr3zr8/ZE4vjEbFG
etkTcAyuGiP7DiVo/zt/CHunnqhiK+j4TPaIGf1Aye/1zBApqn21QKdrv2QSJtlOVA4fl4rz06Vj
S/8GgxVMYpQSHsEdmOdP/z/TLWFwcgxUp7kS1OMfwcmmz4XL6RFniBaujx7SfPQIMtzOAa8RToPG
aiMDe7llgdWY59JeabPmmfSRt7HByUN+6ibdcDuViiGRNTrtsw3znaNvAcv7hIFsdooW8R90d00g
R8dL3gYPkoJ6d+PRuqOAOlZGnKLg3O9YLCXZzGbtgaQJtobS9FnKpfHGoBuznhTgz/7rSY8UUO7p
bPJ9XykKQdv5yUtDSNxKvdHaLTecHew/btERThWm85IGhcGA2IITx5mpow5+QXTmZ/Ab8rgnsC2j
acHHBtAshhUVdXxqN6ac5GXrJiu6/WHFHbhat7+6UUxYFPK9IT8L1055Y0UR69XqyzNe+HRZLnof
IP9RVMY3QkwrRQXG9pCa38yKSqyxKBsW98omracYc1Z9eER6UThvn/cH9feWaMwryhDxxIT3aIbd
3CqYPAY/Xx1uDY+gxMzJ38WAU6itFnV584fCe7qg0sMAfaHKPh2CMtbYyWuo3KjXI2aFvECYE2hl
5oXW/832O8BWbySCFNhmHW92mdNnTelqmxh34Rq0ZfTAHNvd0hvjrL8nm06CK+w7MDVR2x9ExK5m
sSxoHep7sypYFv9hp3DIPgdyQe9YzOK6+3fjYaOp8SHqw3xPgohh4mRRU1PPiM2s2XayquYu92w2
8mTm2X3M//rJl4alDUSZzALpYwAp9XNS9K3JKf24cQhfGeAHS1fDg1wOvTrq1m48MgfrEBPwmvZ/
M6RuMi1i1vOoFd1wuGtJVfNoMWpQAWz0unmwp278UYKYQ1MNa2NoLBllyXmFZO5uxBIqpqExAS7R
Xon8ewVjYZbn3e/2e75kAsT9y22/v2vfb3XJg69NPFE4UBMqHtNXvrs51ysRvmtqgqZPOgSUIo4+
H5o4BXczMOYhIUwRWne1ZkGi4sHduiyoqFbno3fHhx4iPIXML0Ly48z36NdpBCFNFMK9+kzmpl7M
wlg5/rZzioFRaRZ7lIZZTaJY/VqKtsGNjwYx05fdDPi9a2mJuseqL6WFPc8ZjNX/dkw8TWM/Sefg
nvPq5ylNN3IUZ2B2zfb0i007Co/1ZvDZUcMlT+Z4u+yOQF2bhDbkJURV27dJfDws8oNZnmMf+MCj
GY804UtLc1Lp9h363XQ3X/Zrz4OaOyJ18IQkRytdsk8Lvq2Fwddm9uuGHIkBRnYykbUy8XviDZ+J
Y3s2QQ9s71x/ki+37PuX5su2++4GIGPfM3QlylT9XNmDBjHkUtLuL1uboLTKeCPGOKHiB08yRIS+
VucVAxVkJLSB01v4BuRAxFMYYKfd0gUZFjL2j44kQWwQrN+wOJqqIxzyy3z6IbwAxpUUG+XexzM1
8I9Uj6nk/WiysWMppS0IlBJ0S3zjmc9XvAMqanmbt9k+3elaixQmCQcxpIn7ojQzF560tNfFPxYS
K69a+rG7tz1jB9OXF0qMtKJEhhajeoIGgp6Ml8fKbWqB3CflWNEtMpWYi9UdojyIZDJBkiiPmQ7f
WnyNLS7D0GNK5UU/wVNLz+uwKUPo/Ky0I/ICnq/Lrjk8HhXQgTuNE7bFeSLHhggEuE3YO8Xx3oHG
LyFhAkab5F5ST78h8v66nGyhwMCuljRPgJ37sXSx4KeVie09bsI2xSr2tec0y1K7Ffy5rzeP0Y7p
UZ9oenYtPyy/21G25a9MXygu5Ix9ehFZHJb7/e9b7w5OTEHS7DiBWDoJzHPvugSgUCllpp6tCG2y
aISFdONuC49/4XUv7z1tVFz3KMX6zl/l6+na1zdWEmCibBvh4v0Ix1Ktmp/rmnzw+11G/41SR0wY
AJDraDIayBIicP7C/Tx960Byt2gwNjmrdVMg5XmonW6YCs+NWYSVYBL8ChapE4O1dIZCnfssKYPi
caJPrHig7k7T8uNiM5GWKrju4wQqvVerOx2HljMF1axSrFw3NC3uia6PzsPSUAQxme38JShXPoMz
yBo9JazGhn5plTixgaNolHLxfNoXUQrVZNFrO96YAJ6oZXUNn8hpMTbZiJirwacveCObM3TRsjsD
cDck8Eba2oQMX0/8qAXw2o2iXZNLCvcCznvNZQqAWplIKzAmenG0WvDKK7tIqaUGvhS6sEkEBYR6
crKkwS8FPHgzFEGZQfnFGlF2M3w+QMHD4O5udkXLoKO6kC+V/0Vpei/oikea4EFbNROLikLdiMgl
KDzUEHceKd8b7tjNe8MG6CiJPY1D/iND09udA+NAa3EDwQ6bFkgOsjqpjH0KXlwwEL9v7tZtHPnq
BJtr2DAtAJ2bYOskUaXch2qn05UHed8R40iV690XcdFJ6WKJ/oEdpinyUKjfyHQz4BYdA+ZJPH06
D7ITxblXRV7QH/Nc8VF+I/+4LRrmxyfDRPL8VBl1VN7ZlOVG40LM7zgrRrHGgxR4HYUhHqIYq30N
4BdBfyaTrMHItziIXWTK989CJbA8aqwlI2giXMUGatiDWleb43TNEqqAqrTHCqosbfWr/wBwwQ7d
b0tIKEilkCukdYlJZ7r/qpNhYPfXqYLLpONJL5jL7+XYfWBZQtXPY2/ALMRjad41jHbZOs+3KeUi
I3whbQRSUnwQ1/dyx38L+3Ns2vDaotQQaC6YWqCjFC4sqTZuG74J9OxJMAxFuRx80dLvluuaMflc
xljBolG97buYKaGeYjfdzuKwXTOqof9ol5a0u/xagC6XDeFD3+1vVX1NHjNKXjGN6rVnP0AO/wd+
jcM2ipVAPU95WT8lhSV+aljliGOk8qCeDjhSkPrWcfmStn2dQyv8SHlu+BNnXHMC2TN+hMMwYB2k
XCVxTqE7JuEcW4PYEJwgjjxvmCtrr8sOhqE5PBA1S3tW8AXwdGVUK6VEg4CScHsNgOK+Cp05N1l2
9QS3av5j+6Gv4mZrrGa/xRFjypx9bmEGcJ9on8NO8XWd4cI8nCU6ao1xMGpLwX6669w81b4Ja0QD
6MBE9+WRsBzk0g4iXP8y7y//rWMXInQWRc53+QySJ1dUBzwUIDE+BAij2SITz4KNH8nTt9JwVrBf
BwBa25P1DhVKMjBs99yoSNTAM2/uTVLsGHeyA23WaGJCAH6aA+muG+KBjn+K+iKGC2GzPJskKfEw
aRBKqUE1/NUOmlEgSH3oIrRB29M0+aWDqUQtcuGxNvEUg9H57xSqREXNZY3cx6IomtNvIDiKgnOJ
mNrZEzxKBs3jpM8eipZJsp4qBQ03r7pT3yssroxG9NuYV1Hj/EoaaDDnWVtQ9lMWchKoafDfjEN0
n/sd6fxDbubZ6cpAkW5W04YEaLZsM+GeAPQZjhVs7qebNSvdAmj2imYiiIr0lvp8U9UDJqnNDHbt
q03thWoumwf4kiMiCuGOKLVXgLyKhqmFKFzNhxymK6MX7C9Ly4ZkLcMU25Guu3xIybJINlvDz6XH
yqh1UXYel2spBiJ8oEZc4v3d+V3fqrziUpvvmJXtS4jY2D0yH6nTZDpaV5OJiXlvix8kl1EnoVB1
tDBCj3P/DyK2tWOg7sDLn2+k59ctcwGgRRqHfmDO1Dv+ep+ohfjoNMLA5pB3h7q/hvbhhBqE3ny1
8q4xIu2psSvE8j4upLSxFO/oQik5A/MBCvd7meQad7KmwaSW2r7vQi5M5KVxAwiMcXJVYn5DWWs3
9VaaOE77AMprIihUuN5IDltJNmA5nLwYFndZz/3KFr8Q1USgnELkBJdoNwkQ+zWADcDXr6eZ0GC2
LgYk0AmMR7ku1hs5KI1F14v71xeij8yJIHMY87lbf9tQod10NeY8AcJUiYDzyhfnN1T8Nf7bX1rQ
OgDo6WnSZ8dX8eopa+F/hB6pJ0s4DCTGig5Cb+KARUPCIH8Lg2JD5fULhMvYRwvYR4dxZrNiHHir
qZJz3Hiswq5kl5hA/QDdHWeGHuqyna/U28s0cIUdxQoLgPUa6v9YMsCzC+pZJm/YTmCbvsY+ynOj
I0TcAPqJFKjtfBn3djUBuwyWt3UgFix39gTLQtWmV3mBm5QN7Q3wZHqMGbhqOVrKa3ikWA+6hILv
d1JKoTkeJeskg8TnEaCGoBgNAX/uXNm5GvKITmttUaLXI8L+maIrii2Ei1Om1pvzy+8/vQV3ix5K
5XJWsh3ynOROXHjXpacJ6ECyV7o07/a7JwWzs53/ToMyRuD1z+xplLIRR5txXPUuBtPw1jnDXpJx
SvcdPvaj94+KdNIKtXZr36txNZYGGB2KsVtf5eWEq97rRT0TtvyRGLpNfGz55XfRnzCa1ueCLvge
7kO2JArzDKtHyUrY66uQurXxU2lhnfRbfIYj7BhfNON3Bldm6DLTqHWiN0zEvEsZhDNz6/zu/cHC
aNkl+iv5w6o9GsJvXWNbBRLSpZLlo5Dy9XgLyxsXQ3bQGd9OoAdbOm30BEYgeeTAnRjWzMu+O/qd
bEitoFiPcSXliRImqivRyxFSqmVwP5RhnBhO201QoEK6N/J8cLWRLAICFFBtJu000iNJ0EUXjGtI
lz3cvqjvE7Jr4Mq/5F+co5pbTwQSDZwa1dGDcaWt71FIGXpwtgY02KRP019VesRvF/6QV6jMtr1w
rll3ht7SSvgnJsIEGNtkk6hIJUFgzTBz1SneazOodWEfkHSiESLJ5V/ov4U9k2RmrjkPiexDG6mz
JY80xY71Xbqslfm8Dx5H6be/0CIO0Jdl9h4HcpLNqodMFW6HpJAFoNPHDlZE+C94fuYenpTZUWQV
vrUGm0sllpn4XpNhb8AJgpFX+TnmVZyMKahGb/v1QKh5LqQeISrrPlnWYd9rsAM2S8NgbJ2Ko/Zb
ciZNR2CiUtGz47ysi5DYt0nDrh2czSVNSma6sLsAggNUsXByIxnpAt9UUTItjnLoyFl/VUxEY4UN
sFmqfmxWch/epGH6OlruhW+CaqRrBPE9DjjIzVWZmyJWHf5+AFUPI09DwH/DC/f6nkxaKNN+BxyU
2NAdZxH949YIGiR7h3b8y5fVf9qth7BUSyHu4WsHJiDMjjJhYO+Sf2Zwl/94JZlFChL3zt1w/ErJ
RvKd7OmewUdOtYw8+MavDWGmbfixROasrtQl8B3Ae7pz90ScyWFiFJorqBoZB3pycoiGh96C+qCN
QsE0E/azLYBZafEWxLI3fXAkQeWFEe8NnJqIwBxIYSnCez5k1lzGo9KgcMVBJxp8uPV8I7TUOkkq
ajd7NFcb8DUeWekMy41Pc9ZgDiwe/F9LP+W1d/iHUT4wDn/eBXmVE7U9i31dbylBeZwDdALJ0Y75
o9duiexYNjMvW8BbGk1RXAykeWziDKUU7icslPJXpREVmn//YRjiGPLKsYVNs0Qs10hc5+NnBdAH
/sgKcf4JdpxMZmwSLMQNWA2ppmhTYbj6bm87ypzD5qFbbcFMp7WdHG5Ej9BsqJd1Z8QMsaCLL0xk
0+g4bDBc58vUP3Y+JcZjxMTtRnlcwYHfDAwXGmUeQwKjArWtpG81EYC7fM/hXBvt+AIL5YWDC4PK
7NWvfc/Pm8of5fZ2tMK/2dKOeASTywgE4YLu/6HkPkiylW2mU4lce24n0JF2hpdhTV+jQWNUW9a+
dkKxvUJ8+e1cTI1rAqbDFr7tctpyq0XvfKbhbSZmQb15iT173elTzC5984NUxL8REHLHDC3G5TwC
A734TLGLQ+6vwOIa/TQqJo9MKG9E7K1oP77s9y/pECiefmJj6t7Qlrpys3N9P2SiBnq4mh6gP8Z1
Arq6bIH/3tNUmx5f7xrE6rC1c6dmCJD6HflhdSrm8xaXizFK2JlI91Y1wtiWlC3dyYqyVeaPpar1
lJ1yRUSORAssBP4bPyfmve89WUpM5Gipw1tHot2gvVXPWII0K6eCHqLnirP1IfAC/W+mUsGEeYVn
qUefHyA6sIEobXxDDZ6ITjlC8pfunicKDceX0kvzXsxU3/x73bn+7/tUFeEYEcg5VyBCBUl2pSSo
3tlMwDFwijx0pk11DA7FyBnSLUDeRiJU82ZKWLE5uMO2iFeuik8YIcN5sv7I1DZpt9IYyJrohmMK
6aEC+iowo29nT97WgL9JXIwesDEnil3cRayMoIdjYFbyEbhPvLnTQG+HQILxGXpqtAhnaNLzSuuP
xczylzclVlNhxH0OzpydBssmnfKu/D2vgH0/AYPRoVtjyY8x7S+ERo+oyRMYUZXUJiRuzy28VeDX
I5tORi0Dab9GCaw4Lp7697yXkONs+70lQF0s3KmV/7qeXh4PkL4UWp3FiTqd7UPRfMT3ZruZsKb1
cN8Axrijontlvxmy1qyJGNi5+/f8bkP5gfpWCfxvfAqEdMIIFY6hu3wEs5VII5Ch+B/bDL6Ct8BN
aUwB1vwLGlLwmk1Ft1DMXS+CitIa6rNSpFLc885jDzrT+zSggO7hg2l4DtgTUEkJlryjvQER28zQ
kdo/lvHiiOSYznHH61QWxuYTczCO5HcG5I98oJGRGkzEdUPWl0b/rIPxdVaMoEAobw+FtRl7TIwE
E/BrkvDcrU/jyeNPvh8VoJtIUKRn2jDSRIWkU36WWtoofoUFSe9n6T0xk+wZVBQFqH2NIux2gWUr
6mfjnevy0CGuflRCdtAAXaeHqnX0Vika1wQF3JijMavOw1yEESOi7XpjkDGR9PcE+S6VW9cIcxvx
Fo6okUjiWXwyrO7qIqPGfrrx7mZG7V1nBmDeI17rXin+5wLfmx8P5fPLZNpYXuNFCsMLLXh+KfRg
RUAf7ePa2XVHMozTB/Utg7i9GVh9tJckJqy9fWCr//KmrECg3q5CwqamDbVM049cH4LsGMW3/rZK
rsiajrVf3c9zeUNR49rmCRkYdF4AqKFEX9RQVoir+ko1n5xmnKkaofnn1fR8xj8vPYAPmImJQeGR
53ODF9Myv6GPMr/PaB12LN9CPTxRDZRzDa3kRu02uZYf9klhv2XIs7KgI+gLU52TonGFevbwFIhB
R64Okfe477UtzThsWkyKzj5qCcztzofp+PGnakHnoDr75G2OpBajV+XlROo2QoQXfMGMnvKSN7Qy
UlfZ15goiHxqvnV28ElEQTE/gjEr4FAkjqXjtYKxfJDEo0Vr6Y0t1krlrZ4yu/NfhwbYlh8tTDPY
qxx1+DVdnP3vcRLq8F4dkStu4GwnNFG4MRzdkvwpXBRXwAX6DnF/xFi97p284GV0gYnxs+z4Vhz+
BS1hbcf2epr0ah6So7lxL0/ysvlzE3Mymru2VS0BJaXPi6jPo6BqUY18sMERBUhEC8tBM/aed+vr
1N2XyeVjvg7ax6bPLJ0pOUvoer6jPAfkEw5ptRUOJIwsDUQ6t3N5z5Y8+sQCin/1EQDwhk7xv8jH
lr0SYW7UIQXXOtqkjGAzUxppgWPEZZpSheBEXMEBSnb2zTp7GpXIrbnB4ECc3Mt6isDrh42i4ZBW
4E0UcYY0nwHbNfwWQBzJSzK90ser3a+fd3JmS3+vCyLGDx0vwRLECr3Q1Eu+DSL0oUgVSkl04LAR
RTI7+3MLMOjWIKHj2iHSchWw5tdyTwYPzPyHZBBuK4bMoPTn9ZY7kdAbO7bi3ZRutQwrgRp/ocIc
I8vFJTe9Ez9WlYCXTRJT9jTDAKNDWcTvJT+lIhzlBYXbUulj11atPB/IotxNUV4pGnPLGaABkmvm
cL3HEHo+sf6vUzSPH8eVIceiPF1lD8YHDXJC2QWLeETWupTHI5cTUsorxTK3G/+SDy++2KIgH0jh
ChjHktOENqnU7dKiT/AR0whTofJDpZN3daTwaNd9uHwWEnNUjBXgwpRxEWB8py5xr7Elz1dhoFws
vBDhsncYx6W4ifcNmBrxBBwEnYQoT1plltOnXmdRRXALtoUD56n/ltZmPBSF99j7mwu7ciiZlHFk
xeFOXanHHyYir+twCSNq2/1InK+9MeULJpQ0zZCSsyIHQQC0w88Ja80QeKtBHnFZMJ7YiZXDmXKB
hbRS8EtRBlRT3Asr6Ql0YrLUnGcLiO8QoeYXRFYnJm2XVLfegufDfukIH+2NZwDPOx3Ogrtod4su
CcYvFAEmEbzssqwPaOVFOea7gnfoxyakGeeF0/SNSbELLV0mcB9bL2dOme2xBG4ALBfVdwC+BxKe
Z+VwghUPJnx1nHcjJyhwOiR0OR5Ti1gGgOo3zyDY838iipT3wIqYghsOVusqmBz7a4aw8yuALJOt
5Km9/Dr9A1Y9iDZ5JmdVStAJUYVTvs0zynKZs387q4cRWjG7HXmLCCNOo/UjnLDLKDaaGthU/mkW
2sIiykowy06yP3PYodd+YQFC0jZdJBjFLJNjIk0v5/npnijY4z+9Cyu7aQHXRDCSoPbhfZxEJEDl
jxYK+4cRTzYnPA89oQ0GqXRBU5Z487FIF0Dz7uEnC7Y9kQfRI3UK8skUUyS46TSsx+374rJ/H8A8
FbqIq7PYg9XN77pSgSnbGIFC7JSdL3tHevfbablhAqus3mOCqotIstV54qYsj4EtPpjGqoFRj42z
VQ9DxvzlDN4NSPW5991pE3mjO4AE8hdt5UphEEeE0L6QIBJZ6V2U9Vxp2xfa15AgTODtDKPCc9Ys
qATS+munwCRmlQodXLotnc1EJ1eYn2jbGca3f/lH/y4o0enZPsSoCwDsPIqmodVX20vf4vP7XKuJ
foQtvHCMBogwXliva24POB4xvIeL5GtGxLUdapkDNaHsYtZ0UVGnc9DJKFcuJgI0NpdZNr1w4Alg
dSQde+ZuwHmyr+nxanR8LqnOEsXW33cRV138qBRuaKtktYxjVRgZyzhyVFg1VP/M/c4VifxGj9PB
oy66fYKXomJ0kocl5pqV1GCjo/k26ws+8EInIurUyBdlPvf0bYTTsUNK221GcdDjrqRx20+/A56h
Xw92N1hyv6VHmX8Ml+HZnA/ij3624IgJHsP3NHMOMzuphJFohfk6ald67pYV4RLB8ECwgYTskN8/
7aCiC+2gVCegK1JiY12iihgP58RVPKPH8uliweYaRHprrUPH8RnhzxC1qomdZcwr1EGXmojPEzAC
gy4veRdNxQesC186/xMpqn1WF/68FMEGXx2FwWlEqpMJfoVw/Bq9B51DHy6Lu0DFmJP9uUvXwSMb
0K4k0iHzcLwa5DjcDAou6/eIPqyshS3XdSXNHdR1gLVsEqsKnxepddCdCRgSR9KWPAOrCp/T8tVG
fKB0Rc0tXHfdduPlfmBvJ/KM9KWr/tHoXxiGA7/+7UIy66ktEeE7Pfa4BtDI5hg3g32PMnJ7dzqJ
IdjZfnf3UxxubhE5uIL9aFGVPLPRr7U4p8XFouoW6EpwlvQUgORbIMbHyzdC83H5STE05HhlNM7m
CPaOitJt86k+VmOIQlGkjJ1ZLY/bR3gqj7ZtZJjsHPP1v08jYx7darenuIop+88HPmVVsrYccLww
2xWTe74glSh0v1Wyc+tn8HmID3sokMkul7zjHN4JyrIt8nmEU3QBCjkklk26W1foSkOQrkjrXROd
J+zwo29GMv3G8JSgbaR1Ihfahze09f9Ne0mZQsx8ZVz6kxKRUSAPcU85XSbHCYxnJk69NKGo5aZR
5vhbIffg8mX9B4GOMsbscpq+Ttm/p7LHfUMHRewsgdVm9Q0SXTWqO/TBcd68cRexIl8xhl3S6Ikk
0qHJeXp2ycPxfjIKfy3VQ+e8vi+pK1UzpHMXqDGf5kslE7rihhFyrYeXtsax6aB91sfH2jMNNsI3
DQiyxiY52fGarVF/UxdiQ3X0WzO5K0hzvFp6zi84VUjHmSCeg83ieISnUhSaps+213uL9GVxlyzS
Z8UrxHoV4wExxqFWxH48QUB8auSVKnayldEFDUmyotU3QsFv2SOic4uv1TCYrOM7w+1j229za/8n
HwaDh7NZzqn2/2JSg7btuX9pErHCwbwKQALIcAapJWqxe3xKhssGOd8KkTsvmavTgJ5dve0aT2Uq
0womMQHkaRiJscfCGjOItPCB2qzHXSDKDtEJbryl4OHQvkrNRO1NI/qC94w2OdiSGUJclZ2km8zt
08ZPM0vV0dsb/Ta83zJva6oGsFKOi3lgs6djiNdFOTT6G65/C/RWhHYAYxU9J95w5QMrbjDZkQZz
3syC/nM/G8Cv7UrAzkccX+WsQ//+YYjMBw+0ShxEiZVK+st5dJbIv9EV5oAZAzK1sy8EEaSF/8o0
aku76YfBZnbDHMBZnqi7KCiZsFoQPB/6/qhtaRu2Gc8cNz2ELnWCkJUR+lgHXaqR6JQV2QkxVARi
jwCmmv5yMlj2Zf3E0liaVb90yxsAX9VjPpQQOrXpGZeKZrb1kCwlmcIDAbkrNCEt7kCjhYi9cbNd
Ib+ud9dp4NN5FdB3/bOTcsjgkKGb+G+OsQiyod1P8i+BYvlXcrAhNB567l0s5mTE1tOEcDvVXa+S
qBrBScRE6of3smE1kdms24QSAAnB1kQPDms/JjF/9zn5zBDNhP0fRiNGCpfWRv1YJolEtxZEtZVL
u1lYy8IRN4ZHGGrLITG9lLt9QLsRXhKjsLzv7d8MUIYXARM82PolIrSKkMAk8SWUJv0oR5CNZtdl
bSt5cz4whHy9cvHtCGHDv4/Mjm0IaAUWZVu5ky5RzlodyMPSFDVjqMkM9RucAKReC4+3KII1P5QC
5KNqMeNcfho0ynbCtMkOUS4GhgcPgkh3IdiQzP9Mddi1xse7m3nlxQscAh2Ef9pHOTWySBJzQRTz
gOhK6CEAiLKAW+Axvvxg2yB1/AeU7ticduLnosUK3m5JmnfONZ6XlJDUTEYfAlKVEyGF5OJXMrwh
Nzv1wARDsOQ2kngipdGk00mEUsMwe7kPyZ6iXvv16H6cdD40E4XV80HD3/TGOShSc5TWwx5AI7dw
28eycw/UL/jxT/hClkqPTw93YAUNRtCA9uVnzSvJaSuYrJG5pHYVHN6dn5mOlawHnd6ga0ia4MKg
IeglbScQknhVoVMEIDCBzAXnmiWAhEod0bsuq+fYmbrfEqfJwBesSmn+WDZpBQ8PsiuIC4E51yJj
fYp2ddyorVyCVl4vAZphH/gFN0cV+LyCyG5vzogm3G4uHIBf1Yx0Swooo5Wvo7xtY7KxFCw5+9Ws
XW2s2RJ4wDiHJR3TK6FTCPUj1WAJKMiNq2lWgFypLZJdZdz1bu+4ykklAg/mn9N6ooj5+FaJp35r
P8FYEJuECa+FPbtQoxVKkwzk6G05M6aIZhowfKtYtsNCblrauEbWzVdEV+oKMA1NM5Sl8zQGfZwI
Be+DA1ysQkmz30pRnNpNKeGXR5FWeOvmpQ+u0hf5eGc0vCJOxB60lI9HPcCwAeZ1VdMGSkAaSEnW
QrHa8QZ6bjjFfpAACDTkT0zfM/kA0ObgrcYvxxBn9Yd48ZrMa2QuqqL69FLWJGs9noibFkCD6BAp
C+WbBp2SbOsXMqvqaCQdANxkEG0Lu0j8BQJQSpbzg3jnQVdHdpk2mOWVUygaYcgS6hVYaBsINoTP
Lsq+y9bJullgMU8A9zXX3AFAU3oku38Gbf0gvEGEbiQ+DzjRqj+iUj4UuNaB334OBJgxHTxfUuN0
8vZQznlVMjpP72IrxmIraOmCxUZ4H7RenpMofUi5S1Uiw+fXmUZOjgt2tRd5t4jIt+1oZ6jWxFsJ
0pkRW6H5xd8MTSfdI5vnJaGA86nKRFyf9Vp6yfsvuzzYOVPu/2FUJBSqK0fl5QP0Z9LlytGSySk4
CHNZNtdj+xjgv1TU16KyIVr5WJktPhs9Sf8SwaM4V8/13sDBHaPCykR2YJ9W6Yqs4ciCN2A6ihgU
kED1pOATCQy50T085URgjhJpaYhkeYrf9EMX7CEXabcWQtessDwlxgIE058DjHrTSVfKlT96XHDf
8B/eBz+wyirl5Tg49l5MryO40Kl3WllFP3CyprmYyVXzZowzotgC4Xj+l/++5wUOovYPWmr0Dfbc
OsJ73H99UAsmuZykKC09Xpu5SqjoKmwSu7wuhbqlFqu50ds8wqtjZ7VEaVqLP8TuvDnw+xw5D1bt
1Eb531q1g1rbsUDld9gNmSrp2lT4M8pqE/Z7I4s2qk8h4As2LHkiUs+bDuVZBcvtt7tIMk398DBP
FC0HcyrGqVmuYXv54rI/DtkX5xkqh3/XVqjMpQzNKolhV3dAnfHl8yWHyKEibhzbi5ekOhI933m6
E/FanqmUOYbkwVhmf0uERxMwD4G5pb0AeA8w4rzhqDG9m+ahErKPgttJoUtkLqc+GT48I42KG0SX
LyB3v8uSlChQ6g21A68cUFx6cBgFwnjeJMEzib7wGw8N8o+Z+qiq6pZwwSUl8vEqvVkqhj4Bxnw0
NheezGcRsy7yN6X4Vb9ks9FbmmIab0tOnAHUNmL+9UZ3EYAgWndXMQ79sc7XE3gpO363HUhuKqt7
AH5bI1F58QFPuQNSN7aq+FF9lre/wesuDkWmnXbrbCKKjGXXVW2DVrpK6PPZ3lVxdw8zUmeKJz7y
Oi4yKZVn0JQhIijghDrhvU5NOrlMCFcVt0NbQZx4RLf+pgp6LwrQSJ2MXqgT64RtqzmZby9t0+/z
aDqJk4/3vxX4LbQHsNwPPYGdk4yY1pLbfcxeyBsvez3PBgqbuaNmARncvmdlqlmHuAhMI2Loj1rV
PfjzMlZkKdc60nZ3AjS1k/TsibJCSm3AsMhywgwzr503EUO3kRorveNgWtR1YWZKSKiLhCSwhkbp
fc/+TvYJqhlmEjomYp1lkxveyQPHY86DcfEaIkZbbfR2z6OmY6MrMXpMcg0vBjw5iNzzLD9m4pmW
DRkfnr4RuF4DGEXbN3/r5DjDjkoRsaNr+mHPWGLRm8xUxTIk5uf3wEiVIIRTxh7Ly9Og8rvE0ahl
6fzXMxZCGtHaNCuIQREUYTEba8jZV/moM/E07qdnDAu/sge2DDGC/ecS/VRop/0lOBxAYUCGR90S
1vhHH2B8e2j32l/G+8BNTKlabHWAyciL/3wcFQMc5FlAT1GGYdoC7yLpvQB/xy2LWM9Dc2RGC5Ae
rzuCEd72UBSlTs+kmbp6t3J3Xpa7zsxDBqFrERHusYG4xgOIibN49wLR6eYfDd7LbjIv+XTzfdyb
7xfzcLCOwjKXueGv9SeG4+7LIq8hqALW/omdgGXq2/fMcz8/zgsGwYRFdhirpTiHDaHQhVs0NAFE
hsgBtttmOw5I46pjvrQwwvZlVuQCHXHIVmqO8FnRUPK3w0VhtmUFCjINZ9yCIztgpeXPWeh9KczN
hVdipq0qaRNg/7YVY2hxh63dHpiyjLIXG8On4gTepIvdxubtnHBvSxKj2ee/T4Ry4dykrtpm3KN5
YpN73sGhL8LZ+VvRZyYKMSmml6DRX9prPuyBJU6B6RBeXCJa29BJgKh5J1iKSk7L2txZ53BzH9cC
C9iSimNQY0Sx4xyLck0w6UlVZcCMcJ5FbZqqLfqOh6H8mWxnn7lN5rRs6XQFSkdq+qMMusrO4LMB
LusTKxVvW/Z4/M3rJTIczJjZiUyciV/ZzcA6+jPFoWXxRkIbK6ct8V0CM5RtPLUjUMo5egZg1pNI
wy2nCkduCV5g0Ys8vHgYEcBSal+1uMO/v4uUHNKkpREEr7WkG2pWBf+To8bv2J582p7L1l15nTyT
Az0QjjWO631TaLzIq7Fj5ymldCaYvt0tZjgo5F94jcZX9KrFsHPM9/wRYy66meNicT9Wi8ShMnfa
X6xwvHifTdjpNQd6Vpn4OnCiA2G1GsJUbgzkyCdz/PR8XP7+8M+7Z30ncL77H2l7FICOQzWc/ui+
fDLq9TAtmg+j2A03Nsbg4dZwzjdV6Nr78+mSn+j99dN9Z0tvWmicKxAGR6R9g9PEMd81/9wLN3Il
ULGSljKB9U+e3K9BU+mSS0qLmQRZpxh0z7fWBqykrHGPna2cia/uYlMiNZvSh7wx17M65crT5TVw
6JQMjplw1lYhiRgWQxJje9NcobJMgCnV05AN0LJRGhvHmGHbI+KeJCzQJXV6DN4IP24pmsfNX8fE
OBAd3SvTPmdgdBXI6WKrdUEoOWmc4u0/Hs2bIvZYVDczHc33zmFdZyZ8ONoskBWSPC7ywjS6zaDh
4InLUZMXnQ6syZNJeqrG5+mkL+4JrDMoX+OUgAHhQ7/gcTsiFwdtGK0T52CusEazpHUGL1FXhkpO
pwv6dkwqYGSPqFynQ8p0kKQy0rUPUQpWKhAjWZnGtSnsQvDR1rXI6wKPNI5+jYmLvoL0YAYetGFi
/MxJL6qe8n9mKqjsobviYLcl36KWxz/NiFS8KkOB4D9hcEzKmEyFK9aC02+E2tKcYfFnsNGR5swS
B8MErpZSwwQ8fFPPxIzEhDRHFRHpSaRgt1AWRMrQIj5AEVvsuvVk+V+rqaDn8A7UQyjSPLSHG11p
ydR0sBzDSnDzpZ518D2+b9ogzAyFfSB9ucu5ByOlIRjQ34gnl9DDOwHPyeNijbCsfSm1TqNsenEd
Um2+Mq5l17Fqsl5w4vBFZx2LD/fZkxhAyn8aQFsCk8R6lPjnaX3smnp+vzo0vR05XrHr8jJmpMMI
sUc/GZ6XVgek7QKipiJdh7RY5ygfItJZ7TAJ4Ibj3gefGIIjehxf73nmZqh2IqvrC8k1MLrwMnSY
ikRPNYZFmU+WwRGo3A8fBE/5+67TXvfMb84+2UmsH+x/3a1BotLexXqS1bJYgJh/Lh9FK9iGaVjO
ej8InKOEmohTs5Vb1A2qC2uXYIWjDGn1aNX/AGm0ZfA0daARLA0LXMwe1zhJHhbfRlW4B2J0Ecb4
nZSJYgbVO3vzCvuaIZch7UnUchng/tvapwMIGlp0y241y4rfsJdvVpICV/qQKh1h+aWMSzW/ZmUd
QBH4TiDwTPP/icvqiVgqwW2/6GiynjbSmuVsstTPb5yRciB5fHQv1jDJT6Y3mmWfdougCSqOk5yg
KmU2NkHKrg6OD9iSYH1zx/y8NlC+goLPeoht5fOySEBhzLQOLLB3o/0v7urJ5g6sQs8J/agsoLfq
RKTcuPXTkllhuVgaBEj8n4fesiu8Sy37ULnnDJ6+u/CLzI6BrVLBdkVYyk9L85LqdNqscUO4AVcr
bgiAHfOW+M6n5VLWh2silHT9PiZ7GqQEk2M6tJjZh1ZhCGJzjYap3gnci7/9kuNWp6I6BwiyvrQM
zLO3YjUYZSOEPCiumx+GZkBWsov50QJl10gX+cJSvQDNYXPIOd1lUrwvTvIljAmwI9mUT0a+/WjT
KW96VU9ojaAfC/uzHpVt1eSigfLkvwuRno8LjmglSVOzX7Flrno1RkYSMwZVGm6HMjsxxMqRBeV8
fkrT5V0MfrG9M0wD50dJoL3yaQvN4obi/rAG0rxVUYYSuNCFCZZqvrq3GQG/bUhQ0B4MLWAA7nr9
vZkCoEn91d7S4SxoWDqPf0UXZKhULQF++90iN6UXFn/F6Awuf+YFTm+qFrzEFK5cLHdKP6rCCSjg
QTXbmydU1u+4X2y3ElqmskpI0cG+XZhbhdD74OHB/C5n/JFGq6fxGnnbubls8tX/9X3m608hM8Ow
vodNb1OfpXOC4gPdxRpIf23oqdqyKeScpnR237OfF9SXRb/FiSjFcd4+vJZ02yo1XLKQbLuiOhdx
rDNSpedY2Y0LzDng0WkXrISRpqvezNMfwfxlAKsDwgHSmVU4j3Jn1a+Vom42l1xaRbxYkRFbDOkY
bgqVpzzaAm8eQAifS2ASuvnYkztQfDZ8Q2xc2jYNjJJOjdv3gvM+9/xhPg6bruRtTYBIOLY7yEXa
SBvaoRTNPgMiYgndv2DBLcl/pJSPmxlFGdPvyUktkB/CYfPwXb4fZOorf1Ly/gxiBOlNEtjau47C
joT8ozcBV6rxcG6VhDgvy2xbxiaCarMl+Ou1nKPda8xC/iZzuafIFTWBPYfI0DZYQVT6nAEn/KvY
KROAD4WpJbe6HcIHyJ9iM45e3h8RhK8QRq1ub586kcZYjEhdHHZn2bKuly+LwPAVeqHzB0VlwIRH
2ReDcMpbFYf6cLFIzE/g45R3JIsFUdZ6QHx58w2h2Y/owtEEL1qh9U6Z1DlA299I8qIw2LBqsUPc
UjseWRCICoLkse3xJdhqUkQ4ns/EGMRKfVa9qlmooIzIqMQCB347/FhW50nrtZPs47hzKlSsF9Rd
/kdcB5O8McIMWSE2fGXVv1szauDIzzwt0KcNEBIOCyyehmIvJBrJiFbRCPCoo525LnDjUHMpTnXT
vIPfviui04A8OC1KdQ+OWXkNtndn+TTTdwolHcSYVjx21kIKPOfqC8D/7cpGeQeDg0rEg7pXpW7g
uPbCWdX5po0Mj8w9crI168NYoYZ3bZU5OvLKQlBgkcyg/crLqzHHqpLgsqOpI6ZkkLb67vnUWpmf
eUobLdFF4Gq6C3Gz032bQbrArZHAIw7304X3q5fGKZgh7010nH8bJ45IryqqrqEjzqatmo7bBw1n
Ivw0jS244lRfNMyh2DSSZyvhwHU//dpBC7efJF9H5zByi/gESwuxSZonmzSP5DTH/d8c1CATFiV4
BnBd2zc/aFh/Ua48uZfaPXLAkLXuGQOut1zcf8OyMrKhsLUsfzh3PXNjMo7y0hbrV48KD7LT4A7g
mXJKzODXiRfBfaJeMtTDOnd8MU0ODwavVye0pa89Pq/X0XKFLsXg26HF166JdyOqnn8+ntOy14qG
7tZE5UlShgmdXPp8+QkTRH4SEREJGou7ME9dFPi6Hf05QpkH+cat2EiyxZRyApOSJtoesH2/NwB1
DoBQE/dehrcUQtQuEKYFajBOWj78a7hEnC/nyavzWOx+lJnL5Lz/qwRU7FWZhaawu2K7/lK3wzzF
o0jPBM1vwS02X0Cwn4K2JkpPfpHW+fL72g/k4jRn2p6cFzI+SAFalM7nEN/d3djCLIuvGdzavuOA
ZRpWAJ+vwNyS/TwuOENV0BDpFN1HZOYbu9tmbNfVnEAyJAUbN4xB6cFbYjzTXpoxwd00JfuxJLsD
5khH5er46I1DfD6tVjJ738bJYpvl4FQXMTBO2gYFsH6b1odeYQruhRtjtn4RHyf0A4CbLo6KLlkX
4sehkXt9waidKTBieNBtKrTAnHMX5IBAfXz5QVcWD8xbug62n7GnCoSl+UfikVRd/ShXUgr4Pr1u
OTHeVHcGrKIqxrvSsL6yuYnF6ckyJcmQGah6uABbdRGCLdB7u6CM2u4H6id1JXYxWSJCtrMaQ3mU
5sLZy8P2UZPYR+4seVSl5sjpVX1uFVv4UTHxhiByIdiWE936S/DNFIDavgDCQRhQdPAzWirU4dIx
NgTp7vig/Xo3O51JkAXsfIsmOcwiAukSFLF+7sRGxqTOlY78AYYyrcJkom5Gm/a8UilU2pC9ZQcG
QCSIjTMXoGVHR+bQXzO7nSL5gWYTi+oQhAcmALm7s8u4Du8Mk4VPfELsCDSGZYv3AauHNaMWPKAb
V07Tx0r9HUKGIjiehHv4YUUg6zvymEK2j6jSP3DfUUQBs8pN9Kusv/8qUYsiADxkjultzhdcT2Uv
whdQBgjS/LQxyJ3g1fRZd79mh+9fbjsboVBt/a8BcXJywiVNZopvgwtUZmVxwz4L9j/GMsnoo+8y
vwMgNtvqFBvsVIdbngzWFA8/uIzGeMDSYCPrHwqFSCgx86PTZ6HQYs3fYx+WLNzq8XxQF8jm65lf
MSk80BMG+CBeTdsIUmoPmBKykUk1CRqlGZRB4OZQWLsnvSwgzncpB544cgZDCEjh4XEk9bJFin5l
+YnjaQ70+Rc2nOwsUvINyBUNwdfMT/hwjBharb1HGreTqeP7avDOwmZFEGRbHmg4y0t8g38UxnX0
7AsxeQa3ZjaMygJt8aCaoT6pbAewIIGFw19D0pXGqmMLQUP+02S/JLEa/TVGh76XELLUqz6KufVV
Vr6alhpn+tf9cathK6bBMfoV/92AdnFJBhMbx8xiTZdoKlQ+puYeiEpuu6V8FgyUhOUpfFOX89EN
twFdoKJC5W0KD2bimhLx7DLQRDNGkEQ+ffM4SdXyJFXIu4zi9TsiRhZ+/0eT2EE/BuHPBrz/Xfhs
CHOGk6wLgVLOCHXu1Tn24SLOE1T5cWym5N13nvswH/FdXe6qu3Se353FfuBD+KdDW7Z4iqzQpupV
oX2NXWFgc/gtx8JQrik3w1L04hUuH5mpSFLE4krzJXNJeUSX0w3nHF5LDb5FYuJomtaYTZBvZyn/
SvA26qOlfB22J8BhSmZWdp7HwvcxhxUjIHXJpuMV0Ex7w31zC82xvWqR4nNj5wQDevzYPNjAlzVN
HEfNh5WBuJUObv+zWhwQ8D6GLz0Mou21xTK3HD0zNBjaKDRJ/Hbrk6Jt+h5JJcOxeaWoBnJFBk7Z
8ajp2YPgtdHswJQbUimnC7qWr5nR7FTUrftCi66vBCdn0CdISk509QBe8ix7FNPFYo7dWY5Hm+Pa
XQM3ppDpVlwsUCkYC8PNDHoVwAe/X9EJDt9JBWWbNTDj61pqQxGwWZBKfyU3YW1+HzWeSZIxY/Te
EtC9mWMY1KAOkthWouQqYfH9mZuaJROoanTWdfFFYGw0AzdRjK4vU8hCM9TQCSfBIZSspIQO1RaF
QsqGtf+0tMjWoOXnusWmCVycmZqXdwClxyP/k7rd458ocz8uHRpNYnI1UDjdnW1hV5Pt9BZK8WLQ
NGCe0h0TiQM0+NDSkpJ2/KmtVZPv3RshO32ey3iP8jS1WIQV62t1R9W4LLXw1GrnymOYn7Fh0OCH
eG+40Ho3iNTXvIqB67n5gfqkwY4jvJ/ntv3q7fGFQDcZgslvG/4xtBvN+rtAqRbGF/OZEgROmWAi
nrWlPb3Hp//UgNLafQhZD3DEtxK6E5YwrXnkfKwupw//k9zrLlu8B9TeCWk3Y4mg4PVCZBh6aWFD
03rxWV2CCFq7A8olqj4f7xuo683rYypcl1ziQ9PKxeMVVTpV2vL05/swAETuYwDEeO9nQqq1mdXJ
w2UEjXlY1Qx69r8PzC9Tdv6DzYSYntW2VM7rzmyO5MGbfTEYEhxxeGulqArQEFbqsjhiQUYGDkAf
/X7imbEds5JifGBgMcDUL7qEph2rO8Grqz7u4jF0cDugheOtkzr0YPxKBv6sg+le5l5UDl798E7H
cU3Y5J9omUgXn9ZR5OkZ0SDhTCwyupn7GB7VqaxpYflAACqtlYA7ERALSr9d2f7wxdWW6lYhRCdk
U51uUcZA1ypIBtuKAmHPtnb77fFUJtFPu0E3/m6IWNTuSxXo9FENjxl23YnPGF1td++tL9Q59OCU
nyJDYp6FB+xHhmnOdb09uZUCAMbHcOgsn+5204dwgLflDTJ8CchgauhD8EPxCaaDBscrGjg5V+c8
BlvkzLBJReovIgnYtZz1HTxoPvf0oRPxxcmJ5oC26PXnShhqafpO/cB3j3xcAnKyZbj33dxJsjyf
/wUPHSBeIOMH1vawNuEB3NEnjxpfT24DXDRSu0SpRFeMVncabic+vrMZap2U9Oo2QyE9my1QgyRO
QuhW+LoMTpV0DMlswcCv696pZJSzHg5doc2oytj2aASjGHWcPAVZwi7Uagw2MLFwVWU22ynjlH0P
66/ZZSow6mtjjT6Bz5Lz5yJ9kM4znPU6pW5TEqrTdaBV8NhAxvoLa1lc5O2Dr7jMOgQG5SRnW5fX
HdYRmZYeekOVR6Xt3zJC75Ty5YggrmACK+ReE2PencxKD/v4EyQMqhNXU3pnnWxYh7ZccI5P1Wbf
l3rqqOIxz6455MKrrB3G49MJ6RL3lf5Q9qacvi2Yzh7f0GD5RCxEKt4qKTq3AnIq/c3a+DsnRTYP
Ek0ko3VU70q8c4QwxSZKBqsqhb1/CDqnQT6T6g4R/zbq92DpuMroiZItMw0gRS+4cfmxq7ULKqsK
yC3kuIpXDC4iP5IS5Z6SoqQt4MDPzslyg5greUZRfqp577rDH1paDBmd8Z5ZDwU896aYjLrII/TU
sikvJx+Ko2Hf05yvzu55cy2wE0gJBFgRukM5Z+zTpqS+TlyPf2IvikpJuX0dJgJjvxFGnsHBQ6O9
qVlheMU9f7IO3Prn5roKLiYfD7/mCiXZBv34lz0TT4G4aGpzdvDj4/S48S3h7iZaWpj4LbrH8iYB
zNVV9mkSU97ekJkmv2FKUZWW04GbhqyIejg/1RBIOa3CqMpJgbtBDqJcXL9fg+ieH2NTdjXW1Z6k
Ih2uvXmHPedoVhaGkuq9vNMmRvUURta3vUPU0k3Uq1YMdshbkEElbFuQCN7FtfVvyFtJ9eHAzCOg
nlDc/JHaTVEFwZPTNnWOc1U3Tbhhc9zLiU97vlXcoPvSgWj2r5vO6A82/cLhtkkStTTe+GMSuvb8
D/wBE1fedjrHkNCKNZfoSGEx6A32qeUPXZRlPyczlTijBfX2M0OG+q2SBLT9qaTnePL1c35Xe3VL
rjb5U62o6iK3K9/Rc8YEp/miCYKc6+6SRiw3StrPmPJY6yenvpqbqxuJJMAxYnfGBt0QoxaFyaml
OwbeorMxrUVkR+7dvzRYT9nGqVAoP7Z7hjQBU5X1jaoLhdSb8KljdcrdaR5cVyep2Z6itNIK4h2D
tc8utI3uTzMVc/ILpamVQN+wfQAApe8XkEj2dd0RNC2uSix3bIxpHpnEyPcubxa3atK6OnzUdd0L
/6NK9h/JrKGBGx1FOhBUAcjXl1zAJLKNxImPt4lM5P0XtXbx+C4aGKsSm4q26sWgJChy95S2jdVt
wV6bt9HEX0atLPqlx9Z0+W5Hq+CYVcP9sogug8B01wmv49iQYu68My7iCSvF8/vxcKi4mB3fSDSE
T7TMNmN+/rOnDyt7fG45EIVyzXPI9dH4/AYlICpqIeZg7uJlSOA0TbPA2VnNuGdOyHZ3eYHFiID6
I9NyjUeioyWtYZ1fFfZcaUKhUkhDjWdV8O8bBXZM9iIBlS7IF/H6VENyq1I+YjWnXdpKSjEWOfN7
r0OVi7BfZA8nhpCwTVqbwuHgPtm5w29MK+dk9i/sSxkCFBnrxhr7jXLm1YPhWr3Lz6A8aW6Vy51E
N5ry2HZBrSA7Yh1iQhFMJQyTMfSXLG3h2iaPA7lLA9tG4KV4OVutqJHyG473bgjz/Ka/XHitb6N0
fIwFPq+//vpZ1a0bAFZoKaN5yeTUVBZ9XB5hM+wQENszpC447ANymZdFIT+cShtwizFiDd9WigA7
Hap5DTUOk9btBR7OhR2/4D/8nu4tM/wwajklSME7J2ss6DZ7w0iWMlhasqdsZwQRQAo/TCpmI1bE
7H6M4PbOx0kh5XLnwdDqPHRsvuINW68c/1aYGHvZ56T6OLsuJ5o13jZWKBL24MxiJSmoPvsOt5lM
xyaM/q4oYFoCy3AcdhlKMDpvMRpHZqBsxTiL1cuAnuA9NZZQPdJGGmZTssuEBTzhNcibZAS1gZM4
mHIcNMXEsDW1q1dYf6Q6p9QSIE6okj2+FIPARfXjxelr5vuE+pK65kNUzHYMDjG1aCCUbDeoWoqI
bGhlREuWYYyap98mdqT/6LZ5xGG2YjrxtcDEQHtQM6BBi2eONnR16bVxIk/H0f1/oMEdyRW1ZACo
efYyn7h35v9lOPMcIKGwBItqyK2DQWP1QImEWYFaPXzrAENzCdgUyH+RutECXpDYXKLD2YUVvmJf
NJKF0SAh7/FVUvwuDE3rFJfCqJKvoQ30V4FEum+nwuhw5hLv0LSsVprmAoBAoQzJhp+VbjBBq/vU
a3d1a4y7hYuIHf8lJtVzqmmXZOTfS4OCXtItQ1E4YFLH6+cI5/DVg0Q/PXR3TEQlhgYD3PswKoFy
ag8S4wox4h9HQbURgOi2I3E6SyVhP+UZA9ln9HYcsSuk5K3J0R/BcAxV1yxvxy7TdlFYzCrM9T6i
TFN+xSxLreEvjlMAuXn50ACxvN3OIS1kv2fRKis37JjTvenPEB5NmDTYp+ZKsfAvHIXmjg+CQyvc
eG35MSbzi6YiK0VBLqMej+kei2oO6o43HTH4njIbfHUpWZivIM34AYG2mjT1NNDXYv9FhFzXk1o1
tAw8FnmBzszJNhjvUJ3VQDAFrztzOjs04eHe/7S08rWLt42KI/4JIv+ztQ9bslnUS28pe5Jzhxtz
yl8ub8IwbTc/Tx8ztZ/+SaAppePRZw1Ip3tJRQ5kQLv0agTsbdr4aasaUwwZYYxsvxPWwjKdV/5Q
y2tzaiuUKlrxZn/yRZB3wvaVsWbDQ4hgC/xftpjtyHJlGxVO0DLVJvvzHtaFTK/6zLsTLR4GoIZj
4R+LFfsR6zzvyXqydq2eGJuC/dZ7HUdFWWjcN1FCZvUn84VVajo6CxvYOQiFh+MYGx/M9TVHFSRV
t2K8mDo8mF59yHbpWZMMImfedOOg8KLnND9pUs67ZrUn8V/zILCszYawDq6KSLATNXhcoYx96xuB
oye/odbIwuZvOSFiHddx2+BmA9CVJkB9z5+3YsfaW3ZlN6RfCcEv67vdTeTw1U6EooWPAhS69I/x
0NR8gy8mnMUY4QCqQ1rnp5eZ+YRftac7Lq7/mrLzG2DsaJgPKjIWd0T8IyLKE8l/sQY130vdFMlm
SR1KVeUdG6v2eduT4jg16QYHmFoKVhFjV0w7YQE/nGPRyyT3wuJKY/quCrBwm8TxjgWnlJuWVM4Z
F1uBIlHG2l5wGtVbgHxmSEHZ3lcPI2VAkRtiZK/6ClDXm7zuVFJ824xUWQWkR6qyPqMymRcw6wGb
9UX1DggSmOQXa0OS5yNhuzl1bNnMbMQPdc3cx1pQwBcBS6BsCz4YE5sVH1xWuphAKjsAp3bjVLHi
jzNdc+OL/IdDyxiyP+3cAZdz9H3ZWoERNj4scKoSUKZ+u71WwktsFncIRF4P8ritOUTMBNedKwqN
w8AHiC/IGDPMqOYU2jeKWiGp0C9RsrAH2gJc+OAZ0bgNfoy24+JP1+Gah+oeLtbg2K/zpA5BsssN
FpmT6PIL5Bs/Ly/FqSxyAmqNUncS0kDIcnsgaU5yUgW6iJRjhid74GPxTD433MobcwtslXoNQF9W
nLMUevLHjOhLZckQ0pJ2Cicll1G/maqRELyg8mkdWQCBdj6VTmvnZd6NchqTHj+g6ETGAHZ7kIr5
IyoAzgn8yQbZ56GH9ICjnt1F8qrQaRIRO+UZwm7z5vlbc/Ccl17I7YxSnHh8X4MS09d37D5uHgeJ
OEsXZxIPmrqpXwf+0mfqJKB4YjcCE0SweFG75e9uldbuRF9wCNLHEOu9MKy6FIt1ReGDckbbnbju
1hX3LJ9nX7OvJ1bJxIJB7eHKb/ScfxGU9EB49r0Ku6iZsd+O4wrUyBbjyZjhY8jndrKf3VCMn/x5
6GVYkJ7hzp+gyDWv7CEkErfVzotImdWYYqsFUm1OSIUkT2xYUUH0k8rX65hdUC/EFJGeLRQ6NeR4
fOW/xHHB3MLBB+ws87/r6w8eK1smx2QslQAQYF4j5rAcwqrBfsmzmU1uddXBdZVLCaPPb+6uuVG2
HR/F61jMjPgXSi0M5YsQ2ovwGURFbKEBHeZ/yupnLt1XzbcgDnUPcvkfD6/ndvGze85hPnzXQYG3
UeFeR3ZFDqaY0mlt+z5g1G9uWDb/Fi3ysv7DZfrG2jsNa4PoK3uJDeoc/ODbDLmZlgqwpWnc0Vc8
csPs5v0qxSSf2+vGeP6Mh8Zttc/Gc+dgCCZKQ1MX0+UeTTMQMckAhz/jARVRvQWYPWBjHtf91gJ8
xPehAlpdiOHVX8VQV5ZiumjogNl6hF22WBBK76qgI9dYiitR+5j1Gxy0Bk6ljJN6I6pTd8BS9T1M
hybTEWuXtPZHNlCN69McG1TvCui/8Pw04NZKY63jARofbx7x0gXCDkA/Hz3fMILTpOBonE8nRvRR
HlngHVG3S9Pj1zEyL4EubQJdayBPw+13Rrn0ToMqCRaOOhZN0xxbPSCXkgT6FazhVlCx7pWhQwmX
e5su0DStQ+qHEaw8uGrYTe9odE4NtOhkQLeHnHRnzjUU8NlGJSYy2wDTKgVvetHaWVn3OG0GwiF3
OpHnlcZSAt4iWpeWK1F/mnmzuttMSILWpVJYAaDFSkJkORkCfxAEafnPdDLSfnE/884Fd0ZuFiDc
zZhZw6icpeCzo7kDYVhlYGPovVivIZ20oCcuCBDV3tYasYxLdG53PL71dpRTv/XN3fVZOKMjEzuo
F5UcijjJyEJM8Lhlzt2887UZdcxNJuyDLEtqzdTKi/SLvB/q2EmuG7rnPz2UUcb6ozNExjGcBCMp
cTRTUjXdKXsuhM4buqP7L+i9RrWfqnBi9hs2IDAZgIaiR/MBH3ga1QuqCgP+LHBF6UbMS4i31r3O
quDDcUJ5Py4nurR7xwJML1Nrthk2N0lWAtBjv9ENsDttRQsq+YzLM+kBqEc/D0oBjqoQ4AD569G8
LtlJPjfKIINVWh7NVwrEhjrCpugJPWT3uBHaBjGGQ8N87cF6+gKkeWc0PosW2p+bLo5xjwhr6IKG
HO36GsqcNNq2dy7SDWokbHfHjMCSOF192cfpdCP3mRXwhbqX0xyVQkt5moEd5JCphVvbySD/N67F
YKvMaqR80u0rX4mtzwQ5nYkc1rRF5/gOZBM66Qj9C37jdr8SQGDTKbOJVNyAQNjSnapGqelJfFcy
lSBur3MRBy7ukoX833xgShaFgRZCbCijq4J8e1u4CMSl24DnNJTdv1uco8TSS8S8I9UqIM+doESM
MeoB00rGKxWKmFrqQ237lp/ZN8ELRHntz94+P4lI6gM0b2keHjkrAAfbk8K+jxxDIhbNTlOHC8R3
x732r5XeRaBH4FnUHnux7G0LlN/ZaZgVdPxVIUcGCKVmmLdUgrOjniPKQQtzSfX0hqdQIMDAi6hE
jn+8IMu1U9+GQ2i/2xbIfNMAD8oPlZSEj6irrT0w3kUg2AeQ/QCYuAnDEQq9Wl/bOUcx8uwRgUuc
v/W3v7Lh5TUVHl9fGctiuthig0oKGOkxaEdLtvIuU9sfwoR4vYOCOip2Yo2JtgDgDIW9VqDrsMtm
XZ+ZC15xBLHCp+rYEf84kuVThcp/JVsdR/+WJKwOeNgzOuw2wb/WxncRNemX4qnFF/fREGIYPOOF
RpNAbh67MOZSKJ1vzWlCUD3Q+DIVjsTEkaj7s7qDa4gBm3j+r1uzTd6RcWQRg35tlzbB3kFUxVsw
QnbuiNp8ixuz+fEvv2hLmmtuwpZhxDYqazTEJphC1GsxHuVveyPoE6qVKO6z5Jrk7VqVYDxu20Sl
B2Y5cK5bGkJp6IAQJriGGSp8OuT+62JFS2HEI4Q0iYjw686LMEiZruk4quugUP8BLfiEeXNKNVQn
gIFoEX1lI3MOZA7HwP1MbiMk5vhcf4CyEmXQ0Gh293OeIg1ZaExg9fC+pMAsB5aC6qqyD01aX6Xd
nNzIlciQqhVVedT7z72SJbEB5foRFuYrabicFcwz4yXwhIEZ5KcSUZ4/40BFC071xKNCSR0EpzvP
GtDIRiD8l6SH2yFIXSOUeTei7oQTqsIRdevjh+caK91I3dFJ14zIFm6PbHSGUmmIIx28/RMufJXS
GNZsXqSQ2KvHYHDVhfSpNRuIZ9ThPsvKnVoui+HMcC/4JDxgiYoq1tPfGu6b+m5i4f+L0uXTfhSE
3PONyb1yyGHG3yq5PLCZ1N5muF2yvtQHKOhNnaU4zOgfO7MgRumZvjnCsOV3TTvHAX/NWxu0UdeI
+u9hdyJQENeRE5/7YJtppyFj9iOy65T6+PzstqBR/Z4FDeLXjSgO1FOjgbE2q2u1i3hmSy4+h7Hv
+cbLD48qkNqgi+4cSub+3CZ8gfORBjP+a7amZqSWTyhcyrxNRD2lik2yJxzVx9Z0M3ghj01GBhgK
G9heEnSLkvtS7mPK05JUgCKccT8Wd+yGU4YCYr1P7mj15Wi8Qdbn/gpvkSR3LUHC3EqhTRhWF3qt
Cu3KImOZ8PNP2UwEieLISSk37uL1lT3eDBGXopQciZXxyQuVqmPb+czwf3Dg2f+LBknDqvnH7MXY
bfHJxImld6/idM+9ATG0ocxWds18ntnIc8md6XZ2SBs+lqsau8tR3YLzvQESWPtg8Hi7hWZ3UvAq
I5VbgdSe+1wbncxgMbSeXHxCfiZwvm43GGiTM68oem84tVbRB/8JXxW6SulLW8Xrk50or7Umhibv
TsvrTpssWDo/tuo28Yt/Th18FU8LWLr93F8YAhz33ODxQnZifeLoAxVq2CGej7nky92W2gMHnlmG
SnMLpzuRxO5deVwWsknejjkcDuLTRUvBOyp7MsuJJZ2QyiRtU9Fw/TouS5hAZ/3FWNI8BMzcJs0g
o0NXdw3lLhrymsZkPxHUZsa4NlYuu9VF0VYcsovEB9v1VRwaY9cZvk2loe18TZxskFhyFHIGqQWy
xt1BmQ5Ye38NTMiqZRQ9ccvIFaIlJVddeTOyroA/Zg/4Y94F01lTLdSPPrG2/zW9XkTZOq24PGdY
Owh/Gsfcki/q91bxJzCs7hw3ME2lvjy6FE5G3zceTINdnacmDf2zdQYDu5m0E1G2iBPz+VVEBAf3
8WeaXarZmj+jeBihX9wnysxd1EVy2R419PojBWt1gZ57Qs54i5F7Jv1gyFoROLAnksdKkOAdLYbW
DYyTfh+QeB0V1kIhJtflLhTOAEEJ4+8P38787Ldp7876T8dBBrX5Jn/v7XfroX5gUEyIc41ech2C
RP69VhyigqeLGGbZNTL5h7721w4U2zVXUNqvsp9gDLdT2Lk9ohz9iBfeRneV78mQ2xvY7I+40oc9
FSvFiIaYk92pCR53nSbiYJw6tTS2WRrJCi2dhvIBG+qfWJ4X0PNXCvNRC0U1vbcxyj7EBttJHbSW
VLvoPqV9A27hO77tPLyBbgx9oaqfBll+KjTNPwW1o87Sdg+Xaxf+oLihVb/9nI2AeuvBom/svTKy
l3JYgRFPUgk6iYnzFos6dBmYhylw+rlFvHQ2XywVAHeWlIOCYyQmDJOpwPVrsZR+vhg7zacMjAhR
VLbtgPgAejThJSyV5Tyd09qCrcUO9VBcHjdcrzoMuZNXUNSnkb1/eDOK3IuD/lIAefX0G4Z66Js6
y73h+1zr8w/Wl9utpYpzbkx6MTtjSekgs700j9HNcnBpZP5zzjltzOOeTwVgF5riz4sxOdx6RReh
NFWNkW38dZS0r1SHfhn5V8hlcGg04GqzZ0EhcWKJxdOuVEZ3PjziZJc+ob/gY5XPOyfwtfaAbC3S
pyvitL+goFY/Ove8jKGQRYSxxj9Au17uvV5SnmbG9Re3sh+oKOCRpupD0oYN76NCro2hl1OqOcbr
kYfJ68aTWAadPugI5M/bO2Nr/Njqriia5EoGam9fKINZyjjhcA==
`protect end_protected

