

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mfaJYDCVJ9tmCl1qOjTk0TJerc0+CZIKm9a/zNyIQ4axltn0gxS4ecX4Zo1Hni30YBnj26NHIuBB
AOWQWWIsIw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fm/WgFN5BJ8I3UPgZJsI63Ae2cgM6RGTxS5FNhYU6XXXHkx0QJFyFRoU8CrUTLTBjuluj0orlDN7
b6tvmS/b+t2pz/hdtIzowwG7ASfmAm2Rz34QQjDzigPzCKTFoJ3AQFyFVp6APJAEpQMDshFJd1bU
o90A7irB+HRJlROZk6Y=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y9HW81s+G27R4EgUduReRfr2wwhFyWvK6LL9tlnP3yGocqrl4RiI4y+WWaJnw4C6dS3iiGHHmeJ7
BOLahMIyubxysrUfns7VGho/kNW6ikt7VXVZ5L5jmw9yuPTyIBFncC1xqSP7xNaS9k/ZAm5Lw55K
H315o/JmcCyyn5HSr1jVdFPIEuJ8RryEov/1F3wae5vQV+K2pdDVM4yhMeYiSV3rEXBJQCXsB+F9
U7k3P3lccYSLv8P26y2VMgzFU41xdKGkbGHUS4T0+mHvvMFy+vHD9LMvUteqPYdGOQNLjruKlAs2
AHopne8jFhsR31I7KARkwyENb8xzvOv8sBzGyA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
peROq/jTTnGKbWA0WQKdstqCMBnXCQ/l0MNC8U+wUBEgSuxXmaO6sZXlxNbYuvF5VqsLnRWixfy3
wh0htdw2Fg9D9Qk9/a80vu3uBTjVWr4lk8hrLkJnvtq2qtTfYk/OAyM32w2akdkxQ3wbWQ4k1AYN
qu5LIPFvpDfcjJlhCIKstIQm8wteJnd0cow/vDk3S4BJNKAzSiiXErh6GWgVub7ULXmltrFcrexW
PVXlGQKAGU8jNZpJxJZ1WZgcQMimYvj83x1+eJZE2cVzV8Ig8vWL+yju6Io7b1mfyOmpgUuApCtb
8AQsP5qESwP/N+mwguWx7J8Q08qdqM9x/QJkcg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o4FY5pOROZ9YI9RA5p0Ad3kE5yq0whzakHnr9rZ0OajyGLv1cnb96KSQ32j2VgDMft9OzYSZeWbt
PxyURKZ6s4QpIthjKZ5hkZ1dX7jaLHWszkXOn0aHalLo0oDQq0RSEei9uei7Mg0qW4DdwyOjJcD7
0tCjm+xUipiFJ626wm0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Iy13EbSeP18UOZBU/fyz/ghFg8ztq+t53D7w9iholnS1uDKpOjzlQvaeEBmYfRXs5NHQ14Pz3P9w
+hmZDs+uzw8iMA86Fp7fhnCuPzX8/LQRFToaDqPBMIYa6DRqM1d3Ld1ih9i/AYotsuhbtel9kyE1
dpbRQDO6rz2jrgw+W1kKiLC+9RfHxh4rhcUUxHELzdAKk4vXRmckDFXzxZPvws5ULUdbGjwbrHeL
iXS52T7AJBCxom553aM4p0xnK2cy1PSV3ogeM3U2F3Xun8eEJi4+tWr+CR1ygGtAA5TlCtAGBvlr
27svGBQX5xmja+iZxtHHExze4wnvgGrmhq7w3A==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RVccda1v0fDhNCHInFVLDT++HfpYurc6dNEqM4kYp87QHa9Ne4fPEjHI+WvI4PAXowO6tW+feTX3
T/e5eJB6pzI04jJCjK6p/D781dDkkQoBKYIqxJbhmeoO2j84jr0MgmdQYY5cgbbaXIuN5kkFGQSz
Eo3VyGRYCmtfJlean9QS+gf87lkNNT4AKI2eG3SLkZXKRluUCldaUlqjtjKrif8h5fFZYb9yuwsq
fhunSKXAsc1KYi6QHcvOL/gbHo/Ilar3OtapsZn5TUt80BJZAKvR/SwXTTXVXymePYywgZdpaaY8
YYWh/hB3K51qvTWtnQTsDu2a/EjyqPwE0ZFcCA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ay7+KMhXAM+UC1xDUAyP7o3xWwNKph/1SVNJt0GsikZJSSnNHG4zsI8jvwLNjebEEu08CqdnL0r5
ysc20SPKfLvMpMvniIth+gIJXsmroMzwKRsuyL8YirXLf/GY8pGp7aLrsCvZjSURGqBV07M2Hnj1
d6antFfvhNW252Xw3orHYwuz/Lf2G6HLlPpILmo8finQj+mGy/O6EW+tu2HSFoOThajmRh6XgeYv
EtPqisdn40Bo5CRpA1oJxOuogvjjR7R4h19uU7NavRxTlXWAc9v2QpkQZeUvwwZSttxAMF+PjrSb
vwJLBacGapQwB5KVmd1Cw90/LnH5fHNhvEKDLA==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qzOcFXO4O8zN9faGFsurU3eYSecabz3rm5c+LOHjNccH6vkSDJWFpMZsUESSlHQaqMhHRVfZdUS5
lGJ2RK9B+WPWUsy0ZigEqRrK8Qir/Anm/3u5fyCH1FzwryCyo7cm+I2k8+YF0SWIvHVzK8uvNd80
ibPe68fBwOAMylrWShcthBrq5gSqHohNeO8bcRihn+/rRxXxUIg3X5JdCLKA5xMLpnXPZtF81VxF
qBxhvKrrsPRjuNDEcRmff5TnFJffnST0IrV/Wrpgey+qfe34kPc/YnN7G4IcyDB0crCU3KGhkfiq
yoXrdivJtqDdYo5HjSra238d/I8AmW/W9cSGVg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23056)
`protect data_block
ULnTY9iIy8OmQlK70cBnPOIiacJNFCO8L58Zw8vgkfjiTFnmWH68mTEVWqQuPr9qi+TLplishmqr
uncCjGNM4lVgIdewIGakG9ZXKWk7pl50d26wnvyTwuUmdkTZdO0xjDuTE//j7E7Eib3SO312IX4V
JoajewQuqBLr4dIsMxfBlZAILWChncpyUG5ZpQ1lZtJmwwgP4XJB0ex/l3cCflrrKrfVEiWatA5W
bPOD0v/QSEFRkhw73hXQEARrSELFgNd8BuY1vEA4rm1rJgL303JbsOFkqZ1dS+fb2rXbRa5y56gk
N7YwYzwG1aM6+6x258nl+2Ma1zbuwS15pVcMHteeGuMgrZB5qiKTspKrEsIHQYf+zzTvOKfWG7NS
Rzm84YytmOCE3gD9wGdBcAVkv4tz8PyUJaY/ZJktWYtzBKN3SsAsEHyz3Tfj3AlR7CV5cs0lPMVw
KVVtA/EJdqEHgGXCZCS+UyaF/gvGoID6+egeuLXgZBaIGNSGPWKx+TlabX9a8Fbh30vOMIScAgFX
b1F+889mvm882wp7j+WtPeogFRlpy3+XSgWQ3Wnz3bRetOCgBeFDNORXeL+OUe2u3FTQswayw2yk
2GRp4WCiIdaz1WzUNWfeL9v+btP5kewz3t4+ZJ7c1xH8nJTvreSohuNLs7NCRZ2tbuPhVaw6ICu/
fXMM5aci/g00uq/DBZjaEcsxqOILBZJHjbDKScAvaAzYoi9QkLOz5Zt9BCTeDl3P23JWjlJVDyHZ
WEiSvZNNxe4pYQNxwQhxQz0INtlNfBNgrMglI+5FksTcyAvbofiIq0AfruBxLQjwwaEEPhcyOJOj
Cg3u47/Wz2L2FO1tjaZMafmqjwATp2d0D0eMJD7sq8zbNS/C0HkSEycs730vyv/G3SxmACM8S52d
GbjiMRqgG1Ig+BUoyBsmVeLeKdNlMVxPCmk/gIIu+eDi8D3erkE9BwWYpXevHETods61SST76uX/
qaGu1BseY6MZVi/bn3HmS8ePUmkDFgSV0kGZeTN4jt8y/xfCruRuP4V8ogUR61HmtdLXZAx81Yzn
hN0c/7iCsEDoMgTwyjjIKzLMotWLJpjRN+xNsJsqcY6rJRIA2twp941gffvcnWmYfHGmvy0dXSZ4
RE1G42zZ00bNnQjbcdyt5sOe1IILbscUa+dG7VOuXizdpjCDazgeCI0dMUOoZaFXDxzIjfmgQhKm
fbKneUeSI4pa++J9H3JHuH0uZ1ABChZCFIP5f1qfnCJBbT2QiEEfXyfH7xcPiROXRd9PDCxziHRn
fGX6y/iBgHEjofeggun2qOW2f9WIOkBk4I0+dOsilrlWArWnjmGAqSLxt1n4Ke5NKfrG3ZKxsBsq
i+uAsBqaU9yCrB9PLzJnIuiSA2hijG/ycrzfDbu9aERRUNUZF+W71GL1RSy1eSSCfM1FqXYQ5lNy
FsnSps1jjSoXC6Q9jYYuzpv+/cWOWorHiMvjRjqx7Uo9F3BpW6MTzkO1VL6H9qbdrO5oQXEKkaQ+
rrQeuH63w3St6RWiTT3xD4AX0oJ4pNEsagEMYC3XkS2uMLc+oKAKJ/KnCcoOJEf9MFhdkr7NBbSR
71Ps2rX2PyDN/1dOPZqE7DCiVT7DjB2rd+KpdjqjOHJU2HvOkWhNeDd1EMJ3/cz0vw1JdY+y+DS6
m3QcIdNV2ixdzg402uJp1XFRAY56ru2oRWYw/PPJ85g+HFHJFYucTQIQfM8MbMc4a5e8imW9+btw
sduEr8rWlANT1xp0juqmhdX8vgsy6uOk9sfw73vsrXcYCS1TTIMFE2BhdpRxtLRak2x/yxwYR2Fd
Xls7b6zPlRIjWQ/iqQ2Oy0oHSZl+G9sbhMcck6lCTj070yIP8JBZMJcgVU/cv2NUP6WwmP15zh59
KbQwlcbAAguNcr+/uxyah6vu7TGcug0qs66+hqPgR3lo+NXfGDWqZtxjDoyBJE1aSxFYTSrJZtqc
eXh11wwyktw4hcKehZOyozSDOYH72cPMWPxeSv8Nq+hAURNCNcuqMzvVaEj+IMA+2b64YQhm8nTS
6zFjYiFQgzPV9eJ+iubQFrShmMzqNk0yIm49krVCt5/TlOD6Y5kpZzbVwlyFRTccyS5EMdwvaAcm
MUtIuu9zzXA91IJ2718o8D1WyVPMtpmEiXGznlHuqpArKjpgyyxmD80qpDZOP+bwnkQqX2pD64Ef
Ic/Q/GvqqrBjUk4r8W4h5V3OqY2KNSrEm5BRiHdlBiOHVJdkCEmB5ywWdH4pdKpN/7MDjmmiL61m
WeiXAlimRQn6rA8T/YkhSh2nZRtJY3rIJH4/uesKwP2i46R5QCcNRdJZV19IJw19wjUiecMje7Yg
YpSU6Bz+Um2zCcyaJxDSCbWa+3DjZ69YiyjXngBlbebyqja2xmFtecyqdR1EoTCEXkh+VoW3LkCO
ZdO7l6A+U3HfNGRORb8mU429ZZAN3f3cfcT3CZcsHPSS8XFR6rbBkmccdV2W4gl56Q+BRRYhd6Rd
+njSEYQLhbiE4gM8JwHUiDIfjdALvupt1rGFihQz5zL7T8eJQofM70TpcVkYfbQ9s5cy9Iv6WUa7
xiNocrDOIsExuF945sJGqwOT1JzBs0IpR4GX4ZnPppmiKMD/NNWKVnwjItF7aMQGd66kmhRhmDJT
9cTab2cRBe86VsP8OqqmeAzADHXNRPhlYnpdgbJST6UckN0u3Gtsf9IDbhWX5AjmXtj/USat2So8
luim1b1zFdoKIkjxJzpEfwmoeVC3jZ92VYDwGnudYoboaf5Q9+6iU2zS2M5fmlGd/0y4PadcJSPU
NUewVsDsP5udq9Koqgur8KZh3Eru2QQD96BfJzhSKqizl9gUy0HYxmH2wtAqNTHQ/uDkyWlaUab0
M500MBsAEfPfJA4S91Aday2lhy04BZmF16Al33qjzvepI73MktkMnnQmXtXUxTihw5oXGsKni1al
nFjyNGvqpB+auboEBc9ppedBt4ODlbQG3+56oJZwSv8kENJxgAqm1LTbGEr/QhjkYetCIhaCwgbu
AKb+iG9aZoeWBCDNUzHQ+GcVlUqrXgQ/dVkyp0cUiwoLN+r9U491mL6hiYbWLiwdSEy07tMfXohy
WG67vTaIXAVhCGykGLuX/IOE+orNS8MNDH5HjnsQObTgRIU9hrOCZwV3LxTwsIRQiEHMidipZC2a
bf0AKv7C8fRP9bwZN995+3AO0za/F6kbDypkrBGxEXSm4YjIzXTFnWjS8cSNXPm6Buq5YL1IGv1P
NHOVu5B1rBgyMMQNhusfMheB99idlLneFIBLf/qyRexRf1RKUYtQo9RuYB6PE7G05xpLWO8S/MNg
3q50PssbENGoJxO5YZseRV+Ecv55eLlXBKfcWErEeptOoGtIcUbm1oFA4OuAYDVpsQqrvm5RinLA
p9Sl4cAN1e/kOAprABGn3iHflgDRr/vaosyk2BnrWRhllwGs8UKS8to7wFsx3K9gQGndPXnHupJK
mbnwpzhLqvhKZgi5jGuxN+neuWNyo2zpDPMD9V2Mmlaz7vnVNOJRAH/gaq90kqufE606GQzWEglX
wC+UrD6rqNrGmXehEbID/dbtCxfWKXMantfS7wu7l6fPkPou1pcuNBk1+DkjaLrQ1QkMYOPejkia
V3st6gft2Dnwc7CWp9aPtDGlte8LE4Hoc7QVGyYlZF8L/XrdsLrEEFlWtiA4mDLuelfb/zS+arXq
FGdweaA8czDalbsrKus7z3qphFXDJScBUW4zL86GEn5bvT6/sk9hsoBoK3410ukX6RNNcEBBeR28
hNq6YQZ6+DR43XKWisVWQkxmLE/wqIXZPxXtVtxY9n/pEyckSzsOG1ujd+KaiAzLFjjZ2MJ0Zj8h
SgutkaGeaMJGYhzg7CzQmma263BP7Z7pwhgJ6ulH99OWu0FLsbVddtoi0ZmHRoFk9fYmjNm6mB6s
V18oaD8fQJxsuM/f4jB4f2MXys+zXP4daU6m3ber3bHZwtmFEc2A1fURT6M1MdeN/GJJpHMQABeW
qFKNuIK4K355wmCwm9pV1sq7jW5LyQzgAMMmV39Q91tMYODTw6TdNV4cTHGr80JL1w0Pk+tp/Ct3
XTGbS5BTLgY8qPMg9KOdMkiBxfvlJrKl7cTYrEgWRQf6k3S1NjjGCN4C2qgNE5R/r+GL888mA0i2
UhVDuaQ6UXDJ2cX0NeaK2Vyu+OMSbgZVk/f1fBqaWeemE0OUgUiyQ1nK58bdpCAsnS9LEAyLnFlv
swBeRTcCqZzDsjBVL7TPhAjk8eFsEfSnsekASkmSfmYUzjT5Qj5pj/WKva9urbGh+rDciQEcKufw
zj4NUCeRS3kq4L2uyw2eb6gM+xDrHDlntVSBWre/mV/F8bZibdrAtlebX4Kzkbnvo23x4m+RzXzi
67zDbDVvd/NaTM6md1jnh7ghLc8yzhE0NKgX0yZxlk1T1gffGULQyGDaIHTsLZSDzfWcDoWdqWYv
G5c759dyhKMQ2pikV5lufZRYU1fnqafZRgp8YsICVN2tRLksoQglRsETReIYMBMNlIbyivXCL66u
tO5r+BTo2WbEu42rn7InyciUC4SXkR8gMqzMyRxVhBYPOlXJoY63WO+4hc7SrzgN45F+1qkH1Gev
fjbPFexw7IA5FnhXMhgtalPRbVct6SPS+xAGhjGyaT/vEHSQQkC+p6mDLGbbxjQiYzVGQ1c4CB/k
G/MzeI9gh6y8br9xdtf+CxUvmzmXVIVckzVW4TKIHqMc5wq49kNWBp4hN7pNRiT4Z2RFSm0F1uP0
PJtOy558HXKX1SBTZCc3odVHMyrirxieQsn0AUXNTiUQMx67VIn/20z+TWDyoRx5+IuCz8GzVqxi
9UDnfXoHwF8fE8LslmuAG7hTcGEhj0KdLUDeA9V+8BGVQ0Q/Fh7yraC+IXpfbP3Mk6Gz+Kc1KR75
+Kuvyx4g06N4g6oDtIJwkSBn1jWMIdssjkKolg19R7yIPcWHC6j28e91yEeVhzDWCoWjUA1R+zU/
iohwxnljv5oYXNu17mZRs2KZZBSAwRy9jlHnScJZ7Ci2rNNIx02YI6rciHDR4xnM5oEu3bV3zQx9
utjivn7iausx3YNcFCa9aAZ99dlqPlttf0yiBRRN5mCC/OezHExwRsfTAcgZho2EARzaEMH1b96A
LEyOvO9PyMXiasaw3kBVBbwW5eQ+cTaMkGG9bJURqbBof0Zx0xa5Ay4cz+49uI2O/dGIIZQdNsyV
cII21RJxnEkePT5LUyzecMy3HAUEcMerhBfllDLaqOpVRuw5ZsTWDvCK/0iOiw6zxTzdQzQLhDra
9MhqTV77aStC8kYduDAjxCOhA6kqklz8qShVFI3fPuVPRYqzdEUSRkzZ5s0x3tExahoMTJvsrzBp
z33yMizW6TRcOW6Z9CkAwHCKOBZB/Z058dvX/2FObZJ16+yK7S1pSLuc1I/RviBjFDLnnvC9NeIQ
jF7YOnGRcolCaHE8GC+sCmjNrMD81ZG4QBdt8o9wGcZ7pXonhsSf8J3G8UGD+fgNHSyf6dlFENPm
vhwFYObsKlD4Wv88SzGO/KgBVSBIkOwktGz5PzHRyVpUPJipwptLcye7ZVWqjpDtYg+tHb0tDvbc
3Q+rUgCs4tIr6CFoCeb8WBL3bgQxUuMWUwKDCkdpujYChRl7G4760i2ci4CnmHw6fo/R0k2ChEVq
VnZij+2IqKTj5eNd4KXxFGMry5JVRmkqs9ktpFxz7JpgCrhXO81m7+YGTCqNNgwel3QFmRB2IuuG
Ckb4Lg53pIgBRsvBK2rN6b+efsenpCLhfTZjh+lz2k6IUCb5cA//i71uC5cSFi63VYnLVyJ01pl+
iNp0fmUtEgNGyEHrangMZhnU6whGyvugBb9WDfweMLuZPQF4VieZBMDLcF2SiSkCvSZ6qlWxr4QG
pFA3CiJGTzkD/pLok7P3490FHSC2+tpoMSzDE36iwIafB3uSORQPu5MncYcxhWyrfqZsjJEzgA9o
uW2KEN55bvu4E9og8ABW56C7TUp/k13xVN9yfdbl9NSlm9sdYnlyWOBlXhD/RHFwrh/HMxaxIvjh
LrtSzQK1+qzK7RU967g/aVyhCKhtVZ8M7lJuNJcwPIAr1V8uPv+658t/c14JDUsK0W0PKIESzGNK
GhU9WKU6c7MtRwqhnDX9jOpW8pAk2vH/wkyz3A/OAnHQA1UphoUK075lwzYL8Q74FnxNu+DbB1p3
xUMwMXsukzFn3SJWeZ37Q2KlOlWUACRtww5nLUnPaQ1P1J1zs8fBI8F4aV1LpFCU4547RTTGwBmq
rpd7JITRx4D8ftD19ASq56CjUdhR5pFIkISZk1YRX30XYJrvMrqQBvdAaTx/RLysWqtA0HDh9Dcr
J9q63xQYlBHGnI1NqlUhQxfyfP9z1DMoFUsL0zQlo3prdAtfrEyQ71SPRSQsEEuc2DeRW1XmOOmc
187IfgxfnXMVDCo61aX9Ytzh3QbqF45b+1Tu45qOs/CXzTu51oQr5ziRAQPbCRuwx2WPFru04caG
h2g8g5Qi0IF/Tep09MwfuRWQjwIPm9/lQck0oDWUDsM/MZMyr6Gl+DGcMywm4Q9sZfaaNt1AC2O+
0HWBDtwLqnPv3V71oi7D672OcxtxkCt9eTHsklWAhSTiDDSVgLO9MERRr2kIO+rvsSCk9VWXmVqI
LSV8PgJ7+3V3vbVd3b6/PbY3pxKFxlID0haaQG7vQl/XlPDSSEjgp5m7rPNDsCY1MS8pjgaUn7sI
JEhfP9KoQB0lrhAFByO5pingTLAyf33O1XMB/tHlmfL88sPq9Vwi2VXJf49StVQ4iz85WRtosT9v
3UWhpyfg1UV3GM6p49D6RYVbZhehtiCG3LL+EmbXt8N5qKe7NuhBswAoI2tQ47ClGhdAaFKZAIOi
mupOxhspEI4zlN6bXW4lHpo3xs8Wtcu59Uu0jLiQ2OfMmrXOnjzSkVbamUyAqS7Zc69g5a8HSPf4
0i5z8TTClK2YeMOyEdtMouqmMck0XfvLbk5rKdhUtcvPjFjAqzNAN8gf8X7UwcbngiaA7nXxFqMP
MPZqJWLorsEnkQRlNedEQN++qlrv0FoUA4hxsuRaE+eG0KOxkUYYKJ2l4wdTohXIvndUcfa3uBCA
SAmUHIunIqq4hfNxPRpI1mld5oqax1kqZnulfByqMVuPlXYNGKa0JATG9n57hO4gQ3R2lvUefuTb
tyfFChMLZSoq/2P5J+aDK+i5DmXTc4B6Nk9VXR/UKeN6uutiM9wASoqaq6WtCKTDksCxGQM4yed9
2DnLyMipKwRxs/P0axta7SR9rdTsngjzdw21XXtCBSnG7U3ozL1z5f0eOE7l5uN5LvtenGgj8nVv
1jr7Ku5ZqB/JxLixNacjRU+ld4S0YHtoPtQzeRGD3ke/hms6CAUr9QcyPDOAqA3qiL4gjYJu+e2c
EZpGI9V2Fmz23rvMiV4bsmVDFBCYvPMBwgvSFZl3HYteftjj9Z0Zj7t4imFHDirxdB3E04EC62lE
ZEllwKAJQkGwU3rrrmiVXFC44XSBNG+irCO50Bj4+3w/7SBY2y3P3L+QQHZAnEURGP4+x+cXICbL
/5rvdrV8gp7nM5evfdQJVz0jJJ34dw0meW5KMUZV4xGWDMh60Tz2IV3zc+u76brTvsMkY2/Iu+8e
na1sR+7MEDmMeOIMqMjD787Z1dPURGiQeSm+Trgh6rFiudgBmEtKGP3/TRSANX/do3+PFEhxqPy4
/4Jp/K3QJGEluCW7GzzMfP+CrLj7ZQv5Pvk/8HMQo1S8r+9craj5uRsBFzuuqCJDRItDZvv+M3nS
sdy2L0dQry+G2ozfOqYmiJkkvxmMSI0Flee1ud7um+10c4vkWOWfGeJu+Tn90DjU4Raxi4X4ssG4
wxNWRmLk+n7WU5cy8x80auQaEfDxvCzeRKI6v5QXh53mz25JZ7U2iOwfUcaofu/fpVgrCuWY2d/I
wphFTElEvKYr43kGBjCxpuSny0ve44i1TAp6vfFdZWq8dNtpfp8llbmnpiKvYp/KBXTIjOuVEOpx
LkfIxcnFftZBbnyTazmNxhfxxlOxEplaglkfisORrPxCXxZPSM1oUYH/1rrh8BB/CEt8YSViBNdH
nyPW7F1ZfdwLrCjyed0fuHgkj3hPUH0bz8zg7dgo7eRnk98Ca3GYkYzfctKViAj2t1OVasLqGq10
W2VRMWnPmkrZDrlwbO3CEgWNh9BAj0tiR1snQ3rSrGIBiq8LZBBj7/nDqZ1E6y1VCMxDTzxy0Du1
8WO/WYoG7bHTbCvpMK3/eNM3syiOulu1p1VAKf9bg6MeTrJtEJydlR7s8rPLfdExZ6F2tvlLzTqr
KtSf5hqMLWJcwtsCaolXTfysQ51/kiiL/r2AMgaiglZWX2FdMZqJ25h2shG95UUHzO5moo96bcWf
4mE7mutJm4l7Vg2sEGgTEaXsXAoxLEHHe6lhGiQ/G8CWBboFZj5MaAeqAjrw16Pug2nn1bUuTs1G
+qrOAtPpDiF7coQPUAv2BQ3NUbkEV1XhOKk++BcuU6Ed3UqanbmQ3ri1x22SUVC4ZLj7PA63vviJ
W4ZJvP+6RTFY1+BBKgp3z7tjt4VnwmKPe1PmSLbFUBKFmNU/K3XmzbwqoS8FSMg8QATz7bxj/fY1
qrLJ12NWfDz4oBrnGxuIE8Rf1uk0jXbVT74KfzmOP5oHJTPbJYCleFGAMLUjzWdqaA9xc/GTndHL
g0BZbV3XcxJInVTNguv6btZ4pP0acFTarkfXUH4/L8kLa800U6SpNLT60c1aWEkfSX5ReF/v35Xk
QrLBGjEXHKZWFEsrZSTn95tU5aECLl8uQqpXpCWLmM4uX0D/D4opBrbRPycL8txz7j5LBnfqgh9C
mj6pmHvtowIQnhNAwwaQgxhDvyHJEY7baZG/wAr2bkZTh2ODyZB1kAO+M26ygj1t+Thllygf8W9Z
U9fyuoMy8KOR9MOmt0ghLhND8o3BAzd6NbVCnxVtQi3t3unvVJ4pS0CoD49mCEa2WZz9sJOTlzJI
gPjwGjqf6wJ4pSxIeX5P4RI2WV7Q7IJutCtlvhsfR1Ct1Ve+LlQqcxZzLy0+fdlsaJNEpBMz9RFo
MkwY1G29/DHuu4FiE25evtYKUESdoaM7BdUseAnpRvMQEX5dAg7hIsAkKx5uYeE853ZA4noIjgpK
RszLgQLLq2FAu+xJtUprmT1pxtiRHvYGZy1trAUXLh2F7NILTrB8abNJeHp7cIUbKe88FlSvlVBR
Kzo/YKhCmvdxYO4+mgyabXHHRaE3lQf2UldOhMRsJg/+jlV5HuJ9BQ95bdUWSNmxuzO+g5R6JSV7
4IMi6yIVvklwjM1T3gUyM4SaL2AJXgzBEvFWkr539fuRNeyMVJRJU2V2FypzJLU1FrvwRDjLWQjI
2VUtrB9sxmeDNhrNyx/3Z3RhY+oVtQw/vNhlPXS58XhLaUMmMQn4e6uEGI1UOvaY9EjXaGDkodiV
hYJwPob1ZgJeA+C+o5W+ybGNtfvSidHwm8bmiOJmzTSXMhsLbmsFbzvIAVf2ycem/uVUwQLK7V7R
b8n/eSl91h6IANlxmWTqsnVC+BZSUkb45QWeLmStSge0Qs4TAJ39tqiOTmk+lsEYb2hQ9EWbdAzB
JdUeCptJv5LXhFcx8ljpsj2XgfSfZEE3losvpStYGG0O0T/p9QJd/t/7Cn1F2s1YdBmglG/6OhwQ
tqWvbiSLCI3GTZohBetsCacUxmedDG7GAjfB/9ferdlcpI2wdoJcH35pYuM/Uim8+okWq4VGbj/C
8jg15llBLCXZ+54lWhu/wmSfwgi8bfzKtlJnE3xEGCTHOmRO2I0T2aqAuh44v/w1b6ETs47FmXvi
x/y67DZ7pinVErZt1THvUUKBzc5RHZTM/OGWIxg3U4mpcLocdXFOOTvq2pMyryWQ+So4L8kgjlhS
0mgnJ056fkaCS5ylfTOPnLFXHX1oJfaRokKrYrkS7pmAMR8ZedvLjR7/z/eCkt8jEk1QfBv9Ubv4
ZTvYYldIQJHYaaS/o+EbCMLjlcE03no5RHOdg2uX6HTKIZ3Rmvf8oyBU1szUG9DPEiGlNHVgGtLS
zX4J+vLK8nUZ9LPMAn5yjo/xtD6PRWadQ1PqvmXDbANHUPilQUtAzjt/wKkI+2e6pxZ7BZWen8kZ
cNl5fS/Ustzo+GC53bu6Dtkc3u2Id3fOx3eHWrotU2xWPuXCL1nk8RUTW/DGxCbYCFZ2CYXpKIZD
xCR1BEILv756p0Tx8jTDdZkpJmGiw3sSQ6bzUq2YPzFE8xpw3SM3b3C5I0ZqIkoGfEdJqHQiq+1f
pCSafENYOT/8YmRhaJKfgZ3dUs3+EfIWwbDtaIRo2UbKHSL4m/1J4d+5rEBWFhaAgcshyZJq7+js
MTndtmCa/aBtdsQD7VSiRRQxCgeAuToiz/m9sctBLt1TikhkMQf3pS+UBxkseYudnorQOUjdcMrn
9eFANJ2QILgaz0Nu7H5xyAvDbj7ogLbZMUYzLbMUxv09BjKuUK3QJIZVq/6O/yVAJTNWgpvF9nsY
bxFKQFvhVNz4QZ2FZfkE9UmaAZlJbY2ORLzSfel6sqMImOicHlOIKZq2vfgXac+TTwiRmR3pLLA9
4xHM9ToIWo4lOgixJal4+/E8I3nVrEPWNh4GAyqBPmIlBSSF1mP+cYbgBGqyitm3AfluLS4pxWrZ
qsNsPuB0x/fYDmIZVB8m+pJGJZLjxe6eBX0Lm9ZWHjrJ50qBYGsPw3seIG311XVUPRwD1eAKXxUU
SohaLLYP5ZQzKnxljKmRcyORO8rc5hbOL7djbmCL45e/fNaBRbsAAN1CP48IKsnAJHDaRWHvdVPj
p5ldVIbmyU4l1SDfy03AUbRwqbgjt8J4Jxzu+fmJ8QPE+1vngMp4pZ6v01uB3afErXUAcIR5Qvhp
dHTGdqflMJqR3MO9wsAS1vC76vo7VPZZyRmRHGvcO2YBMPCeMOmxj26H1Hh7XKn2qw4SY68qRNB0
Awy01mmSYnNA6hqk2gqM6xLYyPGmsg4IRWLyXP2agYXetm9aMHnahRaS2rSD73EcKMS18DQmci9B
slRkksfmB/kfLlgX6WdwKBZ8tjQIt0DHS9CxdcUoGNiFq8+NsQ+PGg4bnOOXnvSlkI4BWq4X18LU
JGjizkBwVHnEzNi0q8KPFztgZRKc4+Ypq4/DEIhEfNfHaqGfq1WczOdlpqY/6Mbzsj77e89MWPEs
qrcQXJX9Y+tZtY94ZHvIGsGhFBmHFixD8INb9fyUvlctNUlcZOQA6EhWuu6iOfht4vDfptUnzuZd
gpcoPt9x+0vvv2bN9zazpWshfWjsKSnAK1+WnbyhxA0KsVJSJln2TYEwOrZymBixSS9sC4z1H93A
I9GFOaoigfgDWgkj6PIyB7PYtQolDri3Tg4phBesWRKEKLds7vNuawGk+Q+pLqAeY/yeQegVvcEv
5KUfMVNNv33TNubWuq/K9vx1XM/CAP0nhw7QCIJAu/A15ov6IBV+JcVau4YbVGf2pBTBlxmp3OWN
4fBkdDNAfJ/jO155ltdg+O7R8BjHWoRCs9lEjifpxRIjrY6JZ0iO0bWNM5M8noJUQSHlBJPMH5aD
MG2pPBhy9GKhPcn3zM4AF7uSypizTEqCE3IkLSLHZ6q/YEgItXJefHenl5PK1TT05rkIfnU+1lUW
7qM3BVVDOQTkG2KARra3FcT1l3hLtgYEDW1by7Pr1MQjmz/pLNhTmcxkvJ6azSlxzUWwWNpcDhnf
1OKmAyKRJUteFCJnMSE3ZVl/7fh52xxGVm3xY4dtgn7VwmRRfHK2EXYcVf6dKdcdNR3ktrjfoNcu
t9Hh34i3ekZ5mSDH42NN7XPmgu2Mm9ruHDKMVXkgWd7P93HXFSQG1Bo14OsLu8A5MaH1/yRxXtid
HcNFTSsenpN6xdzoBaVX037TsVk3n+sbwh83opiLA511ROZr2eWqFZU3MTAyYjccVUqFiy2aGEBB
6BX5ffAq2IMYaOT3B7+I4cLDCNz4F9/pE4P9wot9HOyOua+RHgV4uC+S0Z7BTDKjcEqywPvpCsC8
Dh27uGqAZZsJ0eul9581ZS9j2RJCFVj3pt4877z8VblOXkkPt9iGEjnzEVZMw6NXxHYzibZ+rzMK
NDHvBACTNKWGsKL+MtEqNCKdXAQLhcw7z5v0PNrjS281SsJHNfqn7ASBsWctLQcsXtz/o3x1AYVc
KARWkGcRPTg3W9GndK+8bBV1YUanH0tsp0I7TRb9V2Vt5aQ3ETB2IEnyqoqWb8p+tEPX/iLT2C/i
0QD6F8czDTgmz+yPHIrvuf9mdOt3EGeEue7K/KGj+sWu0SD3cfD0dhF4NgQgbavmjITe3kWLuHJ/
jDK3EasHUv1XwKGW/CsEdgM2ZKT7HZlVMrvxAS6zpcjZIat2awp3dpQX1lOseatKPhSseMkZeQm/
xsYsuSE6aphJCmlwGBt330pejGdw5JgU/ZsxA1xgm+/+DhRX10+E7z/IeZ475ncTGPk/bT4Qtr9J
IA494Vi8X2rOsGvT90GIuSIczBhQrga3u5oZppZcBmvAF8SrjzgZneD+FV24kXN22YfEjQnpei6S
RBUA9NzpO2uZdN0v+bH0v1e7uJck/4LPkLYh6OMJnfE9KPXOMNti05ZSMtyF8gUvtn94pcpfH2jw
07TkdRSpBQDH3GQLhhpB6CTeyjgO7RFh/Mb6MC5x6Htpa83JVPAAeY8OrlMvkEg3ieMB4WLmx9bi
1FRLBzhuXwD+JeZWH5d2eqr07bjNPIVoJxW7naX4GBS141o9WYOb4D+kNrq1A6R49HD72ehOtjTX
vilG9kicDtTsdNhj1PrrFXU2UGFDxUjpYKB9vtcljCVOHPKlXSnmxGIEPOBpX5l+payNacDWeDys
4PecGKRxlEC5V32+6dBNhheFc4IVevf1IJhhioOse0brGM7wylRc9pZS63aGaplIZknak+JUarXo
rMYwb1msLh0PI6BGSg9ukMcusQFZ2BE+sfOGRh9WWjLrnvuj5+FNGE3a71OAZpnPrRCceXOGz3Nd
4ApusKQBnBBk80my4yPiV2aoENeEJZfD7Wa4lTyWpNf1cZLGcgiPFE0IJvPkCFl2hpoWOU2ob5+4
LTtELVP3i6GZrcILgxNCn9oFijFUNyWaXs3ib1bSNDQIXSHhhTUcUibRb1hhZlLEbPvb9C1+DpiH
KEq10g1bYZlfjGYTSM6g6UDcnJCkT+WM7rywa8bXLk/qnsqgIavwowzkk2dWac5y12ADsxK1dVbI
xVUi85z/0xlyiP7y7arL5O2eyLKtACL9i0Mv2gcJS2UKSAKxSiI6oEXfYadDASRQQtD1CJN5HR1L
BwGzj1ikxmyS57v0Tz7DOcf4PF9QX3jP8uQTpoqD3fv6fL8IRHed3cFljzSnUirK3GlBfUAczI6p
6pW80RenMIc/hGzmds5tDOHHOYhguTedbCNAJaqRZM1qeQkTRCa2nQhzzUfx6itN/G/OuwFfxkgr
vSw1LXVbfobjoRJ2ZW94+xYoG65a0RwoWDWoLUAGeaIndK0LABE+yrbdCmy9x/lv0JiFbYeb8xXp
w+0A8P+4ny6ggdmHG/xlb6EXOJEIfD2YYxCg3B11SIeHAGuDyjwaBRt+VmflIm8UcfI2MJae4FM7
h0B7tp057QniadU7eWx06L0/915RUb2ljHLJ95pzrlEEYR2blRfdvKs4hCUW2b4bVNhVGkStDnjF
On4Mhuz2PWtJyAAhW4DoyMLFHEMfqND05Mc9r6dwWGMmpupP5M4RibU/U7xRRafgoTLRwCwp4n4k
dsdQnWAXJZPdH6vxHllbK47J/CkbY1IidBb5cUPaLZIx8pYZtxH+0c11Fp6677DARzfZfanLznHE
LovM/ZvnCcT4kT1xlTstI/u4KZ8vQ5z0wDVDMAf/YDDKnee0pUgyrgFvEmyW6OmnRtAiEtU2TvDl
DqBUh3voBWEWb7+EGEaplB8O2lYhIMutnxjEXjp+Kodrkvp8flPj6lZv3ZM2EpVDM6v/Sg/ySAwu
dZZ25OhLLwUa9V6YfF6i6t34JSiv4Yzq2iB795UkLXxw7wbvKP8ajLhH0UzFOTAgU+MGO7E4Qc2A
x8O3da1kin1Ve9t8LP+TGk5oiidUNSheHlHXokGBqr7gs+1Jl3Y2WhI6roZDddseIXV3Ay6M7NYE
fyYdy7NwAh2+nNIlwpjLMWzVGwWHvqUUhfkhzaI5Z27TaBvi4CzHWAQZlUG5YsBxg0PSuUX+//Tt
vxgZQla1rsK60fJpCGyFCJrRXyWUGt3RwIscDM+DFKwkdsQntsHpKdWDPYoxv4SgBbyvxFigqEDQ
/7v21LoruOAAceIC1HcJt57pBVv2fIvQoDS+8StCK7WPZUIWK8NtP9LdLQvgAa+f5+/groMQyynz
2UInjZ12OKPvjpmj5tZz1Ly5TPaqZR/3n4k2zaEVywlShmW6UZ/gEa3NeMV0xnORzb+haQbAatI/
fxA9E+Ck8AQnNurDsHXf+fV47zzHDzOah1Qa3ZTdKUEtJxdpw9O7FgkqeqBP0iOE+Ct0lKYDt/cF
ZfYWPMdblhW4v66+AmlSLHVinhvo30/DIj4MP5MzGgZ27EERSBFGZKwOgQnuwIBM8zJMqzSok7zb
cqlHOOInvUfcq8U33yw93X382SNDgcQw+QKGHS54GoFzBP0oe8umuNLqUWoLM/uE9sY24JUtejLh
T5quvXfdR19iC7aleaywvJzH60/UUm43UiKATd1au4EZLBeB45QS30k219z9d6aucgv4DkquiEuL
WPxLqLytj4lZPUfVZ9PBjelMbCnjJZ+SpNHr59cnaB3Q3weK/7VEai/sRxGL6AeE+L97nQemUi6i
3KCqxSowlTO308bRbP1akwGYzbtUs8eYxoj16IGeT9io2KISHLNQHo/LNZEtveNALMYGKYlT4JEH
+w8yWOHFaSuXmOSV8j0nweEJLxGe8W69AevaEl8B3E7RVKvlUUG0HNML4MlNsLF+yl4gzDhMOBSA
BrUoB4T2Alk+yFgBsJ8ZltXFxauKtRs2RzkplFJYeKwnY7yXe8WepA9Zt2C1IS1jG61j1a7Ipvc4
hyU7ZtWzKUHvUzUrddJMReqmw9bBOhsyZuy7x+ZoTqAEjexC1D3Oggi1p9826TB84TgP/EoqzTh7
dAHkwEy9CopP73Op3CsjrI7jmHDtYvRsxtztMhRC/uaq9cBJ7/eSpj+5T3kCdXAT8UW30ouAZxFm
RJF3/4NmQBm7olfT8ICjGDlgQFv07fyhEbFrBkF26qNQtFWujhMYtCkO2HYq21VkLmriOFmwULeG
w1MxlGL5KrS9+iG6iQsqe1ZDXSuz9YoZGiLlmPrZUFVOnQcUoFZwjKWVk1sKngr+oxbMpawS1gLV
OFO4sOcSb4S6BXDnCyFIEdN5Z4U98l7NT3iWeUgU3CBCczdYQ0/dSR+p6qDgJDOFQGbrOwCnu2hO
t+5L+7OxeuKzIyZJk6/NBMl7ps0VEp55LnmQSv+byoauOJDANXGRIHeuYP/3BIqg3P0PnfplBlg/
/b2oJM2I7kjiz8FYhi8UFkOieHab5cdTEobF/KXHyETWgGaj5jICViRtCspKxNCgYr/3puG+emzH
6wQNCpyzwV8a5b4KXhvpMIIz6Hi4UZlcHqbOVB1sDkQLvOqTO4MEZu/XSJ8RvXvJPtAa43AYbMUi
yssGRTMM0GBOUcxASvQF36cEgg2g4yclsyOPrf0xLtH2mYY/pG1JTFiToFIX9Gh8fBoEhf2h4kb5
ZjIp3Bm9GZK5IyolBuXcP5175itXsSx9p0v8/mB+qpSgGzrcwf1WPAblzVhnuczBN8YHlYbERGCk
zBEL423Vkery7onsFndElHU8IeNGw5nCDc+H80tkDWDIJvyneYmFoMBbzkycJdSPVv/kz7R0P41S
hIY9bBtltl5Nl1e6kobbnWPkJbVXhRYgH4ypLCEMYz1qNuVXuI0oJtOtsHI1Ihc3oRci7bF8GQhb
tNypfKI8hhuAS/PI3vHPqDqxN0tqNgm737g0oImQ72VIImYt1ZNuZ7r+kxLXDF36NfHRG862pdZK
YJAHmeiwXyG/6z1T71hRP5m/duaBus+v6nLtRCdwe6440SWUW142i9t1L2+NMx8HRi1fN8Fay8WK
K8jfwTQ2pnCESFRygcgo3LaIIHEKsjscL7r/UhnaJdaSaKj75SHMXkSb6vFi3tEw7VBIXiAjJ7G/
29VwXr9VtptX/3+swcpbNQRhVjQ3aYXq7SpbXAti7Q9EXMDnpE/VuzN/mqs0UFX1b4yZdWNUfLbr
SIhFrl+tXg7fOODpTphb7Lci7V9DAYXdQdkEKwExvEIIIxo0s8yayDnnffHoQBESZsR8RTfn/euP
UleQ7HMt0QeGTVG5LvBCKgyk4wGJs0tIlOXOVab6PEPE0l1IJu1tRgrP7o53cE6GQwFVVe7i1sdZ
5haAUrZosiBoksMLCi/D42ubhvD4yU5ezTYT/FXtraIFxPKIP9kYcb0amxrki3fYIGIPX6GhH2Eq
eL7eCCJXZuh3xvfqaUCJxXd/+QBWyo2BBLotVERPH22KEF+/hZQkftgPNJxUYvBxu2YstIw3qE36
XW7HhENzym4whD+M35ggPllLTK9/IkFiw5WwF4SH8XorOLaHUGYMMOUCA90HeRPQxPUGi/wU+emY
Zva8OXlYN7tShOv2caTSJ/9P017DWQGVf01aVhoSAeC1oZhnrhSJIDwk8R7vdcPdp9+bRnp4KHrc
XwKHM7JM96n1ePQe9givK07yOgpeGnPtTwh2kJbxrN9yvCPL3ieKPgxU1q0T5kQ0CS1B+HUy3/uD
f31+f0v68c7eb4O0Ib3HzZyg3Zcc7MZ7E99a0t7ZCOoZl5NczCI01sA3lqj+wltTy9lvJEQFRtSx
yN57yggpLfPrGjNHzF3fPnJeur5FRq7fKmNe2BrrMQW8pDEQdCFIPaXzVbSVxaBNctio20+9HEEI
AgCPvHjA00pqEtAPhkgDFz+Tb4KwzQFGDMnTW/aKYUc7Qorn0BaypuGRGdTjCw1u9oYNdr3SKEmg
yvVlyPfI0bg4lprBmBf56c/LZlRJhuFayBx+JYjKWP7hxLsPoisG+/41Z9zTN9uTcnU11M109Doq
XGYWE6apIoNk/SkzcY8vy7NvdDXbApEiAHC1mPXuhP7bTIdZ6KtYHbUFADNubsV2xwoN58Nv3QNa
+j7UPz0AmVEYBsPwA49Mw64h9gCT93MWcIfg4QGS4LdxaE+qGTxR7G0n/OU90p70U8kD3nwiTmlq
6d4fLI+3S1gF6O6U6vohZmPu/v+efaRTaOrCfjDAmRSmra9dVGQVIeLjHSqIIPi63mDRw5fcNn1M
tinRoiITs9AU72xkgcOwX3n6TPC0H5bf/evhuBh8IS2wQp7m4rMHOMXdgKeWoJaK5GiFQTb65BES
IjjrMcCydb2RJU44NtvG2RI+ySVZ5IEoEhaQYoO9yVTxQ0Z26i+u0zDQqiIxqDUHZAZ3co2+acPu
H7UUYHxW1ioUHWAUZw4uzXhjNvnMN0QY2dBP2Ksj/FtDKHQJhTLUyP1j2wx/lysBjlsAjLdpN8UH
vy2g1173tjAd8iudx29foI5fSvKURf9AshWtANkT/+dpD5tHxBNKnsojMwaVPKxGEkLbmNd7VCOS
Y6WKRxlrS8/10faeeCH4k4980lWY72bQIOqRZ88ojkP+SY3HJKcgcPhfStbE9SwnMBEKq8crRDV7
LDWhdi6CDyX1oam6aC6waW9VtKJzj2GEwyE3dbC9LOzsHJUFBdDFPZaYh7qvwncfkkljVRKr22P1
+lqbK3AS7eTF48MwIowSH4rMJoy/K73sFtQSeR8Ir5Q3UKbU/bGNnnZDMdeOz77yzFYlpmy04yfs
ceiga7ImpZz6r2phb02ov4x/EjNrvz7eVGy3rWHVvk/uHPIQ5nMkQg0nsRljnSgNDilMDr2FK44H
+TTEscgRFsRzRCe/usdSb5twPNrXNBI5T4D1NQcY3LEsBh6DFFoiCj+13DJcWNQsWrGMUqxEhjnO
WrZxQELXFKxyOsXoPa421Q72dpmNjz6pNLOYfIifALX4rH+7ptau/9DbLQQ075wKoPausXVeW2o0
hcO406mJ9Sa3AJuliLQt1AMQSbaJ4TwelTJNHj364Fy5Cbe277gq9oCEChXi/ZGZSZJYXHCaIbRy
yqYiXl5jPEFJgKSfXHcrp+Ocg4FVOsmNyLUR2HMHeNM3NyvrV7Y22bbNgRByggpMrb8V64+Sz1t/
X8xILSxHFUHgP0OtaBt3mzpqLR6qzfOOh/zPYRb3ZRGZdy1kS8zZQrXjrOTVQM2hXru9eJIn+w6M
CPddr0INZ2ze7diEvPmKosGgbanjDHfbuGlfPIT2TcJRxwqXY2oYQJ5TmEeGpzY3VsSekobiZvM/
ekpmt9UlVy31exKVJTRiCgA2C6eekCOnWQ4DiMCQ7S7WhBXqzcbzNaJQKnw2bHUz+T6Wc8EwLPtt
bcqFZ7OMdBaxH0EIFh/zgNGNCMsaCqEJCWrDbxsTmeiJAaxVavSRLID6LMBKy+iPDYxa0/VGef/N
C7cfwJr8DS3eJOq1kZvSYK/CvjiioH4mN+PrYbs108KcPhEWciVsonWYet6OGRIS0kqnrF2pY6T6
yyxQPHB68r5D90XsdarmzEu/rOMiO6rHeiPlV36cyKcSUvQv4gM5uOf8OzOuTA+DCTcTaAxUk8ct
LtoDUDqZpbRWlACQDKzG75NXnDZigCMA9oTD2SzLBmIwoTBUTFi7Ei9Rw3hgbcyEPKXwJiTuT1Sx
Zc6sPBny3b1eIDS7b3HzpDb2E3P6aTZ4QP+XIRU+fIjxAnvHmsQ91Ft0qvDg0OFYkAZg329Mo0+N
BlwS5kK1rQRzD3LZd2rGNrPFUKnH/cLDX/ZvRoU6hW70jr/a+oWEpSxzi/v9dgkeHtn/sDVCUjLF
dqbrnmJDKG2xirm+higEQzomgBynfgyNl3wgcrR1amJODr0hozu8XFeCLq4AJM4XIvOyHLhOl+Pv
yejPk3CVowWBSJmSidojba9+mgCjUj5YKwl97X24YCVgybCV8a5ENWv6Hh0oyUs+TN9I9kUOm4I8
N+shU7dPsfeL/Dt2ddDmLw1qVr6B/0XStxT79Ojs7XePyE/zu7CA4Pa0YGz0CUPCC2U/BI7MyIBS
Z5e+2j8Yk9ZveMQi4rQBLMLb2A3OoInzESFyhvZ8jJINjGIicxDosPA0RDmU9XAeVw8fJcHa96e0
K6+acACsGEa41TZLQ09dHUooCbOhoTZLNv2Pgunoh5qlAA1L1YCgZwjTjt3uehORmJn69YmdBlYz
JOxB6yvoo/mi8zgGpDjgc2p2QCFDK8Mq7JF82AiSuixmwK5fg1W8+fTdspdNLhxIUtSh6IF0C+1J
/o0hkzz68Ldx0VLWVt1WqMc5AiWUTM6RDbu00louhkNeGDBu/VjYeaXhmMFpqrGruwoQQ7t8HHQj
s0IrC/V3ek2+XEmSbGL+qTCKJatsCPNFpmCyzOWMYPCRXLby1ZjIJDAr9ZDOxm3+mpaCbeks6fub
hf/SzxA3cBzYg6BvD6xrbtk3CHb/WwQ4fcDfKVGV+O1RLA4Ma6PAL4dweWaZYD/Iz8tQaSpHmqiL
hSADXuUMSsSTuUybvE6rw39E0y/xymW8ewXWjO8Lo8uBdzakFsrmlvZgWz3lJEMUyd4L/KU75jow
L9aPSjDBt/TZqmzxRn+1P4ms9gc4Q8Cj3DrZEDepMU9VKRlMBXn5Ab9uw6Psx9vEleLep14ZEOsY
SUSk08Hs9EchtOtFHPwgqfb7435EP3eugai/mkEE91L/m2LScfQXlqLMhx5IEg/SWkOaF8TqGVc3
TlmwKMdnR4JPY2hGOEj+SeiycvrUFvnxgqXHy4psO8oZsKuLK/FmodtV88PbJqDF6S9eb3x+J5Zy
FKZzj/oT9NAG06DrRu/ruw20S8z7DHjS7+IGuoZBMFfS6L8kX+uQot+XvvgCPkWUifKtNkstu+Eb
0dgbXlfVe2bSDin5zTyd3kBRIDPuGJ2KahwN5G0TCFeNxIcZDcWsinyFl9h6JiQO71f82ZdtL8DV
vuGauB3rE69z+o+6MAXSROBCU3g0WX2LcAD6zkUkxu1lf4gVdXFMX9PTy/4bPyqVeoQxWVoC4JJe
LNWAXtOQJjXWX1em6X7LrEAOukz/yb4ykPsEPlWbdvuwPDcHREKJ83ea812gSVlXgoK0SMawhFbQ
ZbNOF7Wy4923CGbOk+0e7w9YWlyTPxPV44E9oKnEg2OJoL85QNY0DSNlZ2Xpc1g+KYALV5NvuM8E
tb+D4tlEIKSu826nWDYtIG9RDJSGObPh9WUWnxbD795gFMhJTYxr6LXX8SpR5v58/MVdLiUqO8xz
kfcfAzoALxsckKGLLd0XzZqEhf7olUJgr/2p0pxZtW2rJ1bKAJTXbaBF1yoSrvjTecrNFrqR22vS
KHlnzHR2kNfZNFy9Qq0eQidvN+oLe+iEPQeFF8O/7Pp3D6gVBOUFFh1rpyK3BuJylPzPYh9RAwMu
pgd2POzCWiRTdiP6ufblcwOVVwEtYCJfjow5uHceqWAD1Uife2EmWe7p3a79/rPpBs+TQoFqt6+w
lmhsuJbcZAAj2ELTi204Dq7ZfVBhcHntsN8NRfdgXc8Ifv3IEXmLNCz3N5KyryLk20/Bej0EaVON
J95zTOQTr09Yfm+TPu7YR4DwLkqnKlLHEEXdZJZWDBXNPZFOqev2roaB80wgQa/55AJf7vAqQMRf
bJJXjI82fb93/IvAirW3TZHZYjFT5EllfLsLyxB/TA997i7KSQl4xyK0y7CLKJrs9t6QX1gFvG1b
j23zWx5LUNdsYXx6KlB7pBQAAQ4ME4Hs9K1ygR0sUJnIqiY4J5EtJiVRAONNZLBfWKsNQ61TB9Zr
wHQdQ5m5VOUGGgyGLh9ch2kl5N+XsYnZY8ZAQyKhUq1+kQN9Jhgu7KdWouSjmPPr49piOMeyqZF5
IwKUbAGrhonQeOFQ7Fn4cj8YzaxqtOQEFcG+Ae4nGfQC6a84Jw1RNzIjFhrAQdcZruO+VF732qeq
tYADwCI/fBxrHp0HBV/igtIJgBe/86SCHiZ/t4BXgOKw4kduYcydbkce8kGek4cRJGlsnNX932bB
V/rjZ4hFlYjbdNF+iI3KXPz6gndsxA7E65J6PwEp8JAQ2Ex8vMHywXvfJj5InaTZ6qb9IDV68ltk
VtgzR/BXZOzwo1a4XpJh23nzJMoEvmxzlKlEJcCR0cAFtQ2TX4JGTvyswmVlEI6vUMTWbL64ep0j
dxCpXBy2P27W3VBoIAr4qUcT0kU/jmKgkLvLgsWcLZxICGAmDTO8Dg0RPGGw6N7v1VZXldXCOXI0
k4Mop5J4wzouByaQD87TD6FgDnVZO2OwlHTNICRP6B5tQkw5wx2bglzc+WThj3sioLZ4mflDadDd
IetTbajQTxU08Hu9C1/3zSEzU8qXWYSdqGg8tkLJteR5aGoaJ7Dmyz0nFS4apqVYW36T7Pza1ugP
OkmpwdMuLEZ6A8N+E4M66HP6Mb3UcrqgblTla3dAcL7u7GZ6wonoEz4FXNO/8w32ZMm8IjYpKsp8
bkK/MxkX6wZx25nzKpALC3kKDnA9htWwHwUpEsbBAU9BFG3dJMfrqeBQEo+pxUgyFDWFhGUqvLiW
qLbCVB/wXVtv68YCDDz7Sz030nlBRoMKQ9UPC3vwivVPqwDHR++4+FQ8kPNNPxmN8V7PZMSGz8+K
NMZx+E8ks7Ci/GoO4Roo7BYGXwxXdJWjqlzI5nrw8qwGqeo56XbFJOrRnEmOJ+7Avc2SDNOI0+P3
EVJ8MNnvJ1LsQK82HsU+lZLnGtR2igaPERoHg25g2wZ/6lEo2+5HCY4E9lS7Kz1Ad4tXo4v/eYGZ
3/DEA5ZuC5bRPrZbIkOpztbzEEgNCLLndclsKcUJ2KM4Y1JdNoZ9OA8xYJltTPwn3Ap6Nhy9SosE
lcid4SDN40BuX6+F7020D3YInzrmoj2QMVn9h8j6gwHf3bnTYJYP9BEl92J/gA5n4GnoXmbw0MNC
u7fUfMiBNhE2AH6hssr6rHLuy0EuMlwCjoV18jkDWO6PQFz6QrP7ubrYUeK7q0gHLqWrFzExWXue
Dz5zkWly+ZVJEsAfrwxCxy1se33mzd15PUCdz0C7U8Pov2aE6SxerCFTHpNVpOSrZ5Oup6355CYG
Mvetp+QDfJ4KdDGzoYX4ujmXMpFbPj7IVex6rHIS5YRZxz/gTLE+pxN97S4UrakPpG66GDMuavg/
reug2jGS/MpEk/TPcs2ymkeCjB5JtfIrbAjD8phyz/PRRa3qgJHK/iYwORon3SsPLpLup6oTnTPv
vO1qeOFuXhvZDKriuhxt8p1vnO3UdZvuwWHEOEj2Rex7hd+XwRj4yaFMLgUTHhnyjX0UQa70nDZ0
gu1RmC/NMaqKbgf8NUqbGbdCbS1IX8/72yfd/5WyRHULHdjB/Na70iy6g5DCzmNfTW9raJ6VZY+V
p3vlWqRlmqiUKdHouzJLlDqS1rIyEn30KBJjRYVSNBlSb7a1HN9jecA+0ZdSalioezlttLUtBscB
fbDaV9BjmAwYk1MFiBEWF7i7z9AOuG8O1NOgW9Wvv0q2B1hwzabujbQRh3eTxEbmlq7L77xkcUpr
/W+2R577CaYwirAWBOnt0B4q/5Q6Qye88SY6eCv6tUAPrBs8ElQ0MQfOJKvUxkDvvPrXulD1pdeJ
04zBPbW3CIg+730IpcMBwOzY8yJ/DdGSO6UwWYYFk50srrWqoSc4q1k/BFfUGhrJ5jh6Gi2AR8R8
ovSrEowulNGj8N6FBNEQmw2oxHi8HR+JL/EcX3nouLbaPL1YHWR1l0VeQUnPlP8HhpKu7zb+8XVK
ih4Pk4DDjt6j1+BIOJYxx7XVzWpTodgaHgCz3t6GSmF+Sy5eSVUu5We6QWxSLwnp+50rNSoPsDo8
u44+Nvnju80jOEtKmV4u5/wAIilw+5qSMHK+dL7nnNkDakNWwjFZgmg3x19YQxbSYncCSJGg8PoD
aVsjJms/fvYqc8PJwdM5dJi6xRRkhczKOD1doAIGXTc9OcnxkT05Wc9D77V90qn7lfvu3PgOOVC5
Wb+hafDTvca/tEs8gmdIFHHtQ03tYUYB3An3XWdtA+uzOxSEUwSZAazHUf715KmjaPQ20uMLJY63
/y5rgV8UxE8IIZcKuhxxNxog+tm2Mjz1wG6FvAEAZthNs/ePgkGuFXy+OvDTE/ulQFsOdtKssyVA
xRxy5f569/68iW42EZ4AJNHeF6GEBMvmlAgPK9M8Wdc4IyoHKG5G0V1C9LK3aONotOo3rvpDhY0R
dExwZe7Ktv9Uju6VYk9gyl6VNMAx4u73CvJ07c0Y6HwIe/HmDPpH1AgPMoOAKzGGGERpjwX6RlnJ
MKHyUZqsaEHVWYAZgewkqlspbBjvv04pwmLUauWYSYPKnBxxhXPemL/+PA7XbnSQ2xU8/Qt/0O9F
Yuc8jwYyXaPldlxrLabpe9FkXKqtQLQIISRq7K109P6/bkORkV2tnFzCGHMNoRaLMjV/Kdnyj1DC
ai9nbVX0ywzTK0MrgI8w1a95R2CcE5y9mCk59D21pvMMsZvSuv3nm784azhBqpNWzF8NWyZXFp7j
9TXDspTZZno5QH4JxxXhSq7t8PfRRd4AdW5k8qAZqImMuTqpECmQVZENTNoaDsvlPgtj0kgEGL1B
HOIHHM69jrO5V0rQdP0agqm4//0gQWXWGgAH5/zlWpVn8spLP9ouvQ30Qtfxmy3ye3MS6staWKlQ
BQWhZXk1YWkISpLOjSiXdS90QlZoHuUJV5V42iuGXK83ETzm+GOy1c1abGju4XnWFoqMpwFMnADx
2i/Ke9mKqLD9uJXKA+kZA55jZiDOC8sBbDO8BoHCoRsDG8SdwrCh/grDoJ/ddH6GY0jefZCcfAj8
ul4Inu1gt+P0ugaz7tQ3w33EB72/nwNZ7rTjb3JE+76/y93UdLybr1c6ymKaU2wLgrQIFEgcDZeJ
8dCT82uEh2TpLPv6n31+lnzV3/ze3lWZF2u3eZelon7YHqfpLlcwsOfIiyaunCnEBSPhdh5WUK5B
U4eWY7Yko9zUnXTph0NzbOiMcYOeNmRC+s02HipaZB0ViIABHkCrg3LLt2OegME08/3CQHiGTXqu
6m5AkJ5foDNWmbM07KUvDbi/69hT7XJZy/Z9cf17aFm5vyUNgl1/IG5HL0XGRJPQhBAJQIY62Tzj
Vip1T4/7UBIKt4OjFdIZ6RIB0XXgbNk8VzdzcC3sWurBV4kAOLlIQ3SpGscLTov0uZTqn2hQjAN7
geEku0anNzl8p2B4EwoRzkP1dR64Q6ED2qid4g8iDKMawZNjHPzFvorV6Go+wZAeVDED/E3gtt3m
LYHLvWZ6alqrspOEdpndNzh+kJ2fO+kpqrvS1+IxMCD6iinlsqGQgdxEa4wJkBg9KiQZ8rNYO9yR
NqksCmALSh79Uc6beIVpvKdf/ZEfEoQ+h1Wu22l5PjlUkOQERbWDWBQswfantKATFOzP10z8R5bI
G+nwcWPny24ujr/VASPjFHkX8MlPYKRmoPhOp20/ohUOKLkghiikq9ZwDXZsgfdNy9Hkn2miaa92
8gxBB1g5tM8muCp5b7tmclNlM6dec+qlkmPdOgMNpV1WvPGHuHg3KuB+Le9GUcufmUPgqW75UUj8
AQxwYZ1d3hVNUThQpd562JMkMZvGyenGmC2i4hUlBlJTeUpySpuWD1RV/239yceB9AeoYnH4MPkc
SKhz9yo8t+1F33vC7yr8L+QN+E6e/pHcmPdXKLww3tpSqwXr++B9FulKM6ii5Jh5A5O1G6zHq4XH
QCa0t2a1Tn18hIplAq/s1FQ6qVCAgztywBEV5iOWgjzaV6oP9v6tDcznzMagUmq0L9YVLxVIynHx
vnx3lfJmhocKila6X7jhhv+VIKKl1h6NlsIAPWIbhH8nXXCwNSJMrdRNnb8fAiIHWw7y78PgEl3b
HdY2g9s3/AgdeXwhLqN3SyD5kX/clkNicQ1aZ4SSpB5fnGgWAP5HynapfffhnH4sHfC0wVwlOSS7
K/MGjocgDc/cNnBK6LaeL14Y/3/A2k/8c4q2vu+EoTD0AdPRQBpKyCikNy/cjdb2A8kOerWhWvdQ
hwrP2cpMiryBYAtyq4WcrFdS8XCvC/DxrtSUUBqxImhoQnekKQbukmbbZ9oriKBDU3UZdOVO6RqS
FesHD+9Jw1y7xarcvSvellLWUe8sAvwcCiW47lunDiyAeEfqTvftyYMn4KdGCdiZyrv9NI71cP1h
7aqy3MZAahYCsKwSjBRlmBLGn2Lho6rDZFAb8K1xQ/sZ+gReXdi/hK+WSyWWTEQOHb98vfjcVMLt
gtmxg84Ln659svtEHOAd67GBChXVsFpCFIIs6FvwDhMJJ8iEaQxYtbiY3MKzR7ve+CD6InExIOon
tofQaUME8CXjcDytuPKxEAxbl2g4d3ZYbkNMu/ZyxfgC3mtiD7SUZemSi3OrQ6gncA7EMh1Hj6mE
+7WEltC81YWdi3m+IUoo9MbVJeBP7hWx2+wOcdRYp5cn4Xy0g3TcGvLlUXOBQnRX/TxT+skSOZcY
oPou6dELIS3ZocImjmX3tk9luR0uNMJZzztZuFZS5nmOW8vsle9tVeRHcgeoHsQSLyoHnQbTNHcm
m5jT1Z4iNuXcuMnP033pLKR3vB3Qf3LtkAtnJ1J2xufjGWqE2NZPJdddt3B8G29QnKsv/wElhLi8
7jpsiizWiG1cEAIR/v3Wv+pCXoiDkQVHKEBCJ8FnEkHtNzBlv7m81SLDpzt0vRcmPksgdgI+EV5x
LIYi+J0TScJyRjgNy5XSGaCuwjzCN7sv5CK8+bIWhWotsaLNCRdb4UhaAMIOUtIkum2Bi0dOv+ZX
AdOFL96N5ofs/vDF/uB/MvTt/Cj81T+l7ZFy60u65VxtlGhgvfLUijL0foqR5Uxz/SVHsPLfX1uV
lo4H1E+lqWhpNPUcgnrVz9KrH7eefuPiN9k7ImnJvJTPFmdtyZKR5kHr3mDBsXknHPrOd4+S5/om
yI98hPS7YcZIcdp+W14eGZqesu5Ec7k5wA5AFae96N3fZQMSOJmNlg4cZvIKQVySwC5tqMLrZghQ
PJ/wLGkOgT3Pk1LqRhKu4I9E3LuN/ntBV1otDKvmT7vGE78VftcG9Yhpxac7PlZX6JhiVHh70HYD
D0rLhXUbgsbfCOYpza7GPyDK+j8WCUTlyq/nRKtcN962zPeM0yuvD+2Z+jJxdnjYJGHsDwcq9WpS
rcEu9X0Mb6Ky8/hvz9HZ4EWyKhM/fjhMNO/qEmkLY+/7uwyJktQqffvGfdjM5zzZ06sTDEIT63UX
uAEUtTGEIlF9cl4psrC3Ax1UPvk7YSzApt7gjfOcgS0ZuFOO38jeClQNzJSAhUUWk4Slhzxny6AD
MJYuDfD20pv9IikqT2c/xdl3ew/BNLiTmz+dUeXGLv+bRQ3KOXQzsuA+ULQkk21FOSoEGrxhDaJ/
68JYJxg4Yg3n54Y8C2bqRIeWgGmAEeim5qQWVi4r3u5qS+FxVoPFR1lV8mO/V1ekEVUGkWy7Btrc
wJiDIQPuO2SmpqxWGi+SEEZaE7wTmAhxI7x09AJpbm70YkuWVU8n/YFtqcbBhgs+ZQjFAUKPt12E
WersKXSNxwOb+wpBIJuwV9jDqzHgq+BcfL1Ks12d/vSoVQ0xm9zRDOhERR2zdU/D4WOPAJAooIw4
snV0CjnAaB0x0lqisf6No9ipOYjqEEzabUnoudFrP28XqBkK3SsUwejdeJjcB2DX7J8/SrsJau1f
pp1+zR8BNPNEAntcKduMXx1PW6kF3vbLop49Xniyi9wKbE4YE5mJBedGbIjo2f18sfOU8qCC3VO8
vLP8G6YTOKtZFCOI7l9pyPZ3aFgqekPNXLBWC8NAaNS8/sv1YzjK/itQEOkP98mt/4zz/cFr+2Tj
nwDsNXpc5jPZwjv2u8xOrFhP7aG/7mhTcXRfNbvlkTjeNKNItQPF3TZdiT099ulB9clUslPy+Fbb
LlU3bmu72BD7XwI+/EeaDt2ggju+u2MniIcUZgXBmyd3mzfrAK5vALkG743RnndoA1E9/nqM63T+
8p2JSOOuLvXMYst8rc90qGbsycwCo/QE+f/J8JNUTV0IPj3fdojPlxrqXVRZPXlnOx+nV7Vmt0eo
zrRfnCsK9R1dxCBOXrUe+QN2z2uLdao5epS5ljQSLxCwYRVBOWk0lDDsAM7UzfI2ESuc7iA1L6dc
s21kY02KO/nAAVqP4O2Lmsjz+5AOI4o2r7zJWs54BAEyxjNx5X+vDUGs5wD6i+YzKzewEFfhe9x4
2FvshWUuoH2t17RjzSnbfIevTAuBSbrPgoL1yS6Ue1kBEbGqZlAGHNGAkaVSvJguFyS09vDre7qg
0Qx0L69I7dCXZmtI/wNqKG14mZGEqJm7wM8PSkfWcUUwExIBVgCnXoG7VUOWA6Wpe+z9lzalO+Wy
MWaJD/oPUal998CbqNAt2Uoe87M65F7ef1EnwPyu3vZcTCjojHJ8wmm0tKroqKAzmNoIwtDvGE5f
+DrlbxsZUB1kkudIOn0wzNWBLZc6uFx+lbwWFy+SJ+vqULEQTyZdO7+XdJ5sSjEHYGWjescd6FrO
WNGY1kMqG85DRGwYc0foeFf7T2kF6ReutnbsTklwQSGTALgBUstD+jdThxr0ujWi9K3XMBPWOAau
rsmdHES7dbZFqDkk8tFQRC1FGSxrkGdrMbfrdU8MzkxsTdnlkAvqNM6HrU94Jwbf0dgqxKRKzw7x
FDqs+IeavPY85Yb/KTH0/W33IvpT9SslfJ1ZBH5bND+EKGsfEA6IFevfGZU63Qz9qXfKJtOVjd+K
pR7y4ix+I0bSN7QCfqNmQrud6J8UgyS5idWelvB8XOx+aCyxwgVxG6fnaxyekUFCgZQM3W5QNttj
fSCcobEbiuwrHgG5eOJQAiqg7wPrrZRU/VnWIcIOKvowW/Blq2IPNYVj53yLsQqPGlXlO7B/g4O+
GU4v5wGm7FymeAlOGHBYNaTw+BD2A4sscG9QdoHfvHSW7KZKN75YNu4ULbVqIzDuzA/ITymFPiKg
5qziVSGeAN7oOrymLBWLhGM/ZcBkwyuxsHLIaXy9wBUcc4lwWSSaoLEyv0Koe8GmjfkyY8oMh4DO
H5KBlyOntN1KrTBb2rkLSkQHfkB6sAnsGZqb/uAeIY0XaoUAPxqWJdE4+RGg9tvcAGqA8I8PzCM5
vo/F7NtpNAXBmTdGPpDyssvmEUx2WuRFItBL8N7vvLg2yQF+TEacj481EYxSFji8KtwdfyuBJUAC
mLNtlDVRq8xX/UyRgT2yATvXtrezyqhJBfSeGXydhAF7D84XGyh21qJueKwzidRT2YvPirtpT+7U
L/y/u415fRyQBuXjo9y0v5v/Z06Zin+t4Uo1kZFuZblYaO8pYQlMworvmS8zT/potlPAQQ9UiNFa
pWIPfrVlWrPzr/W1B3hqtfQ5M2mqwhkwwcQfhksLLV6jcERD1VWWBUB8XLDpNy18IDSmpmb8a6tn
LAK2bUkVACioqjh8u5qY6j5cEBBp7FrE0BB0Gv6kaseBwACnvurEdxhL/xsB7VNlBKH7ZfyS99se
0AQX9ABbk04kDvJIOLZmS3n2IqF0R7KwzN0vkL1k64q3K1OLFTn/jgkuEFgcpfMAJ05Im7DhQhDN
LJf2EtslR4T7//cKJuhGiTuUbSBlDsqHXzy1FiFS3ni/Wzo0lLMxmCQ+26OQ8BhtQD7VfWiR/moH
C7k5yr5TrrNoRj0AzYUlnZAEO0PtEJ2BlzyTucilcITYFEOJb6puj2vbNQ2LGf2mxr4xYadaG1m3
GAj2s06GEKXueA3vA//j6MH+TrvXjgjk4ldAeV8gvYCrVl6bN0VsIAHohVy6xlKhvYrPtuSLKNxF
TSXCOgLqvHWvzxUZbh5Z6YxOJRLPN69OEfaKQheMPafoY9JJNcxQ+4WU6ehsQMN0I9z+9Qbvh0Lj
73r1vBayO8B+y9JlISng/RBifxs3+j5H9hCs1Sac7LN9Vwk24BlOgPu+q2Rq5m6fMGLwFGTXH9/I
PVAFy0cmFsAi7YgysvtOkBV5AYs+cvAhAfOdKQ85H9nAO7p6GYm1xepm+YQGOjyHBDmcEgoLpief
39RsULLkzAV6thUbxhIH/jl8FIGVUO6Oh4h4q28dZtU15QtLqP+nONZll1BavQuNy86i/6Dx3rQn
a97IOxO/Gx+tI0f1i0It0Vwsa4hN+D+IMEiD+YMqbgMyNnt2JpEJxqdoFZDmZzX4KxAOvQZX0TpO
8F7zwHfit+vvHeq9VmIkfG7VA/nwabOkLDbyewkiqgszyOeOkCs63D9zq/7tgznQAtzl3T5OE0mk
NQ+asw1gxn8uTYU5tK/p62WDZqDQEvsI+NBZzsPAZm5aoLmrRXsFZ879M6/KTrxJxVUTBOBcqCOi
/cX1aOPrXgxT+uz21uG+I3VvPHBuEGFY1pTrcyBbnAOrk/fcBRFb/Lwq4Hbg3K9n3LbyUKfSmtdB
KHjvMmp+VkJ+O1omPWzQp8sFynqHo+E4goqm/ReeFZutK7MqtT6NZ2xRvd7AQg5aL/86iy2c69Ik
5t++l57qNMus2bZchiqJ3r6OoQQpmDhxiSh3Q5Ni5h7V9MMpobNlYXXnw+48mxgbE/BCxm3yOQhi
dNyawb5Z35grvvxuhNVBKenVyRebWfUUcJFbY38kavjZiiGnOCjdLjAzSOgH0Ulv1lPa9kzOq1/b
BGgGRWIYSPSixqtyEqDXqmEma9cbt/4lqta3T2rkY0t7bmVXdhTYSi7Qu5iGhzCZJ80iy4Xkfdn8
MYcfhaZoAT3SkYjk3COrMk2JsbWMv10eT0hjb0fFHeIEr02sdYvMwPNVyUE2y304AsZHu8UVBfoW
lj06GrQs5qLHf7lOSHXmcMQLMMp9+9lmYkNGMqMvht/+ZG+oWcQjZP5nPXqYK2mtk9WVN6WnjqX0
vWBz9SVtjwOfUac7f1Z60an3F4CRrRJjn3imbt3o91LTU1Zq0wCpWWJC+THCYGAcNeeSnzLxRB2l
5tpVQRGAvyMgRXDKRAfLe60SsuSMyOeupQK1PuNUpyWxH/UuABTGkYfQq0q7zQR48uhbREWHn+2t
c4G68YzjELfXdYPKhIqC8UdhWqPnkonNeVaN4yoNH2heCJZnCzBD1Sp5qv4+++vF8ueNlpB79rB5
2Myjren1mXKyz5ys32nqzJHY7KCNWDV/7kznQbv0GITINCtDAZHnlz0TFL/UZ4U1qlZUUhKk5Kxu
mB1SmBx3bfAi6u43HJCbhjY3TG9VmE3GX2Zm7Rr74MilL0Lvcp1JXxvX0twu/25PwgoCDN0kUyPM
WkDfY0Yhqmayk4qR2bNptVN8gDjk+o9pHjHZzX2tvtOC+J+p12u/FPqKMSJ61WES1lbDPdEJpUr6
qu0J7ReflAs9flJESS8/xFJK3+83d3n7oLhlZUGPaPqqNczdxGljfPX2W6y9PTmVNBaUOwHf/3aV
L4PZjsLyJOrlYLkFJ5dKwf9lb0b6SEWDtvh8GJ+uVR3T4pxAoAz2DHxIWmoPxYDnazoeJSY9SV9G
1/zWjQqrQQ/qAaxtY0QYiH4ncjGgSQm9K0lj6g==
`protect end_protected

