

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XIV6+/PXm8FRNU72sonnILYjpxjtmIZbbVLNSWrsf17Y2ws1SDZw37iDqiHVxC1cBgNo/dObQumt
yWJq0muisw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZXPA9HFe7cAtyRoNz+yMSPw2Pyn+0pRPvi5XjdJyTktT81Si/ij5SgLi6R0lagxdDco2VlsuCFt4
OL0Tj4wvHy1Dp1ZlmyT/YK+4naDchHt6lXN2dYFjXydimftHAQxst9Mhv6lRib5QRDOa20ZQpskn
yks2LbBSk7XEzudIYJY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bg8I4RzLDMU1lDDWoHaHEhOZTFPFr4IVYc8PI75p6rwLWa+GCWy1qa8WABJB734VvQ5wpTCQEDJd
rxf1ecFNcNhvHhCyE2wu/BzY21WCLI1aRAqFQXE1qi1Z2wDjSCFHJSnGjrE1LDefRxcxG6Tq9XbG
It/MsawBNQzhK43GHNj1+k8zbaJGp860b374HkhV1ZfNQJjcX3XJZ1QrIoPuFXx4Jhi/vjSlVFXp
pw6iybj5y8cMBzzatmsSoxyLcoJGfbq6C8apYs6F5VefEZxehY+hYk0iaREI+yUEx1YOnm0lzVM9
0NDqetgtQD4GK5VbO0+mw0/9k6lrl7kHG88ctA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uEnR/Mi+1UEzM6gOG0vkJoA+Jn3kxV9bb8otdkKTuCLYdJMYTfeNAGMqrDN6fOncHFTG1XMkSv7C
TzB09OOLPZWwUC5RHySY8jhavl3U2T+KX683mdCktfKMasAgiszkXyARiIK48HqFwHJ6chQHZVFP
PHgr0ToY3Xkuv4qeSGPvpnKroN4SGD/mdjKnjoQHGMZuZK8qyq5742CAWbQu7VMown6q0X0UZPcu
1EmiqSozGNEg6NBdiKBwGO1I36DQN4XENNdX9KsMUX56OEaXF2SCnvpLoCayaA9H2EsYpnARgVrs
/vwfUY42CXp95G0sE/mbV+1ahx6recWmvPJSDg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NoPXYyMJfSM1kcGd9d2E0y9DsmmxrbygZhs9LH++zh9P1OAn6hS0Bk8t4Ndb86rV4ZNvh1uF6+XE
APAfkag1Joec7lZ031DktS+E+U7heIbtHrj0Z8txcCoU4pcni4l4NRM4qg2jau2rUeq4Ee2HKgWS
atNnstf4UDlnanJjkbw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EsC7yizglwjm/VQRLhk4w7OZ3mJkXIBqwvXZeGGoI2t8w43A9I+u12UGUeBgq/MHOJNvVYJy+E2x
CC0Muz6vedVRM+FhA7lG1BhtLDfdhf5tyuZ51k/7eDcVeO3IHHvF7XSPJrUQ3MWUinYFQ3+Gsygi
Y5R+qlsaaGcS2CMkG3/Eih5tpkgSHmLV0ktNrQA5e7TmEG0rhv9Zq1LfKnAJYbEHIFNcOJuSLtA5
plx+LBg8QKQ+k9ZVnTJfrTN8PCfGwKgQ5n3P4POrh1PP11JPRcM+bn8OQexcyQJqzY2NV7fLOQVq
cI+aLpHw8NbqgXQRENmxsQ2ZAaG1oapGd13YQw==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qGiQK3HCCFErao7nb8j52G5u1V/rXhGG+ecU5rXKOUf+5W7QurCsJoepMeRrQbXCDAHalCi6YEjP
SXPVc1914DtWdpuOJR9bEDnAtPisBxcDbhjyAaA5GzCo09H3cDy5rQzcsoGiGTT2ezg6Nk1pmUz2
fP/pXAS5iVEWqPpMvSBiURlCFQ87/ni9/RtdB0Uj6TCoM5tkOiWtvD+IVC6HJ7yXfevf56YqU0CE
qkKXwNZZsQ2OGwuT9rL7/cvtRSms1VFzrIDIdrlv4cDuAG5rFj/CLH97nZfGWwZ7B2Q4iiKHlcJt
wt4vxAZVcrklHBSJLO8VzMXOGbZnbCZmugsMLQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VSFFGi5I+8eqPTjkRlMIk7PN+dnGGbWsm1buYkudsXq7lN301VzY6tMFyneWG0aA/kEh6PynLm/2
wd6EFwFZ/CX6b8btvoZd5x51dtWrAg1xEwmnB+ttvr1gRv17BaIzDKRP3nrVwAbeIrguXrfzGUUK
s3UDXw/ik3avc7EUEHARenGpG1MkKjjnV5jUzueDFEIdC1NuYD802BHFg1YFB+51wqGLpBMwLm7h
CC/EmDTGGZYUJAHMTXNrXI7Ji4rxad7i1Rz+hGhk3whN8mhDdU762+MaCF90usEeFK/PE4C7MhI0
3sjbqKNFCjO3MEcV8pp7cgyujSgEWcYVd+eWmw==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lkdsksTGPshZmOBDJc4avUeYc7TNjcff/db8BrH3sr7m5ZC4Y1oBlYsbaqVkMalTZKY9Z63UDWXZ
AfhEkvl4BS7BTXTkLmETGWV28hDtA9OrBk+Eim8hy5x/OQ3KnP3YUrkChGse4nMdIrbWLmb2d33O
1kr2UzGclw+nqYyjAYWpbpYRPzVjkUMp+TTxy9b73hnEPvTwoisEEXB3ubzMq1CGEsUcoQ9+5GmB
VaRWjX4pdAVuuCXQceCKOsWQW+4iI9n62RvZjTfnS8VkElcmAbPOhCFrpH0kt5KaEJodOswVExOa
cdByl8ewewezhdqPRoC8BU6bxXhdis0m1VS7qw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99648)
`protect data_block
lDqw83d4FFzk2Cnn16C2AOzwlSIpxr+19YT8/FTDo0LdgjNGyAjDRssn6dD9dEA99ZPN6Qastu84
cBhdJS4aWmU01OeUrPeUTPxp6UkJvKUL5Irhui+c0O9OO53hf76BGbDA/FwfVoLZTu0ZtVLl/vp6
KML4127Fdxui1vrMSHV4Ha2xxxo8ubS31GkMyU5DCK8oDgMdpzIaGGL1w8AcjCFVWpljxAFC2qgw
czotTp6pSha+XaDJWDWUEbH2Hei3SZHnjL+9BxaQ4JyJyj//g1L1RxiZyOdKDrznqxorYRXKTaD2
AMMsyvZZkIuFYj7LHfASbQFSpAgbLXdQWPmAGwlWI5L76TJzsqNQy4AmssLU8+JEoC+HW5dOozSP
77MA0fm6ot6BbeMNGqqTyTzECWd7D0nf44AFJWLAKDMQjlz3qCSbh5dxVge/ny/2XeuTIwpbyf8R
b16Nvf5jboCRaZx79hACihxVo5qIFuXlipMIzlIB7J98EoDwkLa+zeWPThiPiuMXnxFn3wP4f6A5
1mT3NpoZsE+b6+V7XqHhcaJYGDpl+zn+TVVwTSuoKhQOs2ltfXzwrtoXY37qtR+8DZsq1aN1COcr
iFtmWAN+Z9Il2zaOKUwxtFuuyOoT06eZT63I0A9/+Kc6tgDCm1XbPAsevMHK8GmyF5EocylH0WwK
sxm6DY6dq8Jd2nzo+UBlEAhMbTbahAkG17vh1qUbKLBXHLOvRmB0FYTXB0uzaZZSV2YroWtw32oh
aLLzCy9YqsIZxljrgc6omL4jYOQxd7TuxRGcLEIaCzCVE9+bfSl0D79NtK2AQczPTuQ5N7lnz7cW
NsXwXgyG7OLpLkqJ36loF5LPP44K7ZgUGkalOFaPCxdeXMVYaULWsrV/19meRNW/72o2vwt/jHgV
/FlLuLFShQ36bdpRNXbP3o99/3MuY9+JVfSc2Y5ppqR5IWHqxN/pUf1d5LsF26Y0FXQx6HqKvvLC
7gyD1A1sU5olOVSAKWPdl49fQUj712fznJ8pNwfBcyY0uc9PhXt/nWL0fcN8Ocqsy9Grx28KcBPA
ZskkHxBiWmzXz4QYe5ffgfVQHSocrAPDOxVSlCIuZhcKZ4xevTITGZAOeycLieBWKGLPjJnsgmvG
SntAghMd4eC0QOYTQEP14C8pUWarFcC/Cd+M54vVFmawpIVg3ASB0EWj/jtb9SwPRO6aW6DBXEUT
MTV7iQuFiu4wF93j85ILp8afK5sENeYi304XJ2fqpJRbPUuzAy0AtySFyovchRRpvLJ6vWw+3duB
a5/x3V4g65ojefziZT3eJyx00APcAHF5T41IYRweETzqcTeSIKtrDiDEf5Wk/Pcha5x5PlYKlISo
HRnD1CE9KJBLuuQCcgVjNQ5g/xfvFyldk75BmLB0AS5I8WIEjil1BO8pI7mTLvk/Eg1UU4Ldx4+c
mK6OAMwwYtx5RvPAXOYOXSpwfL3hHj4Y/1G2dFJ7tsOnn/1DjMlur7gjIFtKERbWWmYch915vSYv
/eCwsVsyam9LR89WMhSTUqy/m1G6nE5/bkOQd9Q82hzdhd8aDc9Mz5pX4V8o8h7LDpzOg+YEsDVL
E+cOeL/ZGPc9umqJoed8dXOrOvLDs5gYL8403Q8g7xYCXgV0JWaflbmOsqpjeG4S4cgT80Sifk/1
LkGElazt+SK88gGRZZmky2juz4cO5uBvnxCCFggSf8YnpEMEWTlpOR0VFRwF+Fps7DcZm6C9ru50
AOyLYi6jnpw0mL9NUaD1WggH1bB35iE5g1lr+O2xenQqMRq/ejOJoh4+/Id1WpiEKzJho1mL1RyA
t19yBhWY73IgCLBDjfP2sk9RmA9DBBqxo6uX0BgvPtITBn1SEDrsYSiCcpVCIzFPi2ru7qWSL6xd
IbGYoRCLOzEZMbdEEhprVaHtroFs5OO1SBBh1sEcjzXzRwOPQzJ+b9V0FH0OH/OxgHH0HGNMOTJy
NfsOGgImuAAGiGvdQRwCu/uUq+fuM9Nt8SW/tYjwMYqsjfJOIuuxnZyCMUZ7l77R6Vp15HByUZUm
Iwd8vf9E0mwo8Dw6NiJ/Eq5Vivu2uwvDS+xIouH6YUii87tDMQXyquxXPlSuMI6srNQwLtw7dClv
abvbPdPzdkxbtFzQPH5U4rDJJjjV7yNtpkOj0SNbxqvYuzYoT5Tfmv42EHhg+Uc6k6LgZKrmFlWY
US4h8c5UZOPLYlqbZdOF56e82lLSRqJfXZhSFUQMRF2KNwmoXX6rnGHjBpDmvQ5//zGUTkWTetFF
p6YopdPxr9dFlMZz/Lou3mGodD5aAXY6WRQzh5xx9gEpTqF2VdhBZnVu6hquHqXNi35hLQaDX8Ny
y5Tuezg2qolkSOBfavGt/xviFnqed5QgE1QSEdwXBzTKScxLtWQ36YjjqMx2rOM0dPfapf0JF2ar
/RP21YyCISBNo7Ujn8yjtl5SKTWa6W4bo8Z+9cL1c1X2jp1bUE5a0ugboush1x8iELoIKrZHxFCK
65E+rrloFaA5DtUy3i1bn2GDvxgVR1PsqqnucpYIJtl1UvYBoe3nPpPSVnRw1wJCo5r1JuUhbwB4
TsaFnn1M0RTF1RpVtQDO+GT7oK9o3puguuED6A1NIP38Zw6f+2plil5ZjjnE8yqMIUQV49wz2egT
r3gQDOR76g/w6BZcUhSvEpEkw6XPfKkc0XVqQIzr0ZcwBEUyj8Ixm19ufuPOsjywOg96QrBo/jTA
tiMuUs1QSp5tKdA666wKfryJjfknxqB3kQ8AIVqGf8Unu3joy4sBE9eX1sGFmNXutnJDVce+No1x
JNPAdVwZIhdBD2x3wo2QKPZw7RfSKNS/NNrIi1CVDzc94mAAo/4v+gfpTR0sLHCrhS1VHEhc7KAc
Q6M5rrTwa/Y5w6YvI1XKiyoi2SNTjLmNpHe+Fv2/BPOpsP08U/3LklunB8CXjKKgKGlpkciirG5o
RAAuUZlGIta9f7EF1gDxK7nMqFr33X4XoZ7nX7BMvhu4IMfEJ0ICer0Cvm3k/dYeEXQ3947X470Y
3z1zDnFMqg3SQg7uIcmt3s9tAxEuQsnKqzxAuGttVToRih32ZghmB5df1X9JDXqoD9YyB3l4OUkx
2a8c3VPhBdzv4oW0IEVe+o6BxqCe81AOfck/yvJk94NkhKt7HVeTlZP+CeRRVZxlp6aPmrjK/6ef
XWMaJrMqLDRS415683210GbrkxUeymca9/iMR9mvp9swoEOvQB/Q+8dmGPz+o15xfMIjPqITkkAI
67eDLERwqTJWOC6baIxlTkQk+j+Tp8LRpuBt2NcrCE20qAwvcWB3qdIe458gn0zGvgUk7IRaZhRX
uoPT6Xf6A9ImPrFZf4a8qggwLM71swnMIHvwbUf/aTrg0M0P64s4BIlwbuPXmgKDWJCHBYdh1yFn
sMpRRL7PDaTjGtyRxdcSO/qmCjCB3oTPp/ORdaYxJAphM8LOEZos+w/1ZdkrlmRQQLUbmtmnn9pp
ERUz0zDsYAviQzEjof8BU9+Q38kw2zI4u4Rj6YdXvQFIqC+PiQeEqGrNzd0FUBB3jkdf1wNdYSQa
n5W14WGTFlQmN57FTGZC/iV0CbcGhqxxryXly2r1j7JmwFb2HUBy9ANo0sCpTNGScYNJJKSWUQOs
r8q2T3LqVNz/sm412D4C3sG9UMHJP/uGbQw7YDOjf540EJfuZOYtYEEshMGAIdyORBu0IJmZihmI
Kfi5OPWdR7raOC/vnMXuC3rFSp/JQZ0PglSB1e11WpWtT8FbiTzLCLuciPZ1dCONRdHndFPGRs2d
MAzyf+1ucS8fzbOrAjDkNgyzdMrKLDvP7juBdM6PeI4m0Y9XE5W79LllR0WqehTLozfeGsFmaatr
2qrxmXvBeYB4AngeAfswd4uTUaxNdSW432AVvQ4OwQMhAe7agNMWLuSvlDHZ7LXE3K+zs+9vTKe3
65Z28cxkdALoHyEMZv6bpVM8KeaSz8XrcggOqhZEhvE6oOzJ4ZgHQxZFSPCR1FEURQ4PM/TvYJ87
eUxOp07JqxtM4SE2HSGsMl0CY0uurSYAt8NrhUYnLvWURCHpbRUcp7wbUpwp9p+NsGFoZEEvLBXa
XnJtYVHLgbiltCTmzVHbgD13WwqRbww1nniyUKv28uw/CaO/nfpM4QHc2pDqhHGJLwUToaouvaez
1iga2vxCzI304kk4/gZTMXa21RTPUxdpgFIMQj3WRM9M7PSMYTY/0FBlsq4GceZVy6CGxY0s3aIC
bVnCWM0Iq1lrHUnFV2QvpbHRejyRs01xyvNXTKGn2jDXOI6EDMw5tj+e7aZ7HciGeZVzr9levyIZ
52+w1qv0yHS3+jjWZAKCVophS+TMX+LJqRMg5ZC7YqU9KUELadiPOLjPc0oP/JH6kJhX9TgVxweJ
1/r/z7f2NTYmxHDMopC2Fyorh80ojakKbnItjXswDUlsXcOu/rCTMHSaR3K/CRzCt360MeOLunso
63VpNj/0iSk61olKLMgo1clrJ0m4W42I0UJx+QjKA1+cUvxptIUwx2Rg3HgiJ2N6GUCJa8HVo+x3
UcJuaxYEduID8MD4XmW9LiGUPXBup0StE+SJp9PEbNKVVOn4iSeMK2BOfZQzIB5mIG4+sVHqCDXi
T0EdCBDDVQFDEvA36XzxcYogEa6oh6f6cobkyTQEmGtvp0kYi+QOMFW2mWIV18v4N8UdCEQKW5vV
NfRJhbDjr4xdXonlefn/CNfBzHU3ZikKEbaLIMe1LQUBrPj2C1rzymQrB0Py2w7QNXVuaZbDGDaX
osJyx3jfIBajYwRhyYbbWkwdKHyPko9PelPe0BKuP5Q0Kgv/2QwdxJoeSjrlJS4Tkvcvkel7qRF9
PDP+bLUEdkcEWAZsjxE/3DIDpXfs8hxh8h2qXkO3lU3jIFB1NSxWJOG3v1eSlimKJRFen/Mkljpn
ZFIg8J5+8g8wfekNI5F0AtywUWG3H8THKhhci0qAIJj8EP7+fssz6rgfMj1Cut8S72ILldGhJ4CR
VelQWXTH/nrMAIv8t5Vh+BE/S4rOba5fgG4c0ymIoxc5b/vQeBEXzpNCAaR1LtfSmG5Ow/9aDzSq
l+14tg9PxKTEPntDE4c/aYX9qhVj2f2llYQztBQOpOOi6LK0KpSsYIib6jkyF9ovjeebvJGPvZUr
XmNmgbygKmSX2KHAa9JBF634mTqs5zbty/YlD9PCWz8tCaGjd4dijqb+6SNYBdIhCxoKlGbBJM5M
EdiOEjULlEt03mH3EM6m5q6o6uvKBYIljtTPwzp+LV8ckrtD55jwLk8sXdg0ITMT3bz6bzHIFA8d
lucdVIcPYdAnG2UUrWHK3iHsoT0evcJE8/yCs8tKns8zsDGYrid1JYT8PQGfnJMz5Pe9avR5ekIR
CyzyQbhxbbKX5mijCyJY3oLbys2gZshgydqjmnjpnRhcxcQo7wKIWyj3qhE3MrX8WKEfc1E34Yxi
u7sio1fr8Hu+3kJnWsyvJTtNtuaLVwePO16yeDLVKThppJTKXqJjCGQcvu0ghhYhCHR/hBpdDb7U
VA7IkU/MKVspXlSIfcPm++5SGpJ/qVIBoY5W+Xe8LeVwKrF0QbFgPJKiDxLqbx5ilJ8BK+fWk6/K
xuXqwQ+DlvPTDSwdlGaHvPrVt7tlT8U3HLmyLu8u/HpTyAMur01hyuhMzOUP6Jg8uIDV0JTsF+tQ
kOvThnyg23Y9fVRKN0LMRM6IvU+xk5ig0h0rRHiUiqsbpAhlzDDtT4vH+5BNG+/gudJGy1NSJO3d
B4NA7GR/utMKkKBJq5qUT+dIpDHO275/5la24dnoeUUqKKXZE8zGbn5l010W3xkyn34oNdIIk7j9
rb6UwPJBZmLMVsURBZRlH6AyQ/dyAWirIYnP0SGUcHsRYD3eswV0bYPMaPh7jsd3UxBSpze9Vo0t
wUo/nliPv7vUJAocSV6CPLNcy9QgG/QbzyVjppArdLzxHQz9HVFByYvRRaSfgqAZTOxJg+RcYVJb
XoWYOrYsL1GSl1JQeb/7fsfLlOdKCZIzEsJZTZsgOnfufR3eDRRStarHGZOi9mfk8wiMB3d7aNIC
tZhCPPO1++pl+1sQt/M55NID/cxMQZd+6tzkkLPGBnyfniK7TgiMcGUehLsnX0t/NiCyCcz7aE1f
pHs79XnXjie+nk5IIyRfvWPh3+U/aeRk+sej3HMXU9EEZYmekLFjE1gWev0yKg1XoilC6IjLxajl
0U5ccild7cFAWgMDzjAxQ+9vO+yA8OwjjbH5wq8n4KVw60w1mi2ByI5t0iBYVGvf9Hznk1suAPuc
tAf6In3+o0icSt1Zyf3cyP7fcRLRPwTErRE+o7/9z1AIxHkJGiiNx25Xk/KbXhPlLBFRkg31BL95
dEYBgG56B7r0X2SUuCYZwZbvTvh7PB+T8NCX9WZux2r241q2miHh7TUPpetSl/1ty9jXjzalMsBA
k6RyPhzUD8IX6DONBTfPuwx5FsKR6RmhxjjdNzJr6tu8pnCIt0wOoZbk7Wy5w9/HtlbuPYrTUuac
hS5XfdBgW6Uin1etCleZRaJ7RrazTpCd720fgul8dQojxGvtKDZ+0KKbpApij1SeFNjrHP0QhCIu
YBbHuib1UkLA8Yowu3pJC0OKuMMTvy9VReGDxxbbcYMkHh+8ijZenIweRmCA9A6J366BSOLc13bV
xyZ2rATE+8fbNhb//ryoSyzRE5MTJQ8hVaf7JTOTUbjopDqyC8vf5mPvxoj7nm9xtgT+TsyCq2vv
tCiFRA+s7WqVdP2xIlqxoriSrn2qRPH/QHIU0w9iue9GsLG1WZ63NHF25OIjGE8BRxUlw97dyXZV
ni+PEQxznjMc/dLa0/YM7TlNw/HJQriZSLCcTeemzdfl8InR4p/ieaP2yDbHiilxT/R4Yn80r/3P
q83PPE124d7Gzaqd1+wLA4g5XKYcSQ0uP3gXJwG0V0L9vThjTH1loDtteSyrxSu/P/55vaYk5fKx
+xe057qx4UNDnHmyJQYNP/fu8E/sw83osVDBKWQZE+p6aZYsoQ78lBlq1d5IKGCD9R7CpVoKWVni
RH4uEtPqD+izqOUYEyLEsJZ/LMS99Y0xsnHl8oeM9NbwyIF7BAvzI2q1j8KSH8T260x82Ii+kFWJ
9fAx+OaTeu7LbSVh9QSdG84uC8WdLvVnIxxyo1uQJG3vPtt7/xHx3kuvds9pV9kMgGktm4alq/e7
8dTIRL4uScQcQ6Xn4ywi0GwFR0w8iFQLbR22193SukuDcdKbn59oHo5V1jvxYgIycbGy55yQd7QQ
/Tbjj0OaKkSoudjZboxPcq6BIRHwCy9WrjbAeJ8VNElc1/eqtkPDX6DUepLAZ7Rj9t+Xy9Nu/SbI
4HseUuSRFBfd3zRr1bs1C1lYqpfVdkdgZ9393lSk8VcfJOiihKdtOLgdFRISTjeZOKCLeIj/bzag
hL2GSwlgKhla9E3dmqhtSjUd/ZFLYUYQf7TrHLlcWG2kOrEImMPavZ6oKwBb9ZvrnesGWbHu/FPS
L2aD8WaRIGtisjqftIVDR4for9YGsKHc/qEggQKMIUeVDPuu8okhV7KI5r8fgvoAuPAsMwT6UHwr
uiDApVF6j5Jmc/rXeR/gVGhlG5ZTSBv80dnXoqvOLE4xMvm+qTUOPV4lm4Kx0JX17VOnFO3hMG+j
IgUF6APiijxYT/Bkcg2lVS6b81u28e5dZVMJITrZozToelwgB7OpEse6xYEj3V1Xutpn1sGx4yey
bKar/TTzpMlCmtTKtWFNkcV1eQKs0XJsZMxfGbfY5L/zZCuJgK9nVVuJZQoe3mH9MQ14dVUW0Gtt
UTyKCZGNVyZi3rdi5ZXLdfZh2CzUjb/d9+DSb5dGaRArKtm0vFPPnCFVrT+2kTuao6kRMqPEMNUh
wHvj+1acWPq2efhEVWdzwPCG7dfQEBB2KXtJCZY7f8hsX5AEabGQj0RqyZu4NwwMpNthkAHAVLVM
uWt7jfJs198ltPoE3+x0K7Zs/Pkkq6a7WeF5OLhewCgrmhJkIVvUbePl1T5zPhEWvAJB6d0xOkNx
f4Tl0WAomkX13ztepB3QzdMdqQjJ+LHsinBGdPs6hvjCAnP4wEvjTj+ScObU/SLcY6Z+9RnEHnmR
f5xfE5FRubJMgE7nQDCoqpzDIkC69r1bmVt6BZHyNZY4wiPTh5GYLTMO5xGa5on5Tp8bXorNGGZN
2/Od8MVwYLjCb8bXExP2JSQMddaCrw8WNM6tX2sU7MpASOoUyxv4ZNolsWE3pv8F6ACGN7qp8mfx
gzsU9sURQ3Las9K94y3m6NIN33B50TxdCdj9BboX0/0irlk3Sl+CdUYIfB8pSvnTtcEIiEQwW38E
RJ5WJA7VJkBL9eCCf5bIVODBfuThnKzYplJ86kMheXttn/hR6hLnllGfg/6/Tg/ncsYUMX+8hRc2
OEiDuKA+J73OuM9L/rQezXyDG9OaPpg0v59gxaLrTXGMe4LwTwdNYt0vDRQiCMcgWcSzYy/lOSNR
WBTcw6j35lY3ZbEIJK5JyuBTLULNw57x+jpvhChTOLtybOimBEwZ0xCIXcgD0sWRFiKJgGOtEfoR
vFCVMCRnEwuv14miW/TScaLE3neKiITd22XMDGdqG2mrAdZBzAT/hHu/RlmPjjAoBh7FR47UiP6e
2sFdFW7L8RXQgjuH/GYlc+GWrt5j/FdExzwp0ECjnSvhsxGO9rfcarUSdY3ooFYb+Bhkx2i2JJga
7pelSSg2YJ1Qg6lV+gtTY0YMwq9gV3s1s1G+8gErMu4iY7oGHRLXHheqpoNYY4CahIaAZwzzVX18
ZVESsGG6Ltg7S9FapwDkIrwkM7gdX48Mk7QH9xZnVvH08gjrmCy8jNzvonV+2SkMkAT9RglMaVJe
qGRGz34xRrdhRjowYQubFiXJv3r9GlA8Nz7KRkY40CnNZxdJnLXhkMmGv6wrhvXiiqcAfbT7VY9d
ludpLzGTo5pucdzxpf4l/zLN62cBHIih5pBpv27biTFijTciRjRCF7qFnmTBcoZs22/E99oGriDO
OsC55gmapgXO9eQ7MUID18mqC41etFTioWRvM09mayDi6J/sSVvDavS8fftbGUPjWCJ2OBRTTo/b
c5Vz8z/Js3+bbqB5m7kgQvPFSiRGvmsEujeASUoV3cNUc/H47JXZR88HS/tC/EJ0iBC/XDPy9LWT
B2oUdDuMNlrSCSo/HaOkX9wOCriNBMi+25gLYiGRm5jbuSbc3H3OTM3r0LqmYOqEYEPbQtvrK6N/
xUbk1IBI7O4DM9vQF9nL6WjvigpuoTr9hj4QRHsefgt0AGRxWbsBUe7CkESAabOJDINzHsQPI51I
Ja4iFsYNSEafWLKJ2pJRV+WQFmBtnEOwgEpWKPG9Er5Srf+nv5CeTgeO/XjAmCbEm43gH8zJ7fM1
jqIritRXzOgvd1TH9BHpWoPiNhCOJEkVUdPl+TaxPOxCWmDqeb944A4w56CMjSMaCLPdyz/wJN0C
DnPY8UAydQhZq1bJR5ABuVw/gp6uqcj9nmAW8bupJp31Zleirr1C5qhAMoz/8sEBJmcC2rspHu5+
9ZNa/DeFiobIcBkg5rDA7l1GjskjQO+tZO/pYGKCWAmDDw7tVIGq7bKyyIdgCAR+nMStt2IT3LGG
/1OlydTNoX8/ZSIBfEfF4hrYo69DCiRmGNaY5/YF1lYA7zIRRrT7j3QfpEFL8XedBc/tzZz2hFFz
mUH8mmhaXKcofYcpCwwuCJacm0s3axbtuD/h0AD+smVa1mHrQQO8Zzc44vDzcpDBG9YdXLK/Z14t
JSUPReXhmTWFKvO/coklC6ygPtQstfGdQNI+GfG8+pwTQU2O/VzHUi5VVw8u6dTAUGTl8/fkB0wd
DkHE4DLvLkOeAlLDU3ahTNmnx7sjMZxn2FtocQAImj2UbIdCV1N2iBkGQXG0CHDNK9Rje73EPwMb
dbFdAH9yUNXNOn0LiXK9/Bao3wjLLfmP5r6Vxtsqlm3So9hd2WqRTMpRZ6XkoKMa4NTpkhTeG1mU
OvjylRTM8CuiBcpDLxOtYXJStcFE5W39h6/io+MJJUpA4k4dR7WSb5aQOexsN+0lcwvkV6tZntMr
2WsfIYsML4RwT1mDT1p9JGAAEh4ubuwc9Daa3ZuMkv7QmuYbbeVFsHpP65EeIwDlknio8r0rboqW
BQ1iWXuALWcU9yk6wOv4QdaG/e7x3c7K5SftGhg+Q9Z1LxoY7D667+SD3uA8mLiSjs3OH4eMm4aX
y8NMPGcA0X09vbNoUmf16orKLtiz2bx1FTBVErj6ygA3zRSm1RMReZmX5HGcPnD1+nqBo5sVN4NI
bQgw34aE23GZybwOwaU4/8JFOgKljSaG5K9iQmvRDyJRdBO1JdH3Z4MwwdVeyGj7NWmEiCSKULTM
rGhA1Ime2r+piQukxUxKkJTm5kGvZot+1YGXTQCEadnMcAbAvvNugF7e6c9RgrXxT/g823AFbYJw
pJXXeRewW9OkFCLkjGT9uHbnjXdKYR5e2peGTG17juxUjB4i9BJ6I79I3uoPQAIXAyFpSBtMHCBZ
xoyel60LSGeGY29/VGAIrqXuMRrpKZY9F2mXobSzhyYXzDtgLmeumqPI0aDDLe/SFLWlHhUVWaX2
DPg06MdEAczmfC+z4D3+OLIxl88jwB9+tb2PfPrDBm2n5bNSUmv/8k1mAwUtH+2lbx09FeJtTYwk
ABrtbcWH4L7kjvc0/MRp5hkPdUgII3o5pFn1L+Ov6Z3Xg6VRq99L9WLOl1MAkj0z2pz8TjoWObld
UwUXwgHJ/KvYzLv/HQRzTJO0HLa0ytXIaKhSyC70chwha60HzHUUdWuJYL8yKtKO+aqqiefXwn72
7t5byOF36Dag2ILop0RvPYEavWSkYBHItKNtlxRIjFF2P/vze9/meQHIyHxApjsdbPTb8cUiOyY2
CSpddDMoRka0j88+bgXKltz4+4wsByA/G+PCvh1zIyCmt2+W3clE2v+KewwxgZsbxkDLLfJV4Fv5
otDfJasZSuSihFbYt4YZkrwzg5KAXwpf9PGIKixC9O5UxqKVyM5kQlRSV+sYO6xsELIkaSO4uFv6
XFeGN+wF7BbuKzFe96qT1/pL2YQmyScTUIDNpiclSfvFDPjbGi+YjjFFa7d62ELICKvnYtrNVv9o
ZKQ+XoY2r8Qmfxs2vA4zXaG6tdKVIOgs/6lkgKxPR4MqMH0xpUyvi7UKXuXmapNVzsGATkv1sUHv
O7+q9x3kMIoqsrRYQrI3wYHfLM5t2NG9sYgBJQvu75MWPAW8LfwE9viLuw9spnHytenxuTvVFDVb
WoNLqChs0avP4Cs6X4jJTjw0k98peTVJOlg7D7xUoEfxRYSmt+u2FPjlPG0HbjNY/PGIob89jJR1
mujEK0f505+HKm9e5CKVjtKmTr5xLGnAPc2P+cD0rFg42VcUqXPmuTCwWUhYs2sGXXA6kcTz+xSc
6ehxFAD6nCsDNcxNJykO+VCloQjxC62VLCyw5rgolQWC6WuUK+DaT5t0EPkF7Rl9GcFaTDUwNPGP
N0n5M+3ijAlMubOw036+5ROiLMVrrDb5jqr867Dy3MHwCLdY/DNMFWA4gVI59nf03LpqR+mBWmYm
NKoRFVqdX7hEWss7+LpdJ8WqshnaicAhVCIc5MxWaNuzvkul0towm+yiLgYPXMJsOy1GxMEtgiTN
2iMNCTdfeVVp0iuIgXAEnoe4bZXP0qO6sAnVZBJq9cpdNbipvd5IOGw1ShKmk97Zym/iSZFKqIiA
z8myGFC1+13VUpDfW66JfKv9bSc9sLHfQKRsfVhouXx1mDBZ9sZTjl2M0IA7DRatSkL2vhFztyhN
PKTvdUZkH498v6aCylHAISTfzXKWQI5OEUxLFsII4uH8Kg2ySulbuF6loFMjOPffD+CUXvtD/JFL
AXC4RKrYB21igT76RjKcpa3exm+69WvhO9oBOTI+cSXpPo/MAombwvfUfRQmu6y+xa0OYKbDffdM
gNFUI0+lZedlALMrmh+G9WtrCSBirAOMsqK7M1wIPnllSgzlfKAAIeCNDlaero1A/ViT3G8K35zJ
dOkBAA+kVZMqSuSPDID/FbC+lI3HIwCg08fMGRqOfLbxrSnKiWIT8C2mj4emXOF3JZmNqqfYdCUD
+goXv56UWYYvnEloQv7ZXOOXfjhaZtS7o4n7zIar7UooqhBTE/AGD+GRySBcl0g698AIKhqopQtn
oQHjirb6q4cKPpr3cSJmN4n5rNytZaGjJDewGJjq/0Y005evVKjbffABLxZzVlqmdLERbE1k3Mqt
LQx3t0LO8gfxq+m01u6zDKJ5CspvrGdQYCCWgnV/+7xEN5SNg2Lwku6t3tO3CBDzIa7HXkrlU4t+
T4udHhUbZVpSF21WbHOZASddsdIlsszeDN+/7sAmA9gf1u4ondG7Z9ioSC5f4NTOpUQMZ87m4n/q
Zqsds+/SmfXkgGx3HKPbULS/wqmSmgakaOtJ/FJqKnhIFOAdBJ8QB/zd6ooBU2h96fZCRwv6XkCq
cnKxGWAuKmsrcH2/KsY71ZX+AOjDZGExoVm4trFffKuwHx4xqg0ZOhCcbgsu+MnESN/fQyXYovUV
pBsmOqDe0hI08/kHZwBlb8HvjZ63RdqYXjYygMNUeeAmAf95hjbMMq1Kx9HmLy0wqOZjrkVvfKuh
DAL7aY7TyIOC7RxLHK/kJ2gG/6y84EnELXHD0JV8BKSiuB1ugB37iUFiHL/vGP2FgRfLfGDGc3Py
wzH7NbIgCm9JODSdDa3YzxXxuznLe2ax5s4Pm0iev+DbJsuMkZaDbEg3luKn0YzO5rGt6zP9i5iz
ighd/e76NnhpeS+lZQH86TpzMn7ESoB3xGyWTP3EjZvxFWLE6tGQ/BL4iDl/dJCD0GaQl6XHDb0f
+i77FNz2uFOdbIy1eOkcE36wVdSZLNyYziKTgVmMD5LxhACsFDpw2HmKBtcQJr7OM1L9/EiP3fHb
vPD2Ggr/L3fPtI/ha0xM6fNhcKhUpIgOy9dstFkZuNcBdrLYEC9uZp+OW6b/er4XeLX0nKdFzQaL
9mOw8so7jdHm3LsIVyj245u3GOjbcjE8QLRjqvYcAfefyZcpf7/bXuVGFt/A0ibcwwzbLeEUUwmr
XxS7FdQMxojYsspU3aUQyO7nWcoShpysl2B250M17r+HzH3zkRrxwrbJh2e4VAnAYn5ud2Ls0gL0
BXuezl0oMaHjCzwOa7FuxhAroRqZUBSe1q1koMWiR1slBQgIqzIZlMYjOCrTkySMBanVtcNRmYo2
xk70j30vuVTljGAos9iYbjMgr4K+8UH5+42asdjIxPzfdL39lVSO9By/oYkel4jeuZiEgclupuUC
tPCkgDs8blp0UkenqFP6274xTR37Gj4ktcv0Ir2ZSam0O6qKhuNZDaUB+EW005yzPZHhRekwm9sy
ZhX7ZAPYqZk7Z7gN/3zSNz3TJUriV79LFoETa8MJn1IJi1wOQzq30oP2rQ8HdmVFC+3MlAtFPZWR
mWSRR9Lu+7ogghs+dNzRxjX0x8Mx/uOfEo4J39Zpp7uLh4CGv+h572riTleadXyIYTdwFmozsreJ
rC5FkBFVTDGE+60218IwpptJeXVnLRt0vDumWhpBPW+e1bKVo9l8WsFeoWJWDxgCCwmzQqGIOMY9
R7p6naFIXiAEtIfAHcKKFVkwCwGIWICVYq7eRSD5yJar2IrFoFOiQ638U1qghMRukNVkWatnxJA8
f99HcKB6G9UnVIc/GhqG9Fe5iex9+C8+79+7YJO+861onCQRneW8gQjS2oWHWvDUoLB/x1ghiPPJ
J6NEVOHgt/rhpW3wMpzQqEVUeIMx3fxXO3josM16ww0G4XLLrhFls2/1zLOEQvfHQ9FJJg+sejY/
s68TI7mrvL+wwh0Mxc9KvqrlQVqMy2iZHQhwSjIUKsZ+hJZhBAS74EBaTu2nnjhO5yrjTCCuV2ec
17pm3phDy1LJb0MSPws0uiUO4qPTP5r409vzgrhQQ5xu1gxE77DtfUxHI29z1cr02pMfKg+1/3I/
lTb6wrXkQrR0mAdYsfNHzmJWZEybHPsn/XTtkM2yK+FY1O0UD0lsqYdJt9vHu6L+VTaGaz+vkOlM
eqIvCa+7enG2VXRLm802q6XEmce8/fs+96EN8UQFg9anBGWFWCxUvhWCfRA1Ize1cMEWLykfwOKT
2akUTggsD4WgKwcRGE6KWRLuSndiQlCuYHsbrYFk42XGwROrcQfOdQiwfRhA4vzcm0SaBzsNdPOu
2hZgkdM1jHdIchYAT7m/1mfYuJ+dy6ordbwpRo1owlsUd02K76nfBwAe6tiny3Fkr+gbE88WH+dd
NOPHcZOiRTIk8C9JqbeNM9ZZQe73tHfqQIVURBO5YiwHcNyUGY8gJ02FhODZGQ8Otc1e2n9+URdN
MHPYIarZCbANNrayCsSPUPbZ0aurB9+r63uDRNMSwVvZ7ko0r2sfcB1VZDA0ibwq7K25GKFBVZAh
r60tXh7OHEfRrVBELHuqjwwoTmOtMte7ctPbQCyPr8RnMMl7OQImIEhJQ9j2NQjAdSCsK46xosev
fsUKHAlJMX00268J8GVykoNWx3zBKVOgjiAoB1uiw5v9kFFa2JWBUu9c78X4sGlh+LeqIAZdtSE/
HjHXdnxLjrSwhLZCXSF+bX7EjR8swFizU+gD7Y01jhiU9bdmKLGshM+iRjFWM9vlaXzsfmlLF/fu
SJWEWbhe99iSeDs1tSf0Ik69zE5QRVc2VUkP2crUagQUQwSuQ1zOhbv2IDJwYEWW3sAL6rPM87+Y
py/KioDA1YdxsrNGwVeowE6WPJLi2n7FTC7elzlrw9lyZvC1COyB4pkoeruoT/+xiZllAY0mg73o
SD51oDouw6Jk4KdxxCBcrPdwzDExHtqECDkqSK/XbHApFmTpNn2kWa6b9OfiFT8MWJaJWSh3pp/3
6HxZHkPg8sYkieAr1PlSr8vyNXN/RcAL/At6UNA6X9fpagFdYYmqL0/0pfXL6yBC73RFFDgMvkwU
rSdtNFHx2vVyd7Nc6jDLnI7ofcJsq6MD2JPT4784vNPlISnCk/iLDfLQB1WSVu/tOEfMOwp8O2ds
ss6NpSw+HqMsfz++2qQ78687cmW5P0KLuDU8/hmugQdzPxSbZ4LvUSTqRZiQqm4CurYjM49sNh2H
XP+CAZqSGAzpsyvmTJnJs35hg8vAcV92OSsSlXmQzSDSJg3IGcqKk8RGgHRlgf2aMtpBmrGuzNdR
ZIcYzb2I3+3ViDFzlDSImM5i5BH+zKCHG3eUde6xCvXq1az23JX7kRJ/ucTrWT9c8FPgbwJUj6nE
HOIFYhRKU3mMK27GBSRgRiAyqUTa0KVk4sX5nO76DOWahelfrLXk5E45bZ+pNmUjDD7GceYT/k0N
MqR91W27YuE4gEmNFpEjYEGvWAOWNDGJqBU3Q/zUMzLyxHejnuISHl48kYt/pcGtiCnoWmjx0Eqt
9XcC+IF6JI6Ogor1nP6fHu51f5oY3NsCSU6rW6Wyf3zZO3l2QZZ1zb4TjYckt6QsA1yJNIpnpBrA
6F6/GcSuPUDDMa92Nd8c7JRrSp6Zc/6nrIDWIH6aRDQDNrA/SouqbFeG4RMljimLR5rAub8f8Bcj
7TUafYV2xSpvdp6bSw2S/IMz8jnWwFbGHkmSVQR1CdSKeOqrOORHlOe55D3fPdywqMxIZmXcEGRs
r8sQcbG3lWC+iAjd7RrK4PW0iLAlcTqqT8GcbCbhS6WB877etk0twu5/3ofccwGNtYHn5sySBbba
ML6/OvtJ8bB1W3y9eM1rXXapBQ52ShkBdQcuITHtd6nFzxaLfbCV4vkz3g6Qj7vai+WBU4ln3nBV
+YVI/b+rEwm5jTwt2+PAZGJktQdPCbtfFv0cpbazTjAvHbeJ47IhBCj6qE5qX+OGZnIDZVDRahfJ
shvOMIrUrV7RpExLGV7zkuCY0GBjK6mcwjPstS/Ufoga6Jp+PRBTZpmFj3jlCpu4E18fxNfhUzyM
HDTlwbXdLEjBd7tvvLsbc7RQqLSkNJv0AblZtq5qqIIahGMxUZ1f4X2+VBwUCyfDOw7BPzA6FlQH
8h7LJSFFwGoSE3vZ9y3khV9aJzL3HkQ1OP/vIZZL4P3NQoEsKqrbJiMJcN7ZIhV9aVZ71BxJoh3W
779Pg0qdho4stxQn/Yp7R40QFtJBw8HDjnOjzTHnuTNYqYZ0kXGYFv59euG7zLwe/5avw5CIqUHa
PCKw95rpKBSkNxx3jDcv3dzqZJfJqAU0T2gZQGfHHCY3bVmKqqOvfhsHVo74+t+2ajhKNuou7qGI
obAp95npnnPrQrPxrThfOjEB4gBzxHZSDzI8HTmFZKLmWT4ERcLOyz7Jjn1Kpy5TeZRjYynWWC6r
sjyCPNLz0wsbB27icYGR67hXR03kouLJsajs9gFt8++r5WNDU4i81OG80dRryuGs0j78kNF90D8t
PG9r8P6p3c1S+pV2hYXCzF1+R3ksSkcFAcRef0J36/1TyHTdY/uI7vyomKW7evk9hg77/8vJiBd1
TcgCxA7JP+jiecoGDtDe3iB9JysBx1glB6be28Obhe2WEQVkAWzKbH+9yToyaQIupbl2Ps0Z29V+
FTn0+EZrSYWcYhyvgOpKOJbyiXFCtjdjU+YdI2LZxA5QFRuvi2Jk1oLpkMAdOSIt6RxWcLU5WEfv
N9LqaEwRMbPCCuKZglhzTt4lBP94ZmgD5aZoTRBsbu8GU34qkvxcRVCokSDzyI+JKAfqHjo5YoNb
K1Buxj7qChMfTC57kxcOwn48LUsco0tlOFmmsh/uAQXbDImFGRurYOBl1GgPx+Hq8Q8QB8pesQej
JQOeu/HUHhnrPZiPXbwT4IHzFxmXufgescMXY02XhAT+IsTCutZWDQ3Ro9Qvwk9djBhmtxduYIRJ
BuCTVtdgVnesv9ERjjRC77yiRTXZ0RYHqEWy/9GoiZhvPnmsH6T2PiIExa4Rp4/jyFJI1NWzMA8J
aPmJWUAA02kGHbtzqRc09zTpz8JQ9+zkqOOakOAHSo8YZ/D8zp5heedxXQmNx6Hyny64v5pbcF4L
IBrXmUOSIg7fUMrgIAF0QbwVb6tBzxJXR16NaZVt43VINk0vWmYJIUyFM8fFC1Tg+kiNX8VyYrYm
3AHGb85h35q8VHsIOfGTkkQpDHCiHDoMIbBV3LozQ+fai6U3lQU4wSSEKjwEZFuOAFB9HukA7T15
mFgpG9ey14J6DqVoXcG/dMi3w8/Drr01Xxi7MNbP80gq4lwayWoc3C74CqPGTn7OCcEkb37pCHJa
0t97hi3OCEr+CSCGexM2XpJ4Oj/9eUkGX48TToN7KkcQL7+ROPvnRoAjml4ptRg3MiOTSDu1BHKu
Y1zgT3+wlm+7jNprkVEmXtNFn7tIqordeFO3RkVWofwVeH9aWBOwQpCQofako806rUjdj99fk+hT
auDDucOFeiIMSxx6GcLyHT8YOO63DBqPDReizjTNMV6g0TBEVU7Xbfk1uo8cQWTcRHxSVpF3QtXQ
ntf51ZaT0EHGB3TBawp9xh64tzmSGusX5hr/GOcYYo34QxgJXHb2tInaoLvMSwopSjal9xVcy17a
/ft+6aPLmBWjxQ/8xnck1N0epSkkK+bTSOdSdR4O8OezhHZnIYrUg6Pn4AiQGvfaIu8rGdo55ZDR
YqqOYc/PRPkCu56M3jCfxo5XI2SlOTpDkjgw7TwkqPaxi0DNFJy6e65RUT8DIw0/qymqcTp77jxd
w9JBw3y+K2eCyvezKGT3+G+fd8m0PIy6jHdiY5DqHX6ZRgEW2gM6OVqQJ8kUiavqe8j1eQZFyOXA
c2BZMpmhEWH7I4EluADQH85cPyE/vEir0sZtF7bT8xJ7FSuI5AHCLODGAzw85j/GCZ3XfwDB1yxC
YAGeY0kh+9tfbppCigNrGSyAecm9oau2Wmjzq3w9EbRmP0BTPTHr2czAU55/XEzwrbrNwXy4x7zz
iM3OLY8vS9F9rhYdyzRv/AivgtJuTu65EQe3Aqw9kIV1aKTXLvu6e06t5U57VeOGR4Pt2YNs7PsT
TXTIlMjmhpxFvTY6S65tlCzdeSC7xyoZv6x//Q1L/fKph8izZbTp+a4nIW1YSM+b2OpNbwNkXAPD
0/s+MIlheRzyKyVYb6Z85pVHoczXX29uOwFqHazN640aEbdkKJ/DSGsLV9sDiNLncbS0cH05cpyY
vStAiQ4m+XJRkI1KU/GTWyfIE8xVkMLmTrdYcGF1I5Y+re3377o5t4gywW0dO3pzzf/Nzioi7PFj
DIjlztTGqR2Aue0Msaaf69q/8JyGgu/GGCfec0y5uX/OSJDGA/A0Pd0UU4Lah8HlZTahSY3gRtjs
X02mj2ErwjDp9GEiHJAecEbgxOgwKA30iu8iv/tTzgXR0qb8fgKXtb8LCy1Z2nMCTZc/bDt+fEXQ
8lORxKurWj4QSpRbiqacj8RjoNqWTXh37HEEkT9U+MvdUh0/+NliFIGbu/WhA7OmwwwWFakRdzxQ
j+Ii+v68LJBXUq1U/siYtJBzHkfpFxaAcs/CkUVvrg5wK9XjMmnOyE0uhL18JcqtRfaYtFZtY6ux
9+eMW5odN6fVcucBSQHF+6fZbqcHlmvW5psqEsejSBp5EoHMsp9zRIwYgKG45kbsf+dft/zAK/X4
gZalmpxcH9ap0t54VrsDE1M1BdVvJJ9vRx/2F4af9Vbc199YON4ysbjIQKjlb5ZVvUzmzDs5pfvw
4eLgJmAis0J4QWOaUG3MPBYbg8vxR1kqr64MLuuyiekhRoEYCgXWA/+NsbLzSN+4h1WAy0oEbEDh
wVvNqklhjew69LV3M42R45zb3KBAbDR8ann3xtiI6RBONIei609yDBvpqtNktlVB3+uGss8YZeaL
ytriJLtNwEdsCnxCpPrTstK1glwUQV2UntiaINXZd0dOcRdycLLQ11wC7ptKqB7M4U4kbMNrVEFM
ySzqdXq3Lq5x4Xgw8sQdQoKRoYcD20Z22XBxglCYqzvLtck8NrISvgeQUr/F38kiZ0z+KkdKbGtU
CIKAM4sJ4jIkvqfcz1Sg4u/XTeQliBaGcKbGlIbO+pE6i1z4wWMEVf7dPGnpiaY5WDbPCI5jO8uR
QP/xqt3tmORIb87AjKHflazdVx69p+CUHQE4nUvT7yunzKmsYPxoXHFfl/hjYi0IM6HgNd6JzHCW
Oyl9hA9vQuLCY7EzuWQGAhoYiWz9CaEjlWxVNfMB5Ed3NVBNGbpTtq1qr9GCQY3l7hnVJEuofEYz
VmcfJlFjgjvdCCsjz0Hsadao9K5oPe7g9bFr4In/2MUEa06awSgeyrbnRpWpj5oHGrAqfCyNM2D+
1x/nhzhr7M9tLV0bVSbXlHBfB3bu698mighoXLeFWOJSUWT8UJkyztulKZS17pLvV9OFQD/tywYG
tFsp6FIX8+EczzDddOGHUhc6n4BBkwt4+0e6GcPMSTkUitoVQPB27Cp5zZUB5FfJRlvsqxN1C7FA
rEMarHMyDhc6NpotKQr3z6A7lxZH4RUBD3FJUrX1IdJ26EOeeiUclU5gbPHekFMj8NuaI+5UGepj
e/XOaRhQHXVT9YtqCvuIhqJq90rVHdMEmBu30RBrqAnTKH3nCDPeI/y/LYK/nrBMVzro21U4+TSW
YAxz/yMFjGIHnYrVC2VrmXsV8sAY52nIods3evwYqLbnUrG2Qy6J3GQwfbeA9cEJhYdn2ctevMiL
LbJ2OOQsld3l6eZtiG8ZO69XCs1wE2yXmuHjjmn7GZq14cUaQG/7iKO8Qyhh5UN0KI54idZmvCLF
vsqFAyNHSVWNPqBaGm1ouLQf7PeT5KC8Zg2daOaB/HxByq9rgCL9AewZngs7xm9vlSyaZ2RivnDa
ASGP9Y8wuNhyv1KRLmTw2VwI+UnTiEoOz4jX55hJP73cMVW7drS4dp8XZsPsAdy3ztQoSMZdLxkU
cPYQEyu0dXdGLde0pUMOwDaCM9U8IJcovRVTDgUFzKwv1z3KNfnooNOCnLKiFhB53IfkXukHQl1M
+SNXIcfi0awCOwKztIF2x7TiC89GHxcpdpIdjwTlEAr00mucCXoG+5vny9nBoSVPwqK25qhQY04r
XzVe1zpXUSnz4uJlnL7I0tTKgU75YaZeV4Tv4QZrUEem49RWLwe1mm13NDhDCtRWTAbo83hRMcog
XKKTaxFuWuiL2PnJVt3TheI/yr8u278ogTuYNM0FySkdmPppANw3RItToUB9kho4qPDkiQOndJ+V
ideSwXGe7ZQzWAtjBtjVbjXE/kvAZPft5r4VSPtBIorAUebyoJsPeMs3+Muqb8YKwS6yakaVzVPU
e5lkAxfAaKEB90ZrBxffkGGJyrbLop+seX532POdWYfxIUptDudmgVbPY2x6V8RPLZgGaZwlZkXV
2rynFyZf/bk451wKJV41xejwof0nlxsjMRg6mQLYPWmNDvqY4Pu8ViTXizEnhARKwJjQrKxTYNoS
K2Rr9j4mwdPQw3UnGmbaHakEHOhTyYXMaKGkBhGNptnhw1S1i7S+RcEXOkGA3I44vBml312dF2BD
KI8wwfg4ZntZSffa5ybyG1B68cmG1aPARnP0Z3MIqvTU0po1rFCHb2eyPgcDFSZO7nrJg3gwbKGp
+mVYLjDlyLRtLXItUee38vmKs5ZmG5NNqJDknlVHl/U/Cbkn+vWA3wZS0e6XHBfRiRwKb5ZE4+NB
IgmADxgIPQCznl6S0sVlGLIuwqgr9wCzxdHXq8c8TwFl2BBqumhIgefmF9FWAqApQkkSRNuTRm1N
0csTbMkCV7lefO3NXCir+wKDhyxFZuo6+CzVOGh38G3iwIpjdueQImv0ajaBQMfMmGO/0XbxJhZw
Q5Z/KFF/8a3oFjjqnbYsulgjF2D9yf+crD2cjpjMelFV/xi/14B331yadgbId4dt65/uuVqRpCkE
p/E0P9Z20TiCCszp+CVFxEq0680DgqEVqCsy5w8dll3pQC/nFx0WUczbNiPWbpkOlImE6w+B2fcE
EF/iPL15Bw1io/bYv2BLeGoW9f3n4v/ejneaeXDbkTA0z8M59ePZPeh0vF+MLqJxJw1KxW4OGoQw
kgVSMfMduupCwet0JW+nlc0PMp1aqRZXAj+4lm2PGuI36vCsOFe+Iix1N3MJK+kliRPt/ARYd+Xx
tqOKUcpNe72TIRSXQxYZdguPp37z9iDKpLfYVuQQy4kyFEivkzfL8vfQ2nzn9xp/7OsdZnSvAQ15
wMKe15hTaPBV50IwtLsRavBdUiWRS/3iPq/3wNLOhgqf4E5pCTbezltkWAfOpjKm0WPxH0JRaftg
YN1lDAi1CQjYcysaVq0EDllMtzzxzlJNLt2w5WrdoinztT5Adij7+KKgmsR0+levm+XrRzbdwtka
+pwUaHgzB5nPYeBebarW7wdF00d3ITmqYn9Km21dM2I/betVVcqA3hLQLJncVjJCdhdTlhnAEAlI
a/P+AycZnAYN8wmVDoxM2HERsV3quP4q48gXp6YJO/o6kjdYY+joaAQaACC6h4k6FIun9Upo3gTP
vq7IsI3mDOSQscF606ZuIC/j7zadSbUCRhkRgiTsFA2debcp48x7ilNuoXtpdqueuDHtyXMN5oaL
O9P5/D5QRHjlJcf9yKnnYEgkuTWG2UtqkIoGuB2/coeAYtcpKJEXvTABAdnDHaiWf5uXw/WIaByY
tJeTJCYW/Yw7O05+0fozEoZLGCcn88EhswUa1p3B2Lw/cRQS09yuulpX2LNjSQsbIAHCK2quzYgC
FSKWUlSgxzyedDh7u0pNH36dv7E7DDO72wiE/MqhrCYjK0ftQmnXOILR2gd5bt/CtuNGVaiSemdW
kPoWNtOcNypNz2Q3mX8R4oWEVNIqzQfXTi1s0KEzqzFNTI7ttQIFtJAoT1BTv6S+6UAEBkAjgrcj
JOQPlMEyOmbTP0W0QKhmGgV9Yguo12roaIhu1i1am9a7olVi+dwgvqq8PruPkL5fVlQt0wYQNOm1
dSpnKmiuN6xjWk4yeIZ6zljBeH6+/gGx6m0Av0Zx/UN61fZrO2DxMxaGpfNytserIloUT76Q/3f3
P3yGgidYUibtmzl0nZQpOTsnQmW4PRUSJBbOjjGH49Xrd1y0qVtxrrZ330wDbbCxQ/b3gHxesS80
su8isN1tZplPc0GE98chNcpiJY0Ffdp/Go09syQsoMkgkaSq8VThTRBU5GbdwXxDeWWfocUrPLqz
JNWNUG07KKRSdkqdY+oLm/b4tc/7HbuQ0GNG30Z9ieFCzm7XTEs/eW/8ylHqtyibXThv8b9gVGak
nsIvNBGXbVMI10KpXHO9YGCdQvzry5YTbwbzfdOez2Xbj/Jk2XByLarEmibbU36Kj4AWHNNIhQij
dLcF7bmC/6dc1NUB0AETdTR2exo9Q5AcOZueoQKNLq3XYWqMccpjfVPNzkXPhL55dYHzOSAc776x
WWHMsPW4jkUhu7lYSwiwMgshadrfSfrMieeX01yGiUFh5MqD5OQyy+6UteRarkNV10ratVjX+2CJ
JaaZXKtOcrx4LbY6wByudkLob5U6GZ3YBTO1aZqoPOsTjU1kihVrK1IQ3H0vze1TpgMQAOdzxXbu
kFfmfMZmasL1wOi7QffHIilkqDQ+8tOS8w947wR9WOpAErxXOHQi2aNscR27+wf0baGIQEkzab0i
wjb8j+g2Ma+nOdo/0jDk1rquR1eWLJYP+lwrufgHWQUzsTwICpg7x/sL/8JP1VtpSvmm7r0AUPui
iz7kx/q0JK5XQnSRiXnoAJFitVqF0VH8LsTFT2pVot0TWsBFcqLejSpV5Ma6+fJJPoFYNVorEmls
+sXeB34LnTPbWs2TiGQHLUqeQMwe7WadTWzWokTCXLfQ3MteoPYPJ4GfQHA7mwW9QDJxlQDJZuwX
mZRgqb+/cnmnHD3HjdURaFsAlyXAOBPgyIkpJ/GRE7b42Bb+16FyQnB88TfzILLJHZLbIoaQthlF
BqFOFFL3P4r5sWvq1fTNfqwaWANewHLrxqSFGICUDY0kTLOVUXsoqQ7YmpTSGcJWrOC9N7Dhr40w
86TfMVKWi6ijPprZ0c8CuciGya0GEFtI1NI15Feyw9aczn71MOmwnmter5/jPYKaZlE1VXhl12lB
l9JNzVqbPWkp/CjvfvIFqjBvwTPJGAju64cyoKPT6UAkyMM0FGsW0H0grBsbg/zqLWXb5O79gSOF
J9lF8J6FGA7ONxhcpkq9pbQO22DUc/upaMxO/r+4vV3ybQiMEayleCY0suALFBhtiSQvytI/p449
3RstAaeEVduN1wjMpiJJYSGcSI5FqD2NaYhlD2s+5CA93+27gRzc7kfu4s+ZBqDx+IFSNdFn/Fc5
UxuXZGYwtG0n3rpyqgHUO3fjRq3Zh92voQj87fxLDA5MaJLgmnUX2EaAulBxNpMB4skykA8DHJ69
0y6TAxiZcnJ7Vdzra5fLfe9woMmtXgfowRwwQajg/V1Qv2dGkcGBVQR3zWYuUIJV7f1v59i8zBw9
bMvOJ8a7QjHVz7jwfxuQ1xuoxeRdZ4+mu7rcRKC0bwiP5h183UDrH0WMM6U+EEvBJD/HPQazOlUO
xz/PR5K5hWvq+g+u9lSUj4dwm+6Yg++oPp3pDQDIIFFWdYyLWVQ8a/zQZkCButBpilZll8tf23ru
Rkf+8u/ApjVnXOoUE0e2dtM91lHLdlMB1fMwwNRPZSSiHC0Fl8ZrwLRAKpE2clNQsmJvSEdpZSJe
Wiajhe7KTtVRWA2cw/EO78/0VEYn4yjW/mv4y5pXQ7P7PO2jEwLaRAyZo2MXjOw3XK4eGonCo8hm
6mWyFAKP+QHUiTsDO2ahc4FjbGB+hqbWMr+D59Vto9wW4/9AX+4PR41pRuTlJYxQbO/9qPvop6WA
eLaJn6S2/m5ZE/R8UzUrxWGBE5wDmp9kXzITbRHOK9Xhz59tuyqejzCLNyzjtxwwbEEZRExE7lzt
j/+z6lqvUq+J5r6Z3tdS0e2Yjbi3vqpBLS/T4pCL0rfk0IPWRhNCYaHt6kJVKw7GGsWRQXWW19Kk
WExNDdaiQG3vcmwr3WPQrTkPCi129jEnMe8kxSOg4KRZK8bVlE5K/Gb3qywQV2XMd55vaV9RxIwM
37XivpXhWOuhcwOJoMIP2lnc52PZbWw8EPwpXPxio7F6zvO6a4ZIliA52yUK27Zv0Wx5Y6+BYmqj
R6xkzLz+deLlexbf+3WLlwGZxyveBBf5/wTle6fZaHHZ/7J5SWHs3uKTPIVQqr5C9g7F9+f1XWI2
2NCIcAoSedIctmv1xx9qW+idNpBSB5TguN6BlBTJExr8gVERokqOpFvrKL7gzUliHgYXPQsU66Po
9fPfW95E22H4egd69u5xMyFAz7CQp7sJ43vFT+llOAJ8+KvpywryNyLk8d6P9XgkV3+HV7fX+N9V
kIsnzg71N3IGABhGfFT+y/rzMinTOcXxjpZvZVuzoMLSwthRtr2hDYKcqdbRUn3sWX6TuBNXtCpK
FL6/g1IPkdTyZqv5C0Q5qJ2MhOK/iom+LwT4/fA0gw+li1T3v3926BDQmGCUrShOZLJIpadrxoOO
+J31c/7fq/iW0FtX2jOqjK3HVejuzPCJxotyhQjQnuo462EJJtIEbUIPBYFZOZvmRiRblMarUdex
rDxbPDwsp56tIlw2DMiZF6uvykk9bYN9rG4nC6b6g87MlA6iO46HDboodPkkItT64ssR/P+JIrBs
h9o87Ai08Q863TdQpylhZ+a/ElCR/SeRAWxkIPoqrFwz7yCe9Emi8ioN7LvpcYfdK+NbUUVAqPan
FmaFxifN4+Q+B/H1iypP4GHBtFhs+xwe5qoiA/k51GAf5FuFarSDeaZjT2KqP2tAiKmfmb6Zc6bg
Jb8TtL3ATa+2K779KlDWRgM4AZrMwY5F7fxhosUkGZDSe8D7Ya92d7hHLXHQEcm1m07uFt++w9as
9esuQcme+J9av3hQlUb49kOsjhwR4DYypjlzYgjpPdZ7/ATFh0Zdjs86g7kOZMiY/POgEFGryyBj
ffFunVZo7WN23pxPSEwukQj25kvEUhQAQRJxswSdyTStpF0bUGdM/n1MmQHOHEKgknaOpU7VDrve
lwMSFtzXaPkElevAqEm9+tkjXAhulwKsfjCPnUrvJxTDX6Kn6cbkkCS05zmHUJIzksv0GiwKwML2
VhPAOIe/v6X6OGjY3c8J37jEG3w6plQ0E7l8r28BSChqtEz+WBNIGG2YLokWchbTpK9eHlOwH6Qp
xEwV9h4eVz6zW9UelqtzWmF0OGISFrkm+hcWGww6OKGYGi0Ahazpankw33MLv+NkS1v7pmTqIi9R
fHm8wLztIMh1zc11XH1khDvdBUsUu1ghPkHBfRMzTsj1Nf9BfQFAA+BI8hO1YNWFNZUfaH8w5A9E
PuQIBgUyx9e24AT5eUdxnhRKGqC+/QKvfuvGBc58PqmDhbh6jtb6ooW4gzBOPVqzikUo/wOvqMiS
YXJutKmCTR+kuiAc0Op55NNB1D/c9VlRjQw9wLwD7Xw2Fs8BqbJkZyeoj45UcbLHyAzJSYn1rjLB
gD1oG5qua1x9Id/419dqBRy/LghHYrJMlV6R4Mb+GMHdzgC/mgh2smMefldMLKaUvExbbc1+/bF1
uSePCUTNdckqzlLdDCNXMQUe6kRg3m8ksy3txu4b4NNawcYA832cO5NnJsQ6KTt5vTJBPugVp9AL
IO7KvRLWHRNGWyVIKhIGFUTLRNFEimlPbPLkomTr3Z+wytYZazVolj/rKoJrMNdPjai7pDqdpLJm
l+ttgOJIKh7ZB87GUC9j/Yqu36n4iGwiuPmcaEq7AKfFyQdkfHWrqz8VDiF33iN3pBYQXBg64o5p
S3dzfnRzBxHjk8CbB+RgwGLS/C8T3ueYPF03k/L1HRvkgMmAs6Q1216Pxo8nsgz282QUBwMUQoGE
ZXvVfN258gO0nJE3wuxkvm6Nk93Za18yJVJfJqbWSIdCw1O3yBXaKkfUhVe6HCbgLO9BPWbw3feq
2VObcmHR1lZQurGWSl053gsYFI3JPI38HugfbgLSw0lhMt+o+j00V7O8ZmYQG3h8/T2YY87hCGrD
lL9XegxI4TWCSMUQnTSaTIjIuCpzxqTBUS/cPXv7cBBhJXCuucA6kVMgrLjMZbT4/dwQlB4tP2cp
/KfeIv9HND9YZeLRt8BQmHSkhGLtevoNqANecVILEEKUxhdN2lQR8HjXZoPSTprtz+vKhayBT7Fv
OgLEjYvJDEXSSOK8LeT1nWCmWuUzVAYuFlV5PYJBR31NiRWyHJpb5f9Z/3l3VoWjk/CbDsuTWDFh
HG4ebjhHv7vkV/IFvKMznDKvUfU+Jxu2c+4KU/GsTyD7WMk10RVqLVTKs85HYRTrgUjE5RmiTS3d
jFTuLo/EBXklfrXObJxbZS/yRhbdA55Cvy1ZA/SpC2qQmpCeZJ+L35A+/PqQvqcWNPCNRLcAEeY+
GnaxtqsiZMC/9AEHVbSq15RGBemVWO0UYhIm8puiqQc5gmXI4+83VtqAzbaXpEREAm3GxVS8dtUp
3GTAq/kGvSSWvhUnd6w3IBbbjH826AbrXFtpcrs6C6UIQV5ZASM7hUsVER14aSkRfw+3awJOCmQv
rxRetNwx3+R2oIfJq057M5zILTTTdadOuHWoHMpDlY7rP1ucxaOIMKm2RJwQdG3rMdeBlBn1LWaX
wlvSxWPchtKIwgMzPkpAVF0Pq9WRcZR89qZxHoeVij0Iu094GQifb8qT0qoUurnRCIgk6MuEcIby
h72x8UHOXSoJDqDvXufX1DdZtm8Q8L3nm3198bmPZ2OzW+PejixpF8CGFCnAZeu6R2qd90s7vLNW
Zms4ayLyKlsyl7lZE6unjUrG5FvttCsphLjo5t7rzh/LSRjVWE014i8cOBKJ6UCMp6eeTyjfMKxd
b4K4TePk/Iph8b0rNlgKIZR1PvwK0rwBpByTUcBmp5+uLLCb4MiEPlfvkn1DBpLbO9Sc3nwVBiTq
eBbg8EqYQZAo079GxkSARBN1G9TCnrmllaOauVJDkKNmhuuZ6PY0ds1z7ckqNBbHbem+cxBOXI6q
pOT7HVhzme21Je5qEr79V6CsEf2zYrSEeKQhE+J/75AHzzjydDQhhstCLcWxHYj1jX2Rbw9deu1Y
VrHEBRfyHjY0Hgr0k4XkTj9OQWEWy2CADwUPsDDR6vr1wuFFDSwbo1A9jRrz4Z7NwBr6J3lfFfwv
A9LHeATfWJgIkzZuP95l+lQ++itEqt2dqHMmMJx+rGytK6HKVhMHZmMTt76aJAwhKZ8pWqlJU/2x
OEaA05iy+v5ZxoTHq/hXi8Mwa2UehH/PFCVNGeiSGs0Vpf4J1zR6B0xD+twqSxeSpY3Q73PH7e0S
LFTM3e5H66t3BsAgXPFOJ4oQUWBI2VYcnL+cVzwGr/+hu8ZAkZe32/xNLc1UlsQOEgTJujN4l3R8
BoNdh0gucgo7EP8IMZcKNEr0Vy3yR16V3OBPWqElsp969CfZj0XfP/I9z169GNgOVfFlW+P0eZ9H
mt5Arhcx495IgPpY1NEpXuov7Rai+mQB/SHnzRgmCJruJRLnV+hdpMva5ijWFJsSqbDIWtfNnb0v
4FLnYmCunv6AYaG+kN51DrW3MCxy58dsl1ARUBjilW56RIufmIhUqhV5kWFuiRaOxMWp1dkcxcL2
Gbgrd3uEfvWzj1Sor4k3IIgmSNB7tOX5ZekoNPGAOxRxnX3SY23hvlGFKDGSu/LjT0tY6X4QQtr0
3AaX+vQUROV/pvogI5J6A6C8UELwHKBGrTLjHMRrxNYDigFYQdyBIT3QC+LAOBOLMIDbPzS1nYqT
VYccU/SRgj2wHX3mzNWk2AG1u6miQXQHbX/Xet6/Hgq/yDStijytuzS0hsKsOTTinL/ariNImkKR
KlC96fru861kBok5SIaKY7IE40s6DcrhH2lgBnjvrFV0S5TtITVtnbZqjdMAhxBJwam0zXoxmwCk
RCBw4V6Z84ZazsjJbazSKYtP5vHSpUUA2fbO+aGty0UnKsKx4Y3JjB8Y1/NQ1AjvQ+OVhrjeWnMW
BRAgzGB/yabSbugqOpdn41SXpBd0/te04YorFsfpnVxZjGJFucfgbpOOLOcCFwNFKBw+RZmBo2a2
xLI01WiCUaYu0c+vhqS+emw5IeXTeBgfs+BIc4RlbYvVuErNzofRJkfi4uuw63A254sc/5JCOXk7
wHvpx3cm88K/bKWhVRSKtrJDk9FzLdmKhQRQeL3xsu7rfUGmfZqB5qgZsk/P/quPHqNokA5QUXhs
4uojH/Xeqkkwjz8g+RXqRm9otCLRGYoeqS6745oy7945c5PPVUby5Na2zCkJEwwlz+Lb1xWNsoVe
ofZ0etg0Vmw6QxXtzHveSptvo7KQ0deuHSnGDbCgh31B5OeXsDLex+qSb7NuOQly6Vo3q0IAraUq
1Wg0sRVYvBKP7uvE9dwnIq1vVsWLfuAEwC3vB7QFbIYX0eK7qDW17rFBZK9nQG4CS4mnyYM1gTkM
8XUNhoR3pDedA+gra8GxOkIol1XyfOtYksk5xpbKPdN9UgVjNTQhotWr5PeMLJsA4CYF2oucP/qe
tOfabWc2o8/DlPqbIW+EytSILCUN0gmJibj/xnpxHv1E0S9gVn4pcvC/UHY/891BGU0IOBBNuIes
DwtwOUAf7D0UUOUJKNbox1ePdKTIF4IqzDHHJqH53sH9b/OLduorLZSPzq6vA6nwxwfJzV3Ee15k
T25g2DKGEWDf9Fzc40S9HM+Z7XKpQgSt3I6b0InTWwIu0c80dYtbRfS4/3FHphgZey/pi2eT+20W
kD29yHOI1TdC66l35ruzTGjEGa8SunjfJtW6xTrk1U1NDK5323+F95OGy8qACQYVyvsnEVy67rf8
BTnsQUdBF8oIi8TstkkIl4ewkvHcwQsMKZhzTAA5LFv/9QhtJFQrQFNriQvr/RmALxAqNaf1Z+xQ
0ijVpYUNAt0+e/0GNvKgf9jgXEe0LKBrUkrMAAbChpX9yaUbX1AzfeNKYC1vATMYDoK0dGBMHHIP
FlKdKxoW0sHmG3oXta2E3dAcAEEU9tyPhbFhjGnxh1LmCjIj+CS3Cj5T5/5kU0Qj3bu08EjA649H
LebdPItdKYvaeiRpE5k48SaJx1k2ZANZITAddpNtIlZKWDWFBcN8uAIzVwGq7IdVKbk4j3f0NyC1
9Gv020W3eNIoxqEZPHJYN81e/KR2mXjyjX2+qKbTCnEtPKvKIv0kobqlo7lDuYt/bNAQlrpFUTyu
44tTzm07usPcv1YPDvdDMYWuCuWLj+XNqbuKKaxPDn61btBq7aSmxruz5j5koH9rH5q3JJYgCR8A
+wMs9MIW32jIGEX9XKDczELScPsA/zho5FKW2nE7SvVhZDo2pBbsqVbrdKgh+5ISsRrhIBKxO/7c
EO08/oUjEvrNlvDvnwhHQRKhIzTE4ZcDhwesnxmiB4Ut8j32w2+4lJQSHArNzJ0Q0wiKMRrRj+O0
u9bDr5/YZpOauQY1uFHMVCS548g8XaUplY4QA3aE/Fx9k9M1puR81soOOLd882jDxQuDmzIQmRmp
lR3gMn8GNIaKtowqGY1Y2RfotXbVENf2XRTqbyp+hu3/zic/VSemB8OAezWN5tXad7+f0r7vqXfJ
dlubzME3Zsjm1e4radKkHKSCeelP4594qFTdh3nLyrVrHemx5la63J1HKumF4FZPqzN762+vnJgJ
QPpYfxhodXPZabICmVdC67IGoQtLxl5mXt4GCIZ+rCEUadtX6yBFHL9f95sR+ZbApUpRk8eRf+lT
dca8Vo7kswXZG2bJLU/kEdcnN6FiVP/OcITfTDVBhafWDBqeILSxxpzd2hALeMKf1b8UEt1xa/dU
sMtBOexKP5pMxBJhdbL1lQDoj3Uj8p/8Ii2yq9zdtPFpQTc7G4OVeB0NjFIKj4CtmK6cOJwwmaoa
ssMjZI80GMQzaf3VmvMFEHrsAFBAfkNPrStqNg9OTZBVeQwknMlbTgyzjnw00+g5j3yWPfC/MpQ1
rdjcFB2G8zGwZzqBTK3vZLNeK4HK4whdsIf2MNld29NSg4166Ec+fR3YzSotZCi92ZZ83HNaBFfI
Cxk7zXAgmoQ7PPImylKRqa8W2UUzK7tUTXlUjKpWwhkJNkHQbYvkjTgUzwTL+JOpbx8vuOr5t2AS
krG3veWnfeYzpbAX14ggYi/bEOJnRJBhBlYKdwFy24mKD/tYjHjJi4dDEHXcnle2ggN33sqfHxBT
6DdI4bhSGE38JwIuATFrgqVvWkmWR0UDTrFXsLMBuRpJbNiIeNl79x+kvthdLD5vCv55u3C5ymN6
NtQMnqXysej3dJY/oqRRfZawDQxzG+nQiORhKkZ6SUTPLEr5MeXWtr3ur8uHnWEeywqnyR5Czuhs
OhoeSKN53SR0z5RmuKW5v3klv+Sf4t4YEBpGB97rmb+APjxETBPRDTOJs1ntsP/ElvmNLj/1Q7cR
ONdmrEReKyr27vdg1AvANdapVNgKvKSuOcIpfGJBJS8gsvXpY5ehQZjuskBQzNOATGMdsQqE9qsv
sSQzqfT+XpDPJlHk3pCzjLmop7eDVPeqjlQMZZ0vMBzcnSK78fT7rXEE0ZiShnUvp2C9rJEw76DA
x/i1jhmLDTr/B0SyBP6yJE6E3Wk6/DQh2fzu75n/VgIMNWOMkQ39+w+8rrU3tUQKYSYO/1g2pVQt
FH2OSmWYSF8A57jPQuWH8+x1r6P1VKaS90wntjok/sN9HnJSUgTS0a5BjhEoAz9EfyELH8/iXsy9
qLZOCKxbtmcmRS/5dSacfM4jvuInpU6oIz48N8Breo6ffm+amw96n7WdemMeXquoZqfikSxpmb6G
eJwF47Vj/0JF2OgoIwyDNg2/tlM4YfO8QcT40qXWISoOmav55Xg4YTJKT0jWXZI9+EwUyNW6kjVW
gFX/KYIYF7oT8EL+yA4tNFRhdYO/FvXTA4TXmBA36nxkCM4EVB3ffXMv4h+hAudWREXctnsNrmPV
M9RxbPUQRGCLDKqegzdIIUMbRv8Ki36sSqIup45jwZtl7GL/Z1vxZH95fIcKz2hLTtBY32GshMIu
meP162N26Ag7hFVrp7ttZVLvcCOBgdRlAhN3Hb2Tujpd516mT8yUXqmKmuzGedesYrFpl3+p6AKW
PZH1Kif4nDbWKV1qxa+m2yUq+/ebaPmkIcithwNh1Kv7TbJaA9B3F/Q2zkfhJn2+6QS5vW3q4s2G
bkrxaF5oPBntZ4f7ACTe7l37NvBGIQ4dMIOXyBHKmIRmKINCaqYpRFEDpmP+xL5PbANg5t+W6dm7
kPWEKPVvWgQEaWTM+uOtywIyvaioQYwdnK6Ax2Jxl9AXCTb0xMDPoIgJyiY4eigsy6pdei1oVAQA
EUdY9qimrTpd5Qi0XG5vSmo8Rl64lmEiQ9zdN/BlHpWgdXjrCsDtOKh2E7KTzslIS5QwQya1OSOC
rnImzYSlRatinfzUtF2TUuJ5JZ9oEJjhtXjDD7W3kiboBrTkRe2H6xdwHLWS7tRCxaWX233t3lgL
5OYdBKx4Dr+895Q9mSXLXglD/MEpf4luvX+/lY870PjSPTaVBh3Nx6RV9YAvp8qSQ22eojyOZidM
N2ryFMaMaF1+4cMNGNfIdFk3PcUIVtD1H0o8jithOIMZxchoVKXEMQ6Sz6u7D6ocRkz4+oeSozdo
WyJdlyRWbPb3z2wTIowocJ6aRW06041bNMP5GcxcsHWlP5aZ9P8sOC/JlLVJvYylTHQIgUOrm7uf
yvPdiahZZS7CkOJ7mlGkB7OY7Sns4otIEkOalvQsOK7jGmdyniHp8kLWZdu7llEaMT1F5At80rMz
c2swCY+x11BMJ2dWcs7UWppYNDpjQUv+MMjHoxZf7g1uWsI7Y+vJk3qrmIHLDDR2BUgm43RBd4Ql
R9w8S7OydLpMkf/5ulQJfMrXn98Au9Rm8HkTuDcvTqlhcIppyFSRqwIB/m88dKrCx2nGO4Rj3m+C
jCiKboh9FHTE3Zoet+Byz2iyt8ZlCp7JTumzYndDKwFZA/YIasHWzz6rZO6C5msU4zZMwGKS/80f
DXCSPD6k0RrhrmVqRq99d1sdxlytEANqV5DfQIrhBJ9+lAsJ2kkWUz/v/ngNvl9HjBcO//2PKH9g
+00a1/N8nTrMffjPrJ3A9HCSKtrwQRnA0Na/SxEF2vGn52Fm/Bb4Ik2k28QZLsICDBQsocU0k+1E
wD21o8MEUpf4pS76YqUJbtp7NhLz6YPGEEupPsGK4IN8nPiODEzFqDmVyKYdnS1W9dz/j5r5aDsR
IhP8iKZqeQ5gawgWjJAXHYgT3EWRAYKuMrLAzhLvUQ864BeOYMRRFW4bqyja0by6PCIitsz5y2iZ
WsxdcUOfZPiMDJXmVAGM5gMRtzWxXGxMJCjCPdIomRm7TKU5JaVXwdc6RRXQlIWlOI5kRiQULxA6
+iydgyfcKrjBkmx4CeWOD4djx0dB33Zv89mcefvb7YYCtwrC1vDtmy8RLyuIH3+duHHGDyiy8BaB
UcoQmT/L9G16oT4bF3y9j4M+C2PwMYqYNX7ITLe8vYJl8KBwsGvTd/EdWGUDRpawSGnhltsbcI7/
78fXv1G0bqPcxNrRCSnAlUyor+3KtVSgUZhWxAiMXkasyreYgmBJ205pDgFLuA6QmlAEg6J0yaGG
ZP+K5ulsl6LsgJ2u/8ijIbRnEg6Jxn/AyTxXqn0gEJKzDx47k07uzvzxpW1jrKVRZU1q3eRhgjCL
qSrC8Lb9raJbgeH4EeXu1gabhh/6yNluFTrhXwQuPRhpDhD9mxX/8WwEhZidtVHjgzdF4Ginr3Er
OhiSrzsZCCa5c4rYQfmp8gKlpK8JnEayWBz1qeXNq8ZUFAqiSF/YjcUMFVxnWytBLHj2/Nc30lPQ
bPZJUHgev/F0/kwy0egqdKHArsnAM1HkhaHZOF9phQK58QtWLHx9baUOJ3ou5G/IC1yiGWkOVVnk
aqxwMsnnrEVPPaqS1bAnDYOknemGw3UnQlF7315N3TIYTpPYy0Ty1hfwrHFuITAShHAv0RMrMEjj
45krnQR61zuzYip5Gk4omCP6Kz+38NTyxgqn2Z8tw1J6jXPMssgn+pLIUx5rHUG46jgwvGZVzDWp
1vZFvyLRqiJXc0tgwfD18sWsaexVKEBwY182MQYlpKzEWJ3s+ywHhopn6F/Z5X17JqT5wSaXnd6C
cCrS1JC915OA5dzDkQj3KMpPrdvATRp/gY1n2nVdRdRskhCs6kz7GJi7Zbzbie9yLof9zkob5Z4P
1MysGQ5I4Iec/L0zpSlp9kMkUSG8yRaOtE1bO3L8Tl5yBkcgp3fTGcx+8CV22VKYPgNhyzTer2Xt
sUEAHduGM/sHn0tud/dCtZQ9qjqK8MUjz2LcuOOxXqFP0Nr439RKVJgw61kpNkAd69ZoM/AUSaRs
CivbyLbY6sTlPbq6RoQma9LFFTBWR/CdCTOy5VHVsy/ujpQVX0vknwh7E0u5LonWaFy20I+fUVpX
XkUkVwxgXLiOcPuw2teESFA6bHAztGsemGgvppu9aXQ6DqQseHmbLPX3tq2Gz8vWNziY+cxBVqUZ
joJkbRDWiRY97V0ux+TKGxmxW1KLo7PJ2y+CIf6r20kNdRLDy9XL3VFgqdaTuI8+bdlvrQGT3L+7
1FHfBH840y0Oe3zy0Sx0YIasVlqzdYKFD5bVM2slzDFO3gmvJZLBXWkmxqYXiEdcie09Uewnpiny
99WsR1+WXArGoegOkx7CVUU4LM+I1TanKwm4RSovGqZz2p6AXqD66uyc21+QTS4tlRxJW2idFsab
Tksw1xyTQuIxEJTqgJaiJqb19VdB6QeYrH5ANKe1l1dx5U/S5m/8ngFPeIEXTsXyoBJv79Lpdb6S
XLB1MRA+lqGqyaGJzGfY3Xr9Z3JvK91zeNdLumaRuF0jZ/gHMXb/Gjc/ApoIXnR9yuwJYly8hL3c
WAUpWfUFVJJFvHKk8kiI2bHVe2l8D6EaASFoe3Ri1k7s76CjoFILoyzFlyvTn8/Qtl9cZnDjMcpn
t+zJsQGWZDpXASf7mrai34gzRZP242rjtZnS5DqHxhUmEXxnBklG6G/kl7d+Em7KIDpwut8dcDBM
Qs6L4rRB8S/ay4dp/Gjh1gGjcKWwhgtjK8etPypHcwS9li1Vydkpjk1wKAxhZDu90CDVVD8QcBCN
1fVd618OuXgVO3IUR4cSrptglElYzTXgChaMoIsZ7MBvtJXSeK1KR5Rbi4drHDJLJzOLuV8lNJ5+
CZcHnfImMAqmYvoRwirRbXUCi7L8yO/+2kcBcd5uH1mAN+z5T+KS/XnWIswdM3YVBXMMCmVL7IgY
IdDjuh5sOl+XQTT/FtsEfaEf4jD4+79ykzP+SDlPr1HP5myjXW8eg0zXWodeYnzHqCnOGnjjjNuO
cd8rmEz5n066+547JrOh4lDM9ep/7oh7y/o2RpEBXddCLTN0JbpDC3ZMw/1jPgF1eTkeCSpJ4ZPa
3VtAEMcEzyt5hUoPrrXVVajpfi2/OCg6C6YHV4XaE+7t+NSaBzN6n9nS5WXQV0JAkcwTTchWFiKj
PazoqZyYytJfolwoEnutFi8Li3IG9ndXSTlW/iSr31qNYfAjTR7/8nHJ4g0vatXgaiTVWQGv06Rd
7dZUyTwUX37N7pFFBOa16T702gymURzPjR/MpifIS0pJF2GohRlT1vIrUsPafex3nYYE/CM35Q/q
23u+XuVOhA3SGHpD2L/OUbLHuBPGuYvajYJHqHIKwAZHgY1dshdRSpaJFyXqK8+dJ/zYwLoo2MpM
Tt7IIAtbcDWFd/+FTihPG1Ob6xbwREof2E7eeVYQEphlTmkjkitC8n4cpac7Ni4O2DEzxJkBqDl/
M0JleEizvRGwgMozFXoAdhdEXU/1DxjkzMXQj6h8dB2y0dk0Rs/oTh1bZ2sGE2Zs7pxrJMyywQU6
qNitpfEwKt2GIwI5HMhSaTuXmxIwDMwk+9eIvU667r3flXq7OxTlh9U6HDDozFNXAB+lhk8IF+dd
xCUZielghe3t5FqYchX1qY1hayzL5+cDG9IPhK2AUDZWqhB4nqBMjpynYeYnBaOgGMMpmmhV6aWB
6NraEzeiKOGLuKK2TnhBY+S2Z3dBQxR2p+8Afz5GKWr5z30H1+lcMY2CY1nUODF9YHKp5zYGDj0P
TuCGUdMNDRYMz4MFQcVPpryoyIp8YKlnFmsAMuJol8YvT80vG7kBwLeD3nXycoowGKgZx2lNCXEu
744uxCnvEoR6FCssYJ23y/TtDM8MF/A4JAOpBeFtzsj975A1D/dvDK8FMECKmNkZyvjMinFpTH1I
kS8D/pprzmoZYkkzRyFy/mrQe3olR417kegYZoZMkYMpjGAz1RbEBD8ZLuPVHaeDu/4ZJuU6gDMo
85DzE9zLUld8SJL8gACceDYG/OCKPpyIAZnNcx5BKn+6897W3I4wQzg2rZ5ESSohxm4ASTxU4zYC
zlWiH7f0BCZ86QHMwCKNKLx3InpOv+ku6miMRsnBJSt3PV4/h5Dh6DA2ZxJq5oYLdF7XFiV7PrTf
1ijy5MNnlR/2q9AzU8sVSQD5PsIk17yJvDCktAFYKqIzWi8BK9p0y9wdirDreS43JhV9PKwvdh3t
VuC5EhrKzg+xUcyXYxoC7DrxaP8d3hvViIVaa3fWHcOKuCtPM0rn5vf2eNlRNDPe8B3u156bF+U3
PB3EWSdSfkVPEEmWS+05BheEd1kskE0CO//rs3mirv/92EgttbpMyvCfhNR7kuw28Mt8PrtV3XBS
MDiQQkJi/7hp1gtllBaoGccM5JuQ5zzGS3sgsWVxw+BR7vFWFHzSB3dsTAiVCqkjYWC0emwaiidD
0NN1aW1LEIiaB5Z6DLPjdTsD0tm8S+9wyZwcm1aqcbuM9iofZmlpx9MO7olVEJw+OxE6JTbBOYFH
MnTMvYMaHwwo9eyKSd5ucJW8Mi2tGOUastj/iwNVl2ylPO+dbQTIF37LoDo5a7Bxna8oHWKe+MCO
LYjDnv+bunuA5irri/RnkvO11e5DqOT1gTvFgDjg85yb6+ea5Gm7wP7IDARQlPSq4rcg0Iy7xCEc
8XIXsxLWoHGVj0DW2AJTbHerKtCKzrSLGG1Na6FM8NJicdXgO/OiGOjiF4ZPr14SVDVoMaTRqBhr
YdtZPa+XMH/+Ld6rIUjipZ7ThKtlsgzlCMFfomDJ+7Kb3DFOyBHUqReEoowM/3TjpraJRwfRusJ3
fuwoY30O/kvLx3U0s541zsUBVFrijGL/9PH6tz7zfJILHkEU9kpI5AsxmMPOADlBynYU03jzyPm6
IrlwPxzIIVffhvAqezCfJMf4Ur3nS2d0PoT4suRVW9xZ+V5+zA8Pf9lrrvrD/MKrFZmIDTdx+8VJ
PC2/O+j0byuZ/uAB0s3L789/iPL+9e2ndvAU+4BpUocusH5cB6mogsyTF/jsACnPXxemSdN2EbcD
+p9PkKlpnF8AqFnzzWAMggv8gw92MbazwB1aPfTUgypAgDvk9Wh1PIbT1g25q1jxCsgiM0tmv8pz
lj8StZCNVSreWIpJHUIeAGsPx9d6gSMBX+uScjEWq+HhB+c23VLvJLE9ygWbxT3IpTjOuD/rkvfi
p0ZcBoI9IRiKire/rmqOVtKBTl5sr+oycaAJ6zFFu3I257kyyj3LHIgg2wOpP4vZbgvhh0zR2sKf
WDCOGivN+5H+HpDyV6FKjPC7InQbImhL42wz1prub7Te1XGbXpdzvGLgKjRM2O0a40gYgap2IMsC
5p20U/9Ee1vPVPWgTQrWFwX0aUMK8MyTAddgPEXhKRmvyIrFZxC+yFKG0fkNHt8PQBWwMDO+t9S5
yJjx/Lcai0n2cefJmubaZ77uBhNpNvc18Y+IZxOFMVhiabUglI5S983fy+VQylVGpTBr5+P7xNPk
RdFxC6ZFEiPd9GQj9Mn7HPaJhowpkglRnIz81KeiUP/1mHCh7KVsE9YR/GTp2KHayYEGp6wWMG08
ahhJrTdjNUiuh5EPvavUSprnZURGpi0EsIuTDN5ULKI+1Rt2Sp3IvSPmGuag7B5QE3/0hciBVCm9
yoc8dpIuLmgGXYxbUvRElNMrbXwYVQEMoqilZ86O5esUhqlI0Uld19SEHq7LgGPFyZzym7uJr9+l
qVjQvgMT4kNiGPO2+QM3RBVemO757U2myXrV1hhdiQO77KTrAo8WvV882plvPyZLk4cm32T/Kdi+
CY2MWEOFpZirtIHLt8QnnJcjNRzWrrYFILaogrzvJ8hkC5oyMg1aq2cphuCib0OR9rtP8Ha9Tkk4
oqvwnPHdHaTBxOlKJ12g0NcU6ct42kZEF6JdIbnuQ1eLiXb2rwyUyc+aCrPMr0zwF9PGNMyE0toD
scdnTgQ33q2suvYXyH1RRm5u/YMG5vjyn211BniyrBERBg2r0EKiQJnB8CdonT7eYEA9GkpOPOSr
BuoBTqEYax2WlwuTSAc8FCQi4O7b7P/NALjMiR8wHPTSC0ek+UdWk2nOxbsVzEsEIrIMmmiEycKP
aNvpum2atKl0ItWk99TMslppNOqBkzkbE5oi9y2vyyBcGQVsp3xzoDq8eXTemhTJPhJs+erdqv+y
QwomyGixxmLJKq0cuktfJGH3TJRg5W5JMvUPW2EbVWS/5f3XLrwdK+2bwsVkf6/PK9hkJLpxMEOC
S4BRklZYPsPQ5U6oZttkP9yUXvr+4m7XTa5JvEZPhf4wPPy6fWGc1sxLbokTM2vgWCiXejLC7uIn
Vpo63UKqh2/rKsU7dzVny1D05TB+aUN5p/81rIEK+iZu9cxxw0ps3j8pWpOpKlpwfPhW+MrSO+Wv
dZW94Ekevy2PYpxVpjfxtnXqfFOVGftZDCJH/UHa+Q+pEmUv3od8lFEFevmP5RB9qci8pgNNCPl1
kcauQD81aE4KZdAQyczuUTW6nphOuHac+23QmcBs6feZj6tPgC6NFSjmyI0gY4AI8/P0aMEmwDdJ
GLmpgGhFGPC/9u9aegOEj/hNxeBf4Z7XafvWdN+45pOpdP6TvpmzeR4OxXGikxjySyeJHHIt9whd
Fopv2N1yARnJxUiptHzjVcE4HLxSRJf1gSclvWhEeXSHth664TDomDYV1wArRpPpyx3o/QjGvduZ
BI+WsNftIKdua/GazsWt3qHBq6uGrndVKGqHDprqyZzJscovYjHUlrD9UjhnH/MYmI4nfhTE12Cg
qH/QarjBVYdN4PTe+LVNavRUb1ENUhl3JOifk1RbS1pCvH6kzoPCCmq914lW1ALVBEhdbAyBCoU0
ltWSo34AAfJMgWld8INMABOw2SfqVJsjeOQCFophAnAgWKyoR4JG5aCGJnx11ffVY3f9LpjYwOqV
JSC5OHoTPwaAhCYT6DROAtCu5hZlxAzM+JfgmLG5h/ggbdfYH2X7KCirovTyIjiHy9opo4/b2X/H
J0RKk3EjHqU7fDTr+DVQHqR/22G8qUU8N+mqtkNJWUwcZ2rwrMa7kVI1FwlWQmO4Jv0z1WXvFXBC
uT5cQUDktwI2mQptBWhZvXv72D+e6PWciEkxkIkqiVNpfVXpCjKBk6TlL6mIzFSj4+ZZXmF2/+AD
cNIPg7Pd/ifp3nifq2HDz1Ta9HE6G35hdbP4AHN2W9B3uU9gg/hL7kKOYaF0BEvy75VlwVp9a1qZ
8Mhf94642VhsDkH9UwT5oZ5+8t1QsC4ziA/KbVOdeisEq2GFJnKnRk9C8C6S1C1iw1GbX6+O8/p9
fWc/k1iwGAEirQkaqITTlXsTcrITdBnP2Nh61UfGw4DEadgZHNSs4+PA8r/2JB3umTMuTjKnxW9c
56kqjMMZwK66iBFQ8VkEwyrXL+Q2X2Yv3aFZl62/hB8v/8RFtDDIdcds9wEKJD7AZb6UpMO4QjBV
ZYE86SBiE3SFfjPUmo8HWOv5wLiSJCRLXjwJ38HodjignY3YAbTtCpS7w3/E89y1RUUxzYTK7Km6
8l7VTI0cLc0tGPYfDVescRvdq3seACt2+mTj+Sm0Yjwx/tgDo/xWQk63TWXBZgRc53aWO8Wws/ql
adkUdq8kAEEeTus9jiR8gw/mTMFr3Obgm2/Iqs086RyfY7ZGg43nnDVQe81zgvJ5w4SHBGjFkiSY
pV1c3E4T12oncW6+kJrnCFjPRix+be1SMJBaZgKq2inShFIBZQ8+UrLb4b3x4mw12LCLKNReG5gE
+JJar8HWXNtORslFMqT9kSpEtMjX4YxKQJI+wTIc6xxQl+SdvF++gbAiC0Tm+TQpKxjGjn4snWxa
nrGhisycb4u8MDXZzaxPx8B0ZxR1IvWMAqHqIzzuUmGpv5DZL6zBvakuvv+5irByBwLpBhSY3UCJ
3EOrs1QeieaeGUdfNyfeIR7N/cAAl9Ee9n52ZKqgocpv1Ijdxc9wZUjjgx7ztESRcl6j3jxBzHok
TQ6AKBKs0hGpTKbQzE8jxrbzjIEj58DBfkSrdHha5asgVr4SS4cIf2QpQMEwXku0SsPC0b30zrNS
jLJxIxa3V9HonwuWCbDXBiHQN40k+dvyimWaSfiY9Wrkmiw8nu+lim96o07iPXqIiKHl6xBLG+DL
Rhu/XgcRE2vXuluG5BbGYMeLuVnZoOu2uwXGyRWyCZu3eYxiXewqSInSN7l2F+j6GQ4IYU7jwXiK
es5EHogqL8AqcNtK5EYPj/nU9N+pOdqZvcIltVdutJkMWetfZwcgEkSCT6jUZV9hmJ2LAsJE3/ZW
2b1S95bZoTMcI6T6JiGwfZi0edZ+NCn+7pmYFVgHJi874oy//cMOUvFrUkBTovhwbXuCFpG6kpMd
NajtdIcLtVdqPfOVK0V/GQ+8rG5DNmXUynUhwLC+0Ll5smcOuriSgDdq5XsqbTLNXX4aEsPzknPY
GA5sgBYzLSMKp0u2iJHg1z3DAsipf0wLLoaRcxjHpHL0kywwhRUiMEfEk+fdKLgTevFaFqahOgJj
vEcmLT9k5YHfbtpMTe23i4yWKJ0W6cH640ZSSkyyaljGQpQs5kW+Nkaeqm9ujefqwCdhoc4TQRXW
Pfn67kVJV3OMXABDAftgyltx7tzd6+bA8odC8EVaulqUxPeHK0AaffVmQFQ5zM6WgoMh66LH9ege
RpjPTpaSUWQz/pok9yq9nV7e5QOFqUc7FP0B8+d3IdUYt5gU5d3T84y6TSFihJ/16xiP7eHHx7Kb
bUZK/hKl7puMoguixS3ZrKYPC+jtRR/TCM03juMo7T69MhH0/ZQQI7UyTm0e3uWnaPV4LVPzVMkN
CwBhm5szjQlV5Wg3zi1WZnhXkuA7Za5g2rv9fYHNajMJa9VmkrtIxGaQpuyORh+lAASyZ6AJ1E5N
XkwIfsyuxoPiBkbfeIhycmEJkGXIzMUr3bujQxv6ySOrfrLAjT8F0rUJS4CslNS7ribo/d42YG0/
1cFiXh4ygAvdoeuN9BDmmjTcc6iPYxtUF5jjogQKBGf0HgzcLUDWLss7a/viFqGGP4UUjNjLS5Yg
W4ZdMAn8bqECQLPlOa9hNDYiPA8FC4p60ijhpO9oiZkrsgjTmgUM18Y3clrxt1UcVfIVCZ8ouQaM
nEMhkqSVJrkmGXZb5pNrqFzAhNYSpv80poGHI87aI6JY6C5wTBk8dviCzR0m3WVxi/6Mg4pKlDrK
ZFKRF9qHLO6j6CN1GPwavtetOrQiaG0uRkPkh1QXSAHg3e84aeb5xcu1au+5rjEL4yInZ42JftjM
1AdryMORyzyIkQvFjoFzOogI69XyMpwsutiitZc/nQlM61/VopKVHybFWqalXz86vU5i3W7sndul
KzvghSOfywCWN/OcXA+4cC1wafSqQGfIJK9S5sLWphGnOfhYvgvT+gHsq529nAWAApeWFE/42tSG
P/V52Rzfv8j884TQP0xVRImZBkeib6CEvVUbrof9vsjIdWdtfD79NBsg7hWJprzZ4Vuxj6Y8JcM8
5fovqurX9RPWwqzc5gLTIiU8zGUX0PRpyQfDR/xBR2uJEXxMCYJ8z+qPSExaIO9OCTRe/lNzlvRa
2nkwmusqCnF6C3HKTNt2gCK6cd5htKgpqtvSHhuS2pij9ozHfMnBDlfxpAqJfnrkdXYLsoBYtuRA
R6ZZgQ9dTCfJga8AyHuvGS0ifTA0sqNm+FUIf9e6+F5z8QZ9xUh/7CQaUlJAFXiKsICNgUPqKB0e
qNtoY3+pa/Y9daLNDfW08FOPLIIA6KJKRet09JVIePrmU2uouO18nQlhVHTYDKV8pJMZ0TaSjcP7
r/W5a4DiCZRrRX4U1ysU7xIeutJsq6oz57+G8xyuFbFQ6fuHsci706Y9ump19Rx8OAji03/ufwoI
dyyMyqKFQcBU0ePrVFwipqhyV6tUcNoYpw7yQuDvSH/A05HkbYFO6YnSRQrfjIqB/2xU2tRTcT7n
g3ISxgA71UaZ+2+aN+UTLyXFY+r4przp9Dy2PxVzULRm00ynetqE9VKIZDPmfnKY7dpGPx2u9xBt
mmTFAigXPJ7V64byvS/u627W2yjvJONViuTW9LeXoV3Pt58JWEjPNH7V5kcNNILdbh5LKQ01b7lQ
8eYbjNPdX76jLHroC0H6VnLRjrhdQLJT8UBdNZyy9FCIg/qqNNq9bEgyYPmyXf0ARMtPr/9+DZYG
mIwFvP3I7OUz5HAbMTXA5Jt5YayudWumK8JVm/JJgrWqtBShKvwQpCiH2rVy9rO7Z6nsta8jOWsj
b6aHc9Hi/9XOgU8jRacdBOZ0zRtVO1DVXgSORVJcRATlCYV3+/TuDU0RLJGztVLTkHwl7J1DTQOB
ENmHax80WZXMBEWZo3+L24GWatI9FH4YSR6IcHvCGp6a9yNNZXIERqs8Xi8KCFuGL8hJe1gJFEG8
CxQhyxLKlmUMvG6BWKcrdy/tyHYIFLWYfio2aqyKczSZQ1dvzHUHc3ntCpbpaKSPA5o7i9yHhUZm
FM4OKmL7FDGIzHC2v/Hh1CW/oKozaMj/dl6A+E++2YfiHX3xa0Rk3GbPhSrtLE0tltl3w5bukKCj
eM/psStMjTRZcy43EzHAZ5hfd5T7YpaJ2AFgDo+8r4Rw0BdcEpISWLM7Lh4Ner46Q+P/gp0OCTmc
Of3CYG5aXPdJSHF74zJabOJIRpcDyVcJm0/aIHPICkidxBYXb/XSy19NoftV4sPMusDTRXUdgHcG
6ZTPFoOJkUC4vA4pQsl/JrhXYJDnRS6N2lgfjnh2vZ12gIOXuWNgpVXDiTWcNuoIab/XeE4jwEiu
p1/yHk9AVqLJWv0D8pFwlckc7y1ZNpT8aFikGUcCdm7wZJ8Nhs4G6sXt9h+9XbtNdOnPts3NdIiu
Ap/YiwnO8cPBc0tjz06XokLCh/08n88Xif1o90l2bjaS/7g76ETmIn7FbjcUnIdPXE9xU82xtJFt
NCQr/NzyXdMjFbpKQzpdEPiKrwUt2tgQyz36ThIesVMVlxEtGNofhknxikTlxgzue+89MsinZ8Np
kfZ9a9RBIegO+jK3n/PRqCy7R2T+RvPKUMC28t7ss2hJYyGQClsbLrO9U9YaYg1Mnz233zocaQag
wMFDt66s3O8eoIaIFlyn7QjePJioXOz3RN5jODeEzwlZw2m+vye4bN0bBr4DuFDuznVbl5284d0N
+3TRkq2WI3nzbClryrsGLYGFwjLX1CKVOc2OFLsHwUaYOEBNVwIEDYQVWU/NbN+hRutth3Y22XMq
nhMURHcWGYjRQEtbAOcrzZJUvWZPrNla6j8rhsjS1lG6Kezdw1HMP8JcPma5bHwOlYuitgpX7Hli
Aq3r3hoNrwqeVXwD5+65DVCP+CLWVNTRCjedCIHIeCvSMSil+1HLK9kANQ2Oa0vQYEq5LJXcSlAN
frVJokeUcIeKOvoOyWlKQpXhl3fEHt+Uc7i0PFvMW8X+fnumEYyLsqj5sDkKpxFt5+NXy4Tv2B/e
oUAwrL0J5iasTYDzL0fbDubpMDsF6jlgCycH0Ga4O9oh8UC7Sd6N+dQTomIgiZMx0W8k4BQp+Jmo
leoTMq6735FNDeAgGvk2AQ/zpr8L9VlfHKZ5WKoXje05/P3c+gv1ydpkAv1DJ8ZCyjl7+10K01E8
JHLsXVESlTZRRU90cSSHmJc5jqQ/ajJ8aTcir4cCNmRwRbmB+LCKFqfuVcqCZz+0rvWO1XF+xYGF
aX9pHuNmbKhTe1zCUdCt6CznguabswaoajpMasgHK200j0NtSG2+RLs7iZFU/YNWGhojTVKu71QJ
q9iOGoPHidLIxyTGLq7zy9AdlQXfjAK9i77PzzI0EfR7NPubBb8n6gN8H/bjKHCPoynWQXB7nnaK
KQUCseMxXNuCOChyrlJeCZV1vihH+zK/F92PXq7kuO7Am9XKT/t6vhEhctsFsxxMLnFObSeh2HOu
IGTUrgLl5g0iU+5/wQ8VJV/0cyMBdoMQIz1859bDSTwEI4i9ArRDk60reDsXSvWqnb3qS8wBEnCy
nmo0XxS5SHcs5LDa2HT+XV3E4r4tYE/9XFwdoIX9Ygb/Aumvepwl+uFHGLpFly/y0pxqQkpCYNkM
s+c1SjY5/C+lBIjEMLN1nrQRt5Pog3/pGHRg5rtAwi8Cw8vIhzTSn0fGlnZzX3t3Bos6XKr2lgrn
E3HwDL/owI+liMSHSUjsSGhNLW/G1LUXdqzB3w1MHYTlLNUa9LV7QWAJ/ZI08KoErZDYbhnR7ChU
8Dt5IIuyVlMD6xK03coHP8vHobqHxnyRJp0Dbr7CcE3Y5/QXNVJrtmk2Vxo/EWEjodYg1crXfoM1
NVcFYwzdsv5L+mh7YIINjF/kPhfBEzxLNVwX8lsoZP9W3jAlrgxjtM5TkIfdrXrxSPDwQND8F9IK
EsPTtyJ87N7I+RmaOlPUl98aPvCobdOTunVHfyDskXGKpVJi+QJPAV7tC0f1cjqjuw5HZmXHae1x
s4dxdhOc/hr3s7tyB8uZfrS5nWi0P0Nuxf76wKf+GtdKetkMFmKUsx9ib79HLGd3pUpdrCbiGIIe
TC/4effGhJqHaydz7uSC6CpJMVlUhFzOLtbYIwDFYZ26Wq2nS+8v/mHMJ5Dp8IErQEHq+BX6UT8A
TbR0/J8LwSeqX19GpazlKl3LgzGvxgntsR2t4DSH4VhjjoehleRPMVYYTSEHQ9EPvHalAQ6zAOma
L+Srk2iWVEA7sZlc/G2A8EC2DYyKBoUomEcfFDhHmB+qCrsrhGmQWf9sk1iJYddjRbFx0OGuDU8x
tFfnRTGlImmIJ910bff6IZi4ule9E7mWXBH9qhGLh5SDyfK4gUqVAf9fAgXFajT7OhIhpe71Megg
gJrkX1uyMmDUhohr7bbjWZnXlpJzI0Ny1vPXLAs7bzL5VitQjTl+qBeRAaniWuD1BOg12VH9W27t
4wzYKx4iyZSeMSSgH4seOVaJ7aEsh5nhHqM4D3xCkDe1l2oOvQrLKDJ0a2aXdoGntdDoeAkYQGyL
oT3vG31Y2z5vnMEUCJKJEtuEXYiCh+OzxDMnc3Oaav5Edhswi5A/FSFkLc4XSlwOOnWAe8NMVwSI
d7QlAtjtUbLptkhKtP89G0WEq8RfuotjhDK+ZjEh0bcKVVwMkke50HbyiLUptNIDX1+I62pUIA/j
tmZf9MgFUb1iRel4+AGHHJmqUabaWxKgC9wpHq5Hrn4YvpPdvhMBiKjXcOyDaax/uGZm1lJ6GYc5
zsGVfEiJXNKadCAjkWSWM5ixZFo0hZUoqCHFlyN5VdkG1A6s8R+YQh4u9w1j3a2NyDVCPUcdVe9+
5vcGTo0Ev6WPBIcRez9L6Etm4HV0RUKwR5lc/r50sXKYQn+uL871rfAhOx323yymo9t0cxBXGYpu
Z6yGtzD77+XGgcX+ue39RYQsnw4hOrJxDtP2I46wOt2JMc3pziA8xkEi9R85LPzXswfPXWxzC/VI
snrFoJm6VCE1Of9Ll9GIX6ZNVoVdSyucJgMdIv3BmrqRpNWDTuwXUy+o2bcTRSv6d7/uSdWtD7y1
lPZbupeSQPSA4nYDKDMaNCchFBbHvNLw5SyaphemmCtrSnYeU9v6og/BmfgV1sFZWg8k8kNstOWI
2G2mBqq1npCQpHvCp7I5fqyino+OVrvaOVMy3sncp9rx1bAjTXd0qdinB64odtstx10pDyZlPbEd
pB0eoB0Xadew60eLBED9gm1SBfLLuYCnHNFouKVO1xpQN9x7Fho2UkL6x+92GJ7MAi2kFnz4xe2U
C7rKrC/gi13OKeHYtVLNy0TGitSrEHnaDJVX7Yaus8zJAgHTFTSaDKQ5PdTHt/FD0r5i+wa7VuFl
dwIwKeGfEBAEJR81Zx93FP5Ac6CEsd6RVWCAnRdrgpUhUIbir3J0k3h6dNSXCIg9ydn5ZKohf3Xz
qjPTFvQUsDD1j+cdOR6IEIn31OkSAffpQ7Pp9D9idmIYAQbRkJCNL8FmAmGIoAp+N5sWCnlyaEd6
HbG3nr5btqCuS3gVVmwkYU8Q9C4DpQxyGlNdN0B1OK0N7zJihoQrmdtueoyReQ5ty023jYdxvD1W
wH0PplUN11RdhCRtKyOZkwdlU+ZTvicIJPguaugl3tWwXUN6uI8NUuGMiozEGs2XsogRA9xpAXel
OgN2xwGoc0jGYwy2Of379874YZDYtI5lJnDrh8FYFGjEYvHXL6jNS0X3JbayUN3+UMF618vrv+Do
qzXiPrxChoS+DXYHtrVaDiIgk21NoQZWz2nO0R/04h66+n3+bSXphJBLIKCy5iEUKtyaWED2aZHj
NNt5p5pPggYrA3Ko/1s0177kRWOYclIE8+1jFBRBJ8S73kgi+VsAMXwfeMkNWtRMTMXa6RmWRs0v
WHfFtmazq8YReMl3IwFSv9b/vSYq4AdC195v18eO2ujzgxuGl5ljCTzrC7M6bEiaHyksaIukDEAp
IF2QnRP/3a4BOOemye406RoIB1xdR42x//neBQrT+Dz8l0Zxe1dttKWk5nohAZDz8MhXFfZQHmdw
d6+0w2m5ab+ti3l9+uVVxpxkVplqWGlM01i3cYfGpAGnJCFt5PVau+O44A9w70h9xmQnDCta6iAl
m+Zj6xUbP6h+v6BwQz2LfR1dJKAyrW5ZvlKECRyfOEE6zhUx5Wat+yPqq/wy9xqGzxXZOhkil+7U
I4bxwu6j79I4WKqvHC0IEGlFyfwrq0D9T2oiFKH5iBQiyBh8Pie0dBvPSXCQgKW6+afxtnmHNa4I
8KBlSUxe+FQZT8bVX8LBcsnBxFFWH2RZWkNll/N3o0zQxWrNwOISqIWhh3OoLShuEOX7/6AAcRpj
jOtHsKEusWd/SxXNuIBksDGYrSYxTpNOXzVQkPDR4Ep5kRWS54RlCQP+q0VIEa6WtmE+aKmr0nIt
GH39FcnksyJ8v46huEWQMB0dk9xvcPT7+Rg7YmpAvite1JUx0mY2Z5s6VocbrhToDkP2iARhy3b8
yAm17tzPgk06hQewQTi777QzUKnErDykPzQXOEYqVhSrMH7m71IkkEItXjLKsWs01vn3hau7teDt
/TtxsfMftDwUEfAoCRzSMRIKICLAAfTHEcyNgmQSPHcbFXKN6sb3SvaVXhkixyO6d5W55+Hrf+c0
F9P0ObotFjRBLkffy3n7akGqaCTT6Puydv0XZHPUHOMfSmWub7+ND0Yms13P/a2t7y47tO9GgD8d
+IFAxuT9BWa5lnK0y/9RTQDgxXE7tQhvQzIPCteKRcIs5cOIIRAbYzva2MPYRmsXmgfz5qA8IAV6
8CPyaj2JBRX7yGClkEAPmUHThKNCHnE1L82K3rfmzrICDV/HOdDquu+y5aERoVwJkF7ZHm5ikX7V
VlPAt5g+mrTiuJU7gAPAhPIJfDpv9wRrzBlRDL56bjvDNMip/lfrZwfom8cyarEb2nUOucW4g4wA
eI6Rmn2Bh5w066ZbtgmHZNHETPNJvjpEo+EqdOQa/B670R5PIorLlzNc/FSLZVPpGqp4kVScZ+Ta
/LxYg9WO8qzdNiSnf1agdYKTShSOjqA4ChuzLRv2Na0zQXkeyw3qE2wP1deiQf4YTdLRB9vUQhPX
r80nPcpNVWxigAOVOJ3gbwwGlFCSvmbM9nAMcbVs0uxCGChlmJWhRKp6GNDEulRZtbkWAEZgj0t2
cQDysCBUj3f5tS4cPV80H4Vn2EOu2GY8A/uqmBiy5kNQydWVHQtRVNhx22s96QKAFoO2G21wmLNB
FSDCm+GjobrN3GByt552trhkpAJtdf9e7QJvLaHNqasxjZNIpF7rSPWxj2UUeFRyiUHm8xEpui7Q
teeMKtYoG4OMAmuO/yRrJtFAkIb1anmnN2lgSZaEJj0LsKdMSwAu8T3h+ixuah3MKCEU8kls4So+
E1A6KL2dG8eRRRlPozkZ4uYsN8WBKzQi/Bf0tcdJqYSh1bLPn+cTqvPIBUpq1NPaLCa0FFzbziQp
GTGJ2C9rMaRusLpOwn2zG0R/JYgnqOFYzF7YI+wpalz4GT8zYtNycrioW1/iys4fMD1c3RcXm8Lj
rCqQyq+HdhdRRzJdJrfThPIsA6FrqDP1qubFoXG7WlyNrWTIBfZC7prLONIdnC8QQ25CnlfARXm4
qvR5VvBVTxDgoOgVQWAYIh/zMyis2Q+IYNEf1LJBqD4Ba8OkaZlZ8HIrO6uWcl1zADtlo6gMKtRE
aRn2fUOkAuEJJBWQh1ttBqezKkUm+xR89DysT1f4CqRDZAOPbEeGyGlCPtIWx8BTXh1iFMalEgh5
KXEHXhMaFUfuKs1CSbZsb/t0PHMQU6h4wGpEqtfqMZas4RnkoISmr9r3t7MwpkSDGptbhgAscRqx
yyI+DTRqS2wnhbDU8vBh9nO4OhTozlqLNz7jCabtixzgf8r0/wY0Miz6tNRswT271THdCBj7mBoC
gCYAbU/h7wJ5YaFt/U61woRFaIrFMMvTmuKy0FE4sCkAJskIq8zdKH6A5rg2QmFlceAssj3pbZ28
pH5cd+N2YZMseLXyQWRlovLgqIWHLSGL1MVOMah+sDxwQx2YYdtMJ4k0rcR4bvs+bMa3p1vd0xfz
CjCDtZv7U4YdrZvQ9T5jrFFqTKd7fJcRiTEfq4bQFSOYR9lW8u6lNzxpv7FNxdUiCD9Dbsav/zNe
ctx2P/ysuTG7EhvUZt3gfi1F+Uodr4n8RNaK8gAnmiUTa8ksESnqVnA3P1HRxdccWkmZx9r98TXC
7hYjo2X7zp8AMQl/eWlysGXPjLufCfOsw72O4fDOQ+7+qU8GYNyCMq4+yTemfeRF5aURPGoZGYIl
lgMRxDMHf1wTEB2cYUe53V3qBn8SpCynsxwOBQyJMVDIfxAxTksYa/9FK9MNCSjpzGWvT3rNzVgm
ZoUscH+XQKYC/7X9X93A+9Fg8rbLhFmXr4nzXu1WAYax8sP7fZF2vqslivYhslTnnB1vEZIZAswb
/GBj40H/ujLRMtmCWxN/EoFDhlaOAR/2vTYZTVMb23KcrFukOzQt8dKL7KvQlaCnN6rABieGl3+E
Ghs5aqfXB+lDwfE6Wz3XFFb2nkJNlgk9I29X3O7WmfFXxHuVSQ86HKtwgOfabVZ0ZUg1gBaNKAFq
ztsILDGIxU1PraeuQcT3/Wz7oqeATPpy/CBjZLhFefNdr+5P9RGYpcRZVDyuAjmAJbRD/sMcKHyS
sg2VdA0itFkLuZlZgF+mXTXAxwvzQ4co1dOUgGpyJ3znR5tKQsQp3jwxEEUasy15dvIfoDwTobVJ
Lv3kysHIZJxad62SHNavilZ5MpyJkaLmgsrJ1vc0f076zjTitGLFexnmHNoGcf5opp5RC4l42SuR
Ash7PUgErmOCCuiQr1NrYvlOODVSC8btR08DpI3nKYe+N4yHg5gcuyXkBCmWRmCpC25FR1DFok6+
AeC9OA8xgmVOBuc37xkBoCzmh3bAPseFDl/5/N3cRP4VnYy7bntk7lrVWP3+PKDoBG3SxbcYlMHI
1fbF4xLpRc+OyB669uMPcQw+7Ah0BGe+mEiJd4jtdHj+Gxy95a2HFeci5OwqI3wF78/+YVjgQxE6
blcN9tTBamlNfMdgxws5qfZD/IDkAePrEsbrapfDucZji1vqVLdI0QNUgaoePZf9V87zLjwo/zYc
Veg/TNIqQSSgCy8OqKL6MBguyTLO3+NBPmTqeGCSBP+0NLYF8pwzUxuJ4qTy83/iQT63xD4ceh6x
IrvEGJM4zzZL9q+572zN9akTeZx0o+HaJg70P2S8MErn/J9uLAI9yDjZYnUKvswnDgBZG9q8nlbM
iFpIagf6T1goIasVh00VwjeaZ48pGZceB/wRCCBN7OZpy0/zINaHZJdpKC6kf/n7Fh1O0ChEkDyR
q5FtfJPeNFcrRlYHq3n51TjX7Ni01DPnhHkhIjHExKvApD3wQExyD8eH10u/QjueRqJ8xCZklVwH
zSApfnWEj6AQll0AYbRVcjS8/5rQVdsXsUVSBbB1jiwKVUT6N+Z0wDquBp0LcWvjwf2dsFmQnwPM
q4GgRvouVr8XKuBt10tQMvZ15UvAvij1EdgaB3seso1u1dt66kbAZfGAVq7z4V8Fz00dQEJomldY
6GVOd3qF4gqHnQze95Z2x9UBMcSmUFPEDefCckw+ja/UPM+ffwY6Wid6N0DeQPkqMBbv5yqQNvu+
eci7VnWPDifEvfI/q+hytMQckuwYAIm7VfUpKUur1IHT0mvLjEW3qrci2LPnwqx+Q79eULgtfv52
JmULYRKQP1b3SVnHkg6HE1dfhJ1J24NrBtuT4KMi+tvLyiv78/uuCW8vHRMuZ8CaAoXXhSCmc2iu
pwbyfwKqPfnR+I46+Xv1rO5sL1T5IKqXXLOoWONK7N5A4yNn+b6JUSdQfT1gVFEDZ9A3wX3WssPY
6fiaXNdPcGjF7l3nCRYHd8Z4zWjPKQ+e7BL/DYB2/AGHs+78JEVrZMdDee1ErVm3AAxrGhHIN7xJ
Ej/23L08mp1jXbIHt9baYKpAh9t0pL7Rhx2Sgaj3lxT/WHHEzjzagjmGpbaCq+Kun24oA0ZEsYLr
actkzVmmml977Jyd8oyUca2UySnTHP+ZckI9jRFpjVjT3Lh+9Ptt5A1363lafts/9nozbif+ct+L
2962BI+txy6C+pTp1Tjh/ygHvfU2f+N28FN72SdOzg/QvqgTzYvm+E59G2HnrS2URGoBEbdf5M1A
N876lzp4emoD6MjwYkHriy0s6KlQVAOr+OtKXR7pAYrJVxOELZn6FtMvVYHu6gQxD1X/9VDuu871
Woq+YO9FiMwLtgMK3s0Cvdgzx4sXg6KEohJl7MWW6dPF+WsfapuIsufDKS6aC6jIkEbZJfdatd59
lkyEcRwY2PeHMFTPAoKEKYEQj+ic0bvZ4dWcErk8bHGl6YMKoNXcg3RmsecGxgwSmcsjsT2+Ey1O
Snm0tWA0iYjF6n/oRWL/US9HKZVF8e0YjjLAFoeEYdKjPsTFiPzPQb9hdU+N7Anpn2NKXosfIltv
BKByKlO16ES1phbwdF4l36Gby4ouMShlCbIVRdLRtPxKZ/HG2+rkVuDk5qtjZFzl2IIa0xQTEvS+
h+FdJqawF49j+9jtua7olpxOSN7r1d8GiDbDskVU9ExZGSEbpuvXB8EPW/kn0p4Y2m2qQy2FgQ5h
M/NGW29WVsvLnls3syPlsQsqRoVAb3yhD1k/dCR117ooZDqO49wtGoEagGoJsMvACJRt4qQTQ+FA
jPOb9xuletgZcOWO62Aniqzdne1HJJJVqndsbY48jUeK3LdSuLofuCTjhIBJ5BAKMcptTiTwg2TN
fpZeusjo1X6Kx4AMdW4WY/SFOKR6rCG6p9hI+Ou6DqeDMsRVF6TLL2i9oP2cRF6ly8Rw6Eb+jXMY
x+yUt3bzD61UF1jiXt34oenAmTQbr/rbWbiW2TycCBPeN7xJkmNVdVfkGYAqoeU1wdGZDGkylPBh
lt0oAfLjF/IzpiqIEx4TUX5AmXcMh1wLYtX6b6YNWeeI15S0k3+bNcikWHwTf4mLfLJv+W2TSpon
uQUhcrpgqfDYUfHSzxNte8stfYmjC90JXA83O5KGv4BYWlgtzd1aJexBpBw7cVRMjXnxu7bRwtOC
4ZmWGqItT89FHyrqQu2F6LHkxfcEfcOLz8SyYBgAO2Pg2T3x78GbxMjEDFW7DrxD75lhVxcS546S
XlaAQ83f2ImwCn7clRwZjohX1uq6h4pEnAObN+QN/Mmyc2pZI1OCFGUWIfTz6r2gPFwnB7do88H4
mmWTJ/1+iugnomrbYTyeaGtQZ2/ko8g0SpKXjJteR19bPEpoUxyT8sjVYTgf9QOT/TTYWs9RG+sp
hOqMV+LcvMHgINlTUGhhVA2MTGG4QZoTeSlDZ73HMgElqep67H8vqzsoeZ4TpCpx8DeN9+3jT5f6
jWsRmk0YwyX5zIS2Zn17L4/NF5yM3s9a5K4AdCRTpgxVx6X5BEafzW2Iq6yOPwUu/ShByb0i7pXG
exWSJ1LLPZyJPYNy9EmoCngVYcXzescGdwP3LLdTkOxsEm6JMh/ZMPhg00QoHCDchXYVgdlxBjjH
Gvr3s5yspmo4Sv0xoWgFJcGnGJuzzDy3Fhd5MT3zWJN+Bn548FS/5btmc+NyBY0YSvsBhGSk1zm2
swnEa0JB0VwgGf+Z+tCc0no1e7K2vP7N5sShXebGvmZDJKaLRf3rsAci6S66GnNXnLr3vnolilMU
ICRvkuB9z/ZvT/X24Fvup/Wqepa7JPhR7lQQQkbdbr1TR330oinjTYAdvwchPQo0bgUyzGLbNv/4
ZZnnWoaNpnDGYFK1vQ/zmY2ilgvb5I93geZMhMxjIojIbxgSCzNE/pZfUBxyXGN6NMG+GCaYyL1c
d7aJ9eYiDX0UMIqxKfus1+cI6MPZ3o2Xqjq/La0FkKu4ACRHsM7K+KiPTZATpBsckto18pybJpxY
HjWZbSbl5F1kI8t/H7Od8cJlhNJeOxb1cMFwxwwgjp0aoCy7ISSuY+S91BBmEWJlBpYyq/yBWINz
Dd7tKrwHEt8BDM4CDQTzj3XzAEH20r4/yVHGvi6WTHhFPs3a8vwaGXU36mLeVlwss/Hi/QOY3nyB
aN10pTuQwNaPEXSfAZvSzjEUAqej7PIpJlT7h0ja2PsyLq3HNHEjg0U1XuoJRfoEJk2v8im/R9O3
vK2Rygv/3HOsWTNtU7NlWkcolsABhrsJqu3rhQwtL8TZ8Tre+LSlM8n1hdhvWMc9C9OJoYnQVTiX
lwqsJake58RtkDLKozFmomRJDw22U49OBEAn4/pwsrUxmdi6Z+umRsmaXP/pltAgvuQ4NoF6KKx+
1Ljc8WRIEuUFuiRmdOjyFI6RfgFPoO6AbVBttQNBiMEj5L9ydJcBerqrr7QhqLjqwcaQCirtOEZx
PdaSCr93/sNTyDrYVtPVCyeuI5QLVY+4WzwKKLqqBFDyz8ef6hSh952yWOgV92xV65iXdy5Agzbm
+OLy1byUkjL5vUmwp+MdkgiQ3succMvSxnzU0xmVfNoYcnpsxtjsC9msv0KJxFBqMv3JapYjJiNe
qkO/flNgK9eYEEEDOBUiTRPieoX2zMAhRhK9QYRKcLrPWMNHh9hBQv5TYcp7IbvkVb/MiSygramD
rQJCDeP/mrQkGi7VOiG82sfwhf/8UpR4+uqgWItKpX31RQ3yZrbEPEcpyW4rUkcjLZEkKM6ZjCuy
/9V21Z6HCdZDO/m3BinraAH/38AkkvcUHjAWm3/xk/Wyxcr8KBl9mCtASdiGM7G7BkoOW1m4pfhi
wSF89rAv7VU9Y1ntQiq5ipqGE80AjJvmIxDpZXqAeNSOWBEZJFNDOrcH7PTpKWcNUhKRpnAhslMd
meCI3k+o+zoeaMAUkG3th4wm8XnsskCKq7sRShaV1ZBsyqTWkZdLVtzLCp0Ebsbrky/w18ALPoZF
2X4HxtDuMSvNj4BVnLwMuWt1ox0rPRpgn2tCRM6MYupXj/+juWTmpO8AdrA4IkB0RWIKNwUgJMqe
xOpLbWFV/DzJJDa2FfNzh3/l5zMv4oOlcSUPGBXsHiYwIO60BLKhOntg4SsSgXEFxTENDuf4JKth
ObT47fGf4FLwQwciRu+uE8C9K3eZILrxX9gPCMJ6dhEwIIY9ar5/1BVuJXTo26OgFpYbWYf94PjK
bmcU3cJBSFC2aDpwptneYSt+QjcmRn51co1Z/cj8NMMUvHIvNmJUuqfwCksF18vYG09czG621Zmz
jvoccVVmC64eKIFu7SeCvEHyGbF8cUBmDC0/DhkiLigmWHjQE2Ha47J7YFSbEgJa6MZVkax720mz
hGffHsalIJRQmCf5Wq3z9VdR8Yds10gWuZcKZuSZytJppthyGg3NxbCOVzzM8fl/M9Z80g8Ihy+z
1pf3dgFpAjlxsTz1LB3jBhUyfEZgUHKwhBGpIPu9iVHv+6XIusg/iVoGmwSFkIQ3tzMqvzyquZXy
vcUPidCOcxyI81onbLW4c0rHX4xgUnYvQyWR4t+1vuRdKcuX236js9g765VPbz+KeCsSoSQlT9Ql
QvAqOTO/wRgJB10cl9n0ccWfSQ8SMq5/Iu0mzkzKtXk99VMpbnewy7rhk74rQKm9hXy30tMb8lPo
CwW9OqaAKkIkOAyEkozAfVk1YxWqSxPJehpwdfcEqwkeaKkVmHM2bQUNAyUoPr4U5aWeZl5eJC3s
kP++LaSO/7oXPkMntzCI9grhKJDPAZQEX4KBrGO/0K6qMHqiBiVnuIyUZfVtna57hmOHxeG2pjT8
8RtuH/xXGc0R+x667WJG08apHiY4mQKEy/p0cdYZKZbSKCgdvlHA7ldsH+e7zd7h9iuZU9x+hO4J
Uxw+CnEgUvigdAkeLsx4piH4UowYT15vhP2LL256WT7jRYRoxZwPwmuWbFMTGfSMoKuE/JAQwEBQ
qteLnH98Vh/OE4ouxLnzBq6g3TugK8Eth5NkshSzSU0EnMN1qk1sKjkkNPvZWm5anO1v/Rc9VjPJ
g5skLhjOl5gzztqn9ebJyIo0KF0JA/W8yWHtzoTwTu7kteRmt7YqisGD9egVK1WwXLCifwWy8y58
xvW3I+CKrMxvhDWtMWkz02Gh4oOFNl9jZPBatSmuxU0yQB+Q2mo1uv/SSE2MOBSR4Qw/FSOWBTEe
WIi9QWA24eNnyYuGOg+Aml8jRDWbAKz84akUGhQRbNpHzL6SCA593wZ0OqTwVe9EXjJHBVyWPv4K
vPbD2/15IQ21ABgYGx6dyvzZPRN54dLJE/Cwjn1z1JkwCR2V+XNdoatfhtAc0rIMi0CKdFPSRabr
5Nrz34ElvVksFmUCiNiXSCsqKPxtPGbdjqnldq0u/uZuWkGS8jU8xhEU1DQIjvaot3K8TDOiQSxJ
5jX1T0uZg5kucfA5/2ONpwa0NCu+9j2oCrylcmTzuca6ev3i2B1P/XEwgS8etr7HNldZZtt1sZSK
dPn2vjRRHZ8NTWSP/HydyK+VnwiN11XjQiTR5LeiO4g/W2W3afufctgI/NhczuY6Bl+er8iqN57V
IsO9f9wJv/Gx/ijKbEkItihkF3GuFHi4Q3grgH+Xm7PCCIOh6ueNaLaRInitJat/gTE79QnMe+0z
RqjEjPq9GZwGRPXCKFB08bGFFeMg+6RBsSco0PQx3j5Cv1Z1nNmb9q2MmFBDQvH9IS7rOsR+a9VN
cIMgLBFE4XQIgwq7wZ5TLN4sJ/DVe3N72fcgmeTUDm2ZYpcmZ2/8xgMr49nXFSl3Ha87CIXNg+cQ
6bDcjbTtiSZlGaybWIJiMPVK+FCHrIsG9FBFto/vklrcCUDtY2xfoILmoj+HSibqgvyZKWWco4UT
oUX5IqzEVSuDl8+QuAm4Mls9vbwik0kbLC8TaUq0MXVG9YbiaD0F4P/7nv34m4f8k5ASoN5CG3Ri
LDx9VTcA5E6U648bkW2LdzUyrRSQTja0btcO3JP/VuOHCKt7PzW66QOjQYQ9J7U5gOyD3/EI0dft
6pP79cq7D52SIABb+uoQ77ALjlSEYxbuutNig5nf3j20Q0qNtklWmGlOkwDG+EoV2LOvpUm3rae8
82UVocPYZsONvWGteiJKX/o3c6/Dbl4d1g0D5XxgCVbDdjh5sBMtJQmEHiPm9nSrXqg4zQxP7C7E
sIag0JshyGWSe9iENOHuGssrEEoL/8ocvQhDTK8l6CanYceoRM83J0a7enKycy9An8/Id5ItTaIz
KKE66H1cl9N42jOxGBFQi5zrZh2nNHqiEVvWygbME56G2yoExPNUwkPPjT4O9rScAe2lYsFw56A4
9SpZzoaucBuTDljLzFuqs9BujIoF8lLgcim6r5E55uLNoKmQatsMjdcbkUmW1LB8BQ7H7UKW/42H
PdbxunqeJa/WQ0KnVsrbw7o8EC02NVc51nJUldy+kMKWbSa5AUUNOtCg4ZlBSwhwnRcXHt5U/LNt
2x8lsFzTFDfNmswh0yEsIdxqqKsoFNMP5biRDbBFMyXNQOsXLwXSVDOyFb6SKIpcVFYXFU+4HPDU
67sAQ5LxIBKvNYTSSTH1nKjPL7I2V9R36pVrba86z7ZJhU6jK11mbHVL5t6oMfz+tn4FYlIrNCAY
3gCOTy9eahYBvVf3qpg01ufThK3+/92rijPEHxdnHmyGE9VLrtuDdl0Jw6uETZeimCa5DKk9NFdZ
N7SRgYSwxGo2C6OwREoo57fCoaP5Oj1qcWXvxw42f5ta5WQudroOXCR7St28/dk5I9qY2Jo+dWFL
12PdTSjZLf3B2i/heOh4QvgGNVZhQFqsfejhj1UgFMpatK7s5Q9igDi+9Um99tduLQc64S2eS6yA
tVItD+aVwu5GsYpvnC6YRdHoG+IM861aslBYTx6+AxBdQPk+jQLqlc3fazXu/asS1bm4n6pLiA+1
JTouBFXEDBJDC1XMMONktuhtXgrpxc11bLTm2VRPepResVouCPBDA4IV7P9+i4DLbgUDShsOFs2E
BKWWlk5sLGNPDaH1hmu6+Kk2X4l5x5Oa2Fam+0+IBAx9pjXd9o4u/uMRKg7Q/06tZnhg0NwZcbhe
Dwh6Bbo6u+jd+a8DgETPGClJdhUpCd5I3MiMR/JL2eB7HLXUC2b10XkcpKcKOw+QzylMDtHVWVfk
hE/0hGxZ2Saqh1ni9V7byfG0KhbW4Eo21dwzS5LAyOWteZHtnfWIGF1kH87RDtD/ra7HmojC6Zt8
+h3H/zhxkGrz6JgVOkPOcmnPMeqvkJlhbbcUHXmfShmZHRx9GjTpM585LPnm05rGlznlsOEIGwK9
0Y6ScBnc8fxAXJ7A1dhlZZWMLaR2aUmR4EIOKZoAgekOeVDsz2h4izkpkrIvIyMMqqbGK4NJnvaX
kVwCEB1NwnPTXOsC5fb5DeRI95h3WgOihWEkLuali8S08Vw4EMay+eONe3OfRNBDBzd28RYrw80V
VdCNr0LBV0wUVwD9VwZC2isy3sZKhE2E94yMJd8IhZjUtFKzRbZ9HD/b3nRKXFjWqIT3WXqtKPZK
DzWDUG6gKwUgQfgaIGsfrR9NBxChkDdcmE4DRHVXCANGyirHW2pCu0XdWTZY6wPbhc/RMgiWuLZA
FCSbQwTjDaQRHB0QwkNDJxOp06XDN42KgeGkzBFgiDFcjKiWaTVE//sqgurFR1Tl3H5Yw9eMGFeV
5BIefRi00JMrJGof+HOOsjcznoGFzWUkI5pF4z/lzHEKdyTaXmAqjFRtDeiiuEr9uR4UCBoFtVI3
O9IpaSGSAxLvylWvKhP3+J3Pk8GOIvV6Vh0zwEpD5dXYiSAAJdu8ynpu7aSdzyfjhveQDIBLVIMv
XH1wWWJe6cnhx6D6sQn3YgqMGSbqwtuMhowW6LiU5PNzh13Vm+bse38Hm7rbD3YmHw/GOBdZ/Puh
j2LZA5cKHIWJecYZ5BOXGUnQmQHUCD5PobDPMr2I8KDui7puPsUYvw2fVW8XIOcdP4YF6OtOx51v
sTLNr6cVc//i0revOv6C8EVtH678xRXtYE7MTPbNjIdNk5WOXmejd+NCgrDi8C2MBucbXW9BVp9R
6EIie9wyp9PF/W1y5/vsQkhB6Gir5T0zQHKcCmXFUb2vdKmYuqtulrb/qL1UHVThvjRF+2364WEn
KRW27mhpG42TwpBtO7Bd99CXFsVgS/3EZhR3Uxqat4sJrZc/Foo8sWUbWPX95XVGHbhucOBXUOdv
rTXyRETthefbvP8xA7WmQskFyPrFT0E/QU4cvDFF8Qv0hrMIkK705bkXtif7DN23gej5u+LxSlVb
glovSqeySvvl/9+n4hLuSJt5xALcQvm3p27fuXur5BE+xOYyXovsJMfe52WLiBpj2Kp8F5o25xCt
JEhoTyAzQvwg7UP8TKzBtyhIP+eLAAJR1Zj9De2i8rwaGonMXNxmpQ1ZJY8KAiPPJCDd1pYmL7Xl
SeRPZEFoHtVewfpERXAg8VH8ZF6ET+tB1mP8Bb0SyMXCDnJPf87SKJHiV/78d3A2mQcFf+8OzqBb
TQoxOp8JOqkQMV1XYC9tRgGhoNtBx9i90t1yH3KThovrV2o3qh+VjdwvbtoCFx9p7PFaAsDGUjkd
FtSUYRcbORD4L0QgshwlwqyopjdFHC+UynXASjNCoqSYrP3+pwjM0nhSUVKSPa2CIN0FbWS8Aswu
rjHZjtdTNBxJqiKF3WJ/HFjAZTYbYEJiW9dM+GC3bqc+xnDdadqys2zUI85EDnAO62GPCuPx8+Ir
Hc+BuUGLnA14vnCZCoFTUQGRh49CMj0SqeSO8vIaUDe2QCoSbW6n/dB1wkl0ZCEhP4/xNlCfmLv2
aj0+xTV3PCbtAYKGsHBljkYqkL+/ctay7mjYJgZwfgjZSO3TP1Tqq3ffGZvB8eDOAT0rsU1wFlnJ
T31rW0OF9F6dQ0ClCTA/UqYaUos4OjJf/m4V/B4++Lm8GXWXwcDTcSqBPTAGQ5BCn0ENR9LTUktt
W4rcUxqpLiSSJMkjJrpgNgWfJs5jAHZoOC+Ti6MsI2MTZS4Yw4N8BrgyObYHGfTfUr5SUS0G5OKI
64UodEHrhaJy2kGr3TdudHuGYpu8kKiIx1EPmu+PPF3OCYpZH95M/Q26j3AjowEqeIZnpcVsj9vV
cUAe0foJs3FfP/P9m/B1Hy/PvG07TguBU0tiA5fJKBiyjUfsvZg6qchkJtz0cyIIDLW1g9M68Dqk
OT8v9bhnsrc9+JpkYglu3CUoujIqd5XDVUkqus7WOhbloSa6Y4KVK/Gery2B8bAU2uLorB2c8+9T
f4lDOW4sogcDzXAeGnt2UW1C1gZAqjFk/+awjlHi1pjLSp0oJ34hfEBXtCydExrH9VBqYR2WtYZ9
XuGGjEG8c+qugiWS+fT4ZEr22BhOH/MYl1oL87gKePA+IqBWoDYje6QVJznxPE5ftRCEWl9B9fof
D8pyEqbY/fjRHfnYSCfqkZw5jNIRmKppD6tVmTEfeaaV8AAFAIs0TzmpddJIfqcxwWe4mhzX69sQ
btjtjlbqO7UbdyrqvsrlBMnTHHQk8LY2X8Pam2bIPnL63b8DgaxxsvLFQKa/9IHoiMvmDf5mMbor
Pz8oHeXRZAjsRBJgmQKvUChs3BCFCLMChVjQea8MBzcIbdKLW1R4tq/NWt1nA/YGyntKrN38eA+D
wm1/tro9d9QMQn6ExcrvRSdMIOfGbSb1x1LzODQCph1gemCMIP7veBiEhL4Op21NaIIcB+3vfVXm
Q1Js03uWSbH7354sE6ONnLtq1u4/WuNJG4kPypNsj1cnPoYtRBci+fBFlu32+B8ACLC9QCDZaq+V
3ShU1d2JS3IydF68nzM+j49xMqWi+J5pr+gha+zywBSEn/KpfonZocxY02Ph6B7WBukP/0ydq9T1
NBfIRfaSEXDMATqTcQSH3EdR3C9gjzbP+wBv1rnJQMBGTIdXx8s6H6+BxNwXEi7VcXLkWsj5Nfcv
xyD8nPT0XwgdmnGrUSd4sic3bYB4QIx+w8xlB/TeGaT+PZu+Fo/GOf0Mc8lpAZnPunMzIdnLc8mF
uHYELmwemjk8BmW3ps+AVXx7ly4YQ2eWL64ezSroR3uROP3oNtLsK8qq9ioD6ex7R+9iWOMvNQmF
Hjayt1uLXFns6XJ7Y1uBsl4+HlwgMI6Qkh7sgfrefCaJF4hn7aYaM268qm4HzwiMxXelZ28zvahE
ZPOisZjIn0VL/hjeLfDpnGadl8eyh4qRzWdMHZKYE4qr+4dhJ3Yhui1Tk6BhOcRX2QxlJlrd/Wsf
JDNMx7O0VansM54xzb2wLZ41FryQwN63ixcE4hsKI4MrksS1+eYYtBG/ZroapPMGrtkAlP3odw0b
6JE0e5LtEeVbsc6xHSzlutWXmIF0d+bCZRNs+kjV6JhmtEeBQjjJLLcJtt5jY3RK4P2r0eAcSbDZ
wVREsc2SMRNTjMw6fL12Ua4QTGsL6Hg7PiELYNThB6ez4ZoQkeKsK6ruVSEzpuKx4kPEu56MaKzq
Buetw9QdODvFiUbOhQtLIlbMimy5CYDIG0jwbYi0CYcCvw7c4bga/1+AJe+aePRbaJOig+eJyrfa
qmA40BaA+rf9yeUan5PNJX0NjPbJMNfj9lZBRbxiWCw//58rC6Aa10NnLP2Ll+68GvZsOs+VqddQ
Sy/D1Xl8ckw8pM26t8wtiaYSlILJhj+UNfinG6mM2cfQuBzgo78hVvrr8LNh30Jz9ythwneYZ17c
Kl/kfHMrYmy0sSLiiNIXegQwTd/DsKRv8Hq93BH91bOgf3Ylh+Pmi0rQ8r6eu80VZfl+fUQn+sAP
wjSQcPh3JfxtFbwC/UKNGnSmXFec5Os7O4dXjsh6moma6BtSd5RATBhO7QSBjDSxwyOaZV5rSgfZ
QMP/cEvUCRn5ua+Gho8c40/t5CJBWhtql62+mmLHdNfh0kM1T3t4GnD6hZUlrrMs7AjhLqIsj/dt
27ecsNij37MbtuZjUFMO9h5R07COaCZWQXnviCVj+YaDea4DP76I8f3xIP06usMZ9nBgGgTtmCFX
Lcu+L5LNVDWEuYbCmOLLyJxOPTD6HW5YoCfJGfLSz0JeJGkn0fWI/QIWcRXrrZsCp4GBVOn/Lxkv
hHryRoqMgZBWNv9615KtbRt3KA52btCilBLJF/sS7wXKk9fShK0mJ7rp81lPxhzu+RzrYzZCTlaV
TZEZ2sKu/d4tFjXECuANkHmqLAG16IK1EzFuRnD5YpL2WJSEv0gECi4fT5Ge1+WPAI4bp7iTMzaA
/ohNm5k5xAB338S3YTUOzfZHG8vq2X/8xU9yGzbWVorWfeIzdZDFrj+euB6O4X8/QoRqbmq+0bbh
6YqI15OVszCAw/DT5PZkLtuFt4Bns65YUhQsNH3eN2umBgG74JJHSawC2jdtSiJspa0cFJ7tVwUm
6SWFUJQ5+dZdcXa4S1u8Nki5F5QGUVKpXFVytb2Hr0XhB93mMGmlW0/qeW1fc3mog+xlPbUzSqSX
IlukytmFb0sKMtn2uwoN2bLEUaVe9GeCEJ+N7vR9Tbfh73zY88h7BI2X09ZTTR+IvXPA4uaKO0Al
9JOftlmkYO3TlcLxaeUHQ/FG7UpYe1zuWW/++MLziuGa2oMvtcJVAVzUVQTxrrg0ClH6RggKAHWS
4VswTJiQYfXv+DiKzRwqytVlRubmW68smF+mB5R697HCO/xihMYeyWQ/lf97fnVvTrX2dv9cWHzB
rhFcdA8EU+NckimBuKPMWIgYLfcT7iduuEHG+wCxoMDJjpmmF4IhncTDPBOCKA/96CAhcFwdEC3P
gsoslUWEoDMvbhaScf4wo1u8F1RvVOFCZlkcX3BfXxLeYfahlnqCjdL3io+K1g/k3GLFMd7EQEeK
5bMGdEZ9Jsy5z+At+3/xoUQ47gmBw3HF8TDVEUyuXy61sJHDhWoU4mgaDtzjI94P1nskRz4J7VVk
TjC9cwmzqNX5OqCmE+KnTTWLNobt1rhFAWht4wTgrcXToUuQv6TV5SW0yxsXSnzeKq1eNX1iQSSs
kFdVtAlcyxSxWoGMhyZkjFdRSJCpRWS+31HehBcpRE4Pt7xn6t8FpnTi+Z0WeOUrsbGIpCugJtRD
u6oYu8+ZONmqVZZ8jpokp4W97c8RF288i++657YXjM3ZUjY6pmJI68s+uGebAUm5a7GKJCHBNsiR
y8YVOnjfDMzTgGkbcTKLljK1xCJ/5EVZwUX7lTcFp+ZFpKM1otNf67+dkvbnRd/yxdzkAj7IsLxc
rxR9oR6pCzjShZwvAFzka6beFFCRa9/3eKh4lDuQKxH+5kZUcx2r/KaVH7ZJypPb/BfhKn1OjzjW
KR22GS/xAzcPxzGWfZh/QDDJejjUeNRw44pHLYlbRfEp4uyHEhYQDpO1u3jUF7KKLSfhCgwXCadC
hqKju6FK1xDrAy1a8haDu2j8yj0Xwp5WTJRhZbRf9XWWXRocqFVVB8T1pf7HI1EgDd6hoAe67nSq
Pq+a/u7Q87W4lirv+jTLRxYXGW1tM1rbmUfyKUvUuuMqviz3IEvxB+D6uar/2Rua44vgx+MEVRRI
UzrvOtaLXV2yZaw/gmXbHlnbP/9qiiFd6fgUfysCocKE5OeY1LoLwLIkYMpWrna70t5mAFhAwxFV
OpEsfyZbBQLnk2phkByeiyWuVva4m6ixA094qmiR1+Z0iNvQPSUMLFuShohKV9yld/uzOpMCWsOo
8XPngXVmXO5XDkHCFAxZwKBQtHX26NCtInApU9VcFYVMSq4tuabBivAbrsGPBTItw44YDX5+qCMI
g9rjDRWWNT9lG3xch+19KhcSvKsQcvitfIfOQf7jS7pvsyOCyqSOl/GQRMYueuh4wLpQm2ET8FIN
A0gDO7LVsYw+W2RHFfX4QOwvsVJujZNc6BLloJW7Aaux7ac73OP8XT9sXCP3G5LDmCr32/E9R3lR
imr6uu3QKBTZ/2L2qK1BMrtd9uyqRe9seCK9BobMuJGFHF0g2PdwxG0XY8GRKRDx1T8PzFXWW7qg
u4iKicxjMteJv7ogLvHB+JkN+/fIzybG1g28j/S04yqxK2ApFpvHdUV+bdoqyvsrUVOCJdm4R7NM
BV8VeT0oZXq5m4cH+76vFLOGchVfaP/536ZLEdDo04BMc/0Dwzb1NRHWD5+J3126lnwOSkOtR1jf
Re5JPN51fRzCl/23M5aO/klqRtEEFMxwjWdAKLJZbgpJ71WAA3l43903HPAng8LPZvrisP2hGT1U
FyRU2UAMkOjOeJCMY9i6nKCSZONYaiqsIB+O5CgA8mzxyMW6FPsi7hQ7JtGDUp8ZFqmIvBW+vEKJ
sCmCLwubkVlNtl5xOTgKy+FmLZmba/jevPHu6LGfNmTRgdxdrT40yUi99HVKY/r3ISeOjQNa0G8W
YR1XF1btJZocPSdLozay+8uqoh59lzT4ztWhamdZxHzKlBR6rM+hheokgIl0TCkdBzzDgCsKrl3j
ndHJfejNC9n1b2JxLT9eee+Db3cRkEV19vDvezH5naxzJV6VNlOtdGHH9qBAuwtBGf9csFkeAGDm
642OfAfqnDF3dINZ2Hl88hITIroaG9fr973NSkTryEMip5NpsuoxZSBn57VVBxNJXww4Q8hcyjzF
YJqYfoys9AyVgnsafCQcCWKWMuKMZPnqifvgJCi620iEoNuioqZ3REZigVqJ3e/RTPtDAIpY3e+/
qGcu5XB8Bi0/teE31XREE5eijY0VtYdj1T1zQJUQVl8SLe/t4m5/xvSxTrHOWUD0Vdxi/qzpsYUW
mybVuvVBU6aJxCU2gBidkDRcj4P3r0FV3SL5QUP/STk6yjKYVW+QfYplEN5eDpef85zcFoqap+7o
dDMTATzFz9RJEUp/QNgJWAdj3Om2Y7ZW47iP8Sl2NBHQr2CgaHiGvKNa3fq8iNvPjfhIfvK65Vnu
Z4v1orSVseIQMREqb7K3bx5fabLY6mIUTcHNU0y+nVNredExkcLUPLxS3K5a1GM6+rnmGtCA+yNZ
YRVh/T8X0vHD62w3OpK6CtYo/cvXE5sJJV/u/gTAaRtpdB538coW48RBYOLubrFevtFTzEqAQEeL
1WjTjQTsTN5RCnXN7tQhfKkGoRMDmoXlB0Wj0nIk12uNhUdZE3ooIro5k8kJ1FNRgxK9RKeaGAy/
3O6qtdV0A5iS2TePU+U+OMLo/RJtroAUKfFKkRdCmm9ueTblVHtA9/O7hWFkdVG6k6bISK6giz3l
RzbN9tD2d352I3cTur1pvVwQWMVFdvZ6Io8L7pb2WjyEKhTF+mGCMjiXExkeYV1x3k6tDT/stg3W
bC3K4E5z8T/uOokM4rfcqrdKwReIime6ECNGYECLRjWZt2Cx+6MyXfPYKHwXBeuadhQHXWg4i0Yu
ucdDKa/PwFyQZKm1YasABl1qTeIRKzWdP7Nn3APuCKnGQlCUTI957JJ+djYakZM7CmzIzzMwstJN
M2DCvfO1iMFtMruL557eSoHqvSHaa3ZwKGzJ49s+NwI3j1IAE8ZCCjZp1MQR7zC7uGwUiRbQiMta
duR1Qpozu6uc+dVELHWBa74rlOZjyVY/ySnjf8bu3Cwc+BlCmXyTcwHyO/J+fHGTdMVyWj/UNNFy
w5CGm47bnguEt15UIti578uSvCyg8ronxGBQvI3TcEAl6k2aS0f9xNwHh9RTMdF1hATjUrI9RsHi
BReDPMV0X9nAnewi1pAMTDQGitbLSb0YiCKgUtkH0qephbTc6g2T9E7JndnYQFxO3HiYX4grxclG
7Nc8hOcjfpXmkF1TFwzavXEiiD2TnX0cgdLFP2EerLmyIZvMbQZlR4lfiUrxCuCI/1Pt05TBxTbD
PI+hx/jSkd3r+F3zlBjpmcX7hE3BRoVbkj8KaPgL4FU6MTbl2z4nP6st2wF4LdizIVIsxeolcuku
VI/OGB0Mn2WVz68FjQH0NfQfqC6+NwEMbD9NP2eCfzeT8VBOTBu1CMypJe9PMEeVGoMHY9fe2+JL
a0qrB8L2dc3NHaa1/qhr9A87/NLBOeNghR1flBJ0qoEKnaTC4PlBVUTjn9qHz/ady8CwQWLZkXcP
TcHq0WzfTWUSUyHK8dDKXvR6bbViiyjk3bzbqNr//TP1uh6DlbKf30CHomidfGTxjQGymjT6i+2q
mAYN5Q7n1+kHlDcsybunMX2qUne2Rw5H3rkXrAY2/qvkUW6G7CBdyarR5cHIQ8XljEoJ0umRK8/d
VGrv5444wEdbpYGD4HbSoFwfy1LfKgPVbxO7xueoy4G3MInjHSjjvxk1/2QB2GawDYf/NZNUKXYS
9KOOmd+9qjKUstXhPQyjisb5Urnf1Infcm7Yo1/78wDSTUjg2EZbVGCtilbnPaHH4WrVMi7oOkgX
J01kDP2mY5EJz93T4jtmucO/ddQTjtVnL7pv9KQv9ukOtv8s4uZMdTABi30sziRT7B9JuD2GeRN/
4yP50O5lCEi8Mmz3Nplz43Xesf+akP8lDC+6m89jMsPct1InooNlw2lT6mJ3DNbjbVM+97I2DV3H
On7EDxb/9FstS2tqyqGE/piXs4KfHRHEkeHl4OEcY66ncPURUI/8SKn5SMJM87+G1wjbrUNik0He
W0WCUiKLh5ot8w4fT54RX8OpAEJT/RO/FQy0016uSlWBSW9iB+CVYT+DifSWRfu8z+mRJmEh8/rM
aiXMawrJZnyvxLwch7uBhuq5MriIBi/SCjYxZpCnIfaIK4Dm+lOeSFyaWCiljpZSECPXpY3Bgfxf
55serabW2fh2Rc+BQpuHalwkAZq8uxzW+B5UIessyfx5lornD2ZLHFmH//690GVdpWqhrlnoT9Ge
4F+htzAplLci3v2LMcGXuq0LFrUadYCpXqZSd9h6YxjcUaTr333gZ6XMA515bZV0y0z3AMfbkFRB
grSVIeC901jeeU3t+UXAtVvT76UtpP9akegiXCm0MWRw0gCcfRv7/5vZylbL86l6pDIAqW6yf/J+
CPrgFDN8ELzgsFch7ydb0grSQWnx+VUpjpuB0k3Qm41Xf5l9abFsSo1ZJrcVOVTdTqTjK3uEXNLI
SSn1xFG+q8YUWU3DIUHoFeGmGv4XhD3ELT1kNbgDKo0qhJK680+6pVxadnzxZhA2pmeQNlHQ5roJ
dVU5n+nCeKTVnPw4s/wDmC54UttoiYfOnRwzC5kioiMcYnoOllxC5cpWtgnAdTsqOzmvlpXyyzPx
p1hoLklNLocCdNrS6+Jx5rStWCJmL/B4TUway1JgOBGAWMPwFNcvSpYr6PBGoiwuCna7iS0F2IgX
4RNCgX++W0rsJzcqVvBvUvLx68LMwW+m7K0aOsxQOKUpy3S9L8MeGckF3b/1sy7bBQVzVhtyn4/8
pNFozcvOUZamO9eudzlVYaK80QMqUHn4mcmlfK3Pe3U78M+kugPgYHGmrLbnYHLb7vEuzHlN45qS
gb7fIDqRzdGHMMf6mK/PuvcEP05ok4t3Vt5wMC3kaCOMVT5AOsJL80XpOiPKiVq8SIIjnMekb80l
WJedILYEubCUuZckPPA4CTEuVt8ecFDyufJQAK7WDEgh60lLgHqBFYkKkRHv2p6U9/dtF/76yPNa
UFMj8PkFaZe7YDGfu4FFkjMFqnggFh3j0PrefENtkq3oFDBrMKrDDjNH13eScm4Zoyjo7a1hJTud
S29ITCKU1etKjF8Yx81lihnosc0Oj1PSopuJlEc4DI4axR6cutXZyXisiOf7w9yZdSi3cYBTJQac
lWvIEdDVdYsG85TlxBfw3yQXyDJ/bbVJ8NAeShiht9VpX2FrrtsnA2pXmfO3RtAlG31ymWIhT7sR
HUpEhmvrcWtmFE4FIe0/owbcQILFgyMKMxHoFTJW/wR4677d9IJkzVrhkkNbjiqfwP1q0aVQeNfB
2BnSQ7ppQWuqHWPnCedrAJCefBvxCOWpFkctm+pZH5Y2T0opHWscjIolkkIE6aqVN88X7UNmcXYe
svdYQQ12FWCMoOUfJQgo3uLv3l/HnJWVrdTy+NYvUd34A8zHIWwKW/P5PcPKjtVjfJfzbUzZRpQp
qs0aiSgX5Ku96NUyxF81YjGJFrR+nipIgEx9DUuschWGwLQt8u2lB4hSoFZSEqcY/d7GANN4S9TI
xHsJfumYlI1k9xFgRpfHtB47do5JQ3ny77gbfAivXFz0ujjMzAn724+5Lv3qMPzOP+iKyvjxanK8
Wp0+1CMftNMQQ64bFNcpdWFm7bXToZbyC23oLk/fwZvaBP6No2ttCL7BHhu3vmx+1dl0xm7wjjKP
ysJtbAx4M9vQHqeOkLF0ZuAo0M3RndV08OFiob15qUawhbcyybgveZn7VWOfQ82n9LmxRFD+smCi
CPB0sLXpnNf985Ftc6L9DVBOT4YzbLmmwpM9yjDHvmPheTIHWLX2syKSTsBT+/7DkGOO0Y5G/ZkT
zkf6Be5LzSGLP1r/YThsblbxIDsMkZb9PCSvUaPGl1J+Snzi7fvdf1hTiBjH1jhYWo48e9nsEewi
C5cJebBrAiSds2wq20ywyle01266Mo4X0iVLTnMOwKH4vwMLFOV/6zEU6UK7f6sIH2Gi9vPrGZjP
hdBxqu/JSkBqI+fQZNavdO+ScN8BXSFgPwyrTi4otpCAQBbXcYdtHU1h87H6s7cZf96SiKqX64Rf
/AKVouaL4IA8Wf3j4eAHEw+oN4RWD6mPuZPNUjh+fowJegSJvg2M4ogyAmloW9QFe/nbVU9apuCn
IU0aQjwy3xsKMWwPgD6Xfl+9Lhg2Spm9bmDefSEvy7/SkZoE3DwoudZr5uTjZOjocgnfYiYxz5HB
xFNzf4ZdN6A5GuNUQnSBCMdAOsai9gJcN1gX5wiWSUxlS3ROsY898l21qKGSp2Q+qnPjvm9frJ2r
5j50JXvBxocN5LevK0Yj7NnlwiZDCqXiZrDhDXslc933V8Odz2fQ+y2ssGE6FxGsrWsbSOUHJcB4
XCO7C8rbSHeICSnf8ZPKdU06Ypl3axH+nvkV1C+m7O8S6TrJ2R0q5PHRnfg3HXF6KlNoSXqwCRPu
RfN/kcD47ftS9G4w8sVA9TlV77i6lK5u35hE57csa+IbCbnbYzU+tm1sWQ2k07wJwFVTgPO3eCiE
keVWwOerqOox7YEwgbyNY/iYWWyG/ZPgg3tyoUAK6V5V5b2xUZ6lCAEYL4y0SwMDBfohmzyi/hjP
OkmeC6hqLOz2+Cr2fa9laSOtrVw9bfS75wPmvfm38dIhTggMYyaloE7Ko1f5Ly6UVZdzCKVzjfIO
uNgoDRdgJSIXZykkjj2uZXL1Vq7ch9t+R8O9Dp57E1uwGg5b1+FqCli56E5vxhnGAMoN0SPsouW3
ac5R64uTM4W340iHxdoBID6d3xTyPaOmEzOXuWaob9FRHUkVUhlwFH8oQNQxdYcf8pQLzv5Lhyqj
8294meZy60yhyq1VwAzjdft+5BXDjA98tmEOuRllUR+d5djWEa0Vrr9t8J3hBh+9MMu0VbjrhYor
OAbNJiCaotN/2yKlYSIHmmbfkNtlatNXIvASpeQDxCV7/emi9LXu7mxYBmeCZpspZcIRcrK3WXAl
bLAozgiIfESJ61+YmDWkgpJEkDvPnW+he9WhUVk0p7/F3bYdPoZPerDe74eOnLPLvXT4YJaOZKvl
wYztqK6EHKg1jlIp0bfphQKqP0P3pcVm5V4QpbpgTTAzkGxJRbnDYstLgx/zFhG04MUtkyaQMJ3B
ubZlsjjgkS9mcQW9Plvnyiz0TtspNEpYAKZLhB+qK9JAO4glIFagaDveIhkAAPTLmzpjCSKOpmWY
3FRpZZeGpddMz+MAlE5JhrPQP0LR88SiwQRDTTS6H2V3UCgnozDcna5AJ5oYJLk1N1E40aj/dJ71
f3KPi3HhDfaTLNeuLzUgkd+s8OqOxk+d2RtUNz2/liAn8NBfErWP9KHolTJEdcUHRupYcFg6Gn2/
6SkA+hfGR4kF2OwpGHxVbhoJFyKygUN3CjYixukeXxElsZKWAvzATgu1nDkUrHv15iQDy+v5POZW
u7zA4ThXfNzYXS5DWL1mK1ZTKZIO9cLusbkaHadrIYvjpSFlKBrllGkAqw6PqJ0MmwLZokViYxA9
o0+EvuyBU29FeUCVj90+kO3R3cDn2zr+82kYOOPiLCVbXTh17TM5kPmwmu8FLfynYg5PFIjJaK9w
qbGW3Ax7rJtljX6XN0dIgo/tLTC8W7CK5UN2pb5bxFCBduWLZQiZZ22OMAAM4H7qgV8LhIoXL/Te
dFNzK1GP1ULtE+tBGO3aTKuwpmeHMVD+i+K3ZhTmdXwcud0L2nN0TS1A3i967a2YIHrQpGYOLqIv
fY3V2fO9hFaf7OXxFD+2CddNa7XS5ev0QkXh2oL5he1OXBd1d4AmM5xAeZPKAEtLYhFKuxc1O8/B
zZVkXfCUzk3qaAOsPkrKe2AdMvi4fCa2/XhyUydkVjrU1PtcDm08y4V9rYuFPxJ7LumMBQPkBjlc
WrZMkHJhPideD3vEsYg6ZqEBWTxtaTOKa9J1JgUUsBaDxAIkuQPHUsCDklCv5ozVfMY8PQfxz2/F
nalsRS3QfHSA9zDyLJfHIKgurpw+FmMLEtYUSKQ9RMMh+1xH8Z31XX+5oYgQq+AidbC+VsXcY0DC
YkHiuU25EqCtf1mcUHufxLU8vq4yGqk1iFq59IyG9ZmptVM3KwdcchNoVWnHZ9dIhXQyeS361tSi
tHz5x3t/HP9XGWyE4ZqCqi7e61XtS7CBenj5KjMuB/SAwryMZ7fZq1xDZaF46hGzwgY9fQIDYk1+
eWIelnM5ITlA6SzcKaFVztanVCMyVYWWGAdkZe+Ewhz49C/U8Q27d0eoRip4y9Vvv2hA+map+teH
c39v91T2IqjB5F0PkpjDChQgngPNXTyf2SvbGaNDYeWi8R4C2FoqojUBTR3jHcUdxGiNs7KUwUGm
e6eBQxwYA2TujbXHdoSDb8NGuO6Ply797bCk0og9YH4OXvDbGfnuAM4E2BwKFZvVclhrOwhUo56P
8r0+kJnrGyPcKAEi1PCiQx72rQdpj+ssim0NFjWuvDJuE2fA234hfCGzhTxFeAyWWjXjHN7FwsG2
r6fBX4602CiFOH6mFhiO8QW/DVAJIFFbEFSq5O0m+74GDp/6MKEVYbhexlK8ZlH5StELz7F4y7Dd
QAJv1Ssej3cM8EsLa/0weH8nF/sZkGQL0cqR/IaZrzPRdnWbVYssWUulAph1V4yGwtDqcs3B4DPK
0bkACVItxWpFlf5+B5Upiy9opAz35/ijImLuWpdg6XmOXwdfDNz5B8bWaBkG6YVvfU5gQ/3fVrlF
Okv9zdVJUjh1VK4P9zDQbFni3Dd2zkdNM+cXZtoarD6ocqLZ79c2lVGcebVDWNyOOmzu+wUhYxtW
1EV4ZWM+KC131wXI+spU2cUh5fig4EJqgLQDhBlA5dMsOsYW6Ak51n7kzpP3MI2eORaKZ8Y0Oz5e
VfcKIZM0xbArCAj+vMlkXb+OUaEenR32J0jsrH+5gB9zITh35XiH4hgQjgWVYv5acY0Vlv0anLiq
pAMOQK1n2h+DAinOMQlEpsCIUYKW0ILvCDQxLpMRHJ5EWj/1F7HWUoZhSl42hdHkzsBaI3pw68mW
X21RGiZG6Qwu2j3EqjhWs1L4JrlWcatf+Vd5aiiBWQ1/FipMNTaO1HOTStzXEFFE6pB6ptp9GD/F
qNvvZXsYJLGMJFeOrhyZ4CayleO0ahgtRqrzA+/yXIGcDjCAI+mddnxykRuYiSJvaqGOfjC4qrzb
0ATbJvNmD0M+4JqqCTWqdAWv60y6c6iuLjYZzFI1Q+CCaF3cS5ycuWPOXga+dp9XhudFQkaeaaCG
3BUio56vDNJEpvn53538BxSb2J40N8V2Qm3dddAbrqbEJi4hQCll4MepPWM4wykhXijCsRvYCqIY
WTaLLnqCSC5xeJ1y36/ek1/5UYCd2BUtAM/ge8iwV/LHNRi2HF16zlRYxykhCSt+jJaaKEn3cDBf
4JOdw1OQudqfC4VAGx5Q/l5UgcclZvhPAokYsiN5TvunnGwr5tvtzorZME0Qk4ujAgnQgi3O88pt
vpjU0N2lnTYY+B3Kmn5Ad5gOTKvpJZeJMbEF5FMyDqRshvrqJNem0b7yFteF5BUnxHHFJ80rHtGX
qW/+/VDtYtEHEv9TkctUOk/q7IvkpKNYDMjGgOq7gfZilT5Bx+TWz/MsY6fKel6Pmz/0c9fk00LT
7zVg5O0mx5XlYIXJFhs2IY+gm5jxStF2+U60c7WzHSF3TduX/9zinnvt3KVqO+yKH6iyRnevw0vh
qJybIpICPrAlytj2ziGtp2L0QwtK7hYZch+74Cy+/iNme9DwOp1jbjTe0siw+BEhVz0M8akjNWfQ
hEUBSrLb7lMovsl2C+hXVIOmcNuIUZPBF+jhF1BSoCQSuypAmkoX6fqvwa4AMIC1VYd/udzBVNny
FKm6FLGPScm9fitA15pP1cLFmrmK/UCmrBxIj93/NTM0lcCqbE7TS5dtcLyLCzOcyAGY24ubWZfQ
88U8k8GWHENl4N1Gcnru6+96/2TnCcgwu0LEOLraOpSHSnJbhzRpOSkxDHYPzWtv2LNRLQhUhCwX
xkiV+o/wKkGbs705il7+wUcKRg/Xsz0kf/c9hbMMMGinZgs3oJ6v3EyJ79FpWMII2MnPbcahSmKR
nIRy8grfBSG2gERzBlDQ4/PhJnTX7q/Ug5zhVfdpnA4/MzEdbuSdi+a5H8Lw4LDDYEk7IqV+XSVv
X9QAysH0Ee0SUMkMiEwArIoy09uce65o5CZTmv4gZt6A5NpXc4kxLyBGbqEOZFW3XZy4dd9sm9Ju
LAfmQr7uGd9b5L4oKcmuypZLAuTAnbxsE1TDVAJyiK9X83C2xtnxkM2AixE/A8fWb4f6h0qdB0tj
eHMOUgZDqNskA4IseAtk8elhfX+BZtYquUchX+tDe6sG4yNhEPlBYQs9UpTQQ7N3pjq9Z7BHrpUH
higaub1JBx8gtbkytfL9g6X1TAMVHE1IF+Fldphg+z5czsATTAh4HTKGEEyOqUSJ/jz5dUOdFAtK
2miiZdL1YQXIabMAHv5J8JfzZHvPHbxR5+/A71HHAN0IXKEy8yiP09GBbQhaVE4aSxGzRojkOcjF
lBFLfIXkxbc7SQNqQEqmkR44vs5LyT6hT5wTfC86hYh/E2Xisgi0MH4eFBsL0u+e0Uw47vFz0XFc
pOo4GWJX1evWjL0zJiyzjI9+CrSoVfr9Z3G9l9emTrepkafZOXDU/Vy0R8rWy0e5KyPetX06/sxP
tIDn0k2YYztWdD2kdxJIO4O30ARXXZOvlmQquthL07jRdFlX+jvbS54C7rBxrA6YFTfL16JEi5YR
AZqyFe46U80Tbf3K5znPee5fLHnCq+/9kTD7tqNjiK8I7qqL1PGrq9j/GO0bnTFinwuaSoEj+FYT
bIkIZlE/U7Qn3KvknKZZ/5tymayPdpv1og01lsgX/lopTJylA9HoVEwuVdlFWWRUgRJrw/QqtknK
CctHGyl+Rer816VqElbugZ7xwIkBV7r2l+IXpJvQRZCxTFEr3rBitr9MW4L33r9D0N68FcJfiqk3
drgsD46jVjlfV7i9c/q6pVK9kEJb5TsiTbNU+iTEMRAj9ZzAv/MvIftJEkaRqkA13MFuiT78E894
f3JW7hPWrJ1+jDQ3cxm0fTSo7J16bqF5nz40uzFF3vwBpUCKB0dztheoxCCvZ4EecF9xnJfTlJ3o
gBiuNVTWByKKJ+aMW0+S/+wO2QER0NjNVNH3qDvcetSRm2b7Iit/dmp0zDCtTAswXvjOoQfs2KP1
0ZabY4npF4YZcwAeJobEhhvKUI87bHoe0XqIx+ow7Yxn0TbeLgfgIiB3UovJ0gJ/kglRz2N/jL5w
hPRmOTTFeo+guFc7eZwY625eVKkAfK2okuYjKBm9W6sUA8O5anXhNZm249a6rplU7mOHprQ+xO7B
JcuqrZTP6MaZjinD4tQPMf/kmWCjqbK3PnoA1gL/M99gIjL56CqPlpzlWYPLM6T7kV+8nWKAOaRt
R4tVEPU/x2Ef6CuCqtGoGVeISmP7Szf2O4Bz8M5c6VIepQnl/PeRSgdDctz02neMLqqtPQuhHQHS
ZUMTx7GxZO08K8c+pI2N0tbbmBxGVWG8ravtaIatWoFp2lzOt0/eTuvQthBk+J2sS303igDShmgp
dhsX6wD+RUHaZ+EmFh2hNzf0UCE6olP3F0xBeKxzyyQO7r+JGN8IjSFW0l2CUc/jB2siJHWDVBex
aDYVGtQhVXeJeOouW4Me41ccXqaBLdQ8YMOBDbR2p3MAbLAB7k8MlLWezTR24EnrGiqtETwZW8Zv
+NHsCuKDHdsf7GdDzCGu+wbErvItK06DeG9UCwEfpqSqXMQGKWJGMySQMZwyuHtNk4ImgPeD7z+D
wkfc0kjiOTHcuFu1dVH9SCPK+f3uIHwKDXi9Q9G+1E8McNaSdt3jzuihn7fl/PaKUx2sQAbI7NDu
gEKH6yYns/lFDTCIGdPKdGg4XVNNcjsPvXz71GA1tIv5DRMYwTdTKukQEmU9Zu9XLxRPWPE6VQCg
qiw58ZFjAjKIGaaY6QXgIrb5MLOEZu4XReoORAlfuL3UxH2Q6ktQKNpbS6rq1vwG6cLb9ivZuF4V
fUouZTscnKxIavtXhWZGZaqgtFXjCNLH4jTx4lA9eMvTR3ILYqn24YZ7uXEWKrUAmfzQYoE9HXW3
Y213Ts5cYQuJXd/q5/9t6UsSLJs/xwTnKzLqFLhF+cC/A3jhwJhlm1ppqxk5vHZD0XOu90fHLsu9
C7mNRqec8WeZkwvFkAiUyb+ugxk5xYS24a76sJM+zf7QG55Ea28tVRJYiBdJ74KHhHQNTCpuegI9
oOaK4pyjZ/mxuQUt5HN07Nl4UVMnTn+hF/02HyKUBhloaBh/XtoTscIiTn8SM1GLu/xbDRgWDLRH
cjC5zX0dR5bb+V35JSsrN67YO98hCGXe5DZa82U/jNtp8LQd7DMqgqZNvPFtklFFZIljT/z6s+4T
dhb2K7QiM3tGLNUzmA2QWgXcqOp0wLKgcKNN3s8EA7JIn2AQam29lFqV7GMnUjGRyB85y2Aj4yX9
PebF2ruajqe2Q1ffzQoBPcxv3n0Vl9lzYNffEafj0vWJP7xeIn405FZRyFMgb9lVY0i1HHc6Lvpz
ufH9iJDCwxQfYP8fMy0LP9vXPT7vI0ud4c94MOrll585QCJE3ohuQEDwB1Qu1I97J3IO0owJ1cFK
eZj/5nRvsCLP8IxX3Yfe9VygDpk0xONRyUgu9APxFG3rc84zU8YEFJqQBRvt0xPU4iQ1HIjBzA5V
zAH/U7q+EvDi+WzxqLl9Jt6LL1Qg6QFgMOPic8j+iEHed8YPw4DEhDVig6L5tJUT4a+VxKtpxhmR
UWn8jzW5HSBGtj2rRXh+XX4LWRfZ0TAqyOp3bIqLTm4+pPSW9zWIM/dWzviiX9qoLrLAD50DrLj9
4rgjgd0lMsm3p4ygggUZb3LKSn58cziRAG1tkPAObR81VET+7dtOKlTjgqIlNOZHVdhT6KwDf0gp
fxKmth5M/mR9YaI6V7jtK2lffHBX+raPdHtW4kxe97m/m5i5XyS6ELkb+TJTWmk8/x7tyDNRynPu
fzcLGKEs87IyOFInROBUBFNhhXBA1Jj48Jh1GXrAsKan94P2CVjtPMHZ+VeKotBbChdX9iHnAyNj
HrFu6i9htAHdlXSqRcjicc1jcZr7h3X26qRkHKmvm9dnlkOEfjV8lKaFunPJm+RVx0tFztGRb9oX
j+5/Yxdwc7zDqzVp7IX5eZBI5dGcZH5/+Zedc4AJysoLDa46AHVVUwOE69i5ZGfjZrlvk6RK5NhC
nLNSI9oZS1AKQ8Ecu0Hkq/aPd5BxihuUghb0Ryw8xZ+RJSaZs0ATCzdZobn/kDvIESXdtW2uabeD
Hh2GnOZ9ueP9qtluFnWpHNtqR4G9AqhtcBG1c26nbZqv1L5u7D3TpouLK0lwxfk5N2F40RUvQvrr
vdk7Y7t4ojBJFZuzx7hbJcsxchDdLmC0RWGXcE85meBbDYKXtTLspoYFuGoJIgu7OJUYOL4Sz+MF
PEgFPOBR+a7zq+NawIcDHzxfynclirn4qylq/q0wdRVdJyO94wxNV2g1jGnyNadh6yNfC6gmaFxZ
lAYx5/ihfnG6NBWEAnJKqVGjk7OyfCvp5Q2mYaCh6mnTLAzcQkKMwiqkOfcqarmV8/kyn3ZLpm0t
/CHjBtFJffVZ2EKzBK85F3Peo74mWDw54018UOuEidnJofkff2ckRafNddwOFukbNtmpXo9DbbVP
69akRnT6CXMvuWVTrJa8uhNGyfgXE4L8ZsYrDpgpOfg4ojtI3I9ShaIx/VQ3z5pYyfLBIOUJGhxk
pUmiX54JYarp69bnbkgdrAYpoiNx++5LnrYFqCnXyYnCLM8C//seLW9PxWw1jWZ2i58VcHDJozQi
LOGe4CRLC4JfTOa3lAMHcvTpkUKdurSJrJhfxOUN/VALmPEHw2d3SE4IT2xfzoLwP3qHlGyd469c
curgU4Z0EDlhNFobbyz+ivhQs1C1teuKsEPh0LT+mJEIGCgKUAzOc1i4vhBXTxPZ44OIQM678Tiw
9KnS8/dxuEAyRT3zL2U6deWiFPvDHrlfMRyYPI3Y6xQM6Xrueb3hfc7CeQfLTOf798pG+JVQaUJz
JnG8R3CO/To7UR6+8IeM+8YoSUiitVTnmOhg+VmIFFiB2SDRNByzXVN83gb3UFFh6vQ+iUyzpfAc
s73tzL9+vQmvbHyfiEiLGjgICNcXJkFMcA5Vfep0iQHTjgJ7055bv6o7q0w1TgQGujixCnaP4fzV
1B2C/0/Q7Nl49vnyGOb4y4hFJXrW+yfJuKcUf9Nuyd+tGdbdNEsaGzTXsh5Li1tLexwseggab01v
oQ6nZmZF/fTeMe4u3cd8V38V7rWcto4WR+3cdEDGwRH2hMhU8GbtU/X477GasHKa0BvwFWwpCuhQ
j57+Ho+WiMHRqlW5A938xOLeaH0e75HqrWQiZugDVr3A/RcefVj8Qeb540Y9XIM00hB/RumZHbh8
rnOa8MS4HX6GRRJ2FSYR00qvKurFxKWqa1ojf0x10Hm5qnc8ENG4nWRMlGjtWsf8XO4LUEIInlm5
IXswZZMj8UTp3BYiC8Tll8IVVMFI3XEjmUjK/fN/CnfB6bWQzRX+ZMKKArWK4RYJavFhg8WGrBvW
DN43n/a874s/Ve7rUbjCs8/qHTgNw65Q1h+ysYjCQGIytbfgkLAisOXIwuQJekxfBvbh3m7hFIdn
So/9aYzC+xQfjRKitJT86F/uq5FTMVRQFEzVaD0pugcip9bIBXsoppBvmn/lPZPqtcbR4KkRGsnf
uHeQHQbXHJDXp/eSf/jQPkTFl7OmRu2Wvf750ZC0oEbvRBZtTJb+Wz3rMhkzBl7ZHxoq3EAixrI6
ptK+rew2alR80jcKN21GLoHzBbKLvtalAYJYW7QRebqLCLs6llfo6pu6RjtoeK4ztyBQjP3lEwQU
UAtGToaCfX4lIDyKkmH4kLGmQ96pjkzVgB4520MXwHUU5mlDmq/OR54dzwiyUxfiTaoAyQvT60vL
lh60EUO9Jd9B5xcUd4CDuyb0RYBUy2HNbKhdRhq2jS2Vph4FcBNf6BFD2mDPexa1FxenJ+ozJz1M
EYEaHSAzpp8sIEkNCxsRNu8sasMTZxK6kjhKTSeUafXbBSD9sDvBTB8cYUj47I/nhYKnwvInqD07
1v49XzgeEP3oZXpQqSZ4ie0J+KHNIRAIyqAqG6T90DdbglROXw8fAzrKZJ6HVlVWGuzEOWIDvbaI
6weoGD7K+baSj+M7SDDjiE1iNEloKXtNpvmZsN/JXrIMwCHrDFULr99WCmkc7//MHEbEGZq5VImJ
NICTCtY7DrR1E0rTwj9IU2ny39Muyx6qbbJZCpTZKDra2L9pNilhEmLnSdO/TKMoBWaFSNnzfKTo
0IlC0Zol8rDPAd+hFLCoKX5oVb1GXO9kx9a3LdbfhbWlHxHGGMPxWzBOCZsjM4wszFjK4F1BtuNP
iUwunzzg1k1ErFoky56bj+a8+qzENuLgWH1OQ1uA0AttbXTQmyHSx8WrpbKzf0vLTmA6kNvT1Ic0
fasGeMT2PC7QrwMtZ6AEDCDgY1mXu+qfFzlb/gB6TW54JP3RjpB+h7+M8S4P6MnC1vpy7iAjqS5r
DvGGGsMyT6l49B2QZzsuEBXMSMygacOls5wFGr0ICmQpP4jkzNY3F4xZ7glHchT+syl0vjQO6eB9
TZ09aaS36egArEUvQwUdlPnVQhqBwOjK6H/KfNO9XKdDPDHD1IuFWSyz1YT5tJMABc4EPNvOmp3y
qBSvy9SmXukOPWjEPsiZyGJn4lY/vHbTRXsa2OSt+7Q6vDXhpzDKxqLeEW1T0mSoqr9y+8MZCMzj
6qhWt4dSS7PU06DRa6hvAraJDl+3KuWqrH8aSpiXo3uTJ+OCafLb3W3wV3NMzAznsJZQEfYRW+El
ZULb41xvsD5uSJzdOrsgQPFnY5N86aePvu/uV7Nb3d/btnIxqv/pQVmct1/OeNyuFQju8SNijSBM
jny0td6kkDi3ZZHQx3h5421C/Bza8wBmTsWOzROZNawWahBdbSuFX5DHoEJyLOnZPAPLytR0QYa5
4L+T/YnaBV6t+Cc2IH17SxtpWwMYtJl9HFTz9GCSz83c8UzOvBJaLkKMAuHEyWvxISrEz7tIRBPh
VLLz/faWNXeixMSji8kLRCA+7MHivEA9m14zUgsK6IIbLuEu6dCsXYFc4AL+mCfpMRiXSvUBZhp6
dVylDY9wOAcFpiXV2SrIlcq0e2l1YMeFZxivZQgXtwp9cOaXN96CcjPW3Ewuk3hdpO3Efdbe5y3P
ujvhc/sfVIXK2UxSjagQKvbsPHY6FHwAAdkpI5n57KKano8/zE/w5exIKfcSbEgboEWJqNn2zvzn
zchqxDXeis/JEGwiVltdnXJ1Go7Oyyyi5IvfrsCJ8l2y80KINtQuumjw6PL8aWjsnXzZFQE07Ymc
GjPF1o7F9qbvyU8rS0EwE5X4br8xSHIlJswTbnDJ5aZufEoe9eUwpAuV5txt5UWqquu1OP2xrXxa
SCJ1eVQZywr3sRdQog9BYG+q8NJ+A0+yH8dh425yHm09408Cwg9Yv45YmcL70oIU+fR8V7lxzcxo
bhGLIA2AXCza7iSULcEgIwYZ3rUrcRy/2/5EL3aLX1bHq0N4Kgt3KLNYbm2q+6gBv8Z1+qy/Ksl6
Hwy8u6iDKsdhvHWisRjQp8eD3Vl/LQK2s87W07ndTBa+8VrL4Pejx1yQJslL/Y9okNvmQJKvpGta
mF9uticFfPymu7HUu38pUJqLIAYFvMVb5F/GyUtZkFbomN3JXuai7Y7cYxBIwgddbbB04zaKSQJe
uFgjAoAgDUrPLmV5rbqxORBeoELQ4KXUg7TUDcVzPiZxtpyKeEDNbGmAoP4GwZmeJ+a7udDhv4Uq
upF6xKAI57rHf4HjmGP3BKkSlnFxQCt/u+4qYSBcBYEzUkfP5jPHmUq/o0jCXNevj1tKC0/ShxE3
+8kp7cyYZrQDvqN+YD2GCocGmjCPYrWlsn2bjbCoAVOKw8/Uu6xCJ/aMwsCqr2gM7DiRsK/wgKeC
XYD9qHLp1UZuDLrp8SYm8xs0P2pcx6YK5Urcdt02aYZ5bUP/US1a9wcSWX9HIkHAkkgmw+9DdYsr
6Sfp+s/znRgn5BqtjqTK3c/GyjyyaVfLnb11RKr8IPMccwIQIwwru3LOLnqiVCyudtF1WuyZ8lBw
cUzwvcgWP+SD+oBz+LJVpwbyTVrgpzqFao1VfPSx/euLVk6O12EZu4rwIXz5HDbmMLtPyjiivS6j
Hr4QrUjdSC3DDuoMcqjvcuCygYCiPMtsSJ4VsBWyC7q80GSWM2I6Ld0Gb6tK89UUR4yxdVe9NxLR
cTEZFOqrN+h70782b/TP38Qp8mJLVwmm884WQGcY3LQKm8jQWuU9lHx/ph5hq2JtDgyEyYiq+Au3
zkLWR4Vz/YVFpIQdl5uyBzcrPFXEjbBAgbZ3ppAo2Ij1eWpRRLGIXU7EvBXew4jBo77ZlhLsGNZy
O8hkMnC9+1L9FKf6bi/hfN8O8L9GXcmwxCYq3Z+Se70xM3dxJcvzfxcU3eMr0PXgnXD6WHSRnnax
xbkW13zDK6UBBXwsmQtxXWLnF9/tjjOBrtEnRtzwml5iTWgTsoulJVepCDbHz+11vROcvNI2MlGk
cXJuVwn4l1X+0LW+ID4G0/iR7hfdQIhPWBWq3jDX9Npuk1gfi+8OHki3oELarhQtAkEioi3tnpPa
caw5Yy9Duh0aNvlm2+tOFur6rwe3D4S2z68MHKTPZR7EGbfIiy3OkEhn106oiNS8YM70TKhJ0RJF
iNrKrcJmq1oloS+P4Pi0E6CAFj0GDQOeMO0W0bhDhTRRtwbNSeLpDaaiQUSygOF8jcxTfuzxVgSA
UXuW81KoynJCylVqEr1b8ewornsrpXP+02yzz37N0QbN2nzMK6uUGvQ9y8LhBclmb6JpYuJWwfEO
IZo/f5pnEcBMa15LGmX5nHVgdBIZBoqw57a9EDt0wZPAY5v2xXBcmAf4UMrnHfFFa1tFYyBXtK2+
wizx/bf3V7Ntch1OVlfOW+7LZ/adMY0qe/NARbet21heqYRD7f3k0bc1AWqlEiGR7FGz5hurICZ/
7i4w0G5fAUZeU6v8toD+xgLBB7Royk1FgpBg6iEC+oT9nkPiCFCgM4a07vbCwf1ZDr/tbsawSxS3
UqssURcPbO8KOt8+WL1Ljq9fU8P/w3LH98OZiTJVBxfBlud/p7ZCOIDMm3Ni4Q0on4Mox516ZJOr
RA15ZK/LImdghqvP3OeF6jQ0pR61MSbQALnV+IoKaJy5M58QKDwr2C9V5vZ5ZB01DxxtJed17kHD
xziGqdLpMiKp9ap7BUNidOekj8U9668VU8OqLwOTZHInxVnOFtcOeyy8zOPRfC9JaSddUcHJpXBE
OsNmAW1KZ4OO6Az83o5MyTrR5OuoXmFj7krB4GVqK9SMvhhrmQhLyBqnxe3kiGwvjLKeCxxD1xJf
kGGQGxePIMhcwex/zeJtsN5jJgm8IlzrSpDqSkI/qbcyTebJDkH6viY/Xc4Oa2luwbYPrcfI/2om
L6fpZSSyLTKkfaPGQtZSfU4aMme0BZ5lX8T8bdS+RM4tAwRoU+shXrGFT/EkxzdDsa1hJjLv3zbE
0Q86B4sx8Uov8XNUnt16iL8zQNcLqXZnDAAdXzGTOB/KFAy+7qqFE5zQgEyDuvfqeR5i1X5x+MDa
XiSF6WbfmDQvF9/yvv0A5ZaY2M5K0nf7aRkenfGLLoBm7hFPLBfgQ4mVilfSPI6gbUzES661qEu5
QoKrEAJvTTaLXXo2KbZyR7zhRrk5h2Kz8XB8uH3sDASmxXBFEreL3cdgDnfzK7c+E7Vgzfyn7NBb
kOiiFAH8TcVBumNKTMAUiiCVpcvj6I+ZYLF+hA0OnG0e1W42kUS8nK1tYDo95ItgTPIMJ1jiqhZL
KyxjC0W1QHpreaOdygX8qeBiuc4p1Nhpv/FAwUjPsTGfrYUL4G8vtXIVA0w8v4KadQSTbkjnfoxq
3Dke1H81iz1k1Sb74xIvKPFKXvFIxnY21JbQYALmlQZth0rHkGnDZGDBKYW/JbNLeJyx15KRzMXT
wMoPUJ3Dr0wpMNc+uL7C8yqRi+bU7m3Q/uqMfUK6cPuXaNGYZA07LlqGndgNhF+v1FEdBvut1fwd
dd5vRElnnvo9LBsPMkb5+mzuzf2qMWQKfZHqdhXeVzieAGsQbKDrRsfk/zHoWOyzyIp2sZny0QGq
6QGLIDzwg7EkyGIrtS45Qns+IYDKcvkvL0Yu2KShq8dWrLtONZozyJVfka4JeY5fh5AE4apf4p5Y
sqHL+W6EJVWjpcW/1Ym7D/JpzhhDH0e/79anPSUBQgdW68E+ZqYJY+yKn7bPZ8IyKucs9pBpzCS3
tp7G2oVT8kxoA4Mzg+BX1x3QhrgvEiIAttSsYE7X6sp0Yl9SA6yvgQyXQBP0eq5JrIAhLbmSsIo3
L0HyskEs1afLAG1QChuF4aZfAFQvLP4e4F/0dMpSNBrZWnJssSJBSCu0i3MP+EAXXwvxaMX19+YI
8/nPsx1m61fjw7S26IA6Cq62cO9luYDbdwBo2thMygut7HqNThE5cSObMNfB+ryYVhl5nQykdCJr
ou2VKhsh2/Z9Patf9NPT49R2TAoNwH3HfaLgV1jQyFp8TcJphchGZbXRYkXFLTSZGVCuJiFdqfdj
R1JixkYVuF83xUAo1jdfNDn4QwejD55VJb9RJzMAzUKzohH+X8OlMqPKmJZx7/F95Ir4eiIgEtEf
fCOQkU0zzw+0BdXqhRY7btBx+TtRn69bf8fMRjdntwAW18DucmJxnOvJHIG16/WvR5zdCB+Lf6AZ
madgUkGFAV3YikpwuUojJazNvP0vJk2h2GD4ei2RwR5VGIW4iqca5tHJizP6f6jQd4KFAEnp3fRo
l85f4XapaZoEp2xIACA8e/0itFHo4QWIcJZS8ykZ7Tqt7nB0IJ2kXhRaairUuqPxCwqliUe3HeV7
P5z5ZbqzsvCSyQ4cmKwxCLGmgoMQRSXbrMNW/Luyh1VKDoMhYZbyHYDvcIuiyizrl2xAtd/4VbVu
HHY0KMl/jiaUCurldm16KB9/C4PovSsUc8ccrS1uNogFGt9gjWR3bGAhsLeQ3C7y9hEKa9HleR3F
4Q+N9rC84mPs13p43fOfkzYUFsXSKvFJIeg5vDdfFFMLg3WQGyLeO5fzZCTP8uix0tTbEVinokPN
j7Kx5mfjA4iBb2MtIPWdEnVM/JQ691k3p1EpSyt0XSIv05Nq8bWnyZXrJwWrxSvhS8X8euiZO8qf
CFe+RkCY0dQFRQhbR7VKu52WRJ2tik9O4SDnVIEKUvKlmHI1i9DZUC9sX3JV3R3nHaHX50Q0b31s
r5HM5Xvpcv55C4efh/LPZOXX3tBRDqjZtiRBcAZCh51RF4ppyHojBK4X0EH3ofUCytFwPoRtAVvp
7G6AOoN7JiFavXptxUdB3Igsnb8f+MouP1ybp9zkJI/UmMLDBgWIR5qZyl4XEDggVc8OWCJwOXEu
HxY2uF7ITzUw1e2Al+1Das8+R2gwxYiriNenJgEpQhiGxDg0ezd/881jeWzI9w1ldTF4gV9e0rMn
ZWq7SYLET68Qg5hr71+U67SgjCuKR2jFDt5lr98l15mstKXTbDLmIsqZVREh5XWmlhETR1FFmF34
Lz2kZGlcGU/WXzY6QGZDCL3sO4NTTAWqXSDfO7JfxR8SjtcyyPtcr3pZvq1hiivJOlMdg6jpnEA1
MPM1I873IidxgrqI7qUQWwt6qMp58ZR7Y5SSHAmRmp5iL8eNQFv56GXrXk7OPJhUbIYj5ZVkb0uH
TnOy1vLAerX6EerMGccRnlUw17eRrz20WIoqtYl1+KBjwvoTvX1Oz+NIkucayqmttyU089zOiC/6
+49LAJAcn7i3KtEPgBnXoF1Y7h7O1j3IvJ8hVi9XL8jhs7rdPVk2+8oF/IKKWYFFvAUE7gZNIT+x
ROL8o9CCddF1ril2AUNquNvru+iVASlzvtGgN96Ddb2MwiqYo0Ii1mKoJwYaTw2Lvl6g1oBDH5FG
cxOxofpEvsP894KGhpPg030wuid6zZeEYR/haDL3g7qcH673BEJh1WYZSfRm/p3gkicu9VPNiLiw
bY8KTJtDnC6xFbtZuB+8mzdsZqVgz4qws6tu316giD4XlKMcpFV/7vsfRY00uyg00E058y+/dYCr
RpJqQ4W73uDcXN7cdIbkP6V9bUVczNxBaDbjZQJuNMS3zLkAcMDJpslvJ0z7NmatQI7eDU6VGQzG
RB4C53L7MZnVRfY6jBrk5tfdHKYhivLT9cyzIHqK4filZXVAA4YJl8e8InrKRYl3bqRejYChtPDp
vPCZl9T7/nTeRsB+lsy0XeTjNMYiv9SbmI0tiSazl5ug90QWJ6YeDzY/E0yrQjJc0LjxCiz5cZ6g
lXWHAVyzMxI+zt5aCJ44gQaOGeJ52bwm71GSvW8gIvbTp8L4bPBXda5UETDHs1TfJQUP1ggGvRfH
pMZGkDyN2T6GiqDxzStyNLLVTkbpsR0svFZCAcgm4Swm8cXZv1iYYiC/L6oxaQKzsFTlya3PVXeQ
pq0NYj/2Ktqpqwt44h/5hvINv+5xgI3IcAk2v0QZc/iry2Ua7akT3hzT6lR5b0t9dh1HfNrVn2nY
XEyRD1nR/5Suc13HEyXJbthMBMg8rgd9NXr1gD/EzcCEz+hHqvIWVY2v2RTk9bEI/GwohqL1xAOG
nIiSjKCs/dW+53QAbfuRTuA4geOSifEzvbrQVx2urqRWyVT3WB9fNQCJwq1kZXmGe/2kiBB1jxXJ
SjXeERy/jfW+btZbcZIuOUz0WskBeIhQOi+fr+BcqO/HjD/h+FYSZz70dP5KNjIDCyMMOhMx3Y4U
9efS47tsotuY05FQBfvnXEde+MNidbhezuGYepR4Ey/z2RyaAAfBTdRJK7OwFFigqIOMSWh5gesA
loP7iJZLK5wiZSURUtP7pziujmOtfqSJclX805v3eC+zWF9V19R60A93IKYZAeKStgi092yVnsUN
sRSuhhiuPEo0NSYLX7F+cjmqnhOhN5U5vl+TdJNW1NAn9JduCuEvQLobPhvwBBNkWdeY+lmSS7mD
0HTt07mzeemjq4JjFKHEY3WHcyPaL9T46WWoLKyX812hYD60yoS83oaz2YG998FxV0x4mkQrKZLY
scZXlgQY1uknM0rnXhoWKL1oS5ftqJiaXxMpCO13QV2aUDrOJLaFUHRXXuy2NTaWRrKBWMFgYBQD
zLeOVG1+CCwHxBK/YSoT5sv8xwidBZ7WruoZ/hSzITv0hGm2AhXNcDd40uTbDQ9JKn7f56R8kvcm
Q5KMjiZ789kALfcd6wodVRrJzETYJsmQNfXHJ65+gDM4A+ltCERyAsTJMfbi4hex/NvO8Rt6VIa7
oxLVUlEXtcjJbUszaS6upqMziQRvWKRJ0KIzDaEyposWRz/+SxNttI2X/Ckh432qi/pK8m3vfZPM
MhtAXlWGumqTCQ5jsrPL1qOtm7dtLoDI5Gf9B1dhJq+HRPVS9d5hS48n/VUdWhXrRG6D81Bt9JvO
zdgdY6lKsHFBjecjY77ej6lgn4pMkWVY8i9r7lHbXjYOlKrGR9tzj9ZU7eKrzOggBjy1kwkIKNrn
zJthvgiMVuazabgjjPZKufhpZgJzGvZarBkwYcSy7P5Px8PtY0ga2PR+AHM5+KoGHyaWe/U3/hQp
RbFYzKn9xhjcDBGliw/H5vtIyOkmsl63bES27Zh8RYwcMtfDEAw3EI3Y6nfwv2Z14wDrnVr74Lp3
Z7DZSaxKJiykit0V+wnAO9hjhhRgalIzhW6scvxFsQ0BcRBCxLwFYlJbtJo2O6xUQAp0y3VBGkbV
xoYqkX86+9YJqnt4fghYQpSDPMsxVZazGkEC/F1HJMcI90qw25MRTCsu6HYAU3PoMwcobmyuAPTI
Xce3iaMhoDMc5unfuXoSeXZ/PvZx20ZFvzTRiprQMU/fisn38strnuaHb8Bv8EMyqwPoj0iGQKQb
/oFVva+Mr18tXbRvfDttqvwc461ZNgZ0SzYky9GSBw/b193IO1/WdaHetc7dCNmjdKMyk42tft6I
HUYztt526NNZh8X1dZLZu0O6WCcEy+TmUcoEUTLCzcphesprZhyjHCmeMaDMW2bezj2UqvpiAEAA
n42aspRfA0zBsd5uStCY8NQ/e99b+AWcWVTzK8Y4Y/KnrGFnkYYfdtNgt6W521GcoSz36XCTGdsU
ZlWJI6uJZVngntt45heT6Mx7CrTKi1Tcnv6V5aKBx8J7tMevaW0aATKu705xhiP/6DoYTuWP1QcC
uY1QkaiedPAAKWn6jHo8xoEBuGN438CfpqdrgdG8ZuG+ueiGMxs6jxd6Tp5e1ctngroyB2LKYQXH
MBkhPhWta1TWv8s+p+xJwVp4VhkwCQUr3VqyIvXDRVnNmmJLmZGHU/bFx9gcExllI2Qz5Ip2eoKX
KqbHQTUSRDMsSx6j1znhzYCZeQC0ApkeF8NWVr1eCmQKYcExcYDus7hdzm+CqvO/7QwFf5b7m+7o
CYnFzJlfmaYVEdlvafwZksSalC/FgFd7uLA9ZckGZXhY3XXXRYZaIeufdQ/6BdXduQmJyUFSn7pF
mxt3+hKRrSQm9tDBRFo72D92VV/mMXSUsz1fQxgc4JBtTtvCRkrxIPsAhrYUwW3dziPWGChuB9Zs
0QeETQ3PvAGo5Xc1xQ1EVoYmEjpUgNTENAhYGmEuSFb7RRCYU4mrIgYQRm7EWUsG9tVa/4IONI6j
u2bzLdQccaXU0wp0aFQVvyEx4aojdnCNWmH0giApacz4ngcmSgm8NnYIXF7jJqotj6fwLztMvztx
LM25ipuQ2HqTaphYvURWq1C3wk2S5OaPlrGH1nPNsbinfoZQj+f/cwOHaHbZJ1XWV5xK2sy0+obh
uOjEltEqI6vOjmrr0vjTgEiUHxFI+h/1uIcKOLKUP2JW5mZ23E9KCM0uz+w7JCQb6ml52hkG+1Ot
0nkIUm3ySOv63gg0Q/UXOkwoLqf1kyjF4mLkxZpk7Lifbwzi37FKOphSC87n2OUTTXBiaMWFp0cL
bHH909Hbfyji6/N7mh0iPNDASwmHfnUQ+PnFSHFs8VwSqpySasn3UncG/E4YQggGryT1PXx8M8Nf
Qwp422ATHtVfE9+kpnZmWSh4mSDljD4LTcA727YiOK3Q7mzIuX1ArpEZGuBPb36ac3WCu7kJ2kWE
OIFoGTeOletdgsya4ZTWzl7rQnLapBeFdX1UDTrAItfkBYyxLUv8E40xzdtqlLf4+dJw6OxbFF4e
YC71plSrwv+DvQilGfCNJYmQ2uhevcxEk74CDajdw84d7sIYPvl8lu/DceTeIwSthrb1MRTpWTrS
FH0Wj55d+pZ+SeVYDPwUhqaFUBXTkyaB8s6fHjN+r3NrOqVP8u/DHyjlxdkgYbAWfsjbWSqzEtmq
Vb6QiWoDQ6RdkoX+4BilIwWNd7RtNBQrmMpVpAolsnXjD1t5r5TMQPmTPNKz9Uu8nZBjVJYQNA5F
/3u4Wua+R8KHSgh1gasAzMRoPVhbQWz2wcEFMTcy8Y5hyVj5x/0pKNga6Cqx0pnwUOPnuXp2a3Vv
aCb8qVQqRt4mAAZJC5eqVVxKT845/HzR6P1Qyfd1TyXEYo0lb6Cy/lFpWtz9VBtmDJjUoSPCfIiw
kGUlg8kP/u0brgHMCneAP2l7BWXQV8YA4q+9tXiHjtEQY/inPPVoesQHITHEi8R9+/8xssWZtsbq
OVTlOUkfNoRftOoA7qyB0yQnCjlsJM7uwHMCfZIBo74oMrzjw3IU4V4klalPRfbtzpkYDR7oOhCp
FTmi+3ZyZDf/u6cZUb12Ua+tNpIld5S3lDNIXK5tXDqotv3qwWoMDYGNIG+p/ReupQU2Wehjtixh
bXa3iYDhQnla8Yyr0nh2mZoIz+G9pMtXxzsjbjjBSWRM+pT496vXn4yY6HDF596aGY1VoAhiQIkB
My7629ebn5/ShaKty9ja1sXjIBEW3bSRLYp+H+fl5OHFNYBTVSFEWGRr/CycS+1XNIHqWjXFtacC
6peNJ7kc8uwHA4qpQUQsCcMNSNJxdFCRaMuSGLURgzmgw4Zb1eHEpoimUESOL40P/kW+WVhg96Kn
EodFo5LfEvDJmVeOR5ikxYyXKM4OGngnxF8+8yK9bN43LBe5iDmdKeyLBRktEKL/WaJ6WzCMHuJJ
tFK6HUQXM/oJQ50IfG7hMNfRKQGsRDoW5lw1QGtrWWqm8xtFhwrXanK9H968R21Qw+RoHSjvcprC
RpX5tRJ0jAiaiXUFhJEbC5kyk9eDvMQLdpmnHO+0NnwPVfuf+XkscGPulP1AAwFscDJvzgwAlFGL
/ozfjYTLbC3iE/I3NHj56t8FT3eSBOjs5OS/Tprf3RARYPHKB3V6HLJgYyLAKsF58Xcw3GSAeGNe
zosQtUIHRV14hfyprk1lQ/XnpFHTUAZ9boCjBl9zreaBQCBoKjcDQ+FiwAw0UMZ3lKYKEXGeprPu
5UVFgC60xW5jU66mAbmTv54p63emWhfF+6MKmZdMFZ12LKBUnXRkADCvdsXoY71FrdmGQaj6tjfb
0g/u1vmo4Y4cbXT5h8vvB2AUP86W/5dJDRSUPeBZ7hP6rwvmnwIqZHcV08B943SGt96fQBFrIz46
UhA6yp4qJENfcCAY+Bgbsiw+NB98kL4NL2PzGc2PXpd1N5eOFuiCtVSabyn015hGp0mrqqUR31p7
j61X47hUaFOlCdfXw2wK+N8tVmP0UtXRN+l33GhMcxlkzxwEW5ZH3Q95ARF2gyfv8LFP3f2vkf15
A59fy7OB0UoGf6MHDL2s9Zy4sJufpaGrjrRk2WKte7iPcmmY6EfmUPbSCB82Rj6nPZiy4iUpTyMB
gVLdJ8BN5qYP9S5hK8kXICcuwGrrlWTVeBw70gexLCcWwGE7P8YLKZaK41rClWdyGuo/l9DYwwYe
upzh9ch/4roDZ21g/eT+O4VYPU/hfneSDAZWCzjcPVBFCLcq+FkNfFKg/RspSm4OmtcOnsINEcCW
j+2NGUWcQkpApPo/E3DJV0iHnCgsuLgzvc82orJ6VXZXEeTOaXs79n1GC0px48g0B/HFmTf/txM6
WGIE7of5KlMzL4LsZSoXiN2V8TVl2tsQfApU6rOyD8sqOZIBSsj3Pr1fzDF1PZqbj9RSOYj7byIl
v7z+1v/jM3XueDmD3yqbSv55/o6MDh0vTMdoZF33CHjXK4EqghQ9iIiCVTdi8NLJ2BKCwdRrF0ZJ
AGGNhlteWGSKGOG0gkSR+rrdCMfGh1F5IEwsyPw5vUvlWPeFTP735z6arw9i5MOst4q+Q8IU2lEu
ppHbohEcLIF03yKWFPLGxCcnGrxDW2OSPPxkwbl0KpHkvsaUMNv8DAGvRKQO+PUFKqjHggt/zvMT
Oe9fVZXOOGTYO1bFNd0PLv67ENOQD/anpG2bqBCJ+wb7xKqwQMFLEYVoUPks2BVWf0uK8iWQefpn
no4tkhr3BlZvsKDz9W79R1ET1mDqRLFtkaeNTqURaR3DvkJTMFvVPtxDl4tQVSAREbtgCn3Bbx4H
EvRpELYcbkUa8z/43+5EfP07WTOyKxuVFRHo9nuKGuJsSr383Hmv7ir4YMR5hL21ArqQDGsoxBIp
Gb8GO5ZfsiJBRS8junETWR7GgOtHZSrdfzczBqm57tzELrZjhoo2w/Zv4+ZKRjysz3DJtO/3R1DP
Zwa3LPv67rPLmwVk2EvUDJaJYRZJHHUA7ZJlxdR5m+3JzI6k55IS0BUszzbNp0Zi1gNiHlvdkHiB
jzBX3IwjxGGfffAXt60qFI4U6vlisrERNWmJeWU564HMxvgD8ABU7rCgMm6ncRHYR72N6oc+AKQb
3CroMIdUo+nbHyzaBgrx68xdpXV/HrE6ijTHUfHMGjYrU+8NJbBlDGBdeV4z8xCf6s5so/5fmHLc
RK6UspHpUWfaUSL46g/igQqJjzynLjUn9hFX4K/Q5ITRQ589aoZArLatFg22YPqccUYQKpEu3tea
eR9FlTRxa8g0uGlrIacoubU8AXrHzIoCG98T7HPE6TjUI21Q+PErsHESxz2/milZUDVAtUptfAH9
CUHFyjt+7cdx3qkz43svZWBjKVGzNjtxcJ7kBriZZOS7ZmiJD5hROhaUnfXH9MIIKVj+PPVakuQe
Flk+4OWpDY/rP6KxzwFUk9G9uMR7HFWFCaSrD+zC1TA2YkhUS2ixdPOlEaD37ckGfLyFHVOrIuEo
3PjRIdfj25KrAbOOAlYSanvfbxcgmGeVF/5ut/xIp21rPTT0wak906JrCsu9v9qVESPV5RNAD1tw
w2aeBh6GOynOwlojUhXj8Kf/7IAFVp92sqhlN0dg3HFfs4fTGgvY11CjjsmL3XDUay2aR5X/7NyN
Lmi3KcgA4Dv/fFgWGZRjZInJoPqbG2bmQqam/02jdD6h7NDlQl/2P/r0ZPDF4MW3pID1lNZcG+EX
dzVYuinhg4t9PWRG53LACjATEKKit2rZpq1/nfXXCVqyDczCTzWOW4vCfIYD9aFjZf6PzTK+wyvC
/iEb66G+78rvy2jHfAuidLNKFL30w2WbIUnXotkhckvGKw7mDDyFAklPtBr6H8WrpBFPr3fIfZ1f
IMI0jJ/dsT8uBab55g3dAnw8A1HiSVhU96Qf7MN/Jo2VhUOFNyEjqXI2JCUom0AnD1G1uYavikBV
HRbVDXzo7pwxr0fAF0ZmvrbpEeo8rY74ZIytj8r5UOvMUrI6Z35ejRIFt1DrEbDTZjgO+6owoFVA
Y4fqQzs6MrCOvuRPMRTHCyiAeFHn02REfKGuWs+JTz9TnxushsxkVmkz9boWjqonVpwCqecQZGj8
1Q/4vgKwaNJdbHeYg4GUI3bTYzw+txmjhVJoatlE91P1fPUzbNaGdpOyDrFzJRXk1W89fNOusPpO
uYxJdO2skdD5PkHMA/bZE22rR00zlcojSuESgCwidxeoKT2C0o4ib8jEm1sC6iuTvV6wpRucPrbB
XqLK/mzOldqdzT9AYi9sHzXQ/6c7yak7WoxDc2uWOW6Ieiy+ihhPkZYJH2O4dtnmofVPR2W8EQea
WYeI+CtTK35qH1sOpUvbksLtirmJpa96XNhp9hBGsJIOnVBoVe35+vbpJV9D45PiVafyHpOrxsaZ
fwuFX2YxpcyYtFeTtr01cAXpQMZTU7NSNPJosM6588UG63YN5FwxuzSF6aQqeIvrwhs0WkVsZnzI
u7iVDOWvUiSNnwvz6uiUZ3Lcqi+SefJiMX0B1w2WoS/qNLh8gTc/F5D89VxRbwnBevAIqpvqupaS
T316Cd7gLiZsupPySc3EZzd1j1F6tZtawc0GuptfnF9hQCFubC0WARfcHgxRsPlgQLUCQYNigc+D
oz/zr+OTpeLzBQIJYTOjpfC+8f9tEHYMVDHKzmuAk8EiZ/Dl7ikF0GTu3Wfex4oML/M56F9TurGV
wNTF+VdfhPE3xdFpdpatQmaNeNugrqBafhn/RxNeBtz5NPohjsBLBYHKh4K1owiKzroJvyTwiHe3
dcN21omicLBPI2dPnn7P+l9PX1VR0cCwiaYnhfLNjW4jGSeexUJYhn9MB1WX5X3Ryih0KzzQw4Kh
xHW/My/WlRkKiVoxeYFqNY0NU0shVof2ygh+r3xJFexy6QaMiASyH39GQ2CUFAd6l8AWIHxQVMDR
C7BgEAHUw0hS64kfTsbGhOnhxMrSCYEPGbdxLEvtzrXRrxK8sG92lBPxyDqyqWXKUd/hSMKK0TuE
/0iiVXypdI/QLECTlhyKQUz+1s+tzu3gDRoqPdbmOZpVJvz6y8uIJgo+3zQ1ww2yfP0NfQ374pef
h9FCGjtDkiDpJl/uh6HuGxzBDQe6vb42BE72aQjdkm0V9fiBQdjoJBXwu30+tmNXz+Nn5ULBBkV9
+d5U91hKznekQQD4hFE5l693LzuIxc2bs7fWjlDLX5+2NEh7SG7OOYnEWlwkwXPlP4yG4sJYGo/o
LHa20rWDgfKyAva+uRGHb2tkzRVdAmAPyw/HDsmI6zLOwCVQpM8mNUVxLnh5Wiiyfl8h9JzwpsJ9
ANgsZg+cS6rzIlO3AMi2Vua3dYrg35Qp4XLXJ6gl0IYl5lzi/V6zKNSLEG3lmnoBOJultG+hmgvk
SvrdWG5AxiabrWJDmQ8tbg+Td63kDXp0ls3a1p2PK3SrPgP4NEPnsp+RGaZLotG+zeZKDRXUrLAl
G2k9kW5sj8TtY8YjCpOymbd0p+tOISqWJICPfzKr/ojtNziZ032cuUFJeJ8CTZA4LIzUgljM7Mk+
v0rmfTKUojNi8JLFtDAz4FPEylOjiFphZfHX7cCpsFT8KaoM+Uk2AXfKOcxNrXDwe8XNyrgQKcEA
VYf5+zusEwnEZmB+pdL5CrWB5edTZBIYjBoGjBYi8w3GN+IkN8yZbMfuybeHskeskY8kVt2HaOHM
DfNx/ePSsz5xid5/fgiarg98k+zt6pd/J2ycnI/TkV9H8mMQfTQ+JbfcmnzvlmAR12WuFMClBaRc
2RgirZjcGUiHdzKVpZXuILGdYJl87CJCM+y/lz52oaSF3J4GBCE2rWKDcOHvSN+6g53r/eRQjZax
F2UnUQbLfo48wUgtSOLjwgdHbrAor0ZINk2W3gs/QbF0wBoH24vY2Tnz6/wPeV1YcX/9nvBw4SLK
Rp+Y+VMATHBmEWPdKUQQqwM5c9/a4ZR0sKjJlRiw7R5okcy5eoSkG7P69qfWyuQ9uWKaNLa+fc9m
X4I4VhB94a+MUVdmcwwd0ZrFsjIjlLbyI0OuQoCOO8Mj0s8pMdIiE3dSznMMlr4dI5XMMYh3A9OJ
2VVnPoV24uc0tLot/b08+vsTnfiPQ+LryBHGFGaFWdjQH7f+2exYNVi1iWtE53kHmXJqR3GkWcXp
FB1NkqytesZnnKWSh7aTtotUqeWJzOD8otjF4ESFrPgNysewee2N+P7jZ3c3CmZUf1FCSL4f+unp
0uifDhXS1wO5Uz3xm51O/lcBS3zTZtz0WxYj3C73EH1pkPpKMTvifBnskEMx7lPtvcGrpBco8ept
2JTB0mTU/4MGHWRi4E2meRU3fR5kZ5YeQ3RYdZAg8U5gAKQ424vbzTHLxFuzcmh13EAt8u84ksLT
akkvlXl6/5F9KrNk/sV4TIMwDM1x6ybJu/R1qinh9eekvPKDMrtvTE1ho3hdiSaayg2uaGjdcJrc
XtuRLlC7TvRKjn6SaWLP/dvUU6RSaArp/pQ/TMtb27ArVj3OrZJbPEN7U1Iz/1Vm2Ho5MsUqM5k1
Ba1EV0RnhQQdPnCnc+Rzher0fk7UWc48xFXxKhIi2kEyINV43QHTpmvTM4LhUP709OS6rds4VL3N
NUubwE/MEPNfEjx1BHCbEQeudw2JDINmaTQ5iIKUapr+6g/G7jcu2qON1+710KSsGFLqTRg99+cv
Mkd681mu96Rb0RivAVSiRt9Uz/WkSeHgLjXX8Psc7S1bM6LxfloV51vf0fyylB4Ij9TdjWnxM+7U
sCG8vxIhycFWdd1LqF2cfZZB0QTiTpcsSxb0WOiGQ6QBSjur4D/prEMQQeMLUZZ+oYzwx8XKqYaL
BRfn5CePk16rWnTu8VOPwvh6/2VqrhT8vZ/GuibdLJM+RhnxAvquyp7C7KgvfjhzKZYMiayHi454
w6XpaxIxM0eZ8dWd/a3F+uLMDXpwacSBkiu1qhVPGLgMCixebiBINXu99cnlcM0B+fyKoGoogA6o
2Di8mjDEcka/eVr5kDQeJPe4vVE89wR9WYGlEE7IBtmMUq6DDjXEjXv+NhldiGhK45PjoF4cUw0H
EeOhozB6y1rvVCBefMjQUub/J6xX0lNLHEN46bWk4764Z4ntTgSg9DCd4NYZjjCQe2TLPjG/bkNj
8lh9ZGtRhZuT0i4OABb84u4dKiK4nO+0RBN7mcZ+sUGCfdHLYvQaUGhpsegSrVO6m+qxOLSoJo6U
gQPPbPQElyOQ8Yc76XyOhpodLfQNXzHvTUfdL1oZ2ZmanjzvDk/gLRijKgh+SYFBdk+sK7BlhMLC
HFvc9UVHQ17O9S+gdqBTELa51/yKoJGk95agz2m85YsjU1/RWU5fo0olgvJGJ2rWQBNPzCqFkcQM
+BxTho6Z/a1AzyYQbArHan9f7CfeM33KG6/rxrSSo7I7VIcwETTDH24Vy7wbbtzqm5eCEE7GlNr3
9hJ5sZf0KFvO9uBdWc4aNliv/i1iP0NYQAcOkdAxLujlk6RsG7/C+TKkF7MK9tw+IeNrJXLlA3Rm
HcBK2hN9ai7fr83GNo03ZJ7bJShdjHB9gGyYnuwFsS9OdpGimuj5Tye4Cmu2r3EYlKaBmLNWxFg/
Vwhx89vf++Wft0QKm+eng5F+Wti6mlWjMsM0ChLCyX8s/zsY92WN/NVFf00THsley1pzq/ntBJS/
mjyRlWzzzvtNiEsU8OG+4dx1N1GBzVnCQyiQHaijTgXn4seNoabxZJSMcS0HtUnsVn857OkhK74f
LvPxBYS7HYzQN5C1RbvzqXKIyGdeQ1R+uxlFbsUyTSRPoCv+OiCREtA5fBBAz/qI4ZtgYw2hcnmA
rvUZoXjOQuGz9JHW6u5RPP2L3g9EGbcB5Y2h3MtxQ7PR0r70DpiAoXPYEWA0EEFdujcwC1Oiche8
/NqoqnswfV73Dh/GUxqZbfTLTMQoCsno5vt6TW4Ks39aKvk7djtYYuvCdvLP7onrnU9eS1p37Eq2
fHMRkjIkACD370KDabT+2Zg340mOPc0OLsH+IrKiLvbZvG50zUUl3XudA+0Cahh0oUFzDmrOmQr1
4W5D4rwmEtTEMNSwMLzSHihzWb/+T9roZU08Ip1zq9clrvw5PoWe4VdYK8qXlaph4tqPZ4ER73QE
V9RNpXxngxXWmhKPCsazWiyTgvlkI+D4TvkKaP7ybF9Ln+FtAtYl1t7kpkVarHGE8tuyEBgn7huM
ifzb8OGk/3cK8JEIaxjxF5n22DiOKRIo2TuKXF5CFwcn98Dz52u3PiQjeENW4TpYIOsn54B+Fx3T
Ra/66qf2QecaHzIuJiI2ZGJoLiLYC5kk47dzXDYnw8UqejYwRgjbfdAzVZpE+VHj37OESmbJCZuJ
HSpE0JteegAH6v+9KHj5LEt72T1tbEhihF8Svps1vJrXk2oqxe43Gc611V7E+LBZIJpu63qdniNg
BOIbuoQvMpHpdL5uFOOD/tNftDmti9UsqyuhWZ7cg+vhnT6uw39heTSyPk2+8wIUi8XByBxDvYgd
svTyVQoBENXVYSsr7GTWMINY/5jDfTtW7untwimZhX/Gqq9WSpxEUcIJ9ckCGMwyqrnZoOH31B0q
M99VnhcZQpWzqIk3AcDpz+nuAZhYejuQStXgsUqR0llNb4nLOw8T164Q8gtXaSnQIX978X7XsFrr
jAwFLVyKUEFGujG9QSCptAMGDCEJaV3msN8rWTZUfGYV6v62dhezYYjtmAXa+9t2UERCzxfRKM3N
CoWW6IFljeSjERJ3poS+8FKc9y6K7jg0rL+lg/8MZc35bDaCB/I8xU434V87mHfcTOaAe11VSfbi
rPQbf4+6VdHHgBUVN8WiHbMFaHSn+BHDo+mx67W4QcAUHFKMydgYglaRb/4VfIqw3OFg9c5rWSzp
LA4z0V7bvSOfCMjw2h1PP4+EuJ2FripIS/SLNtn36s+7eZ989A4Gl0o+6tnwCYZs7PZuee9GrbqR
ImBhABMP9vCjAeAddBJsHsj+V6jto21L/mS2sw6+yKsoUTIEU8tRL/vatWGrxfwOI7yxA5Lb4nHQ
DN2duJsMQkWYQKaIt/FaZ38ouJepZAuAY8/tZJk7oDkHG3tY9KL1OMbbEdRSxaw6/eX6s6rGjf7g
+yRVNzL5satSuq/RmxKgWkCQmYDNVpOEc9BUzGEq7L4LlD3PU/HIvE9PfOAbdIx/qGsOVffwrhvn
3HCVxl9ZgI6w9ftkknQ2JlglWP1ZbujdcQpefODD7uUicGAnuTp8q3n+XM8eR9rTCeuGYE2ysjIv
3GR73XX99zgScBQWW2Of3SsFXI3I14/0fdkzRSD0WBwZfbB225vw1WVBp/PkE3JlqrvzNfGa2U4M
j4j/oMbapE7ABysQNzSjzh088KUFCA6EETuLVIjlo7cTv/chQdiNkiBia1vaZDDIHQGqLfY5NIbX
xxuoKGDRU1R0TeKQzv87aQ4D7EMdSceDL9O1MCO+ZWRo9hnSB7NjQv56MgJHX5huJNPhNxz2TI5l
ndCLkSl9lfdsKbOuhyM6jfBm8K9WFF0B9F+CJI4CZiqtDXapjjkRoKLg/UljGdTtkhXYDBSwqnB9
4rfIVcAO0plUl+bFlvzE/h4tamOmDNvuXBvquKSmlXsCdqk2GB43hykvpmJdRFTMeVJwICFi4aTG
ywB5IDNocjLnIh7ODETG4gryh5wNwyHugyxiAzixHFA5g2doI9lsNcq+rXmgnNOvm5j16uQtGXZv
2JT9QswTWssRyCNj2t5UWBHQ45bAtSceM7TzBEhvC1fE/+r939xUA6Qvi2elktVL/yGZ77W4fi48
TTe4kliXzPyjkKxK/BOn79sP53tNFIDrmVgJ55TpadutFevyKCDUJf0pjBjZL2yMaCeusZD2xEiR
yXWZLcmei0L902w5wPH2LXUydrfnAK5az8GX618yHTckq5JXLhF6ZtJNIsYeUDVinrcYJsQMP2RO
trgZk1KN2SwF111q0wQxNK1rLQEz+KI3+nKd4eUygens90IOvxKKajOwQKQlkcvLxSbOmYY+vcO/
UBuuEt81ozdXB2E4t3L5ODIcqCPcVQRMpCpSRwBilBhGHQ40TEv3mPcaImUcZrGd6QFM/5xBFMv9
yzGB8rL935Rw3MSNcbK8KWgcfuxr+xh1YRXXpXnwWP4WJ6yi0FnIXSLRu+PjwYayWZgifSz9i0pG
xlFeRnEyBgjrR8MAuRGncgdxSqVBbo1eSxTx4R3zr3+4cTmUE+wJkMNGquhpq8Y3tI6wZ2+2AacH
F+c2E/kCfkA+AR/yk+B5sKyTBDcAIqAANPbNAD0+IFa5EGSzLp7h0s/rE1AAHaNHQBKj9Y5LoDZF
/Zz24KsJLpMQj3MM9Tz1z5ckQr9bGdpv/f+nWVP32l+BhPRN4/dSTJosase6xCFkO/uiagGKw/6c
+aAA01vid0DzpLbpmqIC2UJrzA7tt9OEZsYglcLi0ue/I4dGzLyGumOR/18naq1cr2a0rF8X0a/9
F8xrrbWgqRgZ0rAytL5OBUfGCaQJpzzXg55Mxg+Yhdo38d673Plv9cwSOdG0oPHgMQHKRv4oiA3K
QxD8EfMcsU6UDEv+G/cnQjcYgeq68UrNVnl6b9XH1w45SGolfMq9VqrJW6xBNfgLHXPGhn9TmF/m
OTHWgDZof2ib0Yyc1cw0il2pTaRB9tG7uuBNOdm6YIXNKiAn3EfnuJOnXBCsCAJWlNUGFVIOaWqd
AXE7mD4/PNdbB5ThGDjB2MKNBQ+yQWEx8Cge0FnfzmSA6ZfDobnA8v4bofKgVmdKF4SCtggFLK74
JrqDThyztbAeZDk6/HWXVIjwy+7G2rcXKuAeh6mEsYkGMaLg0afZg6L5AoiUUq1F++UHV2dxjUHc
6AfiE3ANS1Zsulhp+hKZoYETklY/+QFcmJjfrUYYx9NN3k3FCBa3Kb4QLEu8Cc86v/cCDxdYLDY3
a6XVgCc50nqTWV9OO+HtGYLEnxo6tEYky98mGGa+SGDNFrhADvOukgMzCkW5qs7+b92GyMDT1tL6
kk7BfacaPCeef+1S+nenlBlaRyCQLJyKG015fRd05+2BTcaoXrsujvFK8XIBn8tjxACa/mrAjTBD
3eIib8vqf231sIbgAIlA1ildqTIgsoMWOG+zhHkUN1zPsWWXOcyH1O7KHJlowgQJQYGDwIO0qTQJ
XQkjtpp69VbRXrqsM+7E+Q3G/BqENn2gIySkYLNJDkYUAHh1Gi/HljX6JButJuen55oT8HIL3RPT
5xbDwrILg62iZbtcDCnAdz7Sx/L+rOolGeS/i0sPJEFlOk5BrM4y5fPqZqGbm0QkqIMv+PaqPRlF
i+mrqbdrOm76WCCxtLF1HQ0Tne9XXry55HrxPAkVajzlgFY3WWo+yOCHRQjegq+fiv8y+3vDZYSM
XAZfILBqOiooH/FnHPvwCA2qyboPbzwdxY4F6+U5rIdPCe9FxG3B7L0pC4FMS7AzrDvRG64PBTbq
XPqTwYWoyi62JNMOc2QOcIlMIQXrDYF+9XDDmXusvtLNYgt0QL8k/v/hB+fdLHDGG2gq9d89lyeU
+tqFgOrSU9reJxkcFPfZ2YoHc0q/mq/iUuGtp99EWCvxkaBHrn7dtXiRewrtdjNDOUG8Ghk/B/A6
yawS8uHzLN16U/C7FHxWiw7g/rjt7G1b25rhF5YVBGCOY602nEKXklo/4+jN18q6H0/BuojUQISG
xV+5WydpE+2YP+onVQZ2DeintgNj7OD6aVhwVGyuAfgDZQDMsj3A1H3o3ENqa4l5FI3RATrJOgvz
UFYxKQ3byHTez07XhCyauDDx2KzhO95Cf/ZyJCUa+Aog7jsMo/opOfWrDwu9nzUTDUegtv1VqZSZ
VKiVq0fjR1s8FRQsiO+bmsV+zKD3HvD6m+FsEEGM3x2VtC3r6ltWn4oq3upbKr7pIe3cOATUmNHY
nPXzXY7l3cZezjwoxG7VruPU/025bHVbrnCcymFXHQ7Vx2/AJAh01K4L7VjE2wO7WRQk665EjfBX
u5C2yxKx7D4X1V1ZRV53azonIknEwgH+je65Lf1YJ3upFvQMT9nuGFA/z282IdkpxOpRPOsKv2EP
/m4ciozeRsPSe6c+8uQN5/ltJLJ/zjzEU5wcR/qVnBMCabfzHkwc5wj1Z/2hTiRhBK87n/DOwgSm
tS7xslku9Ql53Ca30H2Y0b0sljuQmUTjqhurT1/z93dBAtle5NHsMmi87Z5kFmUx2TMHX31gwOdA
tWOs1mZGqqfe6i/QNzRRzhu2z/vtX8oq9d/HILOlArtzisFV6DBBpHwwC9LypJ+UFJyL4tZVHuf1
2wxZLP1uG1hf55dcHXuubajecEK4vn+Eo2Te5kEqOFIEhdG5+XNh1RrVxho3hUWwyUFZVMm6SW/W
cAIBZKqXxfmdfCxhLvcel7uauvS3clOSihSnAaCgiPKZFJKISI1OU79F16mOR6uaFJrjmcI07Brp
kiFehkAjiH+jfMnMoLSxGmBoB32yiWvkheXrT8G352dv3DEUj2kOu7X4rUry79j7h1vNdOsQ1n2b
vnxvbopmSX1H+eC2Awr9W8eSc4GMLRH9WpbAyLyD/Uv5Y4Y24HnoZf8x7ujkqN3v9kpksa+vm/f5
CvDWaFq+NVbE9BSoRQ+nOH0oHOduthfKBZbksE47T9Jv7qRYo4Oh13U0z8daR3GTm4zlsNCZ122a
YPEberdRZllYb1A+o37RjApXXZZD2XGNt5mpU1FRiC0SB6RV59c1P3TDf3JqVIXgPRMjWfzrlpnt
aCMiSV8AeTNzH8jUr9Wj9thepMKgmO7RsWvQFQ1fUTXb1G+OVyQnp2ux85e9K/qUvdey1ZHt/WWx
abgvJsz0AEQQ6S5SLE+uCABZjQ35TyTu9hgZkpx3WWuFaRDOhXOUDTOnCwvYTJMvYmo0t1YTpUM+
ufNA6YPA2K/uy+u1CNXQJsXFaU7HculDNILyOFD2ZkSkbl+CntrnUD9WfkbBMOcuy/HJ4WmoquoZ
c+aFq3pGJ52P4yFq2WLEusuUzcYO8iM06tuDreM10wTBLbyL3ILvxWn7i8AA1Q79lCexj9e8mJqh
b5vc9dhNdC42b5O87bAXvC8qccdkHZpWKPOwXsfNfgsf6e+vlF+TsmlKn+dM1ewHCXIQMzzaAHk9
40t03p31ea1sz2QAXSP2iuLAJmmyjplCAWC1p5HVzhmoA5bEoghfpQvfax6bkYLrZlan86vxWCRf
Zrpht21OpsSqEo2kRISroTkmtxpJ3+lB5gn0zmGwuXDHR2LoOHn8gXGvSOKKx/5vj9mPbd0Y3+uD
OSu851Kg073HY1sK7DCjpaK892iLErtY+cNJN9v2bdlc72uyL0qAabNj+IBPG+QR+F090A1FKu9T
g+Z9jHzPpnHxoDA1bitSFNAo36qCb3KkGis6RoTW1JLmP2FLKG8TvZW1XXIVkNYebe+mr8YwY7nu
IylnG/nj42hWjzmKhc4VGNMdPe7+ElSRRR80uZSvwZSkPREErjW7CJnhUJR0uxcdM1ALHjytCWN4
36fEnmh8c1uLEmypX7ZRpy+JWUkoNAaFe/Ks4sqO/gj+q8lNr9Ok5CxUk3jl/P88fT/jmr+4LOQw
WxJsY2y+N0uz18Xw93THUadie8BsyfB8KRHhUkJ+hdCqu01XLmNokcNnNKL03SBx8h+5QEsIh6W/
MlRsxmuNoZwqIPqGWvy/ekzkDGHrzuJ2Vihk04oclJ3w9NqghoM4E7H6BmvQTEPdSwP2156y2vMe
LTqXQ14jHdKnhEmSu6xK3cOe9dnWFjw9L0mWCGVsu2Jm/tCdi4/RkWh1eknspQ5QszEGKtEaNm8m
+p6kjjVJ9LcAGr4ahdte6sMwzG2bhd6+zHg8sgG0Kp3zRs6svybUrM6SitIrxt0G43CgvyETsxm+
+95oYtVeWsfVADSmRpk0eA4Zd2y31xY2wxh+wFPQ/kcjCNBfAzSTvRBZawsiHpeP5mf7j81YafwY
iaOCupe+sqn/1XXgG/RI736hN95pQignmm426k0PhX8ePT1bPatndoI66pKoCoQoO9DUxKVB9cIm
YMKuGuiJKqMQ52km9HzqkE+MiQVSESmFi/5g7sKFySfHMc6FZDObJv9+ba1ZQmGpO6DweAaCEC9+
QEOSefmzqUe6kaNEjfm7ql+S2kK3FtYp3gZraz0NG+caXHnWQqU4fCg0N2229XaXq+oxEprYUqi/
HwGKm62HvDrPCNWmXSR/xTKrdi2z4ULtvOT/g2Ost/NPE6/Aq/Z6UHRXk/et1dI3FucYeQU9TFoH
SBzOxeZB76RffsCbT67yND260Megvfd6MOfOUIunG3CKJwq1SYxBilHj2F3xqBNgmKWAx2+pZXge
py2usocEy1CZdpYN8i3yC7ywloR+S4uR89zduVcWMbUzhLZ8yur2lOhpaAlK8wAyjX0NJK0c+xyr
pQil0bXyepMl3fglqDjpWhbky0v5GYPMIbdQV+cl+u8VuqRJjDGcfzRAqLTjUeIGPeSlcJ2/SXXn
9F9Qn1V00ASopDGLc9CHVBl/qMBd974i6E4MAUB2Vi0xw2k5/sfKdHGIQSjCDec/CXMHs7l1b+iK
apsgWbdV2A7c3O1W48QPpjpMgH1vu1VWOqkaOAeaG1d5ehw5L33N0/wfmuw/BZIBDQhQnzOBZKCh
edjtxP3VCbbnkqol+3Xte0BHKMw/vO1lvCLh7yz0frPmOqfhswZMUrabQsNahseFSQCCw2+K8Hxn
xNZlPLMT+9s+V8i+IuCUDW1HaqnJZAXKONrdS8yc+PAB1ad8EGSR78k4urTYGcZCffxR+7xuv8Nj
/L7Wv2NYSqa6t2MFPdGxsxe9w/ef1j4G0jf4Ittcc/JT0TreLRhL3Zax+9CezmW/vpD5bzxUIFUM
jfZVivZFjEvd+LuaM2Arg4hcjB4HrfEfY9CE16sRWGp2yd/3HnQDnIyGroQsiI+zsZ4ROtC9s8jA
Iu1ubjBzy0ALMhELJbXD86TCAH0XOBAmR9ojngWewSms/AKzMle6mfztJz6tqVgny6SUZvIlXFa/
O6ePNpetgUUPgWG7H5Y23t0clUDVYUmQeUuWnLoLIYzzcVIlCSd1gBasUHuqjkm1nckKGiJxPTB4
49+amgzV0D9nNz7P3mNxGzEKhTFuvpmRdG65OxWT+GF0HJdXpBQeFqpZa3LYRhgp3T27wQxpS111
eMOG8CLdS5I4A7JzvpYA/XV2PeR/llbFMfyVAGZuBB82lKogrdatMGaBwfu5RLvhAGoysrVHyYFI
fAsODHEjpv03VcXfa3/2QzdBhOZh9DzdEQGWBS/cdsuLrx8PHTo/8NfDw48DrQARKhAB6VXLyEzG
WVVafNdfB/A+uG3/aP/cYF2F+OHzQ7vyugTDbKAtf/KZYeYMqLPX9h+QXDeHnBp+PykIsHaQa73E
3WTTvAaRLpm6Rez9ArCwqMdXHvLu46o3G9OpwWZEVnIz61jJHs1jz5a5N6SQiBumT8mzgT3B67HA
q7R6OgRH3sTIyunsmAuYti5QHM+V4gmu5OsHub/C4MEY6iWOR3Cc248q62I+LUXhWSYMVvv28rwz
jPuXm/cFoWkankWzzUuwJKvoBIHLTyR0YTV8soOqALbP9ORIqSmVql4Jnexo1pis/iHNgqj7SDLW
CAvkblGQk3G7NVrEsCdu6xSBayXwemJNiT+HdYhjhjc48lpNWrpERZM1oL2WJcuqABSk7i75YG/d
jEvYoRyo8rk1Io8g4cx3G4xrxyq+/PbEetSkGttHlxWF3FouHk8X2jvGy9NJTQsftHZjf358o02v
/J41sLxCubvCiEkicuFf+Oeaow9nZQjs3hUK6+xoxkk85tsnHALk1vrr0Uz9gBNM2feo6NgBiiVe
Cx4pDiiDgh9zTgPEW6HBF5QOCro2LZjyHR52oR91UqhZdnKmY5mM8sNNXSL5XVmeUHlCO4rVgOH6
i5tHLvp/RK3311Wl2GaJwu1qK3pn8H/oydvpcKeFCNvamGSN/O1EZEgAhlhd/abw29SxjdICNERr
WS0C3EvPQ3EjRgB0nzMcuDOWeQdkyGOTz4IyRnxwiyiQUdIiDQGVb5MnNcShWJdzS+7uqOybb7HR
o8kf3PWPeL0xDU6SSTghBJ0CA3+yEfqva9sbkBO2ICfNfyb4PDdk+ma64wPuCzzzwc+UWtI+7NMi
3afgKAsCMLR8OlbJDhMpBX4tiAbgdLWJn6EqWNus1S0udAVeNiaeoozqZDRRo1w4yqyCFxBaAZ1Y
PDk+v+fYmjO0wfHQCmRsogufSRA0Beie/c4xvc6gQSI85+H8mPQstR1vWLI6coF6Dnm26rprsNs3
/+wrpzTpgyXreP2G9lyNplXj04ccfQOKlH7BFAoTtoLf1etP6ZsfISqZaRa/K5eejJ+Z9sZLy5wL
T1WHJ6RsZhILj3bEUR9neg5Vrha1zZoxmduREy///2rZmPGxQm3l3O4UwzJxhD+FJHfjqIayKT/M
PTz8vHrtaCuW6JoUhHhnMH+7+OCK9dIvRxT0PXkeq+kfpLJLiK0nGk5QIh3iN1qZT0MgZA03zq6e
IVL5uQMHeL2a3c9QBEHurC1IfCrZ5dKgvRJXA3S+kx8vqMcU3YbEkaTpa46ALVMHqnfgw3zrmLOX
lysVd3xCi8Znb8oW++peiDUgVVDkE1fQv/CgkY8kPVjKn9ZOePsQKH6knOy/Y1SVB5TZnyFJbNPN
Hx0/TDzj3RZetNep2AkxS0AtiTtpJenI+iIYnZyWXBySlJZiZZbRFmliwHxuonYC6YTn917zHIBb
SLyNjQmDeHB1eTSNCcyJ20jXmlbMpFhXqfTPCA43Mtx9okdvsmI6UbGu3dgWVz4jc4g5WwLj458q
kDsex/tCV+w1O2HrW5lPUb/yrqq8GVhu2M8kHY/+cAywagYo25M8Gtob6aW8nzspRgnf4cTDco2u
0tWa8/nBdUb8gc/zBdMYUr3mrtV78YpIqac/ZGg42AZMgIld55AnsYFn/xFIPfedv1dwO2J6m64A
5BglLbCD79iZsYINrA7W21kVfXl10wtNhUIAgsalIGYa7btEQtjIU9sSOQRRFgCn8SJzBJIbKm0B
1BpmawCPQ9leUOo3iMe+PTNRD+PgjamBEigKebgTKBy6qGcOUkL0Epr56cEZQQb6/owWJQAPm2Q5
mI2y+8Nhv42LN9gmKvuDTzYAmF5A9xnyk7HAxWxvCq7K8kA4uJbo2f7ClCIW7rnLHsRcITTLosjB
5OC3pWHubEgDPRgRk3GIlqtIPE+Qd0C/FHEzm5+1N2Tr+jM512uhCIN0aqTpI6jaksxSUfYw7h9i
Zl+wE8G9Db40XiSyzo3bKjNBp1Qit3mHalGD0nYDDbgb1HGyQS6XddWMuF6qFYy6yCREqDJVcrrb
hCLWJssYnTyOkyKd22CHD53VsQp2iZ3rerDYG1fsmZfRlC9Vz30qBP0KnBj+1N8AggO2PGQAhfH7
DnCF98VIzVzivaRy6DCIXJtAKHB76eFaq2152Qp4ilDHYOjreqqUctnWkLa6Qvrx4dZ86kl7B8rA
/iTs8QJRPITb9e3C+p3+Uk9Txshbm3P7bFAktcfA91kqLLnFZsKAAB7icXjDvG4RllVT5Ee6hPtB
XFQqCR5EOSgs0jVDbQEbIu7mbYkR+z17TF5V4wZU5Bw47jbmXnJOwYdK3wW+4kF2yE2fgC+OraVP
Zk7/I2+fM2J/mvohM85nuWm2f5D2ZVECTUkRoIW1VkSgShssh0fnq5vYP3zsm3+PiZ6NtvMWfhy0
mT1t01enAlGJR29p5abhR3DM4KO+Kxqf79LtMRPzV9szQraXDdm+MEHzHyPrALUMMYsTARcxelLh
xfi2S7ndyxh4iLvPXVQg9kQiMqnA1xjirSWDnuNC+gicAqCelnxQAumppV15sbdlsGZGeE4jka/p
fT8zyYHr1yBnvZuY4BWcwhDD/+tvs4xQQ6zzyx+RsBzCqkS9y6AoDGBB1yxAIgDSdf/ZCPBbI1YD
J68ebTdvhgHeSZDVCS8Ile3Q3qV86sIzAN0fsk5Rqv9vuox0DSrZK9mmBEv8vf43sl9Yj+oC5kCn
CUYyT5KYI45ZvaccS0jX8bjDd2JMLl65tCrLANykF0TpQ+/fxIXKf65nCtfH1gq4l3yjWJssEFn4
cDCNDfto9wMsucw5YL7LeDzKfaZY9fVdr4vsxH15wgo6uf+7GKRAPRV0pDtmc3+Dhhzr3ws+40mN
b4VeQDH0HBomjpeJSOCE6k0vv1YTN4QnBHNSsQ0rRhsgjYjEiGDUAHUTw8VUp3B+GtXG4ttd7Wjp
rIFwfMl1kESov+1t43PbJUSPBjn3MATQ/kAydOkc2cBLTGxgRR/ixRT6NvpReVDRgdD0rZtLMDHy
02l2a77Zp4ISqd1pV9ErJ7k4zZ02NVve4GqMzfiYFH1WeQFpgn1m9PUk54PC2RRKpm5BcaQ7wcLf
+bQP+aGFYDGSHlcWylKpIbz+s4wqSC207+1VZ8KaFC7yjfFWimTtAkxZbv9FoVtzXBqNgso/E41s
lVjNC/GF8mZN3lJgfUk8MkQuKnpMtc9gFxJ/GwHICN0wZN8QKjMnfApXDyy3z1zKYk4UwMeqh5s1
VIKRyO/YwK0MxzYVxMKPvrts8smxnxtkotW5413LrYN+A1iCxyvCwIfiI+QsD8k3kPAuFxlWp2sV
bkkBBTrt8cI53BuILA0qWx5sZ73IEFEIY/6Ooizf+bP0FeqcWT9vcntWCODB7zBvDuhtjB7QW8ra
1MukL1kWx10B9IT7+x+zmlamgtFQL377nnFirGvvN9eBFEpoUO5XRZhh4sSb5LFVoinoGbCMxD9J
piYIER+yObOLvuKmDIRntzg4gbwf0saxkh482Yyra0ti+XjoOrVt8CT5+yUYEOAdCM/RzQPEnQxY
8A87IAIc0vrOxx5qdwz1LWO2XHGtjSF1xNbNvoCYO0ryFg1Qu0w44gra2qR3gQPbJL/yjMYO4STw
ZshbiWDqf52umjnBB/0bQF1HfvntS80pvbzLrdLCx823ROdaG2rv4GAAolt/iqk9jnHRolu/4ndR
Rbyx5MmhfO0ZB0XbKOprYHZBVy1g55Img9vxdrP09TkxwqHVnwtXTX9NdxtQmPN7grXcI0u9St2o
ml8Ab2XTNG9GzCdfgOS9ldPq7RQcX+E6/5P+iHtX2liBywKIufic7Z6oghJSbqPwcNOiV9K3AUgJ
5LZOzpRDC+fwOpFdJhmc9guuVfiqpG87ufcbAqNVOqSzdzGx+YBOyyN0yu6FNF/FK6GJDgwE6RIN
sDyq2cLcFxaNpP2gcz74S7tiif/LqSo74hrqTOlpGhaDXFMUZ3Vh1tI1lwtLMTC+p0nJ5KZfiHZr
iTCKZGTtPyDx6pPJ+MqlZUqVSS2XpH2wwqU2iU7zPChfz7f6ulo6wsBRidsbDxktaoNeJmHvI6Ku
Is0f5kvMNVFpx/aeDraKReCJSsmiagFHltIGVWq76M9mRqTUWM90Z1wFeKRuudrh46tDeYrp5pC6
jpEwFlFCfYD6ggfN0s8c6Gx1VrKj74YvfCtWOehg3z98QEG3rUQ5jJs7kk5Rstc8QXSGetr1tE4A
CojPdBOLvlzBBqzIUHue16Py8C0ntmkq08RUDfYCceueGvR1rDNOyv8z9puhiy05hef5WOkRO8+j
f25cI07LjeXSScerChd9KfpIwq2TE8M4qK/hJKEY7HOkia8XnmXWXCxN2uZXo5ktonCbdJ2h3N4P
P7cNJiy4BFyTsOxCpVbb28vLkJZ8LeNg4OutpIjJwmadgFP/i2cCoMtT70SoZi6PCUWRbQqTCkEC
znsZ/aFnL5ZqW0CY7u3rTgu4BjatwmhO7JMJ7Y7GLfyJ/gfmXGL3WPlRra5v0sNfagMbSwcuZDoD
R9LJ3lnTYfGGTVl9cfuNkwQwgjnOG2bvw6ATigxoPUjqSVXEfJFwjNQu0bPGHjUzVodmt7toKDdh
pSPTAr7wi2BNVluHUx7jrJB4wAwhzMJzrE3lsRTxD3bVoaFcZlHipVW6QVE6VpuaBhoaK/R3lf6D
ODa4u5FuCR5/FTT/CzPu0pFaI2w4cUYoWq9YrkhTqIIaXZVnmDFWx0bcShxnBvmVF0aDaHid4oLM
JPvAx09Vywg6bmn1LOiwTrSQpTzEODV2VUAaA1bV6eRS82FiR91Qkri9afMlVdcIZmOmWKDODO9H
v2y7uLL9C9RqgF2rIIPGwOaXVK89ZMzrpvi9RjeFi3z9R1xTV58IwzxHP0BENICWENJvJa/YDNF/
ki/OR0XeuW9UXnS0tosLacdSbMM1F2JTfLtl75blvfQx3heVxRQQYNU+je+ZTwtq+3i2m2zHH1LG
W7syD7DArUD8e0vtOwtgu0ukf44kh++Efcvu93ladR2LZIe/+QC7CSrUQAIQFDlWNyBn/5GcYI5/
601+h1eynMKqtJw4126HYAyqHjqvGIetyChKqNGisvFEggrLUmgSKbL9Id1ynpr3+PcC9M8PfRS+
1KheGFQXLywvqe1Qfv0tAACv67gr+bMBUFV8gYS6zVuREFhLqk+Vd6nGtHFT4oBpGEy3LqhYCoSr
PEY/nOFvBFVuPtBF2FR/vqxonDAvUfyBrvVBF6NsKBMZ4FxLmVu48T/yUNI7OBBG8arL4J5sBKgz
BmQ0x+MomeA6ASLBsDxYR2KmBpUgiS8XsQV+Jpe6UtgTpo7nh8UDvCZLz8dHwGClxuWc7BCokCcn
3uRoCg8N+Jw3MSH2T0Spo2BXF7tsKO4IiJuXtOHLtJ+LQqQEVxg3Udy5e61pk/52b6C+wF7EX+9z
EJU9JzwuJAQOU+Gx6CxeWTnFj9b0lDpizGGtdInI0kVMAwfSBpZA2KBJS/eLNCEBY3xSxP3sr70/
46f6UhWcDZeX1WJCI/52MlVvaDrDKu/OSurfgu84/PP1gRpvh4BYQlri0W+Ksp2GrZ2j0etQqKQ+
9164Uh0WQ7smRDM36AhCADK/ZLQcYthaNzKANjefz6a2/C2WYSjEGZC72Ulr343MPuxr9/foWo2v
o0APV4J7H/o1wwNoOQj/0RT1vsumDw9e6Efhj7Bu385tvU6OFzVop9OGPdU3pxWGx0+RoQlvasc8
k4/s+3fMT4xUBIrdbv9YVrR9MT+7qMMopMkfzBL3eXr5i5/a0h6pd0ePuAX8/HGGR/ivjp7vDBu3
Er0ynnBUZzjKVMDVPuVkXrh0OZifjULRY15xZpJGwCv0IbmUMcMRGYAFywDbiJsJt2ead9R5FIHi
yTcmYn7XFws+Uzbd21PE/4ppOdS5hdGJx/w0bPMI3c/ZuK4hydZwlWQn2XlvMZRTTnd6yuEayH9S
r/C7sNCc8tcHugORFiLtGjzzVT497gFf0r798qF2Aah1DQ1lHLg+5Hv2QslxExE/hFgylfsJi3s2
rMnXSrPsC8zXUx4FB3qgKMsrsbcCKUk4PAs/JA1yvva1h8C2M6MJqb8Une0k5qzNXmwKqqOu+jTr
ydIz2n9IE/vVKxSjIbBmYJovSh8qNJYCl3it4hV100RwTH2CO5SN+ZBT02xaM0qrm1pJGwzor6qA
vvCwK2mUR2XzE/LhtI4dzpFTN8XMTowRv0FawQNMMbKM4FIkni/NTKNAm3NytJ5Qi/pIwkUjO5U6
y0Tbspc15z/0m38/QLY5ZuTJJ8XdDGkaxoK2YweI8fxV/2bVInlRLUuY3FAZZMsQjvnZ05aApHUC
QlaBnfK/riRYRH98mbS63zuv0bdASdp8pAyopuuKYZBZBQftnkC3vi6CtSxYIfuuQQL79/5gY5Uf
JqivjUi+Zki4TZ8Hm/7b4RpwahdMEp2dNFxkvbn4a8iPxs4Yr3TTTwX8Bi0atDOznpapWOgLXLIN
0id+FWC+KNDX5wAq4tl0D87s5WBb6mfnfIWUMry/MWX3OFXCiSImIoby8WuxkU1nH96CX8n9BoHr
1rDBrLo3IYloBbKVIxjzmuOXwjsVTvrUXH7/267asmIPlvRLVJTlCUGWq4flWe8rhT+nPHSIuVUx
5DIkJZyxefx7/RIxCNpZ4kbwQXPWCTp8KbcV7VlJWmtIZfIPmMGHqkZ55JtL13n4zFGq6SOG1xGg
MF6wzeRnZehSzssQcui2iwifKmFl716JwkylOKnbsIRTeT24eje3X0quJMMxxjyntG+9Ns0fmoNH
D0LG7f6RGUCSXjXu2hCatq6ewv0VqA2UMVfKtKMRcOBCXIMmb3pqyyKFxq+zh/WPbRj5CjD034iK
7mn8bLu2wnEmL2Nob+ARV+aBM9XaLKmqwYQqiFXBjyhlKNYef8bBTKpjAr9dnuh+BhU1uRaYlDjF
knVvTnkEZDZ6cgU16zjyT7vsq6wvL5xGWhIbUoLP1iBTKOJWXbb7zx03YYRtq5ilm5PwVfR/avU0
YWZb2yWsQ/rL19cVVwtkxeBO0K1BJWMz0/XQr2/9Ath2s5RgBbYiH1+qs3nCpGou8Jn4/wUDOYYZ
OSJ/edRZiTheBHpcazXYSCJmlXPel0EIaO5sa5t5tUfe2HZ6yu1pjLlNEAHXz6cNiHPHpQXmChBV
zg4jYhwnqvWieEpEILOd8rVUzzzGoAADSSb/QIX1xJsU583DhEOsVdsgbN3WDjVucHAY8CH6JYwa
8xWTdqS6FQmbYiz8t8A81kwo+tw0Q+974snShoYlcj0dwlSRkKiVhpVxOjDPDHWposO+EDq2FtQ8
ukkq+U5gdw8F1ZW9IPI8OXWef7bNUyUlQDMPqeJwu0/NqW96UDQcmxFht/2ZsT3Tm04wLv9YJQ07
6oHS7Pv8+yTFw0Ykuz2aj9uif2ywB2cazBdtJEJD3ucszntYYw7DI5mc8WAflmzws5ZlbSfhyEbz
uTmTeLxbKf3qQ0hnImOtGBsrMNM9vSduocPAMxg5PFXX4XCZd7BG3+nWMIxQJQ/JBX58o2wZVbBY
JFGI3/uZllRzXnIimywUwhUbUN7mXdf6C3IAQKSEXyuB0MFbFJey3aTx7k9r+L2VW6DHDl+SBhiJ
0S+OcGFAet7vdXcYcd6A5GZbWkdDfcZaoKkU9jU5aA6iYsJvXY3YLx8CqVbzoxWdBXmVLIVOZonK
KEeliKejsrqYEFY2j+LA9WaoJfop6xJ2xv07AeYDOlDZq5/HAomtcXbp1+TFY6GiMbjWnDegfCS0
DWXWAtQq7fyR0i9BAd3o0QSngfbGt4M1J7x6GNlLfAFXoVYJvkweTECvrwGLSmJjAcpQqcD8rK4c
SZthh1Ndqj9DXpuO9YltuDKl6CExOx46Zb2IVIm2PCE11iea/8Eum5E0rYff7VjFzeoBbb+fv/+A
ELGD9RdrtOPa970oAxsuMR0RxfoDCNAEvHWwo9Dcr7pZov+btCdUZkmWXFahI66nC8LU39skewI8
bJf+5e55PQNWjQSDwSrpeZAlRrlzX9osQUBDvdae2uqzHIjsH9yuSrtar1tY9DEzB1AWLCNiLoNn
OY3BhkXVeWBdxiYfu/Va2WCQDCytMmQMJ3ihSVpP+g0NEM+2pYKPmUYiCfW8v7iAAafmpaoHLSK9
t68xuMCI20XUTAC7uphPXKfmqJAktzLJKrhsGqFcFdxezIfe9TFwVPHfgP0LUoIZ/lFMuWMQgJqg
5bMW2Za7dU1fHv2gKbEX+uSLEAtpw3CIHnkl28gf/pX8A9Umf5l/qrT3eNFQw/ue4Nz62rVLFSiq
MlGB/5Yc+uSYTkSFA92/u41UacSX2eQe2v2OmapE6Dsu8vq8WQzYJt0rvJl/Z0S6kCb4g+h2QlZW
XBtfWabBgcE6LWiE+mA3bDTM7vt0vx3PPxejGunsk4S7WzaHaWauQYwS5kl389eZ7QuyLfJyHFT+
4CXRXi1LpPGQuOziF0acVUpXKmE2zC5Q3MEILV4b43lArXn1hGHiX9UaB9WhRr1KHx2e8WbP+XKn
JXo46KMBSS7x7RWr1UjcJeXKil+rpiNCo9etsLN0gu12V3vLCMIgFqPiXMrwCURvGV5p3F48Su4I
SfRHN67qPltcTXuzcF/72k/4UMWJ/ioQxbm/64X9OQVh+bsjHj2OU4lX86opkqMp4iOCcAa6aGk2
g5YPCsRDXX//v7RdTF9EkpeKY8uybrfS/N92eSO6mskRDPLe6Ei4GG8PAg/A0SqmWQHzyHsgRGve
AyC2ZTU1OqCs4wocYnWVjNAW5PSQAWMOKzl89uNDkmjLd9nsnYJ2BuMnxxfkY2RiCFydHHdi5GIq
jF3PY13SsT+YSx1iQGkuJp5DSTXD1BmFVkd4pBq//J9DRjo60SzRsvWS2fBTqe/g2uh9RcT4Prjc
W5J0Xkz6NXiJlsz8MZ2UAcFxisQK5q97ylIkHIeRY990ceypmkCz4lCQfwm4n3afSoTnNEq3DZ+I
pa4zTACeBCnnspMsnCZEZQDPFv8TAaATscgQhDx1OhqyK8FqxuJ7CZn7ZfoMGN5jXU6Rof8AJxAX
4Wnk7XtGPafE/DyRls45hcJRD/HByykebcdPRs1GpBr9WoLBeNDxHZGDHi3aP0tzYq1+tvAZpL/x
N/urkoTWA9FM77ErlBRaktegvibX9QM/m68WX93B81dIo7wZLB3LwJKQbPPckh3X4DyU1KQmNoTI
EEIaDiefWv0sShcYG0B0GN5w+CMpr+LrQq+BQ4n+z9IgMrBpClLwdofnfofil5cQHKFaSI+2CriJ
x7Ls9D3DDUbqXAAF+nMZNEXIONXJrsbzdYnq6qyaoRfhmcAH6yfzdQi4GiTawkaPtPI56BtaIFvt
98uE9yyIF2UGFZYiO2XEAdHe84hy3SIRmiD86+cc8GHEAuZjwFOESDfPUXOmqXK58wDku25g6xQg
+zZpyR97ZsxwCDN+kpSzlbZ5Lp/ecWxWt7u0i+PAlgdMPZEQ1zulWks7eeBIVdoLWdj4Y407uiZW
t3HPEJb8oWkGr/0+vsxZk4D+YfpvL4wDlN5yFCj44PaHJL6LSCbkguv5tLu1PSRRmNzixUXy5mw8
w8ezxL7uIT1JIcCxcRO/twnTjL1Ng6n6Vibb1w7u2sNBfBytcTK3ybx8NQc7Atgq14gIczlmDtb8
B+Q+TiyB/lDAcU6kUjvR3wOOowgMuME+3M3wWkerZfoiZiLhjGZaRRMdGKMDMlw+oAG/G+7ohzAb
yFIOXcc7Ykm7hahqG2i5kbXKDStwyGHrVojaEsZVdeE9/1EtSuDOb2l7xH/dI4H5zEbtoLSTSqRG
8KeXxBTtkhlYeUTc4W9h7myv3Rq606skoKSn79UUVfw38zz9EKXkhrcnqlEf9nKNiQbekMKRAjGC
9SkB75FXwjyWoguvojG6blMqLKlNSDpQ5xs5h/3M9dDItrFa8fL5GfAcLgfeOALh7S/806GivFrR
65w2n6nU/AQv03pehcB5UFwxD1UoZRUrSb6imgdPEKq157LTU8r7hPya8nCNrB7859XdD7gj1CcY
22c1VSrvQZVKC4vu6s0hoNJ5WNUJ4Fk2PQxK0Ki0QVZJyPom8cluycg2qske+5DIGhEAqwZiGmyU
kpAYvng+hVQ7ejLYGDz6pCzFmYfDJRsga6O436tFQI5gvlwGeAhics8Htw9I+ui2Hhig6MztIRJj
XhO6szOwFghAVfduA3zmYyHJNddmE9+BDdIE8tr331r039+7TCLPmnY4Ij14hEpCO003Amh036bL
lF0IoN1OeLhWinOLnxePAmOem3tBy/Uj0XDggG5tmmTWeeVEefNy2T75saZvbe41CgC4JOSDZT3w
XiQvWZUcBt7Pt0qGj7C5jTemAdl4kPXq0TDtOBO7tvgTk71lGoKXg3Z4RWLTRVDsoYgn5vwzEegY
1CDbj43nBxImIxWie380j/BF2BZm2HLslKrsF+p6bAaoN07npKJ2TG1E96TkTSXaGizxkLw3fmKn
D+p17D5hZfHcO44JTfXSsxAgKFyqCB7xWX2DHorRTGPMBVDNLVyHpiUV7wq3YeyyhXV8yPu/Lpvu
hqo2gJXrER9olYUswuMnfOBR1ktytoEgLc0TM8OILjWvQECWNZK1Hw+hK6Yybjq5NVvUbB3IF9ec
d9oNxgPrSNX2JRDJBLca/lrnf6oBYIAVDx8i89irHrpmOqMNRRZ8jeS1ij6uwCAdq3dCHPrRXWhL
efN8sOZsykFPTUTjT7r1wJFqWMi+Er25S1abIcuWJSHy7l7z7VbDmaMn3fgqGHUAA/V7NBnwgJVB
uJ223Kse9E+meM11bko/yZzxWRJQlRnSG5rC/hm/CJI1X9erD+evlWwH9vH6BbZHhX4Omp/deiq6
zpd1XXjMrnd9rpQd0Pg+nxFX1CzcAgO5vMtpVKirVO+Z/JR8+MvradHuLkkWRtYLLZhJsc48XfVs
68RWplPM+Kt9+hASRhIaXw8bJJ9Ot38k0bWkEGoFMxiKsOMdZ9O/yBBx7yRfB6EGavGu0FpGO4tE
tB0jOlou10ZdBOkg5xGUMWp5cVX/fvDur717VrA9m1334SQe1JC/f/M37Av2sFXjjCcilrtVhwje
/Vx1J6UGM+NQfwFoMZTa4Tv1AG4+tEsGgxpeuVUynCAw/+Jlln3vfCu/819SBO9ZOQk/eHspJvO5
Q+VyL87sPL/DiQdndM3FR83Sr0Tczu6CQWMBrNdoMuf6iDpF29M8opZF+0LBza8MaTBJhW6qwLRi
pBjPLX91t7xUZWN2aA+HEiMZZLJAXIm/NkdJJX/znit3a6LzesYo9vEpCrwiWKHyigvCRjpVh2lk
5m/M4kHHJWWpd1dVt9ckLa8xFMIZmOgqs8Q94mz8fKSPxn8zjWnC6cqT/L3uzARHCUqTovzUSddy
tR66wxceoHHiORDGZ1nM6l9EJexZbod4Bd5XufbKXhSp27sJ5xhG7FddbyEZyDIVqGrycCch8M7U
bWgHRNItUQTERhSs0oF4XE1m+Jdo+HsJOjUhRvojnRO9UKqfdMjbR3k16CLwhFhIj+4AUUWyREeQ
qND81uPC+L3m5J2Stds4kMtkhBR0yJlmhJ+3b0rldJ8A5aTWCsCPiwCR2Jy8E+ugitSQrkYa8G5Y
8A/7rGHBDVv9tIuDKryZSP6FOEP2bMzPVws5yRxIBLG16hIXVLQF6TRRiVJXB/N4ovZgIx+NT/Qe
jtMnejfGxkp/+3yD1CDE/Axes+QXCrTXcDpcwZ1D7X9K3mn2oYmXOyehx31exqqtlQ+ww/Q/pCBg
NHLaXIZWvBW1WPPdT2CYHGPxvzSMuq6iH4wcexm4Z311/XdXAcD81ttI1833TSbLSv6GzQ78qR7g
wU6NBFF60OHsvYWZcNh21KCBAsArrbSx51hFCfdYwMUG51xup0LrhEF3psmb1SuF3y8z1JpZ9X5M
HGzkvLXu9/iEQKOyE0CkZVWaIdcpeGfKJeuR47lMAy1kOA8EkQgAvDLMjyTQ3f+8PC9kMyBLCItZ
A1isCRnG/8hnsZlBkPn/oFrshYOjHjVOPwRcHymhcOvEnTRUBnTGnGLTo7snbu5z2fI7MBptJqyO
dWN6sbtVt7OL3dm9yLSex3uXuSxZgFk+idLoDgKuQyoydYBZrKFwXeL6/2tMtX8FfzLQxgnjMlZp
Yz0Tq6j6VlbXnWnM9XSwJhP6fInSLmJy/Aq2xfdg5b22Uz3Fq/eCWQCyEexvkAcKRztGQ18SWmdg
mnGSGklgPfoHHp2QznK8DBcacM/ol2zbxltD+4XFY15qMaCEwvJaQnqhEOJcY/8NchMhl+AGt+vH
WEePVD3qBoDWhVUq8L1kzZ6gWOwRkJE9L/3X4WMCiuY2IFA+PvEryL4/G2E6LkRTOlzYHxrtTEqo
x8Fc/8cZ011CVAfkBRtffcwM5khTMUzyTuTD66H/xl7d8IkU5S6O4KMI7SyiBkRNVOL4PXY1lIIL
CUs47PygO52VUhde9Q67LtOoGJLQiKPaB6Ynh59KafL2LE3bdjpWWXk3ubhI3uqOfHlv9zev9r+i
FvVnMN2NVqOUI/AYCeYtYC6ONtH+dqkTDOjAityR/y6c3h4Fr+nyov1UobL2uqcVgZvF5Ij5n1M9
WlNM9HL8srnn9u+6vrpcbLZ3tHekPunOmP3m/z/MW4bDEr/TexD8PYz+v9HM6e/842W79FO8BAIa
qsXRyDMht68po8LeUp9jzZ5NVYxGhELJdigjfgtpMxiOWWm2q3tT6TrqAvKHd2Lx7pTYMBtaCNrm
KjlRuiWhVT/IFRA918d1bCFsj41ARWOZq9UlgBlXPW4udrR0XWgIDBrT3vfJSPmYSfZs8SagiVpu
yXpoH2wNNfD63mN+G1WcgkWy9oYohL5s98s6+IpQGa3xacfakfPcoXm2yGnkuhI7X+2ARZ2a5s3u
uXW95lbIdYT4UJ+n+MW9c0qxOV61OsOYofi8JlFjSwUBGrx5YQIUieCgaO09zfPYg/BKpRwUqVCC
HeLIoL6WgI4klau1+cPT8DYS5Sti9Z1sYmXt1QVhWpqRihoxJ4gyOn2AF/i75YLxbichBbFZRw0U
eCQFf7/Y2sWERF07WDZo1YS+JoXe1aQ1vZDo/DuYxKWdPINMS9gaDQTmUkvXoUx0ZtYAxszOMizn
dMkUcsw581qGme46qC+7Vj06UYOqGNRCNV2wzVvc1fCE8LUsqjtwoMK8zl3x0W5VuK6lG7f2mJv2
39uBtnwKbf19gKM+q03mH6DmlRZdepcVuN5H88GRhSWKf67lT5moUqssOLrJcp9QCoViLZf0oLQv
mav77acBQp07TDJ5MNDpIg7WgKCQD3r+sawRYGm/K+avcWo0d1EaLem2LHj1V3IZvMQJ5fNKR8MB
nSX+EKm6kdqUUCcM1dtG3WJ3I4FhN6kIjjqzPrNefLV/wmQ46syJ9LWVOoDImctZznbDNgXMwV4y
5EOHfnn9d52DeBrpa5OIlotzEltqXMbW4Dq7OsQtVHxjpMoXknZfg3frS7GzpeLBIwF0XS0nTYFr
3UHsKQ3PuUgIka7xoDmFK9lCI7fx8TPCdcNz1xqenWNA54icufIcsnhUF1tOSFyz1hZNP5hC2hku
9LrB2foam1j6yDV18TYBAnkz83mirMcj3tIBCkHHUqChFaLRohjzQgUCd54TOZsdbpVeGaSuMqXU
AykZcbt70OtbPTfP7lLcs7OdJZHaDVoJONpV3byzThpesFeflJiz6H0gHRRP1N/wTHEXcsPaTAFF
fA1az905byBKdr6BzMB9y3wiWV5W7WuRBcjAKVln74QDDhkqB5REpUgT01RQY4SFiE/2KO/LUbmS
p88yB1QFAvKTNAMFCz722Q5ZXEyOJYht9u0U8/3HC1lmfxASFK5b0qqpGZBikaz1f6DDeuRZw96h
eEfgXwr2s1eTj4F836jxlVYDFuJo8bTHF/Z6oxtKCR1Y24tL3SO/C/lzvV3Z1ChWUve6lqoxz4TK
50d8/5Y30g5fMZ4YQcLUtPlpOw0todE/1z2ASvSalWgMp+yenmKnCtuIl1hWpDaGr/7pE4UdNO66
zsXC4d5Y/PJiA3kdzIVn3ukyTBhMdz9Y+/mNXFLgp1pFOG9M+kC4j4EKi+Pb4WaPvod9w+cIsSH5
Zz+gxYvutnesO0dp7AmZNCp4s1C6MWFRvkhH3QgE2A+/i3EBocc2e6HdPv3sEDSMKaqVQSCrNqHI
xJ6Ifeg5xsGk1gQ5DU0jCrhG7WSE/YmCOw+KBOejwvQQY22K81sYQh4nHEc976iMSlo7A9quAplH
lv3FvAJu5nwXKXXKjyfTASk1eIaIsDatdUSc4XwXcEtQFQ4os6o72awxuz5i5oVOsmJComzpJRQV
zpxNXkK7yf5ppklkPFZmJLjrSO5l9jiH0MlVmLz9lGd8hfU6IGkiTlmlI5HctfXueLEJg3Q6jDF8
R6QIRt2OBxvAegCME3232Z2DvDI77R8DpNNbkrSYKd94HQOWPlc1MnLnF74Xlua4k8L6DobaAkmN
XGuMC+R3A/oWIZz68VsK7xWpgfiYUGl2okEC72+3LFAz5ffatYdSaEByTufvvl3koPea/a3Vh5hM
YNnqOC0m5rw/zGxi+Dv6T+ZLUNRpaw7UrXNVYDqajOJMd2xBl9QHI0TP3hJFVNU7+6+ZvV3SWUcy
iKPFEjxQiOUITrZU0earoHnCZgJasg5W3gjQ7nGBkf18mMI3UuQePeOoWXk+xgixNEtpeWXEC2Lz
ol9QqaMOqi9/gBa9MBIXajc4tCW10m5m2dpzIEBIG632mQTWcTZOn4xYxQr2wEIXRa7iCUa5wVCi
AZh82GunX7BTKwWeeBsLu4kdlc81tOo+YqLDPvk6O57aNttYsDxca2jWaFeYC0uw9eBI8Ub2LGIw
lm+Knv35Oo2S6MwEY4Pa7i4z/N0f/DSQ9bCRYOIgL5uepUi61v3VaSr/YAYhKoCE71njEakeUia0
1MPZn+CMLNwr1kxVQMTvdsq4xtwaipblhQs5tI5ohim793IosLmrtbCvD4jbdwMUAnpMPh44pIuN
Ez/v14K07BtnSParmOJP//gy/4wJ0hF9FJIQ53/tE0l0Vubt8rD0Lizto57yZjX11rSQhmmDTE6n
rWweVk8L61wuZlLxu1pHAY/sfx04A2pMNVxgXwhRQRSVmFl+QuBF076vzgILIiFLet70ft2uykr8
ZOxqfwdYjtnO7mRaW9QgwzVGR2UrBTomTJKQ+ky6hsB4Noz4zLFFALV9JJ2qv1SaxmFqN4SMXX1p
1D75y9wODl1NZdu+RDFxDAb9Dr+xYO2ePdGzxotJpjlbbby+Xqmx6Xx3sQUakVNi7LBu0Cu1CHXQ
Asw5n11mczeNdxsENMFohhoeyRITpPDQoruZgm/7uzrjtk0S5goLeiwlH3/7YBaYp2NEQlv5ssFr
+MZTsTCWL0ABa1XP1plUjJKp/K9vQMmjHEolEm6IRzBvi9XNUjzkEj7HnWkOh35m9HzTXAZ3bxde
zYWaCndERcIVqXS5Lldub26uqp27+/Byih/x27UBL/KdOUfJMMI2Yt5CuMzWjmgvK7TSJDdVqubG
JcgAOg9RjcmefcOMjt8tLgefqrc2wo4ZHFaMTIvy1AcGEvEXbovtzsJFVgOILbyTNqSH3XxD/2Ac
wAHm3R+VRn3SctnRFYN1PNNPUOk1mAws6h9r20gCi/m/2EB3uC5yd+0LxiO3XRIqGWXR+CC5OOT2
mNIXvsVCXKAQk2j7za+FxcMrsvOmNMXUMX8nQZAp/+ULToSoKENYj++ygeGyGiw/cVTT0wTc7is0
MP6iynqJso0EL9CO5Mnu0yfSCnJvI5oYlSThal6LbV6aiV/dIM+9CHv44gle4LBoBuKQvjJpfTe5
wip31rAMs8p2Aqqr63e6mNEyy1fmGpFILrvuXbYV+FxsZspcFPfp61xsjM5a9C6b5Ho2zhoXIl4C
zQ+qFTH05ouoQ0Q77jj6poXxjZTU4IczUrp0C7KXp3XjNtkqj+8sKKz7eKNHqeRlBsF0XL5AWuqI
JdJjOppgazgzOYILq1OQiEOSRmE89ssm2rZ0rLR2Ow5dRsVIvSGReaL/eAnc/GtwUGrVu/m8FYto
7UjpRW9jl+QtCnYa4pIYx4MyOEpbh79uuEhvAnqu0RxkgMMqiccw+4MNDOfMLUk7oThHIQQ0YgGP
JmvATwlnPWNKoQkHSP0fYo+1SSRkxWT44J4dgCgfOgVTlClH3OdPHrovJqwwy1tJ82hY71Al2jji
NgcpmLEi9oTwGZrzXdJicu8xK089iTNScBTyn6eLuKt2XVYsOE8E8lQYcS1obuhWzWO5AHWaugQ7
u20CLdEHCT9r4z9puMAIfMNDhsnFRpNgsgS1u2efzo+q0o54sWAkvQL4x+Owu8HPPwybp6/oevjt
CX5gn1BgWpObK8anMVbkkiCdtS/+LAI+pKccBluRfnKXTVgtjaWBnKMxzS/H1goX/eNDLsByqLbm
UETlm3CqjhBbA3/xwJmKaNg/WnWcyjstUjrHGJF2SdBbp+bw5o087Dos/+j6+TdgndFVN3ltqqQz
AcqfkAHaxI24Yaij+nabj0L/EjUxF0hQb+UUD7feeSIqCGyXebkteKzJ7LVH0RycYq34anUiqkE8
cDLpISCpwYf39FR69HnuqOhMK1473Pg2UpR2XSdCjCeCJ/ECF41OyV3RJuhbfgT+kW3iLUPlV1bk
RShbRX0KPCQY+7M3r7j9R0+qt5/JeqYNF92zqfX1JHD3phvzK5kzj13fJki/bjBeEKOdi/CQRifz
oEyvjxVEMxl681NlBOHAIRG8sXva5jhb0+dTXtS6OjvAlmTm/jmiCJ80GbvdN2efzcHZ9yu9dDnX
l5GJVn7ynp+f1wHeoLYncYtMPFtu9glVd16ymnTL7T+ro6PNMANxgQp+lm2rsKfFSSxI9fNj3J/M
rxk4oBXFgRM8CpMRd6Dj9SDWIgFuqdLgkiUW0NeqqtS6NJE3W6FfJxJun1YBmTYSLdW/kyGySLtw
AMtzIcZLmRKKQS9ImEwJEIUYnugTUEEzhbvhJRXwoIarmyS3EQgFX16vIJDHQMyzSIqIHKs9pPwW
hcaggMjChUqa+YiFQreKN0CmTkrPczr62TN+mp9Q2O5u1w6abhNukHGyYt2A71Xc4fGRUw9aVegm
4KFx6g6FLKKEEhnyG1Rs7y3wTuDaEe0u+rckHoLV0i14Oum0wweKHpT6KGRVGneaUkaOrRQWAbXs
iitceGvmSYMcTrDNBNP1u544YW4qKPe0D6TlnJF0dPiwQmdIZKhqlHLUY/DTfq+yH3vHvf1yW7Uz
JHYBukSEmhfe/zRuRdHl2DpD63FujmslOLqiHnMiqAVDuHe+eAZnUy2+cVRtNOK5F6YE4cqpJQpN
CGwMjf/LMLUCeGT08T4fJVTSKsF8dWQ5QPRRGH1SKqD2U+0elO2UhwcC8T3yHk81m9YYzSdE7qA4
bsWZZdnCPxYiiJj+sa1/oLPRB6ZsS0HWJy3clexfgtQolWE1OYG40nB2M0NQbSWQgRgHg09+DJ3o
XJbn3437CVUoV/cFqvjhD5IvwgYoVDV9I2Z8jKt4Ay0DICbjMett5134ZBrZgqRW+kogRSyWHKFr
dBra1Rbj3E+SaQEEBt7GClo2MMnid+JTYTUEUux/TZI6tONo48graDFIhXupZTQqfcQ5IrCwZ4yW
auUsvkXB7y+J1nCYBbpftYdFYKYtTsurFKlmIkaSa9JiELcO/TC3yySc1/YVdYWPavWnH9oNkaHf
j2mUTryOmoHKlcMONjwHX4JKGBFgREd+k92O6XFA+fzuFtqzBETPKcigLYQ613z9AiRZKOCjpDJj
sMGimmObeUmXGG6qdaQh2FmvZ9CIaY57yi6rx4wo8h5hybd11KIgtcwcwkZONl6nDU6vxtxsWpZp
4RSZqU1W0xUmfyRzkvslrNipXTKc0rvXT9zKSxXqfQNAI66rB2FYSSbCUp0HNHGrChO6f+NGrq5O
STewHnenZ4vaP5YaFeOQO2N9w+ZwyoZnLcuG0hg2FRE0WNwIwOyX2H5eKAKT9YruyBevODy/gqjH
h01ZDCQY39qEEUm3DoLsJkgZHpPBZgffLYwJ66AZ1lP//CG7eqKg7FdyHzhsHlDnmdJEuVezr5yV
/xb287pMVn1XUqTOlv7/2cBt+z4Io8ZhQ8eT0hqzDLCbWz6ueW2McJfJ72HyQW8yN3KxiPqIuzZp
/DyzRnG20Oklz3qwoSmTHKm6d5jTzqDrzym+HcXOrfUHjtS/b81t4XZDgiTaWAFta3XJ9kcDNU4m
+Nhl/3CAnaaX7GRt7o/M/wW3bym1JOvBFLuiCXgXz8xzZSw3qnvZQLB/gkE0gmaXkj5UPCdExBGf
/t/owVQQ5WOOzzbYEr528vGv5bwjwKlIQ/HliNzxL4H2QAGD0wxISiMQtH8i8Zl8UCtIp98IdFxq
RjHJ7Pz43RD7jOFNKwwNAF3LULaiKM50QlUKLkicgAmp1VMeoIgY+EaOVILcpJnhbPHzfeK/2lHz
08907qWl+q0GDatNIdFxSwyNiFqBapo3iHPPOquh5mn+1NLZXczYjBopFptPMIwkZ/FxbunqNLJq
Rha8Q2XHYKZ0P7dOgtYEgGxIgEktCFHirmW7TmMqKrG16P6CAgSYa+L3UnTTeDPvjCGcf8VOrLdt
LnaHu7X/tMLey4rrKiljGYO5A7ZC7WFu7SMArRqXJpysQWG8UxH6lNKlkX3p9jX13V7fwLaxDode
kQAK9UVNHj2bXKbRDh0+weVp9zZa1ob2qVjExp0B2V0fCzaxMvU5abpUe+c9Qy0uC2mqapFEfGuw
YgaS9I31mvMeS5Vp+4dbL2aogc6MgCfH0y/H34j0httGvACR3/9voC2wJi+3Qy8zCTA+cYv+MiDX
ulEycnQtdcqcQk0i8rk4og0XhCBMUYB2eswwMDqhzvt874j5iuFyZ5mFiBlfAvdI08Wl9ARzRfjo
tj6mBGNtxDVQVTP4HL6qpMRPpjTEMLA4vREq0yP588SFd9QqeOPh5I4WlpiE28ZiT/PUN5T1HF6h
LvGgAkfiEYS9J+5BWd5omRNdfOcdrPvOpYxDG6Nhe9XqKrDeY5Lijz8na2fiqbGqkeytXw4oam5i
XI+Km+dENKb30HeiPuoTs7/ondxmK2Pwl7+qHu6B0FMivwDuaWw6ffNhIyBhPgYg14IprtVWkhon
qfu0ugc1xyL7KNdk1/rMIcK85jEVgfWmfKhbvUoqzwcsVPhGOf05xdCBLFwn0yTxaj7/uSo0B/wC
BgOE+uxVS4GFYeUUTU4SWC+XayOiFHBoTsfLzlGdrftFR812XL9xSPdtql4tvim9fcOY1sN8khjT
9DYK20OpE2rCpOAybUWKdB9eVaWzFMc8/h9mHQHcCp3SmFFb80e1z5X/c4qESFnIgsxcEsrtqyiG
eKsb9b5OveLlevqVblijFgGp42cQpO5C+tI/sGLIZDhrWBij/vrBpAag0l6POtMOEsDkYDOpifiB
W0d0qCtsZPGVnn6GBfNNw+cflNVAjjbrYb4Wc5XBBgERqdenXElOZc1FFn+AVvTqMxRKD15/ZDQp
onqhvrVn+Qhez5k8fYtzgofX8zxBoxOY/RY6agWxIk0TM+S0FQZcvzyBmHgxNYBQjgWV4CjuyM2/
H93Hgm/mVCzKI1HJM0vFVa0RPQETqB6ovhbEYiDQgTQZ6fNdLJ0QHUVXfBSB+eL87X7Y4ogrJF28
5EycJh1MPD8tB/7+MAoefgTkXJJiWOG3UmmYmhSG4YtzOOKX7rok8iWXGU0h+MY9K/EqQs9duaQk
O7e2kn0bUi8kv1ULc5zrW61Omlg2p/hPVKnG/hgHNGaQyofgoS7L899Idhm1D6Mz+Nc+RDluZgUr
eo6wj1ThGTcwmijhhhQtthhOr1Ob8kbIsXKD0fL7kN3YS+PBrw13XCgBIhXhycMNegPd4TjRAKi9
3X5iNMggdFb6XYsQ7alQoO21x93BZSGnTSd/DwXhyW97YNr8zIBITyhRs137w9F5Tm00VGqex2cK
s6sQDIN86mn5pAJIdJg5I2xG4pajHs5MxwJVgi60vgVipOuQNOTTpH3i4wjLjQ4zzNePOrAz4pz4
jCKzBLt4bFjAUiWmrHr64gWgOkXNRj7X8uRng1UpAEbnvb2DgerUHeRvA1yiu0MEPT/S5ncMV93l
/3OMCmThnPiN5pXZmjaZs1JlNy/Ou892HQjBSW5UB3Q18RDkVvl3jE6rrmr5oxrmo+JpcWgfwdDN
QXX5QOpLWE3Yiznwpo1zsEfRGElte8IUpm5+FkNMU7p1Rr3GBgsYhuv7BNO+N4tS/e4cqTSRdNrc
J3LC3K7U2ghNO4luq/YUPHU/8ZTcQ8ZuEZlGfV5rJDxAZQv9lYAaPL2KSc2dBbYAwwYzvG4UAfJe
5ci2YbGvAtU1j5vTZW79cJAnk/v7sLgpc1+mYWPjdM9GNAHs7j5YELHttWedOyMLZXyTNohYlgqn
HkemIzXzhZYGB6Ghds1lXyxk3tFIepLO7ufVqMdplmp0PSOzkRi7Ugemv90Vk3vZWDmM4qGhbc6/
YKM+iW2lbyT5EB4FVHXMbPnMJgkfb6iJ3RTCbPjM+XcOF9zOinLTa7Lfv4rUAH7yiu5QR2K0M6nf
Ikpf3X3sixXxecSHEjQQ7KaSrkUc7EUU83eJ5p4i4V2HY/Kkgk/l6+PFEg1yteWAzrhQdvfImsog
VdmCcbHit6LCYqX9cVI7hO+tGcV+UBW3geASfggrZrGXLaxBYvsHw5x49f250mouydM4VcLJcXNk
bK6ZuMgHT+Bp7z0f/KJDhR/m+zoHxyXkIk0/ovTq9TYUB8PPEQu+9DHgb+cC7kSYQ1enfBgs7boj
puKPuBYyoBpYsSwD8ifviwc/Mj5yVr0Wcaw9bd+3Mk6iLwbTE2sBe0gHaNUlYbED8CBXaF1fqlf2
VX1dUcYFPcq7Hvdvv9M9deIRgs15TeULPf3EZltKInQaXxshTbI+7LTyR9RZzreFk7KWSHIs9Apa
wGkcPLURgILPgbcI2kAiCjVIIq8096f+OKsP91WIuDD+yWSD4pOH+KTwu0qJG+Y4KORdNCmBL/C0
hOEV8t7m+R7zRN2P0ybewAjCTfmHvX71nJiJ9tWYgorvqj7DlbqcDXOPEpBE0rT6tWNFG4fHw6A/
ciW3gLBnbfcPGcVL+XRbowRVWhGOSB8IduKuLiPCI999olXG4X6fqBw8dp4Z0ayEkZ+GEUDYROk9
FfJNsw6+Y+KcWiHxRbGM30eIVD/PNcvlmgvL6+0MLfvmpjV1U0e/yJ1FC3FqvYrM9iC2z2AYj2Tc
6+mCTqzxEzTV643oEW6HABhD2VfYvSPz6Ob5B9B166uo1R13wqGi/uk9NSR2Uaue6eaJ3eTrKlPU
xy/ohKyunhEh+jOMNWxxjFn/laqGsvEgD53iTfrcw3Hvch30H67gSQsZXZlXek/P7J7rR1eoETiJ
MI7Na9UUfnE8iP+071yew6y6/tVsOAY/VaOY6KT+dPvtA00gRU02rXjKVy3uwnra7b94VB0bpn/5
URY38lqYwfA7GiarWjodMzXdzyeMSbRbVZnmYMqJu6YRywDOK++RtwRekppopM/FJDqRL8Sh3z8b
cCU+P2azHlNvjhNN+3YHt0P71fL1M7XQAkENIv2rwcw5ojJlP7COpeDePJyCldLfIvOEtaA/l/Sm
St095tYin7r3jLi5F8SsNVFPN6hvqudL35KOOjglHtg2n4KxsSc7DR0mtkFC3SiNZ/E72bLgFNju
RQlSTaJsxIbfd1dsoKO1c27gygUWAez/k2+2ejsy/zr1/ZMeIURhJRLMRxa4XDVBckNGYoDZUx6L
jiG3OUvTiDUpf6RiV3vPsY3TZ1+wBSjEGbDUTUlCNuRjLncoqgR8rO/Mc6XtG7A29S5GcX10kZw+
59mJncabhf8o0rUJ4wJGphlo8GVuagL5yGIynSWt4R8sNmeWaVJ4noIDw1QcdoOo6vz8nFtQ1M96
9WHMV0zj9tQgJry/71Xr/9h04ewwVE5uYs3J6+umMTfuMGcrbpAfhO4K0/LVdQFtiqd9eWwK6POa
p9heTwefpBbgHULTMXDRO7iI8OQhHyDS4cpsJ9dkP3U3Afo2WLVNa5jvE+DDApqQIjKUPmXNH8du
GsXBuE8bWlsVzmxPsPlOyvLTBFlfIxmrLzMj8ikLQpOW9gfJTV7iG7KsanLUj8JS3Bt5ogmxckvD
qyFwryCRPMttvdKhMMSWphTUoFJAr17m4GSobPgXdqpTPsttCqL8t3doHU84gAQbeAQfsLG5ZdKi
W1Ysf8wl/brivzIgmGoM3xaH+F9TJTkYdpyalFvorb8WMvMm2l5wv+Rm4LuAiyou1L8yJGm2OgXX
DbFn0PV9UEuIyN7g4mKueRCbOHpBgBchJny60VaR6s+kIRwIsrlPuMlg7Dk8EAqQrwcKUJ2gzFem
A4X8eCubZu8pVsnbSgAG18NX0uRvhz8ib22NVUNslzk4K9EcrO1Hx44DRr7F3OCr3PCKYLHxzhb3
JOyu+mO7R+MlkNe4V8KOrTPCveZNyYRG/tTb/74e3UeviIkSo2sCyYKqLWL2wgTGtS4zEM39RTxv
E1y0/9/5Vm4V9i3+wNH/X0Y8/V0tzJ+Qk9tw4AvyuaU5IiQm+HdAMqX+/oJTcXtmWS2kG4APz57X
FL/VFANmNM7GdMDFX2FanaB+kYN+J6Xu3ADKBcRZL0XD9fTN69FG7MfMTEYb6PdoQZc5JkFJzHGC
LfaEDmFhShWKeIgNKnH+Vm9if8R9Li66+tieZsCejHvd0iUkyF6C7yaIBNSt8y6Z4knRbM5fSMr2
VFrVAiJk8PeR+GNY6ExMGifVFZC0CRQqgMAWU08ZuiJlmDe1V8qHkSKhhMFZHbJHecF3UhL0d4nM
rQDGLZG6jFShy4K40efCVLMHrvf9/V8Tf6JrSZ8w7KI+se/cqxLtRyzbBXcAX/Gy+p9Qp3JeZpqS
542vzVYFHd+WW7trKEVpf5ARYwbIad0D3GotPGK9OxgkrLkW/HB6QZpsylLUBrWa1gZrfmcSyB1G
yAw1BhFh5bdV32XClCvyDVMcCsCm3ZqYxH9xQnLsDN1y/9d/vkh8QLFrLyDzUirNHTpUsEE5qrKH
UueFXJeZ0QV9S17KpTHaYdOgOu1cZH25oMCR8/vTVhCN763IaCxIS8NooOYiCigr0QWK0rByPgjM
dYZZS/BmJaP2Auem4iD4B50qI3Lpt/C/LRlCVs8MBiWGYXho+Z2faaz9+yVcu4Bem33q8m+tl3pi
rPkMB0X6vYlbB7iyao40iPv2rvASAPN48GorUi1Ied3r5Jdni1prMRaZ45F7Pg8ghHJgeRxHzBqi
0cpwYZh8YtQCz6qAPQDbW3e3Gl0KcVHJR+kdgoA4tR3yZ34XjDBBUflA7Bd18lzgQiaEY7TIVLYz
iLrtF944QQnG+7kzioGs1fZj7h1ZHCWxLYTknGEaElLAbGhcWSdE06JNYeb4Knu7bi7CcLf7KtAN
wK498k01bARNYZlfEj8s4KoF6kIAjzs7pd17+P1bpqWqStsk5HZrQxPaLWmLE/I/kWU5gkQRHG3I
6W329dQDaFDJ3p4smUiyrJRgn2qYC7dlBVwMa2yzsxUuMDelrla2LUE9G2dmRR+eAbNkKnDU55HL
e49MCsu9vKU7AVNtrFz+3zd/Eanb4b+ZgP6P9L2rPpG+FSJJKSqZZsnk/MymKuTH/DTZfEXw8Yx/
FKe6pNhTu4v5fbXvC7ov6Zi5zdFBdUopg8DjICn4wuzZld2fdiyrVK58GoAo0erU/xrkjUS5YNkI
9uDqe4UoVPZ5AvKSiScm13/VyZifGfrt4PwBl8h0mb+y/W9cS81kpEgoK83TfokSA3wO2h96dOQe
+2LFB3nDjzfRku9Ys1KhQ5k97qp2nzxBKB83thUalL+rwTq6JGBnBuuRiPAj7JhsXCuh9xLlEo9w
l2vhppY+927e+hlOE+M0DIoMNOkjRTqnTczMGtFLOK3CKeC27SCciM0YVPSh4RJvHF/f4mBB7TrK
O9FukKBmQ+ujIdv443yMIPahkZnBrT2UMXwNsvRubEMJgr41e9+Gy4ZR6AGW7wcloMsnIPgWVqm1
40puXLsKJD20JwGmvjsEUJjwS1xC1xx/5W3hIqFexPIBiTgl0lMlY9FikANUrS9wXHIIF9/MdI/g
MplnyRZyDbx4OR3kKPJntqWCV4R6IC47xi0ROeFMzVY0oJvpu7UbPKdjMkbD86Nyn0lSZ+UiWcPL
DZAq5S7+1IOEg39HhFJvEUk84jMcxip0h5bMyr5PZ5+nKpYYdBpvW+8oJa5AjghKxidq+mEik0yq
DfAMWfXE0oM5Qf5Ubj2xPIdW0ECbtkj7ugMqR491Wx/VyH1JIaigYTvTMbzTKo7gUSPqPoQD1xeH
RL+2jvzYcdi3LtBf20/XkdprIwon/OzQq33JcHUohuCr7DwmAEyiRzNTeKZ/9QhLAtVVjWjSmqBV
Zn1qj3aqulQniQf5uqkxhD8xv9zNkUHb3ibPfcJAjlQJef6uILwhnUpgjOLRJnmfHHd4BQpc+xh1
Gt/75H3IJvUgtcDv1XhhVJfw1QOFVCaBbm40p2pZHOwvVpCpaEbxBr57AzUZZAsh0MY78K1R7hji
YsEZkqtj7K4oUhIy+yuTRoGhABh+d4dW3/fXM3sezpw52T7deYsHg8u2DCPq+xt6DKDNXF/Pz6y/
C7P0aIDOnad5NNZbgLDW9VwZxeF6yTkG57KLNgoYs2Zts7DuYBU06WI3MWhotBBKFTHP9vcxThKC
BhuPHEuTW5cHlVn426oBrePP5/9/5Ll2hGLHsavZ10pktYMbIEA85v6BjDv/vhzJvLRUF1oxtV2p
mFXxDUImhbXuHRcghoJS9b+1FqSunJfJX6HixqgTegD92W9v1TNva5TLDqZ87O3R3Pj76QNa0RUl
5j4l4ODIIsin4SOcELH/5gw6WSHxgANFUcdT6xYX8SXRDcDWTAGxy83vG2rtHWKqwU8Zv7osLIfm
BSi6VUEPJSorP6hyFNZsWXtRtfxLe+UPMEbUjLBXCHq0zyl3CgRb/vmDjRabU7Fc7zoF58WSbTkH
tmxlYUXKgkqMs8k3wQ6D0OkNeHPtDpMRalX42/oCifzE/i3P+5BUbFhwnhqD6sF30+fCJBZHtZ8j
EsJ4LVz7jvDvuu+SGUbMqbCMMElDYTRZGF2+h5SojxJk3kHipABI3+O4WSMM/wmwnHo45MSwoELp
2hVM7z6Zx8xYOAH/oqXbtmxkCsykItVszIleMjhD0lv/XHPNFCj2Yu0ZWoskZSU9xk9MV0eYal6Q
LbykykSHmh6ktHOR+BahgFRxz2KjFUSjL4N2KcsxTbsUJ0FGMSlPhV8xuaSvm8A638f9s0ARHTaA
+NGi4FIU9PyZp361ZD95yZlQaILqCLpL/a9U+xmzx6g4WLUpOzR1K1Gz6reGT9ggp0ScmEYJXQqv
V8ToJh4KqlYHQo2lpmXigxF6ucZ2qmcC3cumbdIu0VTiXs/WFeDNJVoeC7b83AP8Wq/ZcsA1o83y
3qDVYbb8GU3hnJT3T+pQaBMJ8lq0LNO/tRgtRP+KKu7cbTX6QGUuaeboNpyYqHTPqg5id+4JH7Xd
lTuh9SXyK3yk0rX0trHSt5Aze5HLDgLrwKyEDvJfjMl8ShfdqYlWX/QvOtqdro47o9mMakCFm5k0
XqvHgrevLo3F88qMz24L1t7/fPG9wL5DPvRQ3LRVBMPNE+3QBTYDkguZUuNKF3sJc4fjEt09aagL
q+8NsKJniuTqHLjRMZRx5z5UPULf06b5FLdsTwEBANvIirvo5dF9kdW8R3OlMhd9ojjg3RPt02h5
jGi90pWcrvAviG0xurMnEtrNDfIIA6eRmY5oH41fhH69Syk3BMJo5i7Jh4shnK+eOuV9CjbAi5RF
JhObMHMELEHJByb/e+6WbbW0vm9U+2a576fSbROM0gbIy3DV2Aw45o07tXrpNOpXmIe3yBsBXjTs
TkKNiGehAE6OeHpsSbM0Gxyxm1QjxoFuABRd3GAoIQInoesqjB0CsX0keuavqAbayw+cVfu2EcS6
EW0pPZs6YAfqDUzt7VLtXco2a1oxP+4ww7ybi3+vh2orLGCwoCose1U6azlxFwyEID++WjQFU4ax
XeSL3GY+bHsFV1rdkLcRGseJVfXAVyvkAIMlrXnfkw04oJM2pV2IwCWJiHe0b6VSI0Ssy8SsTzsC
ykrTjRtBo3MQT5jr6kKfXqOdP0bnKZS+hAIk9te8eVKCf+FrGJ8nTMuahdZNQ2r9h5Bnq+OZbXrz
Jm2xuDefJFc02seqaA+8AEdI71DHSJ7O8MSW3oTKeH/PECp8MBNdR4AxHKUDLsnXjWxBu8M8IJ59
FU3Mb60+S9AWfKTWYxZ3YbNzOpNbZAdQoQd+pB0bmVHkWearEbuCqd6FIab6CQitQQhKn8XmVt8X
A6DKLnIn4RA0Zow/ATQPAFcLezY33k37NQ+vox0Zd3iGyERs+CGq33VeCMK84rtIYcVB+iLptlE/
5DvFYw8tTvrlGEPW+Czbnhqabfi8TXJ0PL8q9Fr/mpRHCY9AAErUid3bytG/pJ5uIh7naWNsn7uI
RoBpLDi4RlEZqDwjUWzk6LioHfkTWKu4lGXLXw0eARag8fi+NFE3nl8BIscolr04LAnZUgyCgQOQ
wnAPxNt+vllWCc33ij8kG8fxlJFcAYZ71tcsp7CTP5tS/4sKEuOt/+baoMiJ2jW2cjJd3s9s7rBp
/jMDEJVH5iYzUYry/udLV6uyDjv9y4A0zJ4Sll3p8qSwNMcry6Jgy8GxQ0O2/xbnYoWavh7wQ670
QCphixP/FSdEoqiJWBo6k+SyXtZVRIFJrsSHUVfXjIKZP4hZUSuTTYekAdUsjEkbMWH9W90kpwK/
VSs39wtmKLPwx/SvJt/cRO7rd7gm8SZGeOkUOzHDFGecYxQx53Xz8YKy1DpKjVlfH3VVAAgZ7gxe
SNAHMNKRHtg9aYPaMEC9dVWvRqFs13RjGf4BwjPLcXrtoo0k5riy0NgelK1xJeiYJ735+bqIE4e/
xbavbgXy1OZq+eg3gM2gPu9Wx4LCXJ6nyOH/qUFvWM1G0gVjVU8YfhTtvllod74IzBdMUlbQXrkS
aJlrzH44sfv7Z2nTEHkEXEexrlJ1EeonUYuzJmEAcyF+KF8Rvy1g886kWiWRP7/WM7Kf5MQVbV3X
4EvBxpxHiczwXhtPt9HqaBQz93X5peFgLUG2peu/Pwy08XatfsmD3FbviZNYtbZRvz3ptZIMKrtr
BDTXODiQl/xTl5Sn07InmgYgIgvbYxQ2gfs4uzaIY5xHsXBoi2QF+ELHdyJTkxxMzGcRsIMRQfJ9
3HcoZyb4NZAU/NYgSf3jLYKLvs3v0aiMBfZwhzEv7ntmG83J1JOUND9H6pX7heNgvXQ1P8yUES81
ghobzOtTZUiYPsNzw4CpA2OqNjzn2GihLBONJCIKl74e6IWTEvAgqocXlcL/wBkm5/c5vhPZbrdb
kB7D91A0B7ukCDN1/3aUY3I+e0B63LCSeR/G4vcH9Xf44WeQYwmOfPg2TiqLnVVF5XZPvdVq44Kj
gawrPGQhcwgk2fTYY5YG61ABNM5ysT8amQxMSUI1kLcjYnPjqScSAxVpLlSuaDjY8qAWVnEIZ/q5
vRYqktiGet8y5GtgI1VFJ211SOE10cfHyuSbSe/+qQLC9ajlimU0fos4xOI+xyjnVI9Eh3NC50Il
K54n61pLjioGkiCKwDZ62g7OTLm2YvO6qJzeSBUf6H1q2vUYqE+0uAc0ZtZ0pwJTNKgFjhUXREFr
ojkeCkvQdANUh8+w7oE+iucZAxHKd5TywRcuJWI1u+G4VzGAC1hK65EMP7ZljMnBCgXYRjlF9TCM
FCtvxfF4t+oTOiWGlLrmEtPzuaClo+5k/jwRLu2NUTOudzNCiSbgzj3TNjOouemrRBMURysrSSU3
eSVDq7ZADwKf5VjGX4+Rly74d7pDgUSeeEmWjBUrSTp59QMIRr1KtVstYw5o8wgRX/R2FJhH8F1K
qSZnCYiLsEjhFWVZB/wrQtQxzAnYvaU89769/2Qbr/deEq8cOxIdoBlfJsRUOCu7OqkUWm13N1PH
ATFeKk7gftxbYEm202xTM41Occixuzg17jiEBAjlp/fAHBo8nP7OjoladzL42LTlkc63WFpbbMGq
b2iydM/+z57TIRilbeqL7bZNTKmBFjSVP9fMjI1EPrfz0cfPlxiZnfoEi1xIs33hz/8aEZGBBvte
ShB61a7ogoZ64neKkuCHwHR7V2DJDCTam8SzKDIsM2HCknQGUW/dD24MijeWkaSocSLDugLEMm6/
VunGNfo0jx6jlq5PUUdlaOOcbzYVSt9KnoF02FED66vMSMC9SALkKiM83TdDR29cEGKXQi3Uxytu
8UsVboQ3kdpz0HRRCzOOlEHYqkO0LrDkRbSlG6sE9u29updbCO9BX2UQ2xfUCw+nw4jGWm2quW6E
URHx3Jg+EatkrLo79opawgXYZWdQrBjNPJXslzMQRGmz0CkYCClryEwAQQRJqUW8F3Kv8uYkaYNC
bB+nwRyDVk2GAdyoXC9YNGjFhWnQ2l4YV8fWdx8kXT8N27+h2EIQg1HAkC8VJQLzMsWNATo2lJcM
sK98txOxiEmnomOY75+8yFIU1UHPa1/tEZTPRlWAubHSWkFyH2nuurTkqh9xnNN5c3M4VphrUlkq
P6qkTiaAw3J+hLl/d/YWWu40SRsE5vWvmMaiPGu8o2JxuziR3Zn55t9FHxgznZsHKbg5ZsKeV1Wp
zzYJA5rU9yBAujrTklU8ic9h2V8Dk5SXry3+mZ5zqmyYNwIFoiiPupEVL3zJacs/Un80C1/AvdCw
SLahWXEBGKfE2G0eT+Hf5o9TF0fSHGVESlhW9vAqXy7vVHbmY635l3IK/SScJI+uanuxwmfRqZzk
tPMUcelHJ2vnWYemZ9VgO6mJV0LOQHPyaliGJANq6IaUJDyd/aciiPdpOFdR24XaJutzNc213U3Q
uiBqW1VlPDAq+tVosWQLunGM7LqzENrHTJeXdl1kXZil5BOjtAPPGHscr8zU3BhbRuc01fDpUfOB
RCD/o/LBp0lv2rmdgEyaB5EvBcD4qZG5c6MMxrUWx4Dtz17LELf4DOsCgE4Wy2qe66kEoHbnCOTB
upJso5PrY//EuinTU4/tzDhEq2SL4QEwrIauYnmPkest+wX8+4kgzWipbIQmSr8Du2oS/NtXHvn9
OeLiV6/zEDELion73X56hODnZMJc7SGMglN3Ahv1vssfPNMxCSYGVuhHd6ozNmGgxOv/DUphwY/+
fo1HqmdlVIATtqG333292+y3e5swEyxZtJ9vlIAe2tYUgFrdZa234dICey8nCpTxSxs5YhzOONZd
bfc9uNdtADL41ZvrmCzg9ZiyCRNUM+iKFlAb6EC3JMyvjE0FVgavZDw4nAelMXF6fGlw53u47g7z
rfupWhFFgtv7gnhFnr066Regz7cGuhP0G8A8kO/fY5KAWATIcawktyMBD3hUIveTYcyLLJonSxev
mnMgLtCYA5UZLKD2+azDF86DcbQC+4bU31uAw/xR4F+dRdcNV+ke4ls+9/4s62CWVUSrzm3XWRJU
3sdbZWSZ3ATHUYiaJmK//lgilHWDpelc6/zccVKOAuyJUJNkaaElJUGbu6xM6POl60xsX8ly4P8X
O7+OQKSa5PCyroiE9Gb9CwceK5B9nyj9LjOwqihqYMMenuxqQ8MFaeIHypjHoqDOOy86WbXvspS2
HZaPG3V8Eiw1gXf2tze6RatgyHi+JyHc2xyLY+FnHOIfP9QcsMk3LZTHVXZdnnqeFf0HO8H+N0Z5
xkdqy599CAvFJaWTvGGSlm+dhQhjF5tpPFKO2Ym0fjXHZiBWg6PzAo1GRG8wtK2vv3rATlRQQA4o
VdGh/lyYmzanJzPW8l5KPUnzeY051MvcDDoBAfRJMvLgiX3enlryJ35bSpGnSbQtae4Ms5eGalHE
SD05evBzJGpZDTae4AalqZ9CyAbaf9IkMg7HHLTVMBz0FnLFfHMJThPBVdIuinXfbAoWiyvjlWVJ
Zn0lZsiHcYObXU389Q8Ti6Hd9JZNPssNKfFvXEN081aC4B2kxPbEgBM1dvv47InMDfPSHYF94rhR
lBvQPzXM9MOFtES/qRkCqMuGJWXZuV1Md5MmoSTK6FbsN7UPB880hCS6wHNZr7x9L259/qQ3TQwm
wThaWajUrduQNWRPX9SFeA9AzIReQ+iAgLm7rcqSd79oYGai/XDd0nHPIde54EfvnP7R+vKkkwBB
9WkiKHDb1933ck0sow8yUB7+rz4Ah+5KvCvAPF3UQO/QiKx5Ve/FjnNNyEJZSKsffi+PuuOd1UkV
GFooxQgilo+P1dy74Vp39CKw4eZXE2+j4v8D4GAcksL7HdhyLUj6W9Wzq/nUrN6uFKJkFAciCkn2
2oZGEe3C6gqWzMPvx1A2/R24pFwIChF6pq4jftE7CRCYkPxZElrmmQgRZmacoaC/PX4Ah+aKon0T
PTualC0fU20/sFyKix2l2P/XxvChj3xez8UvVZ7l4GW+PEL48ShvAX2SOu5Akvv+JISfy7a50Fgy
RSccCXGE/L9KnNd4DtjxAajCh2g3RhbSo6cepbBZPHwL4M4jbDDaAgEBAOuan2pK9C7Ga734ab2x
MaulQZqghhJrNJzgsLASDAH1Z3xTSGRT05HyWJtgPk3CFN4rwyEV6nPslJXtGdjC4y4NbORjFehp
MSAhb3ZepIj3LcgU5H36c/YxVFk2hWqgHluUOnn6vfW+AlMC8Cg+AIueOgQquAwnTlG44mgwEdR4
OoJZvwZ4D7iU0JlGQSAue3rZ7fw+mx3uxw5uaKk6Xunn0LwI9dkycadgaPi6q2PDhzh5lK/C3IlV
w9dTy4RtBuhifBuy37dOSD7uIg1+3NVG8ug8LAN6boyDQaEi7knJHY5s8gTUrh7TDh4OJ3/Ld3ag
K3SKbodgkeEgqFTSrhxvpo/KZFozASYVx1iAH5nzStw+GCfzDVyTrTV345FPpNf21RwMLUl6BBmw
y7jUIK5cgR5eF0Mz/K14onnjJGL3gZ6PLpzOmsD8bR5imZIO0GtjV6VlgRmEs5vKc0NGgArgSgal
jzX7ZqJY/jsN+5UO6cQT548mOwFb/bu94J5kdhWE0R06uCetaNZqoRIX2Ij3lQIC13b93X+zTQDM
pWeTKN8Ca4dDdYC6iFJCFubT+dNA6LrWc4/kwPKz3n8xSc0OMGfyg3TOKDg5oCEawVIrZlh+pntu
5t8V8AVDIFDTVfUH3M/Z5rFZ66xiFvSvHgoO52G6qHglRoDob21ct3HkpIFBeuhDBitGpngq7D+p
z2We29fvl/dMs8cXkv0TDbe+SRkQ1ItTUajQajYfTmsVofORVF7sjn0yUouxojdUTiwyKuSDLhfr
/xURde6zgQqCJL0yuE6be09b0XypEdWhP8sCPHLx/JBuR4n+d66fRTVa+bkB+9XQbJ3M+Kse+MUn
xQvMsAfFqBXNAszFiKIajhI7NtPJl8ukAmI90i+Jxgb8wPWFGGIs1gpaj1ZRgmXJcKHqJWqzCVlk
NSccSgQn9hqrvq/jEXSqxygjxpGuegn7kBJ/o7imbHsMHbM2DvwaVoxs6F104gX6spt3terIP0Lu
SryDU8kESfcI/LCi0O470LmjFNgDErrqmyo21E2yQD66vhcPpqfA77G+LWyn25YWjlSZg/4iV5u1
92eRN5ZW3XR6ruZHd26Z9U9glHCrLOtaaYlHn5bEBBl3baElTVvUd2YnOdwJ4nnik0on7KG5izF8
sk4OaQs0GMtd2XBGSoq4r+JPwJFxW+vi9iGltbKVj6pM6gADeUceHZajnqqYVicFUUMJLAX3gQq3
GZa72aKkKRrYV8At7i/iOmziYU29dibFqKz75CjDGawyzqP6+OriXFrtvl9tYk8nAW4/ZB0xv1b8
6PFl/wcJUn49q9pl2CQWqml4GVflBCDQSQEJXZKvqtYIYwQ8H+yR5nV15UcLkN4vxWkaLxhREaCG
ts2vlwCsW3Fpg4vYLoK0ZecH8dIkv+vCa6syglbR6hrVjqF7aKdG5hQV6BQxdhO1ljs6tDwI2OJh
XGADc+IG2TojpOED7DpVGIsOxTMIUbuNuNgHmBZsRNqzXj9IDPTD7vE+Sy54QwKKzeC4WrSERcPT
t983M+m2Zk6QfwD0wIMBcqd1la5I3Bsexj2OTb0UQbBgb6h9MMm7bSqzbu75TI4ULefagJC5dpT3
jQhjCg19OWfYtd6zlGv/oRY4kcONxgmqq4cTbelTOoSSMsFg/yie/istn3Nb0LX2dN07g/EerMpN
ik1YYhlxCo6eVA8hvX7zcnOcbxzbJ8xEY/zjQ2ILh/aaGMJJSmdPz1OntLUpz23RQIpZtTTHBAYA
BM0bvzxzKL4pFObiGuaFmWNFdcTT13QHJPov1Rsz0vBRVLD1uGvfIIWzlIm/Do7Flu9QZ5g+tTxE
byyz1RHEgFWORHZCeENuAG0X0UyL23A6PGj5HuCa+EewQQamCyfMKmZ7IPxqxb9wVjf7TfuY9hpf
O1OFTYXedlWG+jfihN8LoUSzbIUp2OgkOpyr951H9rxndvJzGC2uNfPLXFNSwu9nWpT2aHgS8AX6
MlDaNGiEVBSojL3CoeKPpa+8FbZpejACTiVEZhnTc14Y4bddYzpSRzjKAXyzq5tm/EVIOSxfT61L
/+Y+Tr9D+4un3KHgZw5EDRAmjyoYx8Iq8tUvQEjFj8Zcpv+STdKz2NBKLttV3GY0KKDVckCTY1bN
k3lWdHjpCIvXHYM1iGi0z+XtA75oxouQahwfMmtXa+3L/hJbXX6iidvvsa8qzJ3B0GA7jZIv6PDh
2Ks7q5mVv69xNeRD
`protect end_protected

