

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YkmX56Hzp6zc9Cpn4dNjn+cZwcp0a7rfSO40z2OhDmDgydIK+f8dJOUxvulgF6q91Q4mdI5THu7T
aPHMCl/TVw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fuGWwt65aqpsijXPYQKf4xNDFqs7QyIeqFdDTWTkiAVBR0LW9IsI9gFpldYOIalAbyJdgg+vAbe2
BW3cMeEdrjzBPHwnFO6i0+xuJESX0JaE/5xqzXi4rdv9rbwn1ipdH+AmDDahtLlTiL+B0P2p/F4A
qiXHS8UnGmSwzsE1OiQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xBK14xUnvjBF786OWI9tF8dgHJG7CGw2bU/z93WYm2fO83KtfjwrA7hbJS3Qvci3dGdutABLhN/t
k9noi7Zlu+PEA6HcaodQyFQS1sTaZzBx1rC615e5FFmwCwGPLIGT827+Q+UWuYQ2CLjAgkPk+Afb
xj2gCYPJa1Z78sjE7D/8y73RbZHg1czi2g6CMxrsZs1YXvZI0V8XKtq3Z8xROxmcRipx5ZMouPvA
r/8WnsIIlS/3WSb2faDRH8qN2lNdnHBRi82mDS5FMLFJIL+SqwY/Unv0DYxfZ6gfk7M9eM+Hw4Ao
qCa532xALdvmwmU/o9Rtm9pn5JKLKTDqgTNNXw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
amF6Ffk5lSq3BWtaDISTCd1h4GTTleAqwM6h7zDrsJtYLGJ3rwqRfAJJof4EbJrNpG2j0AlgcNFN
xvyuzT28bAEdj5+gf8Ze/hfnSFPs+H06iUGXXHaBwCA8u9LbLnWewa2j+d/wZtHsBnCQfaBKYJ82
1FSbBFrJzg6QAD5oRImnWaooW+BjX7v5bT5znd1eaZd6FwCN+OPgR3iR84MLK+toVSaex98Qgzyl
2Gz153m00VS0eqVhx4Rika8jXeRzMCLdm+jLcRjV8UmI53N8k+UjV2SXrWKVPM1fZ5nHR09Hg2gH
BwETZW13E6iGSXZWPNYFQ1PR/gsW4cTcifeGkQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bi5yef2ETUeuuNYvxcwCI2Ry9v2sI93c+6LJ9VHM7OEn9gJVXm88Pf1MDjkB3NVumSdLRCQTqo9U
fvj3dzQqPMoQAZNV/PwkzDY0yCk+iUlYAR90lJbalZBSdnrF8FLjJCr7SdvD+WRQJc9D4oKBezYm
dcy+Rho3SBK8r+Arx5M=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YZnidInB4F10zk3ElXTvIRDB8d2w1Wgi/b/rA/DJDeY2V1QckAlNNvPOM2NcF3sWGaoC8rtkMtV9
CJp3IcLj0l5urwylLRoQI9TXO7xMsXsekwAFmYt1ijsmio7UZYH6kmq4EgcK3ua8dLl4J40gaBaC
spQHoA9jOWjXDNkOD4tQ7iKL9mPuTvRTbe1TySO7/Z9b4j4Rju8m7BjJWRya7LsI9+7nrfG3zTUf
DWy5uSs0UoXgI6Mk8QjAFJ2bX9qwgjkqhgvZuy5qFU//x1E5xj85T0nNSRLZwIXUjr4itLyzhwyf
HYuvFjjL+rOiyrQq0EWaKAi9hrK0Le2bCRxnOA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hkdrbGr7GlXiTl/rFffFMB5gXsDqvhPWH9fAlS39AMy+m7ijia3G0/5wjHO6ZNGm/yuTmZRCTHdx
w4u7snT92L4bPjmaGI4NGoWizChFp378yzkDk5sPcrIJ40fl/gbNniBbtgoFXhzAIwyzyLWuLzXS
pZ0Zg5TeYnqaFmyjsXWkXThQ+hbpwb54w+fkGDMu4q6lsx4aV61wvllN8WWkfH5dYGD/Ze6UIUaR
sInWgwXjKWJl3twtWos3sNtIJzrSiU4um2md3N2bI0NvLk4sONjHryu1tIKQ28svBZ3+ZOEcRYWN
YJGvWSpVAPaK1Qrma6bvobEb+IN+VJPzERAcgA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dsxVpfHRBR8TfT7W2Y1zGAxARhKaa56bkpyUEJZXL8JLA6mh6SWhwPTGmK1jeY+spltqcv7t3W77
KAIaM65CRU5cyYKzJZP3PDam/mK/qS7DbQDYq+GbSQTOD9bK9qwbI7VF0M+WJOPqAVpMN3VBKbWs
HtxVlEBvx+uLiGEpaTx1HEr7KMZvYi7Iw8TpbPz9911lqOxZnpzivraSRt2VDQsmmZY96nuuTQjj
tY+asI5lxKjA0wHd1ddDINo73/ScMEnmfsOJQTaqQggnqpSoLVFvQ5ZQXz54jCM08sDyx0auBpQL
1ss939Cq7WR5hEMnH8B1MFcbemm7hv3oraO+7Q==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TdXZwNQQ4MYnYzKg5OUj4AXvjjO1zxA7Cmablx0YtDpsF/xwqboUFjcDRckHAG6jOGkHbS9sMiqG
vsqxx6CfIHBwyhyT4Tc6uYs4X92BsSmAIQOWERGgqd7AzFuIBzxalyLIsis0Iq6T9TIi68MHf4Ve
5iWfRGAFrV8RGPP66eJAKnkTQvb9qUXQraIQfQOu4ljYg+r9ird4eNrMsF4jewU5okvymlkbWeWl
eZSHSoFhWvwGI0VHSdoHH6hwlV73zsfQxcMSur6d5wSAzw5RYkUkWYdXBIkDzooYeVbc1JjQURRe
ODWm3jgqKgw+igBYag3HEfZjrpicmMffAbyu/Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 558784)
`protect data_block
7h8uQ32Ypd/s/syC9125auWy5J4bjJtkeFSVGB2hAkr2iVQaNbjR4djSKan50uHNB2UQGZeJJBdM
Y+3jr8KWxqiyubRtr01m2KgJj9n+fGi55rz4XX+oWTC7XZ857XVJ2wO1x4YTuo10f8zfMD51/wjE
i8pf5qCBn4pBlaLozY+Qxs5M4cAtKgqf1TlwDxQ4bBoTepUiLPCfPpwe6inrhWofE0q1oMfoKUfa
3xPdpIyRRmgGd3eSC+mfpnkzH7cXGthJfVcOu7ld6ntQl3OR0ZpbBK+K7ob5WZLdKMHF8tFHVKFT
u+eh7IP/HAtFpDY3qQ1HPLD136q4BmHjL2IfSrO6Cw8mdIkeDf9d4djk8/0gyVCll4UJbQRRTrXV
8/B+sBCmB94gs9cJUcYLkadYEI0hnnIzZWiY9mkOJlDn3Xk3qJJsTnpFkwPnpDLPm4KOs1ZPdwr4
75pu1YuWull/3LcnNJRu/H9IjqFNwfEiSQ6oNkKib0tl40jcpaYb0ms79xv7EOz4W92+wCyizhkb
C4JaTNsvp+eQoRRtfVeKuX3psv5IDYwh7o8XwjB0mOhgnchqbpCyVf2fDqA5PNFU7/pMYf+f0x2S
YgAcr+1HRXfQigbBdc5FafjsXphEPvNhjekyFtqi9x9J2D//ezmfqkDitcDtdCOW2Qj0JiI73nCM
LIXzqS0n2beMg2xLfE4ktTHyk9qW2k2qmi7vU6qAcGBHbmmgNjaOG+MpmEGFM5CNT0M1uZC8dRzx
VDLEsKF/GBr2V6yiBHqBQ0yeRufOswpz6ItZrNe5mG9Ci2PjaqkDTEBq/0jbRmFAMhh0w2P9I1Wj
uMwVa5uXsDkC7YGNlzFYUWFph28Q1Ev/IuVOEQOg+N3mn28v/Fg9W1t6g2zsuK4fsxOBI7rOAKKm
4HxF+Y0D/zuft5p0KY3aiAXCk90IDhicBfNTMC3TVFcaswblbQUlzfvfask2Qa2NGpFP5c6S0wgz
DGL+NxLTUxHvHE1Ajw1/MbK6oBD2HHm4jUvDKNkcrOxUSUPvpkhmouKGFlsBPtvey4PUUV556B0q
GcML2sZ8cZM2vA/S+8o1yEuobkRVSsXcfWzWQTHbwV1ENkwaK6iWSLH/0VrtE+NLXKRZfJrypYjP
hTg6rtIbDc0SJv/dsFqYPOKkwPrN/5c+Oy7wzRlnrDHoOFBddyGzYSlb/EA5qGiM2FcLdflRNcvv
9aK+wOw8HYxJ5wfgAr/R+KaXhe4ZFJUJmByWyVFLvqhw1/9bvwSiUdsWBPjf/XBaKKE/yVeVw4b5
Nf31Bk3z0KTeXLlcyHup/N3NzgHj32jStAMj8wWJeqEDHRFiMW5fZG8Bnb+ClyZS3DR9qVCUBDQT
Fh5RkcA6lLE/AsqM9hIHh8fbQ775FUicicKJCn7UeN1SES0aO+i7vmyAJvIx5oeE71SnUhJ8u9On
5DJ2edPNWENH0qJbjHY7IJUPJ/SltD+WPcLsUqyF/GNnTqhm2FbPNme3gPRJ/otl+i4WxysaBDAb
bclIs7L878JCvSjE2YLEeTTmZXz0d/NyJKTLcW5h9K5NiolGKX307vcsgGOZWgbVII1ALb4vtkpA
qvCD107LVstOS0ttDuQT57i00Wq6EDx3wD6hD9r72dYdo+iQABkrQGz58N1qbaytS4bt7EaWMde3
+bC7cwkw0DiT4fq755kHS1LiF85LJmP0ywkDtHh/2QgksGe9KBZh0u5vJkoWH04cp1j9kTKGYu5T
srRwePiFplx/GIrhuKc7hgYShV9f1mFBXJhZEAsemANTrTVCo7HWjasfGLTF5YmxlzcMiyaKk3GY
eKtJazcVITYcCwO6AtjjNeOgiiCTy/slsTPV/nRMZ7nksm/CXaAN1zuPZIbj60/II8OTcoe4vAk6
u+/iG4zxX06MWn/ONzLnTBtLdJZWqagCoLZ/YikLtrLFcBy6dCSnp6fDB/xuwYYuBud13ayoW4yl
gWuKAWKusg1h98RgU5rKfLzyv+74QvTLVaocPGsezSNGvkkH4vo9Ef4u4ge1G6NX9kgcX/22Ow1Y
siJX9PbFaAh6tPWd3WnKrwnWiL6EVlDG68e+o7LxA0nhsWXlZIXsPNgnBCUwWtN0Lg16lFUt6Oze
L1JPYI7q1u0dsWjWgKc7i9PCIGRwbG7g6ua9zioXWDwNiQhcIkxLf+h+SDjyeyA3GaP/J6Qkl7pp
XI/Z9v026VSQCUXNcGqacP+YxMHsjVLR6zZHh2ZCyIbBEHfhNeEl9Gr3v1mk8xLW86htNiP6dhTd
dccWvapoFPpg40B0XA5CqdkzbTL349g1TkAHUMGv36tGTBeg2g5Al8te+f7Cg8CT8F5s/FfFbckm
rSN7PD/IwpfKaaBvy308XcLSNp5Kc+0E/C275+VGKczQceTkFTnSLJbHmeufRbDfdkaagLRWoHDf
RrvVoGFoq3vpEphzjZIDk/n4hKzwFp+ev1X/y1DccoE7PuZUnIJQqzuJbFQJLpkVa6/WoqJTKhbG
AAziwiT7RrnvLOcDwJKD6NsmI30ZBDzxkGuqEjorp39zowxzGHMMmdoJnM+8qNoAd+uQ+zsqr7tZ
ofQBLer3XGoC0p5nzdEfu93T4VfmBxGNJXgow4isyAt/z2HBNvtHNYnoRfZl7E0f0Hg2PzQitDYk
cMdyvOt8EUSvVaHE8EfSRPwVBMnZDki/WYiK+TBTmap1BEnC38KEnzRQ/3/mqXtcFY7vYy5yZF0m
JIMj2LIP3OHmxbo5iiCrdlkSPFWOpLLJGeRiwLtQEfLPJ7SZGOIOg0k5fQD0GdJ3llJ2t0XYX6lV
79OSaU+MLSy99PZwA0x/RwNCxoghB+s5bviUIxA89Qa1QjX/CV+k4UL5Wt5XM8mGKUVvXXGq5WCs
/zdI74lFV42jentjgG8sh/99Us/ESOd+NSXLYmD/TqtaYhA1JK2yLhhxOhP2VBZEy6yXF7svYbfG
oCnhnc/C9PK2/FKCmeiIabXyJ+bp53zJDigkhHHz/zvjgLzkix+NuSnxnKfqZWbCrQ+V2S9VNk2H
EkaoHPtRGjvbuKcSuMZ67MKtTKmcEsFjBllVFwdGg3nNZygx+Sms8jeEwIIswBbf5Q0oOMkhp9IK
rdzEt8UyBr+nPn9HuY+sLfgR+OL1bO9M8A1ouAbdunVnWo8d8hp0aAl2mrZuroPW5F4XmI3Zjnaj
vRWrmJsboYwI2iDqTWsX4qpVVpBogXLwwa7nbSpG8jnIocTRHCM6UXYVxQVVyoyNydBhrd5rwdT0
2dzrCXNanCFd2t7tNtx435efxslfHQfOo6rwqEB/CUY33JnWTNqaAHkD0eo5NmKoGQtlto5Y1BPn
Sna4hHnpB/5pNw4w39SC4QL2iokhRsyDOXKUszz5VdoBvlm++MiADvvmzRQQdfwK8tS9y60EAlrE
uhxQQGR8EKYmYc5dd/4GOA1f8Qpzl130ZkB4opHE6D4V4jlrl3JRZ+LAsD9hWGw3csXLEnlXOXZw
E28OdBmtmBFtnSKjeq2VfeC5xQrP+JSX5E35v94WjNBGDSHcxAx3032FepaE315QQnIvqAjdtXps
M3+kZ3RxNFG9NfhCHyuHrLnoYayFafdI00HA4Sr9fCNuqjFJ/+RAajaBp4NquuwnpHqls7LjJFBB
kCBWa5BWvDufB/onUahhxveYo5CZXAE4DD/++GpHTLXwdbb/aMAWJt+EdBmNqE3sFbzYs7HjEpL4
ccL93ZFs7fVAs61ppuNkJLaFcOzL0UG0Hh/mNMNLi+NgdKduXC+wmX2Jmu6YQ6hSDpZytaoDDRKJ
UzVgS2no/+WLkvMLVUydqKxWGikiihPutWaQ7GXCE7yeu9M9BG4ERFQLinYJOyUQJ6UY6D/1gqXa
EvQwecwcBYDF1Lhl5Y9VO10XFMbje/r3UTk+U4SBn4mI1008fN/1mtBiC5vKZDUQI+RWmKTYPL80
j3xomNhywf0McbEMceTbZXD7zRAjqOuAuQrg44CNQ6a5HDcR9l6ufk6FvPHDVAMOEGXNEMUkcAxb
BegwL335Q4mtOS6GRZBW69VfSl/NlKIijyfkIMasmCFvcX8Rb9ay4dew+JhFJ8w/tcXfVwGuFC29
W0j/oh6zAXGFNlMWOiPaWWNmDixbVgxhtDcm4+ASyjJ6UT6CW/tzAvvWFOQQFRYtdlFLtKuSGgCz
b5xJrc76wfwLr4BlCsXW+Sz8HYwKJWZf8NLbriikAnj8E5+5weJinhSRABB14RMq2gZVm9CYn3w7
DoX9QkTfHv98+vANHpakdRtfCD4DXqD48GB2JiXYfBunzJKXMy9GTUJbOp3YcmbIbbmj0ZvtD1cF
1XRXa0ycJBHOvEV3JzuPQdl0j4zSlMPBHGypoU7JjiPxaa0CwKtwQorQbkhCW8ayRASBnOFl1azc
yMtgqmYUWK5hrLi5PqW51C8OObFXF7SfJz5qG4cv+fIQLy8aspyrJR9wiGU2fSKFtKECNFFy2wLk
/R+uPqqmL4ttZIcQkAYUhNiQq4lpNwH/zRlgdn9wH5/DJLx3yGr/ixcycvci4BJcc6Afrqm21WjD
nu7z0UY7u5WbqBgUFcvR2h0pf05znyqk35fVxqCcGdJcyqFHTN0Za902RIchRdJG31AMusQpLPJ/
4kqb2qG9inEt6iS1axknc9CnvR/MSA3Og/obSwPRpGXA1i4Jh+pOQIvnN5uNUxp94yC035wphpjj
JnAQSKdPkeaDIMGIBUiLL+pA8AYv2+u1NRzLUQwDFpUXkzkA7k+WtgX7i1uzT1ME/yhfOFNpfOxG
HJHRrtqXqtsu4XTPPvpj2te0asuKpEVcGCB+M3KJPIZrsTsukPmw8bCSaHVYSLLBAQ/f9jqBmRxO
dWWS3fOA+tQewdrnLOBIk90E1qGnrC7QK+nopLMazZqxVZNRGLvjqzfV4VNly/F1tW1S2g2ob82Q
g35qDRwCXIeOvaOtHCwQSKtY+QxOfdkmw1Nfzapue9ztiwixaHw9w9/YeXKSm+JkDQoXDLC81Ri/
TBTBvDOlZMnGXjVO3PF1NzRMgz3GZ3qcYGkn7jtl2M9uKTOM6Qj6POHz4shn7fEauCbPRWlPfIwl
dsJUPgGjF3FQkViqHionZnDr6fWD53QxSFhj30KfhcAdTt5hZcQz2oOQF0tuGILPELDr1TEBa0W/
m5FxJLd+njruOmFE75D1UF6Rn/NX4nrL2AnQDS35k4LN7ES3a5xvo3KC/fiOXLB5b2t74CKcdAgm
YMLkcD+ddNPubk9y30yosV9SgrY3Jtk6NIfwu6mTW0jQ1FBN2PHYG15J1duPNU+VIR0R4e20/0f2
6UX4o76f9RMZMA9UdGqBxZjO59zy1R+5j7K2j7HwwZqXCVFj2qZGJi3gzI2AQEvtXXFNyCrKUXFh
qEoUHpKXl0cNKXq+D/y1viCuLg77AvEO9meDgz2BUSqmzztQoDAi375fL9vvxq6u0XS3iOO4E0K9
/xHP0b7ZHsAw7hodFcnz2BIWyZL8bSLOPwbangptyPZNi3VICoHDUgdX9uaX5PgIMmO6lgVeQulc
4XhRx3ztlrgRsaHgzPlIs+XowLXQBMMZViqcnOMDAbdcUsFD6Esdrw7FTOtfuJalzsg0rGAsnpzT
oNakC1/TGKrQU1mLbvMyVOE62moVR2NhpH4O8ogOMfUyDZ3JBqDPah/qBGlqYnMM3Xe/k91KC9A+
jXmwqXSpnR0lyhMfybVeD+OwNmVayrDBUuXX7H+FrrFLD+Giv49sfBQzb1kQ4HppNVn+ZNwCbFxX
IcsBtVxLfAVgvpcgoogImjVyS6CiZbQDJZ8j+LFzgnOoKUVb/eDnzOfOG5/GUStGNT5Je834+zJI
MRR52j1yyhet0tnhdrx96HEIL2XLG1tSRxGusJEUx+4OItoBqcvwAHQ9H4VNJoS/E13noPUhoeQf
N8yFNTqq6kkNXREyD+ZCa1oUCY6lOyRKdtLOGqrieepKzP3vWEb8jDKeVDzEb5vSgx/C+3GV2iDe
co4/otMvmOMlfE23KVN5IUKJmZDVLlDSBCGgnwAsI7K4p3N3EnvXqC2z1Fl3CnAmxRWcHwObQJQj
+awTypXFX9A+RGzAQWiETXSyhM6vzLzu4+M4Iqi2KSXf9faqh0G5Z8tN5CyYA0wVe+6khVCujqZn
WhKCcA2jedmBVr2MlLIQMGXRsXqnRu7dgDwlvn/lPRoING1csMx7eFAusFimQd8vr5tisWqcHR22
Z/Qc6ZOkB6PSO0haSNcPtYPfu3l+tD1lrn79/YGbPtJlJNhnHtDdHTIIgrAZC93oxiEL4dc7iohW
v0PgvEh+GIcuhAUn3I8gy/GPAtsCc9mN2s6NvTfCBJIVIlvoldmWs8FsX/2i9joyNLcXSwLirFJg
/9tGJKodTyVN7a0Gd/Yw9MFCQP5xrS78PCFABm7fwgHyxLn0BZNScRiGeHlcWRHYHeQCHRMMuVGk
omKyG0zUxqz1cGLbVBslUbYxOBmAg4SjEE5E10Ng/j6Taz01B78lDKgN5nJWZVovMuojC4j1tIwS
60otrQPW1gEKfQMc7jyLe+GY9Py2Oj/xX90oX689mXh5q7Q6zg2CRE2Cs1pEd60xg1LzJQe89HcX
X5ZCqOjRJ1WWFwFv/aA9QzDiyEVm5t3Wc4SMRx+Eo+BlLM+rKd+4ry9nX+VFa58F8L5dYLebFQ6+
6R5s5EMATi79ju5qPjXXYtnRCpnBpKi8lWagDForgJHwuJ+LKHTcJ3NZliao9amFRrEuz0z/yowb
GGNA09Cx6wy9vNEL57Dw/G79YEphCndLAiq4l8NFTqmwyZqpN28s8GMSydC6vCMmuBJi6KKpI6vo
iowvKcWOi7Tl1kLQImQ/9bK3YanorVfWCYDLwKsOixtuL3FXWVRMtlSB0fpGGexaX8IVnDWfY3cb
4cnUSgUGHG1Tm98/Nklw5s5aJiomHhNQNn7sQcKyF40FqJGf+1Iqo5cTQZ0TQrcMbVjy8id8BoME
Tcqxb9LKkES4MmNvyhqAM/JYl8ALn6FS7AC3iaAHbxFYViPxP8hfm8lBOHQW22N4V4Sgtu1e8Haj
IcwHLx5Z1l/CgL5uK7LvvIEhQ+p4lIxbqok4Iz4X2A9XuzTS8xis/cNKwXOVaskuJ3NIjN7nMqzF
ZDtrXQfjWBLj+kUcRFZxwSZpIE4kZx6LgJgbsFzprnSSkkJSBR6FSADCSMDEBs7AR83kKqgJ1M4a
Go+/ysyx6I01YWiT9pZwpe96ySNOp6mOgxXpTFoVBaFcJw66gdlUhY7PDTWaUoW6VGOIXDhxI6yt
NHvUSMqwJNrVgqj33eiWiYt9+50vVAFDVfFOeoTWxGdcZmRJsfPjQAADm5tLhRb+PhCCV7eXhp6Y
GigaHhUFILefZRf3tQAcKlly4C/WZIBSW+3cWtvHubpwVfV4I7LEEudc8TZoazF8Mj2IW6y8i+9R
cVsZ4M+jQCkenQ5lSpCZGfzCU6TOk3jXPHyVw7jNbPNPEP9PDw83XNYngfJbUnQD9AcFUG3dX9uR
D84JRNhkl5iZ8MW1mr3BTRxgYMUMPHSPyK8jHVB3TlM9UzTtxiAEflNNblpozWpmAt/ju1JZGO3l
gACRrkGzRgYJA04t2wRbaDVlgc0LjmR6Up9grlEcbfQfGsNPAKQniEi8irCT+q9tb/V/JF64EDUH
/qRz0PBPl4Pgxf8Zibts1ZLU51rv5RtdqtTejkbObLTQxn1omPn0ltmzXg2ZeAsGgclqI+l4Qd48
v83XuoCvzu9+vAK+nOISBWaTKq/nLyV4N7/8mg38Vvm8e8rlz4E7Zc+sepd83Z13B40rQH7b7iQQ
aBIEXuOzDXfjKRYC3RCVkO/BEwKP9GSxr/wTIocTTbKgsTv2vPeY8H8+P1/ufimn8l58Pf5GnwwH
0d5oEIaheJjqbBKIn928SIRO+AeY9qh5QRZyMEGopgnWNq1cP5CigOnAJFkTQ+qa1vgbf7EAYYct
f4JVv4Va4FeEqkbP0xzlpYjJBq5YX/C90mkZBa/TtfiMClw8+JHA+XiCIlOfwyhv0IuiZ9m6obeF
zwQ9dWQxhNwhVcGddtWBiRkAWNDH3y212ua9FAOfTPsaUbPXO2NdXy5DFG8gBgyjyHex5+AV2+zw
szAhO3z9A9FElr1r1ewjHcrFGxxoWU3Qs8Z4hmNTR/uMBMaEnGiXNdnusN9jZonHqfaXEo9835OT
quZJJ+xevWEpKkixNR+ZYkGIfAESCyv7+dEznUocJe54GcHrrCs1XjKO/zX6qSdtYsAzjue7AIDP
22uCqysPnj/y88KWdIIntvXhF2z7FsHjgTyAJ2gHFYdQ57FSpBj8zuMq/1LpFybi1D5V24GkCxmh
goOiXib4vNVvG3hPI084G4+RP1ZT+vTkQZv19mg9Ai6Z9MZJqUBKCajZGVM8g1q3/7lfDSG/fsNy
fC3vb5UY41waNMp+NGKxSfyygqYQfZ9WNZ9KoZqNoNo55j/XqOdiYsUSGxVoaTJhAER6hqhw7/F1
rbhEaKg9E9r8+IeCwgcWVOD146uZpby2qdzDt2MT4sEMBwTTsEu03qlsjj3ulsgS2VzdKgdv7C7f
vBROv9puqnm2Ewk1bnJSto1ue0phbCAnHo79vjUfDhoVC+Wmlnxjv/INLmddlvF2OwLHup4vROxe
3pE11cThZ9IqJegbmQjPmKmgF7pMM3x4PAMkQ4ZH/ITBM+pEfd4FG5VYOl3mNtsLzg9pTiEIyWUz
gaMvPFxe/V7EVfKX9FF8f3WA9G9835XeTXpmtxbP129oPe/BGX9bXpFAdRhqCP8JbNdlM/Sk0Q4C
WU9NcssqJJWIyWqnOhK4CHq5tSCnNOK4tbzMTnolkgD/migyQa6yLJEF+0nJYxiiQWFNO8UfsMKJ
IGFG1bVo2h6NZA3qdJCbeIHAgOcfZkar9jGMj50k4E2n4RC8rkcVXP2hrrsX1iSHQLr54Z+nFAFW
POaDlQMHfG+FOMSOATK0Rxmk4L7o1rzdjjgymWmLpTeZEyVVLfWGpz1sqfr2qmNUNbKODuQ9uabd
HUfK50unypp/5A+vk3Ttx2HXrqwQHjwKZAoff3IbdsGFGxNH6F7W+bJrxfiZ+UCVe5l6u5LGH+Z8
QmSeJWr88RpEdKEvmMgmuhHkOyXV2xaDMhRjpnleVvYld3Dkzf2H5zwrUJKtyfjyS7hGzXmmZcZi
i2SmPEml1dLIOpugUk1D/9PiVK0W8x3bfcqCaWr+IAHjPp+r7qYC20MGHoHIq1pizy4Gc+S1x703
Fl++p+mwu1GuxLmcHKEfinGAqNqc2R9I60Sv1oFtnTt51wXaG+KIq3mMjumdeP+2NgTfv9CojTQM
iOea1R04+IB1FQnjXUTQ3f7EZWluyEWcsfRIDXTO+PaVs2C1dU2ZnMvyOVzxy7O5wdPfxcruphFh
/lwrNQkwZojbQGHDhX8/z5rZjhtyeGnGTh2TKtVNSwOSSmMZFBb0dj0TBs54quNrLHj7JCtUH4/S
0zxGUkFI4x7tx0B4afDdmej/xEk0xpEST0Jdasgqtfgy7wOT6uR+xe3tSgO4nZ/JQ8qt/+XhF4kv
ZsgJ+v8JWldhdFZgP36s5yPjZ7aYAHcyPLnaYkDkggisQAfSrzd+X8BNMbLtStoEg+lkTdDCdO3z
P3gCg4h0ru+9MN9mHCY6Hi0yA7hpHLpDI+/WUGauXm9T7o1t5jtygNpcKEf3j9mRQ7ghqm/XPkCY
iC0KI0Hs4o0s8Ql0kYoOs4YH+mYflv10VvSyHV2a6UH4Ln22oINoOYperqubfiR9tkOzaoqmObvM
9oBv4dVDAn0vMD3zxypwzt6VsSZyqCMS3BVD/snWqq0She4frtSkDxwisr4GsKdiKsaRw29IaJwX
AfS3eRX/D2d1c5ad40apojp2nrTr8DSVc/v8+Zgj2tU8efyx2RkWxDmQdh1uhZwexyFEGqm/3Ukt
q/Wba0PCx98uYemFTrZwmjdM4XOsKBDZQUi/PErPHb03359A5HPNLCYOenlTTNf5AIw2OYo8UPzm
U/Zdr97732SfGg0bkFSOU7F/hooh4hIHhgWp7sAx1XNmDKym0y6OTC28bxcsOj4StAQ02n5L+oMo
nvvFKilUNzraohXUmtljw0rdeXS9gx0WwQddWLU7YFmLsVrF9+mn4mrjnYcCt9DbkQG0NSp47X89
EDLRUMDeUGUh4SBhdgSMRTUIp3pKnQBSXETdD8GRFsBHfLku4m2qVc5SoCt6hP1RRmIC4EpHakqY
Dfy2Gc/UGnuR37/M9aEfuxbFkDSkDm5IcoQ3UnFd6hAQ3RmAffnzWnB2jRmOYYFPXe0C1l5n5gNL
XtqFS71AjGkcUsH+QR6k6i9QLLqh1jxoFL/+ogVbKRiPTdVYngOTXol5lghpNsvJjDl1xJB4+fjP
i3BF1kF4Q2/cQ4qGc+t0v74FzXTTtGu5AX4YtZXXTSRAl6mP7d+m0qHzt+N0yZ+joWU5p/+UHLAG
pIPOnclLw2K4PEQYDevjPZ/SuyNm5BgWTI2oHlU4468FEuRZf9moyMekhF3sk/gtfdZtEoXdghmS
9Dr48Hcw4HQrvDH2q8jl2jNJ7NxeDpmcqSzCy5AMSKf0WdaZNFdApeqF4ScxdNuRKJzw/b8tHijN
IlOzE6do21CUZZmKJvhBU6Dj2++4LLwGBzsfQO4IzO+UQGmeQgKilnTRgCcBH2VeFK4Daq2715S0
8GT6FPTmIY4oTMzkzlHZrJN1U9r6OY2KY/ibtx1/Wcwrf8fWZap3WtaAW/q45soQP+iXEVSa91bd
6GAxYFvfSa0QNElmTlENVmA8nOyyJ3TJEDLphS+ZtZSDN3nQyi62v8x9l+cLLH8dLJl5JdWWi1mi
rPgM+gdk0+xMrq6R0/oEc0WwHZ9bdLBKqyX6FhCT7wrWw6wUcQoWFTz/sMP0Ojng3VuB1j9GQ9kz
HwFszi3qkfW/xLQ3C35QxFG2dSbG2jySsyrbzxqFdVV9O02BZoR4bnvxunFhNoBy6enY8N0mG2On
NyUgpk75rlEXlyrbTKbg2sX2hlYMUcbONa/DYeIqkpbZMHUWzty6c0/t7aK4j6Y31kN448DfBK9R
DEcPwcF8Sb4hfIOGIz3n71hxHJl9FsJHX72NlSY0YyNzDd6eNJHOyTel2O/W2kUlggj384XCe7bT
6qprYpNf191oQU7A6X9cv3DVIRJ9tHbdnCDXRpwiPtxEdhuTYz83NMJ+JaW1x8i8SctlcwKDdv/M
rEDNhpgD2ihvvWRDunrAwGYbZg6NjAQe5sWCaJ0VZWB+jEoNj1chzLEcnP/DQ2akBGQRgG5zJHV9
map0Fq6IbYtNXOHil7W+Q1beW7wAztlCtOIsNWyNAzj7i+KzlYQraCYYypdIQT6ZRTTzo0Cwto4N
qyHH6/+HG9ER7nn1WpDc4GZaEGV0GfQMhvaAFitQXOz4hLqoLyG74F/jJNLoguH+bCeXoKDQuz4Q
TQeGh+jpX4gNoubOjWoIgj2UjzA0QeTIPAio0S0rdYDDY5YTEKMgNxOti7uPx/vUD3qEIZXUHWp6
c1EA1Mmu337TkE9MeDxtQ2lRSxMFINahPTb6TyNOIlmE7gx3Evn4WJ94n822k+RdXtWD0gnRxDx7
23Q3tjf27YZmg3waanDMVPpF+sMjQ9M1oD62UUqV0WbUe8JYy6LXvo1yG/wMyeQwC4Z+QLd2kSTh
7TBSJn4Gr7YBf2yKrhHmaqsRfLcnebVO3YC+a95DvAtcE4jQKIvDPDib7Yj/NY3cCPgQTRFagXRQ
fKWoF82nSjT2iB0mG15XpIlXHbEfL6TTmpqbJ2Ujm1TUqdnpIFRsmrXd7XbcSG80Gsd85L204bcp
wBe79ym4PG6aZ4wfWTa73o7PEVG4NxjW8EOkwqwa1XYSjpBbpJW+/z0ppWyeqceZYwVTk/aUcU2i
kn7uG17HfIucJ+/AnZMUhX8O+6utvUyLpGfSSuWpuKo3XObfc9EqPnUhwJCRFG11sMVvN9WpGFgi
U6T/rvNnYXMxX1ojfoJbbkJU2n+mqMFg6E42IP9RtuTxK0WZNr0iHi5ZAuqB9sGntPnSPzqNFczp
iQhWOjVCSIrfrycVfemhUCdnoApFRBvtR4bJElIRiSJFfpaxf83SCD2eQ8B1OAkRW3R/Z0L3vjc9
EI2LG3hchcR8l254g03Z02CnSn4RVK+nuopflMRDdEcb4sgoT8FW6quIAkcETMng9mjrHKequ0Y7
r88RVg4iStq4GWtSegb2sKO2W0GMB6FVTc9YW3OaOoqpBkDOMNDBi46wcXMm/HKwbRFBi1ADr8Tz
tyJ+d4zDFIm6eTbHqFpJbX9vJVn1/25NsLUZTzu50L2gqHJBo3owERiACKdNN1+xyKHsK/PArjwU
GIa0AIOBMJREpxBWhKeK0CjCDU+Ci86nBqwPb0yyPu7uPV2hDJee6YXBi8acts8/1RA1UVCfHjUB
CFjRnO/BqpDPEiKKY8fKFRePS3SYQeF3b5VsaES80w2FZ29YX3NmyEDHi+QdkqQicRZPljCFDhb7
tWnT5p0gGSOWGXoRvlhq/PIvLyJMiZV+Ukp8qKWmUL/w3mXERjJW4XpkHx+snVixfItOBtI/WX1Y
YH0ZrxfqMQfPfiKQt70PscBKS+VWvxxqUPFmQubqVWzeInzc6yJ6Ya8iAK3MiySbFGu8MtDJxOQg
gRsRO2QUjrbmVUJb6Jvl8ApM0a4psrIM7Dcu0zyjgUoJ61m2T0HGiLL2nyuqSi0W/4GHdKHx1h/F
LBR6rW0u9vW8WtKPhVA16+Bt1eruDwh0wP68pewf+12bosFzak8LXX8AO0BZaa4yGEUA/hGlEGYa
YYxilw5kM5zDNc2owWyvYwfyw13NA4wlYLqx8qphCwXD/Rgf83nmoUIeG74WGM/7YOCF/3yOneof
XLjSnIVHnYzG++ZjKYZwWJjkAH+FAEQ+Y1fl5FKsp4vDQz7AnsM7sUPqQ6SB16RAOLt4HHoK46z+
rK4WMDHnaMqWvwFKbL2ZX9k7BJ042qzQCIcgOLUMjjxQrh/iWzpsqGfYNE15ij2v3QySIpykkrQc
aHwNFQGZg0jkn/hyYdBAM+/5T5ATmcyq0ojsy/Uhf96MF0AngdbhACSuBeHlzB8/y3Ut+VrHu5xY
Wnp81/YsZ+JlfhQwS/lXFgAgXwtMugS5W6qxz8lPOMvTh93UEvAYL9qEFNCf5GtDIxY4B9w/HWWv
ZguXZX48/T1diliTrHT9+P6lFhokpJm4g6kZppLVJbcq4F3wiEYkP6ebb7RNPc09PN1C6eM/t36Y
Lttp/HpFBVpz2TZ8WvMT/Mzvhr6QPmx7ivxjr1a4SZqBvtZmEuOn08yn25pEElxpHLyuT1Y1XJA3
zRfA6ojBDGYmiL7xBaZwtN9kfQYcz9GO5gzUjx0+ulgJ5vjQluyENYShvXowKM28DevULT3S1DoJ
VFwiLUPBF+1vZ+wXiBRwXUktMllTjeNKdWCEbbgnDbMc0Izan+MMAOZaDlFI7cncnetbNERzl+3D
j7cVZ+M+xtMpsWlp+ZT4RtYWt3lhxgN+sqmMcwf70oluXeMru0UyRMpWvSKU7mp5oSGWa1ps+QUI
DSP6BJZQ9ksm8VX/c9MM+75ExHKNi7nG8A57rMlG0X/KwoapIzKiIvTK0OaNJ4qs4BRJNt9f7QsG
CPqh/7GuF+k5w+XZTOq83PaXes8IgHSK2SGXk1ygUP0JLissxyWj0tRLiEiz8dWqVjfcoWETNBfe
AXrrglK/ln0K0Dktf9vEKCW9Xd//fE803toypDAu1PvpeGM63JSfgZjYGh+aZoPZlglLyZeQStgi
TFn3clpBaUTatdudEnmVaVBMKnNEYDtIvQ5JBvqw0ScWIH+Ugtz/FKbMnzBs8/JV4MQR0pirTa6u
HDELJhgVOa1yQ2tx1EsLRHsZMPq1Gkf5chHJGeY1Py4TqnV2FYH6g3Qs3U8qdWYJjIZfP8oG42sI
2RytpBZEEZaCCSXDZBrouCYSR9iON0uLCCagrWZ+TqGvSZOwBw41DMH6QyPFsXbmMDWQy/cpnWUn
tm9M2LHpmZXsU4z9jWlPIZIKFzmqgHMLfDJWxOU1XMpFM0N8Z1bbKRT/HJxuDsVeLV9vtDllb9cO
IANDqBSHBMiJ60PPS+v4JmDDlwfnwmzDnEJXxf8CDaMRQUjpLFdG+L8MP75h6goHGhmnKC3Xsa5J
bzYhh77EMZ9LMZKb3GiMsuq3+Ky7B4QqSlvhr9Ay0BN1ICnjfDxloK7hj1Yu58OuhBKeElQ+e6YG
PLdiRWrsbsDn4PByse5l56Q0CLtF/X38MocruF9lQ201hq1u1dNaDHoeooxF3nyjf3dFo9CVKA8Q
uGev/ZYVnFOCgM+SUP9u4k7GfoZx0IgF3Y9nh72yv+wycy+NJGalkM868X+8T2/TX7pM2u47Ry6/
tFgYkXUZJ+am3Dsvnl2ldFxUxcewvgT28Raoyi3wjEMXMSmImDlsy5lH4AXCmM+0ryWAZjF8diQJ
56DaevYTlotWstpQEGcAB6rHWt28bt5yXjMamiMSHGH4oOKxZ2Q6N+MVMIUHKvavAwOWoDWygqfA
HSPHM3pmvC2qzdtZQ9F6BB3pm4tUgUF3H9UVftFlFRJxHCIy3pyuOjpARzWmIcucdFksUzZKhbtB
CPALXrOiZeggjK35N04BaqbLpMvfcOj/Sp7w4zM7QU1sA5dCZNKM2TnGNYxPCGjVBMQy6mYh1/Ad
tJ4CHlSXxqQAdVmeIzwCjQg5NF/q5l0ODiEbWZ9QmIqnqbC87QUes0DVRPzmnETxUGw2Fve7wd8u
WVR9u7IXgiobPzvFjUsVrkVEIE9RflauNWQqqo8Te4ZCkvz4zBl0HCuLudXA7293lLTQW9gDY3Zi
UhttQDMWHHPvmfQJTA4OfG6WYHoK8HUVM7SSq2iGRs5Q+ocEv14by4AEMujWTlMoKDxV37vRXbhC
QKQ7bj2DcJHrfvbDQ2vy6dttxpkGlb/wdkGrGaTpKvKMV4b6/ZxG0rO+FIddM1C7ancDqn8tKIyT
noaiP0zmgEUWVmrVydw5qk0pVxfiah6f4A1aYlUeikYCqOXVyBwhKW8G7i2bj80hv+/UetluQ5tu
uhGjDFlUR19pHut314vuasDaT76mierSsWpKLdMK630rK5T9tIJX8iTAXBlwXIR7L11XxFBOvUt+
c2Cfn5Lfe9ryci6ZzVBVNqHlq5wKcZnyymIS81L/oC64ATiBa6BlyDw2tktsUzYY6iyfPiQwM568
yYBU69q8deLoIByi33eaXXpNn/Qw5L4K74luXlIZt75JmQin+ZKXzL7SjnCDjC5weeoXEthf8gLr
TeUjjNXJkmcrrRYGE9lFJX8FhZhMv7iJlyKslFzMPdsxCFqC/NzMidzwBxFLqvZVBli++j7H4h1J
B1z7N23H69D5MuHo/0xgOwZM5bG0v/fKrJ1vzrPtMhfKQcpdDhEhq07LEK7JcNEzaok91AhF4hFQ
4JlY25blRcSy1kTvcFDblY/XdWV2ShqRjXzV9vKOaeZR8Aj6/2eLI5BO/QcPJv0NCMPNJhT0C2Wr
eVbGsNKPl3bN5SRJspz8n4wFqIz8kkvHfW5xnB1uerQ8U/ZRO7vGRXfXIdc0lShMSeD0KdXQeqj4
f1MwbSQVPO3rK5pcsA7oic724e7CV82bm59x0o88uKgSVShf5UeVB+FLQrgDWz9k6yxTyolCtlRa
xVYOfSiwvESzcaknGzMM2vm1sRocazAHihek0SX2R9BnJGt8bTAXEWMlp9cjKXevRZ7wXFZKNge5
xnM0lHBtlTIUVLs+i5M4aVeQXB5cZ48HWi/vwbTQPjBbwp3nsyV9KkkxUWHu1Mc6b5vjqRYqrpTL
zaTC027O+oNg7T8w/bbp1RyBdAOBSLDwJmpIk+v3v1dKDSaSdjX3WhqA14kP4LktS5ttud27lpf1
sBC82xW/CM/C6x0YgpK3sLezaDv6UxtrqsMze0SWyYhL90sX8kK5WebGf+4dy6nXGeeVeyeCxSyd
iBg2MOe67ObVGYaxL8IzLlX6KE25GiZaVPulO/KsZ4cDE4keZNpA+OS5/eG/EzBPY2OsNsy0I8qH
wxMZ9s3d7LjOXc2vcrsGxhHqVG9edvGSurPsYWFLQXExEawvGeAnxUutcUhM9htqzZ5OF3J/96ZA
rYhrg2eLyySAikeIvuBWmn6+qDLxZUA8hmDOpJrZZjXm7eFp98NSUNVtP4spZ6H5TBRlvWsG1+Ao
0aZjrOWZY/AobTBv95Ar7AcHlt9S+4MY7uPhc6PmsMtWy6INyFv6A700MHxeUTRHSnALvteMpWZ3
DBCNklj3aaOL2dKBdW2oqA9kfinV/LiOU4hK6vt1xOTWw1wxkDeJlgzEVkoQadkC49HpWj14iRAc
pI+fCCD9x2h1u+4F+hcC6+Ix19oWOdEdoImJ33Zw+WtBy7gXRfTr97dTlKiw7+dm9p40nL4OP7t6
GlsXI+JTGQ6MAhatZsUp3rFphLQofS9CzcU4Bb55yyqONo+mjnmgPBS48jJwfieb4z7H8EVmVqMN
Vw/bbC5wgBtwC38m9NoRxyxeWTCbfXJZhsleNo3sh9nddD/Ft3EHis8+09r94Hn/lxEkOOLQGBgo
ACzWe2vjQIcHWddoSgUxAc/utrlFHP8WoZ4wALPbrXm+A2jriDsDxo/Dtb5BDDBdu15dFgO0Bo4E
T/G7vMb+A1TD+FIiqfZIzTReEX36adHW7cgPZAVjJk/vkhEIJAU01/eBhvSmes9tIFP6ILCFqqV7
btlzSiUSt7EtyOstRtFxvX4zB0prrl7H6fvrsau0C+PF63kF9xG/c+wlAnakpX5jUli97L8aIik6
6NJdJ325BglbhOgQkER1kQBsrHNWhXLb+ZFbuyuy4lRb3dbZFMSQmMbDwHccix40H6BkWAobLpHH
c/owVqKeFiaqRJPCujtLKYnfbzNwiWUfNXw23Bo0XE6IfGdkpALyJklX98wez4e+aB+bn5H3EoI+
OGik7qKy+6CddU9xFh4H9I4TLS9fNogF3cs7o60jllXJBVNoFwV98jsrzWwQCZm1fTaGfRfmbq1E
M/QGIRWNmR+WDHJbbfqAbXOwy7ZZgVgnRzrt4pGaZ4zg8pz65R5Wok4U0oTWfmK2r+mafANON5u+
rJ4x8KF/J/PHHPdXLjKJy6qP9YnK6ck/CIXB9l8tN2+UdMyCazG3g0wkhf7BKirPjPYEm4zwpviC
F59dKVpzsF6A3I4lVqA+t7fxU3aXQCHZR/POi/UGsdDY3kfyDLHs8YMiFphKaE346Cy8BhCguTHt
wSkCKOtdBoFKi+UYwjmGlATstL0ih70ao8nusRy5gIQ/PP4HJQkAqEeuq+niXszjS4Jkpmu+uKl0
iZb6rx3+P4N+xx4+uMBZfl+SlAuC6gPnt1h8MLTSQ6FQLzYt5gZnkFgaqs9fOltjkAwPRwa6BiNQ
O317azRgSHWbZufxXMlQfTkmlbv/wB4da4c84cVpGpcOHC8KMEOhOQcRYCJ+p82X0TyaD8wC/4sz
awFSrKSdVCfVeTwwTwKspNlbB4DSJ8jID9ebOfaXp2n7sU8bm1O4Esi1K1JAUxFRooeJQW+TrNxN
7EvvnPpMtY4IWqXk6jRB5ZRNvUCWMN9IKFk9HZRwGciSvDLgLDbV7rHxFTTS9wnMLMeK2vqvSJY6
ReWDtYvfi1X6cZa+eEUGEo4e2Gf3r17peXUCG8W8ZbW5WUrl5oSzEIPrWP4RzyuEBepy6mZLx6MW
G38499RyuGZPqiXDteJbehMjbYR7m7P48OUkAQh5YgQpCteST1H72jBazt9x2pvEI0pwnHmYc8qz
eqc5KFQjwJQAICXlwAAiEGGqC7QFW2TZhKHbK11oRIwTeQwgBmCL6c1hafQyMF6bIwpkML5NLe8P
/KfvUp2MnvxVIJj6BOC0Zxwt2QstnnaoAw0oTqWtaBt4g3EcNJB0Q4HfbqAa3duF48KlvqvrrNK0
hTgqdWbQyUIo+/4lIhxdlpFPEkdVZzvYdAv7Ar9itlm2+/Qol7dx/+hz45Ubxe3gXJKfAYAnht2/
w2c62UYhfQjL0KEFmTBku+tvVkgQkZMx7E4H4pV+4hTXJ3YMAHkWJp682nOdvcNLPqPqemiali+I
Yc1Twy80J6HufcfuwMajITg1bs7U59FWtkpd5TX1lrxaC0CMaTeaxV+E9T/UViIySD4MRhAGIwHh
VUi/UY5r5qnntRvb/nRlrvfoawjsBB28PUJjnj0BQqw/Xoy3bTfQysBAyQNRPWSWDNch/rg4NJ6e
GHpE5hl9XQh5r207ITF89mKMWeGqBX1ml2Xq8YhQvXpbRP4Xzt5BHJ6BTSzosuc0XnPEUUqI3j64
+TrmoU0cV1mLvqi7LlnDE2U9OtAqDw5RP6Q3OQ5SjuCpOX0zjWSo7CxBR2xV+yll6FgO9sCKj2Tt
3n+YpdZDY+tXSYTaoR56FqQPaJaCWFUW1a2UzawYCGECj9du7U1zq3ov36Z6GIRk4Jggfp3KfrsQ
/qCyPZHP5w12elWnD9PGEF7qfNfLFtT0julS97pfE69G3dACYQ8CtgIgF3tzXRD+fwNqtXkVx4nJ
3/kapQaxm5qRsHgr2eOqJzoHI7Jfps9Gz2ktiSEGhFVRoXTKc5783kuWW+Fk7j++ABel3cqY/4Dy
jB9gVfYyuLYv54ehB2J3hqspk9Cv4cwZ+BtX7Vu1g+ky2O4zfGmn9wAtG75iDsqHcciaig9ecriR
ptgUn3ZUzJkmlkqF4pSZVEeNTmHURmGi4ylbE0DeyJ90QhkbPbNepaayO4Yh4cH6+wFRfG92g2s/
OOgn1LCTXRy4L/CmG8CLGTVOoZBbPAltwd7eezlFYXtyPyWh3J3mXeYOzuyTFesyyUoqK1b4sMfe
onZZfYuJGt+ILb7xl2QEq0s386kQ+zowukk249Fir0uQNcafCcPKPZsZN8mjbQEZ+fpDeeQ9hAwg
wfjil2OnwSB2iiFMd6+I2eXGHFHIb8UGJYGclMqkQTQLywbCKGkeZS54Zol+AcjnzVqN3NgLB8qs
sXScZamTsrfl5d0XbdWkKTMENhzvIzO84Ea1oxIUV6UfP0xOLrMqkMQmBo92AnluEtd9tNEw4wk5
fMvDqiYvnH9cok159zWQ+UZNfWzLBMXu1KrQkGw9B0dKpBGn2SdcRVMX/pdPEV4W5tzr0pU0XC8Z
qKNWyOIIxH2PNzxci6s+fBMnSWTSlbpzua2fPKqLyE8pxPuGfsm90Nz+6ienXHLnpi5cd2CK9qlP
JvKngB7aR23Wyuqvg1Ldv4mMK+fxBQSwJN56U/L36RsFWhC5GsO6CBLD5llXA007TP7+VQzKI6vN
YJCi6fbbU1RbuZlD99b9WFVS8rdMKdKtSBU39BAiBPZSoE/iPB2IGzo7QNgTxDMn/+YLTn8YV0M/
AE3Z0fwiC5/EqpfKPYBFwL7K0Po5DQmrqZSc/qg/DtzhJQ01Tn7+bkJ6ffzPuBp5sXVdMRR8vZ10
cxKfjqrZHShPZl+8xbgIypc3YLV9p6bIGOGiXHY0DXVEc57Zm/24zqFoEA6y05lTZ1ydc2OiWY6n
oq2rz/2Y7IyLscW18hNMW305i4XbWwfiO6JrhyNq6b7ayAXNKMEmiKQETt8LFC3dggjUTLCN+FjG
ymhQUGNvrde9mTiFcpthBCbLkUMYslr+e/qtx8wuCDJ3719UxNQhXNN3ayWe14Y4CvBoQIQ3if4W
kwZCAnDBNqaIf76Lwif/RXfWDMAZC2W1w4sceEVDOQXgmCm3jvAKcY09cuvvROhSy1JFvWrublno
MrFI81cKwp6cgsuZQ8tlFVax09unudwu5CzQBM7zLoe0Ejmd90chjDj+7VWHWDFa5TCXVQ1hBHmv
vPaRNkKQL5xGLnHaSqjFM09xEWrVBRSIzGloLoDw1nwcHrft2efTzvoXTPzuWseWSaKLWtMTQxYH
Q4Q1etkTHlllf5YquruZQCO97Mm6iCTLXjwQMwl6R1VB0ZTF+ezOASD/JYuQ33oZW0v87j/jRyv3
4ZY3txPhsLyfVlHqg5SY20mkdJJ1hLzhAPoYNB8TUBflaYJCQVXDxybypS6CKmYs0KfaAOfvii0f
pPVRO6PfHkBGHFjb1rTpOz92jTv7c8E21LyV1aD8r1SsRAdMj4iTP9gUei4VTLDhcdzUlIDYu7g9
tK/H42jf0Ra2P9un5H+LqiOZBeg0NJuZ0lPILsX93sgjJq/EiMsW3SrdpNjeRuvL/4OiYRfhrb8V
cCBAUTR2cTxXg+bDu78xY7VRWBtmCw8da/JTMT/e7fnpdwXH8Il4Odt4PrYt0oCk79f1QXnOzbSZ
9uuTHwMI1ZlLAhH1imEDL+2PFcTxp2JLuf6bMTFZbzfDA3/5OACw72CRNaUmNsrB3+bLqdvwfEwy
bV/gd5J5CeWBdnJNBp2JmjT1SL0lT/LbK6KfJQIRtbNBhKKlw3uJcV6lU3/X35AoMBebErXgM6SJ
IsLBbXpnO2uRc4OrRWs5XWDA7PY7Mk9X9RQ0jqcPx9xh43U4jYREBJwd9Bkx4S1xcgzaIquR0Yl/
tCnj1R7NPkhH27H+wAJXWn12NbK8HSEqRQChnh1DrK2tCDJ677J45qeLnz0i7JH1iKoQNpJq9DZl
Fk+FHMrGum01iIRpPvi5BqlbDaAZfawbHaFubYH/mOUHtGy0tIq8GzcOlYrGNQaDejzfqrTnfVgP
JfjmmmL8YPMO/XqBwJ3C4UwY9ez7llF4w8XJLAaB2flYujqYVDdGHj7KFZ8yvGix9cteGnKxRQud
UXHKrxNamy6PZF+DPIDoON5UkB4ECL5GCIQMKR2oFWMdQQKjitPVqqyk+x1RE8ai3HpNgRkEU2LY
RaJEYJbzOuCe4aQRj68D3chG8FK+xCEuutmA43WhJkOazh4k3DUeGE1qOwV5gBqie2eixMWuz7/s
K7mZj+47XdLnAyBaelfCEfBvTR5mujBVm/rOWeEhyM7JGs06Xfht8uxm0T98DhoUgtziYD8IrzoZ
P/5zZE+uO0Ulag+ECmjvcn6BLdDREVJKGNL6SrTAgIKYNE7A2BbpGcEUgj2wSFbaY9nF4IGoKMJ0
XItXhHF9jmlLKxvDZaO86a6NG+ovGwqv+jNva89+dkyExn4LUmRBPdUBKSIBuMqIK/u8K9TW2Myp
xRIry3ivxrLYozhThcYazQVSCF+EusTjv9tE7UYMHna534vFahbTpsTg3eGZFjgTdnUFGT4Z+JgK
x+vh/INFAatTMcFp5zt+hKRKJ6s1d40SFAljqnZanhyFvvZFuxrTLproOqMwmK+XSTQiWPziyqir
/v9pUJ6YzM3hL6awlSXZMLmZd+ogiIAfbKO44kv28hFIQdsQxItZWcJG9zLicMg10Ha92KQo9eJw
ub17ep3rtPxmI3N687mmYRNGPChRlpFIDBgbY2QEM8dnfmkFQCB469h1vdzNgUkdFJ0pqjiu9gnq
OLYs/5+9+ureftPVTXLM8eg/Pr/idhBCLJ+bVJ0PDXRwvYSdBnEmEND5FSLj5zlQOu+Fee9tsE1B
oLNpJcI8tw9UpIrJF3BygzoEIytPftJiaEMKj/PbjGutiBuNbguSRFX0s7fCPaa67tN9B2Ud0rdY
Jq/xzQcl1hXVGLiY8pqSi0BsGLlOvJchBj+x5cICDZ6GKYkdw0tQ1Vz4tQ7Hk4eCRoNhezH5Qzik
3ObZArhXBC+bX2eVYQFNSdVxWbj1o8SBSOFE8hjZiJS/Yf8s2oW3m/UBXgjkNkg7Cnz7n1J8pnsO
HqpEZZQuvC6GsAgKULs0ZH7ZJfeVoDwffrsBABiyvNAVYAxAOOaNPVIKhzMG886Mz7fvOjpWs6GG
SOeU3BJDBTxBFKNE+U3jKEci/kk+wg6Mp6E21fu82RDodvL8ZFpIepFycr0PE0McdeDpjQQhmsq3
ZwOV+FdxdVnY6Vb6VrVT3+umkb4G9OYzoTGN343bArOcNjrXrY3xEqUoPxSCYyUg0r/HNOw0mMbY
tAOmjE7RlNRSO6UTcuxidGMbVuBKEzVj1a/FMe8EywVx0gIDDfnRC2zQ+SzL3oiuUh/ca1jCkMzr
N8kIe7BexE6PdtZztYZmcfCaQsT5INEtxujkVXChFZWiD7ld34tFGT4rcsgYjl/pMYW/n2mHjxMF
9nS2ZhAxxFh4ojbFjCLV8qBQ0ZxFsUcfW7GC9AOS3vvW0XaoT+eh6V4MEmF+QOlZddHXvIBOiKnE
Wag1/xi7qSWJtWbRKzF5vFMQUV/FvVvURjRZu0z1S8rv+D7PQ79wR11maakaq9o3yMOApXRwqY3T
jiFr8O7E6+AZIuftR4djZc4nouB6CFSG1TaXwuYwWr4t8w3daBwDZKM8Gvj9IZ9fWcKHzx6yp8ul
+NrnlpuhvDQT8U89JWcr4zEhhq1PY4l3Gc6yalhl1jqIz69vQxMPXjGBttaXDnBa7KZRjXnt7X9M
KqcunM5F0S23VWzJf1BOVrAqB92ITjjKGji8pMjn+6UsPl+9tKQ8WVLrSzigIDZKmC5rVJSfQQW9
xgqqcrYKLtoQwaY0fjINpDOJUeUn1TMGtkdHbGJYCEeZuk+1PPXV0r2WuYWZap2EnZFVnC/ctyJY
FXKYD9TAt/sUr8qJJ7wMSIaOQ/FxaJqSSVjzI279kAiVysZEm/Gn2qO9BUFiV6uraiR8A6pY5rm1
VWv8ndTKW6ja6NbKuFKgwPEFICIVkP0/YRp9CdSV6FEZ7AsK1HyvdoEwMl7sGcPLmhglHowiLrJp
PLnSbigQqhJtvkzyCTQjEhLqtKfsMc/JY79jaP3HbWDeajqSObOkF9Atvx9XwJRChgrFXATKICO7
CTSn6zIY2lLAOjsTneD7G1ggeuceqSop5KQNAv4wML9TYkJmeXFXVRuwcHCgnl446p5Zs2+HcJ48
KKdk2pPf4y3EZxjSQZNgRbouY+FEGkEJD3BwYnVFFffTp6ed1WNxYKYbkE7jrzVIHc01OP6qG4OJ
Jrri2aHyTqGhU0y/77nnSiZ33O75zOSe3OOe8JAXPd0sUuzAiA2TNZs0UEx/rwHoDg8ShFT0SUKH
K2Y760iYxPOxRFf06jKhEakJRKaw8sh5dLNnCQd8DsQkJ7TTcY4J72OlzMTEF/EoqP2BAytugOjZ
fcjhX+oFMLoXCOlGtD50pbmuiDFLf63wXR9CUsjY5xQ700pA7h2rEPLxRbL+jqM8xPawa4BS+mJt
lGHvho0jRnk7O2emws+kfSQla2wW9x7WLnYs5Zx8HRDIQpByGlgOo/NgZ+XlQgkfOATre92F+ZgF
QaYOSNRAIQWSRBkTBH+sy3J8RQ9Jfku1jHgL+UxPVBzqgW6IWVx5ivkyQIeNkHOJTH6nU9PmH0nA
N+z6QV4WWe+czbWlYMj3ql28jqwJDTFhmkGnT+c6NtA41Pxlp0l3PrOEl3J1hbhSkNOSDJMG+XZF
X36XaShd9P2xPQ0mZRJSZgi5Ut9mT5/sF5F69tVxIwo/aT29sY+Uc+zUndPYkUX8SzBxpqlP/z4E
AkIP5EvVMUwCFFZRY5mPuK9iOwvgOZBSAoyNZVJIfVN7Ik0iO9ZOJegmHi2sYaPPm6Ez6I633HSm
uE2Jsu+RpMntfkixC7w/OzbJ7vG/44qaenwlFi4oWQ5qeyPkAacVwEE1Me8pmxHw93VkBkNjxOO5
jLZmM8P9tojIlntJ2Vgh3jTMTOqBZxVlL+/eB6TpdUEsxcl4AAplYtfeWYgRwmqsc3HgWzMHgyib
JQP5H39tVhehRenoGmQoMUM2FB4zp1NIwuPmQuULDmPpnIBV52cgsfEJjmQu9ljgz6GySaIgH40s
XXmpdr6hmMrpYds6GLoppX5hczyqrGFCpdZaHl0NAaDn6hqAjAQ2rLkGQkr/vgU4RHv135zj0Occ
PwTcBzyWXNTmrSucQ7mbk5EebU4XT6kSd15ryvqZuHQBxYmHKIGfZigbjW3lfEiZkYT32RS2AgrS
k3iOfxFgys3WQsZBtWsFzOlpsCQSKcZ5Go5WRcCL09IZi3R10IrK9dVq2CGp5ZewmMg7QaTxkhDf
MEbbzmG8l7g2zMGhv5yB9ZNytlgiZHUg+eKxkmPQZy+y08V35Sa7yN1D0u5cO/3BD2hYFoioQLDm
S8RUvhHWGE1OD/z6ByBLXEJcmIn9oBW1khCZGuMqm9toZESQAb44uVZ8IzSNdFRsZ2O9fXg6EbB5
c51MyHfCS9yucYlxbJu3aJ1A3qmjS6s8eStRW7HPXRnCKr5oDQ3LY3to7VCEC0yHK2O63c0ugyNq
d5l/CUdKInQiCe7SaPhcxfzWEKOWCztsAKvTc1Xa0agMN0b+NqoaDLXigbUtvj6eywAbcTwZ34Xs
Zbkkbqz17hTZLeJ4famT76X9AnR4i//diBE3iSpZ/+1sB6lRqnwbP2TfmbCfLUd83E2I7T5Ttbou
tr5JjYaAP+nkk/ySgK99NbjEKQrk0dakyRepGrcAuzq3q2MAeh8F+Hpwly+R/O8s34k2RfcNF6rj
lFVjrED2lL2duKCDbBICqM4v7/KLyxhJJGbTO3HH8FwELXztvaCS1kQxagjabtgidK8px2YwXkWx
x3u1bgMdPWGVXT62xX6T8TdMp8R842eJzHfZ9irmP6YzPko1loYv20gFg9CbeD+gD0NPHCHyCnGO
RDIHx83yMAyHSkub4yTY68S5EMYj6hShMIeRLbXx6cpnQ1Z54Ug8SH6M03bCMp6dQLliaez2cGIq
FlUoQaTnV6AeksVHQgz6fh93hiRHJaEfZIWg3yUXGXJDdH2181tcZjf7Cg9RX+sozho2ikw4u+Cp
1DQX/AF44vq07imXUzxjhybkTZxgKIT6Z4Gm40iEmT4RjZ4etYLxEMM6f2E9nwaxB8i2l0CCfTuc
iOi6AD8yWXugQYGt1un8s9BR29z4JqcPZzFphhaIuvEAwmy77ZzMDEiui0QfrxH+4wppF/zkyL1h
GVLuFeT/a4LeRkUz1MR2B4YebkPClPTaXAU5VbE7kyYVaVc/seeK1diOl3bcQIdzHvfPzUaHo0Bd
JiF8XX2xE0OoT8CwpSgzOvzD1J7GcujQHYkvHBTFPlAogO+Op5i+a9/wK1Wr+5tGanLMSH03FjMy
z7EwsF8CoYsyrLpUtFk+9VgoWBQuW522Yds98GmA9OlART8e2obz73+2EQD6Mtf/0G0aMeCdnFZF
PaWUOU3Hro9FweFq4LxFLDn5yeEPvxNhM6B3ySyLsD897N86SlGMpwkg+RDzhEjDaVDxKg9eOIj3
ujdIaILdDM9jAeqmVOkPCeGXNG4//7W/bJ886IvnVOGd2Ue3XY5Q+rCm4/AZAgUMMySLRI2ilFL9
Hp2wZcoY3WeHCUP4yg0qtrOKZVVvDjAYLbfaHUsJCHISNE4jJeK1V35GdxAXmKo9r1ZIN4tuOf3B
Z+M3q2p+K9QiJ5FyMFbtg/KtPyyxrPmJt+nVQ57Wdh1082CHNar0ajWwAVjND5hO57HkLBy2bOZd
aS/r5Nr+wOau9uP3idGV3ksW07k6oeTk0q0omWZ+oF35YB3Ay0CcBUN360a0PPS1k+CoZyxlSWNm
iq3gXVNBja3abN423XVsMyja+xMEUk0cT1YaHxJfkd8LxNmIcvFnrFFg1cK2JDGoy4m1M1BKCx38
RwIZpZ3pRb7afxaX834vCR89katoiLhC9686lSmjLw09tGInUCtfK2UXtdGaw/SrfIB/JezcLCOG
Gke3PC4SNWioJ6VHRPzaq0ufgTtOomcFtfr6n+3A0t/CARJi04pZhDqgzc2cALG/VP7kqtvMBLPY
2xHYAHOyS1UhP7TUYzBCZb3DPF5kVMixqVGma6sw0BonnsMwzIPiih1/BSYnCVN2TgMUCEJsiffO
6V0yC+d7LtpM9NaVbf0g2Z0lPydjLTYMebZ2tRoAHuKPkbXin9DlFbRuMx73vYL2SnPUgGjgUFHS
f0IPttYFw66jElFMQ+mt7mqPnRV+4FghzLgbzckikIHdIxLJ8YQSY3LlYiT/ANMHKWPDwz9okhUd
4kPQVN1tFk18emYwDr0BhXuBeJag2xgCSU1NvrJr/+ErGz+DZNo1ZdAMmFWC6RrB3FZlStk/XhRe
QMMkf/bcmVBcb9TAa5s/c83tS93RGgT0MHa73+LB90dk+3PJP5sxB/nHjxWomxgE8ojEnngkTS7/
ZsJhNzEVtv2o4CUmPVkyfAd98tz6bhJ9DJabDRbGD2WzAqq5z8v8AR7aTHcWtoyvr2T1ux8OHZ7C
1U+Kqo95KDMP+c68lpdSwfbyYr5NUtuc4AjXITLpWX3XkM+Cu6xag8YcLqOdBtbDRXx5DYi8oT2h
FX3mbN3MU4Gqdt28I/ObJlvt+GHulAm6PVY532zWGkKhljgbL6TtF42Lprh65i+PWghyOtBl2YM2
WvbpmJax9VzpODVAbRf7fRCTQrhQHWXcXSGumQKW2GK2znLfuVr9LPPdZKXj5WAZVL2ly+TWnvBp
ySRBJAw+N314DHbRa6nFYcmyLdlKSCroLrf2fH5l+lmt9fgsB3S4+rTRajLRzSvp7qLSO1Ctzxmx
5kGiL0IsIeGMWQMgBdymyX1XsC64tq/msFCfsGHnq17UdsAV1ZBe93PpwvX6auHT9sk0bvZvwVvY
CUbgLm2Bn/vqGiVldnag5AI9/7omt6VYk4OMYPvVb7CIt1gFxX9FQu/lQNF5NgeRivDNpkorq/Pe
fb2n3vEl/46MaGNckPjHeUBzHtALJcpfxytSNlxGzxLbmAxX5rJNRYl7asY1eI4pZMCrb3UA7TCo
mK2+Z7HQzL30FT1SsmiqGG4uTymKhhDSe89am2w6aiM/yx8HWzHDyKfsl3DtNu0OobAEZ+vkmAb1
qbmAQKpuCfLMLtWb/DtXYZx+fkYH+/XG57AAD1N/5dQf9uMgpu2V2he58rbmfed2HqLpvDF9X9f/
9PO8sLmq5MiDJ57ajQ95Oba0QgxPV9oMN782IAkW/DK7xFvyg7CAFZR5RA/V8Gqo65CmVfW1rj9F
cNPGwri9Xn3nanqE9Cf/ZkPSz6wIVVynX2WE9kvG2rJXGjFiy/l69kWBFcEK9fbvRCyAhB1S+69X
pOd592o51GVv1EpnsXKiQyb2GRymYKT0DkO/ovOQ142qCB8c589shTnzcqExYZj2V64+iMwjK3uJ
VMo1ZG6THeJDvuBarGCkAOup4ynCZGWOrgZR71EsMW3ha/JcW32HLbXITPU53U/IEqmd6vlXLkjw
nUeLQ6bYSIvV6i4f6pomhHqxXimC2FQKS5jSCK7S5wOmytI3rRkKDjVu0kN2qhaQ5qw3zQY2zhGe
AMO+k0r/NssIiLyicO69asbQtwqx8LCnOHx83tO6rc/vim39YHK3hXNDTkNW1BYbNM2wULPcMDcO
S/tTJQ65zjEP6D0qIvSm0J1xhgj/HIajfpk4mzOX5JLiQ5pPLWheZHB6Gd78HxRso2olfjAIagWN
VeYXR9qgUMWwNmAI+MnTIryIbJCm59vuENQ0n7ZqyhvGmkq9vzC++DHKokCsezaYsURHpVs7gTYA
roaQRbl+TynFNgsb10vmgnAlJbU29jWtH2YH6xPBLBjbToK1C51aBDlRY9msp7wY0n5okAo+vy6Y
franLaNrDCAx+mDOfUe/ZAfTjS9WV3242O5ZEgo7nDlqj78T04DuMqyoEl3AVOm1JsuXFekmVVde
KKEQGcBonUvYxetiU6BlUVbWU23CcagbjyeuuIwx8c75QeFk7717RdFg6qt5syrGxkl0maB7z9zk
AsSroQ31D3KqnYCwux6iegbpQ9x5QC5GkotOfb+84p0LG+MyXK85mnrG2METjj2CfJ/WBR1DovRC
KfjOFmpDo+i30Vao7OQmRFSCGPjcNL0iGUJYhWEBUB+ZKP/2ZmmitSCHEkDQUb/eleidGXIrjSXs
qn1KUhSQ8/iXuVnQ0NDe5LNfOs0WPRVX4Abcndc3m7wUJ1mSYdhTulT+90V79yqioytgv2U1EdSn
kl7ILZJyqfZS9+ENeZt6MZqoXUw2qERwcEJMIFJsJXsLNsNHXLHjs5tLk4oY301xMzZSq000nXL7
kPzxXs8LpPiEJNxkOWR5wOCtSYeSWjIbDTPByPABdXBikr3p0QVQjcAl6OEAGUS0SutMwfNF295/
AvW/pNbEcN3gWGAiHpNB2O95JkHhdSIsqAwOFco2lAavpaRIZ5xBnrF1k5Ga5RV9XJA8bSlxAfzG
vmkR3MUqmK3znlOWNA5jLDoC6lp6eaXgRwiT8V8leQymFoz+q43zIRBnPdqGD55hE7YrKZykr8np
t9VnBvio43zz2WJNIbDQ5s6n/Rga0ha15hLmVDlBB2g/vXNfPqsXSSFLxgx0DYwcqnimvDaj1ioO
8NrbTtsIBqOkU5qpiHBffpNHSEVm5g6v0l3CFwCwazsrFvu0/t64gPEIuyBaNItproy2CnBZPy0K
zinTQjO4f/1OnSdr5HN1a3thqnVRxXEvzTDJAJaGe12xZ3HbqNY6UfF5aD+HZTC47vZymkAjOBqP
R+P0+TS+oQU/KKsVyKYttP6W3GOYrIhp5ovkhA1rrGJ33hKn2/66IdArsWRZKIrD2qsrdx3UHto/
jp6tCAMZfBzbCzYAsyjFGDyEbSUnKleA0HQD/dw/P+A4EYbFZF2NDsI8eQqeBKSZgFJNp7BCg/Lt
AwTC0v7nd7D80U4h3eN3epBTadwYGwfhsgzzbnv+l7hmnkUM1tx/wx2QeaNaMRBz64u9PKTZJdME
kt/VCYAQChsBVS/1OVeQe+VcahqM1umpNXPB5ErgJ9ZbmWTYgiZdQSnug6ZD9JKB4tlkAFsmsla2
CNlP+hPl5ClTc83dE82KLaPDJbc3yll09RV9F+YkysJxrs8iv0yxiA48/b2D/CmVcMF03sUu3fPe
K35dO2x6ZOWDYckAXj5huwYXQxbnP1A5w4jjknImwbZmeOxG3zvjO1ZDWpZ8+zISF1mSRI5pg33d
f8/UrfUSh0GBdB2grsk0MaC1bxun3eiMGx1xGJQdYusbVfz/6dLdPfYiUHiddduePDFK8Qxw9Vym
jIFFukhdqtWzEcX2d3zovTR8uA6XCCbOJtAwl9a7Bb4lCwJJ6USImfv/eoVhyl2hijyGslQcMa42
yrN9JSnqQiUcYrldV9CdXpHhvXoMnP+je2OI6G5QXuHEZ7vNtBi8qIhI/64KnfHrWzPPH35dP5bh
jtjS44nkTyAPs3KCmSx/oLt7I2dqQNOjDD0tAmNscETZNJtjTOtqmH1sLGiTnw+P8cSxU4nfgBTx
ctnNtLYkgjIBKe6jsoS6bmdhqTZzIctCxpNc1r0mSrxDbl/WPTgrpFBKiwt5xvwdpFCRV4JkjvZl
oYaLtI5dRx4WKmcWRS9q727wY7PBMpOGlkMMzMJAsgRujiWrHb6zSHkwgKjRAUArihrFpMx+m3NM
QwbpIEfISxkoM1F3VxKeaiikP216HP3FWMFXxSiOjLwXFXcH1KQitgdEbyjo6jKPxdyk5Ly7w7Ez
SS/8p963pHpR8OC9z2H+zjx02FarvhXPbtXmCbziMC9Wp8DhMQ5aBFggk0paM8d4FX7vC1lQ5dPQ
sm1pCwUPKjpwtLuBl6K7Ncjjz492uJM3jslcdc8tVqZCy+8aeZQIQNRm7p+63+113hUFJfn+WFeV
qvHK63xYGvBIfd1pTrzeZrKJyQXbMRtMzndF9KQHFvpyrE61Ay+y2SEEmqYENXrMn8+e9dT0lXNX
FiAypwsjR8YC6ulsIXGVn8id14nYXYfwcMrnf0PASje7cX8SpD3IVmsDm1u94JV4e9sp9RAlNhuE
BPnIJu6C9ekwhNIJQgE5CMabQ5ZjBtYLi6RPzFzWRcSNPiVhj/h4pKy6ecQaLezOo7fAe0qVWCwb
JVndvxS/npV7bJQ589sBSO+ivGFx80iNG/8veoKBWGmUt52JD7wZWPkJSgSdsDeCQbTeSRaIm2W5
iG4xpuzM7oNe8ap+G83xmH6K5AQNypBEvmAgC3vRNLWHUX9XL/fLugKqA8CzGGPe6t+PzhzvmM5E
O0BPEVqDfgnw4OYmy/ZorJ20yYFJ26Unbyj/ecLMGxs2hVNSbe4rJJ56RkRowxYjf79vWFFDdt+r
w6dA+lU2avOyOC0j8v/Cj+K9IV1/GPjinVE2ZEu3M1NTN4V3a1JNip5zPNh/xeOO9zqryVWP77xt
moWEfTXB1izBGgPSz1c6iCY52hBDzdgT1wJzDXCvUien68GSsY2ck4UvslJvQ+eDbay8BYtTr7QT
psI/IaGOAw6Ue02lOPXZSdUIYCB57ceTII+vnLep40y9DfM+NLfOL37lZd6FBx+jyFidZUEc9W+a
ozG8KBmJYfxDOgyPcDgYZyeTTkQv2b6JE7uxi7QuRRZ0AC4HXSkvBAF0A0hZJGKctErk6luEpOZc
Mo6nKtEitllarPMPwiaibJbAkv8lPTgYtDnqCuyR2GueYQp7db3wC94LukCBZUExNUEhrMXDpVf6
6j7nlq/fUk1t1ompLrYvHoo6pnLg0nr25HNyvFuGqiJY2Z7+nRUnKFJujVac9cIbSrU9oGCzdvnh
GtDv3VymCPZ7qu4IrdDde7dZM05XIuEhoDBETBJ8dSHAMCYlSEpXTYE0+W40XsIAxprVbcIVyD3z
UMhP4gaRbeNwm2b8Y9VOjTFaoxr/6isOIx0/h4UBcKabVe/Kq5/hY9U0D9QXD9Ij0H5H/vAc5Hv3
xdYmg0/6V/W/VbMyRnaEsjJIOkHWAa6dtRN8MVpVm0NRBzzyGNnp+H2If2zpipNZtJoSYfKwnvX9
FxtyZasliYZx8PZeooacZ69CSfI8gk9cee6Bj4fUiX2w1JETNXksp0RZcSMIIBI7sV2UcvcO/jou
BkIEZSFovC3v0uU0E5JTTlfZgD7nou6u4PmMq9wY/MMZzPmtbLvJKYAXQRwkCDslFLNyAOrdzrI7
kVBeSdvzzlB9ikPQh/hp8ycY+Jm0Nawr5P7c6YRd8Y+OQMFj4yJ/RmuAN+8TATxBkW+OnA55k55V
BjSSUNsng8lYK8M+F0IcyS5msaRoUbLugj3z+DOEKhA/7slno7RMSzOQSVBS/k3Sk9ADUZnOOAqx
qHaOKszoKWZq1KwSD+mMLWH0Jah4/LJi/ThuxiIHBNvvpi+sG2td8DSLIwDrGa5hZ0ATS0t+FugX
1RrBOAHvSowoPHEazJjQIkOCocbbA/maUPZ47j5GIFO9hKWK0eWFFVkcAjbYUZx3RDXFWBb/+B+3
w+1CwJxqCa2XwX5A5z3mym+SLX+wxZHUh7dgl5KoSTa3xnMhUmQxzUvDIDl6aLpQMXr+lycQS/+J
Q2pOgI/pOTGmdIPmwyj0fh3a+iFMuBkj3Gkp2yVa4OqEy+uBuXKC1VnmiUMJRFpMSLDoihFG0S8W
ffss5lba0zpsUoVbXf7HWZL6eYr1VozD6uUZHVH8ldMeAYnj1XX1kHprvJUAivNfLRXHLcwMi35B
6ERevaOFAlsNWAdXSF5zXPRmol6Zp5quIX/MAGluum7OWZ4RE6kyqQ1sxUqLejQqxBDQQkbeL6DU
g6syp96iqLIoNaCixZ3qc5+6bVZejSai5uQxQbd305+bidrhqK33E24vFxdv1LKceDu0Fu0nk7os
wncG5jHkitdvHHXHugFscSZXhlta8q+WyYGg9xKJeT6RmNG8N0vIq9DlHXQTVUyYAJL2PyM4O7TS
4BkfEwPKyWKZi6iJCVBUZoYp7cqMU/LAXHulSDwVO2SuJRmvDvZjgToV/4MpT3GInc0ZmKNNxn9a
cr4GDusQ+x4sufqqJoFBRbkjW3fj9AM8v2EFIQOZBiN4D8Pm6+MlvE25Si+JdFC9PzrZReJKmWrN
paDVWKh5/QNKiGaP4EY7nnIYlXs37yurMziTHmQ7l0YsdChYpBNneM09Mj1XXb5yS91rSCQ6N3pC
gZeORhIPtd95pPF2VHJNRUxRmMAcrQ1oACu8icUQSxIVOrEnmhMvEMGvTW0rGc9x8G4T/GbCzae3
6raRJe/VblGrHSaBKnKJhdDYxcvjuqpVMyEdAYAajeYMsBo3nw4dbJKDVgCxkPvGYmtefPHzxpF7
zfRAkBJZVvRf+wawOGr9XWuTMSxxL+g5g2clSILcNJwX1136qKxydTRCQFqiKctCW4pRm7uxY1Go
N+ZQk2vYlZk9XacHvABUhCRmaWipCDEjLhnMyeaiarxwnshHnLFd6nd3uLsyTSR0evbHxQbUFhjb
tSuq+Q8dPTwJ7d/ZiGsB9PmEn9GX/pB38OzcHnV0Dd8M6lYJKl93l3aDU5gK6ZOQcRrnKlYVdFTn
GCD4gqy+Sh87S22qj/zPi7WNRxvH+Gc8yZtcQP6/X/7aI1BXplXCBD/1KVYhQPOXG34FSRJETnA2
45jQCcXQofyNTN7BcfDlA5HmeEiKDheYtD927y/BW+Biz3TIFPj4ySLipE5aMeH7kAX11NVsnJre
0ZIf+NzMUppWC5MrZEHGKHBIFbE2K6Dw5kcjGsv1UvyT8+sB0kWVUTnnXtYuQkRf5cSZeu26f2xr
K5j7EeR7GlNFoZ7pRpdmkxlO/QYriMlTdTvn3BYvAIh3Fj+W+jHGHe30yFLB5vIVUHXL3lt2RKn0
VWeBmt9kRhwplwCbqOmc6Ha19RIII1gzuoQKUhAIZp9hvUue1+ehcb7nXhld37Y0UwgZXpOzxIRo
uBi9w3Yh4Y2BMTETAZeOblTAygIRFVZo4bUluVXK014v3lvWewtRXsPDfYHi4t8B4c3fwy3hwRgJ
4vfX8iw2POtJeLPCc/whbpeGDUi2v+dTzulckjTW6JKjNIH2XpKvYdbbwseVYpCh6f8sutnL7bj5
hYb6d/uG8wuH1y+zltRz0I9gasohFKtZQa52mQY8nwi7UuJuT+ROq/HJ+sg7HCxf4nthofYptVNF
hhZ7QWuNIDLUSy5rxX2b9HScLhtlstqELW6DCy1+hrX+jG4oBsx+3dEGx8N1Tnp+UjHIyCmzvr6W
MRyevJPEokMplwVG0Ly+11eLje98st4pzOOgF6AkeynrrtUCtxVtSirQ6z7mGKaJOXxQzF7LXgVP
08Tlw4spndButWFbT7RfCXO0bscm6YGtdm5E3uBnSLPfyhS+1PsrpiykS8GoL2FMb2TB3VBdkF/V
iWmnOjzVCIkYoJo7pxegPnXrt0sr+apFYt8uNaaQfnyBzuN2YouLF0+bwzAy5GNvGVrknx7zGCRD
nEYkooUO+8qHwOLhQksZmu7JcyAlLchaamr1uiUMFKyw/zQJWT6CMTH0k1TDG+uJJVg1+jvDNjQy
sHUVhhNk88p6ZwSGeQslmpWg3+FpWboW1fpGmxAyU+JGoH0V7uv4fpV/rxDSqk34rLKhBqrSKj57
4IWIZi7XX6tOi0Jsyrwuv+5XwjFYISdBnuL7V0vmlDEsauFDA6NEGiqZVBO/36titxSHpGsRdBUN
0py6JZTC7Urzkl2G4ckC0V3/W30CYCzK/6Hm4oolDOsRX4T+8OlSkArOjfFbrxs1+dzawQrAcR/W
c1DVE3/PI23vXvvFRMhadzF2LLRLuAEnYZqOFM7C/39J2vUiw0qW1vl4uF0wIQz+BqPmccLqwSe6
tCIMdrAfDVpTsff6Ci82LMCAUmuZwxy2JSLfZNducSpD2KmazU4tjmjEUWiybKiBbTgj1lMG71Zj
Npv1z/m/xGhOKoMqus8I6q0vZalYAYNZGethNC0OxG7av4id4lCLY+iI5QPVoiBT0StUqF5XvODK
OsLInUfobxFoF8reKxVUORLIEkWAih+QllRya25Tbc+2h6SdowreanSo+eOIOVsiSSsd594xgq3m
+Kpfu0DgDnIrdmt5auYgH7bGKMQL4LtaKvZSvQACT+VKKKKIS9PJQYxz5zAMYjYF6tb6N77f//Aj
+/pIX1aM8gjELFPmS65DPEZU8Ah1Ni/udhg6a6IHzj8hRKKs7VQqmb/Z2NqznwISzaGK1aSJWcK6
NTfUvuQ9bDkm/xE+/D+hoLF1toHeYXyQAbd3dONmZEUkCp6IJgCGaxk49UYgvqGmkmGhxd2z7T8R
LHOnqcslV4PYJN1eHmwi1KY09v/YR6vuWmVqUDbJZ+91HTfq5BG4PH6QzhMVuPoCskCb1PTMavs3
6ULukuiDuuxUVgo6mvuHrAKuYUy99CHvbwX2WPQYhPSYmtXNgUHAMuGnmA6ZoQFxNEYKcbK6jkVZ
keUq8Xl8o8v9XGWRsFsrxOQLRnemW12/YwkK+mmeBjlWln0DKWg23FORTBGSiAs0ZK0A/xOpru1H
ufGE1K9i2DcotNUPvMZLHPSiLUm8t+Jd2sULzr9rd2IUEzNhWrhzDeISwHMck96sNTXFQ8hVMqMN
4aiqa6zHIg+5KP+xjgNyce5NrsvkbiWbMe9ye1IgKvUY3IPgAEtDf6I+MmxAwWJt7yj20L+87rvY
KPvkgYCf7aHQ4ZtnzP0Su3/x3x7MafB/dqIEpdFDYLV/tGenwMUscNdFdQpBrv87+6gw7CFnPM6G
ZS12AAI3hBGqd3q2OT7L/wKeKdN1l501hbXeOpXVu2AOq4jCg74G0rVXFst/+PNREwc55FaoLwVs
95a50VlIC28NNoOHmP4nP7NzUWnm8mQ/3XwpItQpVITbbFi95Rqg+4Ge2AhbjivgUYmSPyUQybxs
oGaok4r/GyAtN6oM6ThCFBq6qy/36ZfOvGQHyZh6myRb7NeGfTrHcPiPt57lhQU1lw3lqhmSCzf3
OUOtBRSmfbuLvNVjwmVqHFcOxE2NMHgePPVqpew5mg8sPthI7yt8LVYVSL8ApnMkbSGQlow6hQkZ
T/7O9rAUGbBC3fazmX43nSYKYvAY15NCU5IcHPU3WbL9VHCAG8ZTeeUuNsdTUMXhsZpVzHwA+rR7
YPLbIl3BBeFQlnn8sDU+5oBR2skScMKiu6zMvfk4mJxAgX1viX/zpN8JUVASl2allsM27OKhi4Dx
slT9fO9+ZN9+0HaPs6RGhpVosovCJwPGzIZ2cNVo8MXJA+d33E+baGCeXxayhB8ojMYSGb3EkwvL
GQsLRWtkxyeNNUsKUwWX+8g1KfUIJlPjgTcwweB4ZHiL/+auwfHoWO8ZgZfzpn1VVRkMRy+nopKY
V7xJr8lxbPxPdsO4mcktnjLe6ss6zVstJlnqbe5ma3pNU3SIQuubG48/NeFje49tuv9tJMmHiNA7
2y/IcUQkHQOin1qEcWm9N0F1LeWc1F2OybxJTnYRBO+GblYHaBYPuElSV+2+aAMY5kB/D4dosR/e
KQd6tMGtVf+CJ+wnRThkWu5sA/P1tlmxNcmhmITP4SRs3EmaGpdJdhYR4Tckw2PYb23cr4YXIOJt
fplV0CBRiywoLfd10FmLwKJhgXCUZWPVqtmEDntRdxPD0lWHD6kRAMCUyL6WB5Q37tWCtNc1DAsU
1VWZy8bPPmViDrNFsVCh7xgZx/d8NMIEwbc2gsqfcP9jnsYonPXeQjATrIsopRgYz57mclJ3UR47
aMhzgnWx+ClB80AdUOq0FjpHN6a0UtiK0Mtd4+ErpvwyBYGhmV0qt3PUI6KAX0UG8Fvy4mxIOfd9
q3S8HegogwTCm/N039w6zcorpdt5y+x25clXM4702Mhq/3MJ+tKjKZu0ntgG4gMHzefyHRzUyF6V
eePvYww9SErLnj58ww3CVgzqiDjezIi3CylB/Mjm9Wq14jYuTgJA7cHSprHBdbd6y2CY4qtCbU4Y
c3M1N1jxXVUSnrzmJZyVjF7S8Sassex/HHfdYaPHueoTdnDu5zlP3YId38nWR4ZLNP3apGxFV0H2
qc6PCiHKGo2YxcpXZjjvv0UicdifcFAUp4UOZCcvbr+T6czIfoUPbTsrAmVdlbmhoJPtLUpxIr2p
XChdJN8+NftscUmSS8Z6kZPOF5kxpkgzfxju21zj4GPPQmeNv86zTwrb/wC4p/KAlHFHE6JuRAwB
JRJv8hXfVCfNIEZ+UlkCKBvpoHjflq2b2F0Rrp9yyedBsycayBYPnH3orCdadxqMFdSLjWXc3ezi
YVozEsE3sKpdVbIqYOJPy0ups/+OCZHSgbVOaTjf68Q/l1rji5CY7KStIC572jtMUSWFx3C/v1Ta
HQuMUf5GgHwuRlYI99ghSnQw8IqNVYQ8Q79x5qAifxPfO8Swao3lN30o20TlTWpFk85n9KB07DF7
TcZr8Je9wWMvmApj/dM56IxPtjEu6/Tozh6Cd+AZ4CfgTIE3CxwwbZDA4AkLHKs9W/Dzt7vFf9Ou
wyYhbSCEuGc5YCiPGedwwb+g5rpeDEqGUKQJJMJWyb310xGcJEF3lKLAnsEErGmAN6jjyLDWmMuw
jfxdojYesD/a3HH402yHvSrar9xiZD8W8u+PDXlQHUZiWkEPME+mJh0pqmBL5qC5rzG66VCuXG5G
p3tOti7wq4nGbxGBCaU6eSFc3d0WaC7v7M4mmEUPw7a+AtJ+g9/TKovscE77EzGSdz4sYqm93CxW
fsHlCoz51JpWhAcaW5coACNiYjKlLEom9b1Tisb/5ljSXlNGbqaAbxsnFukP86w9UTFj26GS2UF7
sX20W0Czmh9Q+8mdrO/8G8riEQT/zgDbhzIYboCB6v+Ea6dD8+RygDkkJ0BB7G8Efm2qlaFXOrGX
kWYF/gAD++CXQQV6wdcK8pwKgZDMQBFtqsp3YSbo4sbhLcIwuLMHVI1rYR320xvFBmzNuw8zUEWU
NsolljBpj3J/xNQvWylphnxF8OWm1hvxSllnRyTKD8SIgDQD2vibjVsq3ETgPh+e5XrzeZ7FZ04r
lwPvz07Rw9d0gdPrnQLOPeFjVyz1pdXQz+j5kRGu/ul1Te1GIqff2Ox499qhX/BI9i1OjoT4J/kb
h7DBatcMrEulmVfIL8TR6Rbiqge/mDVTbNLWqXOgvfyEOqaspvjcOCb4l/cL7rp6NeD3OMkwJnjn
nc10tZBNwb7lE2HmD9TDvT90nbZTUdPJ9H53/h7Gp/yVybCW40+bp9p+BitaZhA6us4rfxj0oDki
fNF3kJYubrsgv9fzkDzET7FkfsR8oWtOmp+UDJihaSABOPkw2fHr7xZiQasS5ri5P5PuCZB8/sgI
gy1ZsTFrcVgtfw/3oKxRC8W8rkgr2XPJhrSADDCB3ijjBaEIl4u6faw3JeP1DUbYHQZZDGnOzN2h
ncHSX2TGzRFDJwknPVSpOj2tzZ2RXhPr5M+/2JDe5Hbp1nGb/Xz+c+IessCSZw3TO7Duvw1WfaU1
9d/ivdhuyxI1H7Cqp8/uwcnb17zmkZDpGEUxPZPwQBCSSa7yvaT5nq+1uQTypIUnZMaxDXse6AgL
xHSqHM8eV6RKC7J4x60qUieWLDhue1WjRTqT2jiaH900Ix79BrYHC1UurAuH7hoIfQbYhLYmuz3f
jxBYsbcudA2r2emBIywQheQY1eih/nusw9r50Gft50375vi4mmLWjEMTJSjrPmKSLHLVz/P+Gm7T
4dYaCzTx/Rv+jly5NEjiNpaflG4esPEDfFNbavL8jc2sz7NfwYS+/qzcnQ+uBQS3X3np1NVdb1w4
7boTxlnG8wkSZDNN5YfmB9jHgx3t6ZCH5Nlo10mKjDw3PtwrbHG8TeHKnJ7niej8hBj5837bvwWU
x+bHtYaX2bfSp6YuXj+PBiGQyj7UQAklMsTSXI0mKgDEHTswDm6xIr+iqvnj5LTP+g9Rpp3gsizn
oPHG0eIO8FPfn2Ab4XT1kmNmZNWDavE8PtnKdxl6h9HkGzuyG5K+7txTFMqJ2Lu5ZWRQ6v3TqGJM
hJQlb72x9pG8p1TTJekzkl1ox9HUY7fXuOeMWLXd6N1SDummT1M7N3e58PZKozWeSzrmhKrPs7x0
qi9fyTcDOx1JehCmAuFILtcPKhINOFc9vSsBzF78O6HNk4P7s5/oDOzz9T9bck9JfnX2G6Q+BDFF
yAQ/sWCQ/LNvWc2iVyb8TxLxprxjHHskNus0zN9JzUkSueMSrVjg8gJZAchfK75bNrkZn/4Fd9h1
dCT7MtkgBDbx3D4aKBubqdCsYECm4sT8gLHbkrcph9tHTt+E3Ubmq40vhy++aHbccx1+5d9aSN1F
tBTC8eDCfnFJrVeLUTBokbCj7yV4+jW5hc6EzE1KvIILq/d0IqQCcQFAScJa+yNOhYsH7ZluwDiI
4Opqqg91QxKPzqatRlO9bBZyArjRHTM/Q0lzfTzc0jUmX8OlhKzwKepiNUvFeXDcXpRnP2+yzp4K
ghOlMLF2o9+oE2JqY5ZbXYallW5mg3ACZ7agd7r3OSfxhpIFSbf13O+M53cXXrLkwAGrT913oQut
bBJnijkKYKt/5iGZ+e/hMFFPzHB2hNxfrVey5Plg5ZcjvyWKmBrH0mDzWowJsmmY7m0p0DlZqLlq
4XcFwWNye727oMGSo3lwcPBlEwWA/PnOva9c1sKlgTW1ElXuHcR+gAn+coedQ2dW2D4D+3NDdtml
SH6djQynUbapOh1mOYqLn2gVvsT4Q1vxg67iefgzViuCp7TGoJKt0GjZi5BWGuwocAlke65B7nd2
w/KOs+9PZ0mp7FiwOC5S+kO4gsc/pam5lxZGJoYJ3zR2uZIyHFD+6zRAohC+ESDMzcJdMqr1qxjF
OCnSFQQ3waFmi98AUCCj+7wxpO2iz7lnnxKitp+J2KHr6WF2ZYeBZl847T/OXY3ztEwGF3gieLHd
2qynaOBThnMQVpEiOK3QR+pbOcl0SWN7sY6+CBZKx9zaDANFjxQydTR5HC1GdZy/9uN2NcfeCzCw
fRTZkcNt4/DcW0g397Ufiiq2pITwVPl+FjEjMOShNi0os6otwexTbxjWP7Ezs+Ns0te7/i5PdcG3
wOnxRxXWh5dehe8nSSZcwtxvQ2iA2c3Dzy7Z2cu1ww5IA1xQzxJghHgg7KktjUd0h+0zkXhl9+U0
BKF7bwSw0FGl1q4h0FamEuuAwuLNKR3CyPxjWt5nEbE+oMfem2+usza+ggO/47wwMDX4Xj6t5Zg3
+8odNOfvs66m3q7Na9vTGsOYCutAmBENsDnaYgOXsODeXwWf5OBaGgoUucSKEu2xdxJNAWE9564P
QI75Q6FayH+otK5FCbHDuNQ/U44S3pb9BMeJUecc/aN4U0bqnNzDuOc1FTrxGyamFuNEKdeDyqtn
vuASy7gEeh6x0VN9uobebaFnK+jNS0Sh+Jld7WMexFYf51o7+11VsU4dAxQgFf7JYG3jW39cXGmE
o7SuTbf/zti00oo2Y9TVT2e9Cpesa56kEBt7vCyBlxnnc/wVJ1dWawWFY9jhn+IFksJxy66/rbF0
RGOe9YxVFA1mgtWMRE0iv/tlLd2zJ7xk94/kIxz8k81nzukC7/vok9tkmDiodSXY/IMbae67CH5N
oPOEoRMCwzBidmX8Zq1rxM7LRAjA31ARbLAfn3ehR6hrUcnOfVNOs9DfoJvxbUMLKtbLTq2hfC/O
jAQf891I3Ugy37qatlWR9UB4SHwWjbGmLcSgi4/KiG59OcnfXqcrCv8aoecOEKHMlpf8APpGhfeV
pquuIspW7c9kYGF9p9kdd+RverSeY/R3d6SbhIy2idfwGCFAc7Qd8eI5XU7Cr0BfBnsEGC4tYEia
Mgu6ugMDwwqTnz+ZrZymS/vHlDEE5wxL4si2HGzvkfiqoJi0bymqx/aOuXedCNYJfl1ljlfnsKiw
yTHdjJDEs5xbVOWmyjxClMTSwAvI3JDtEXzGxLgaOs7Hy1O67IZ95ukBeGd37NAbwP09MgFJy2tU
l1pmc2viR6NxTcfhhaDOIzWZlthefoQSDJ4p8hxc1WjXVH2wuezxbqAzwznXsCFdKUt78RAF6L2a
U+n+x+9ExKyksMv5ZDr31bGv0/HCFr7uKmhjXGB5wqcr1dvIlPg85X+ezzjLVyVEHDSH1PId72by
ljOFmtksd6nvL46Q8Hz1ohEog2FxNr7bXPW/3HEenjTnHpf88jffsZlQb9hS0iMUh7Tv2TqCp2Ef
TaKQhYTqAHgJZBcsHLcaP4LCNKHrzPiTn4F1V+HDg/D27909suizVmClkITiXpXLTQNe7dma7ykm
uoJQctw7qaxLcLh+hqHE3C1sfwVDOSiDE+lpMiY2GhmsVg6s0rvPdhKe32s6+2msbmUPQpgU/DEO
o2DaxpptiQY396NtjStRVpmnaDPX9azDdXLZaGIIF2lQLEIzDHAsF99kI/GzSHkPbw7Hlwx3NkXc
KIiLNhTHNJ7wgJUqUK5LbKKt8cEtzNY0m3bff+mMD3YZRJAAKYbBFzPl3q9K7PW2Y5vQe1VjvHdb
8Rfep7Iz3hBtLDTCCtV0KDgcPiURewPBQzBg2vLPuYMXo2MVcF704QwEL99DVLXuxB0Kv0gzqJTk
/wepGn/5SAw7jJ0Qz5mHA8pj08eFn12XSOQ4ur2rPkent1oMHBvVW1zysR1VFnwkaYraXKEuIE9H
kVb/2vpcx2ob0O3ZJQoG0fygxCxNIc6skBoTmXkEe04Y2Pk8dByn5EgnrUT9ORllWrdsLeZSwdD9
x4kRwrOho3X2nGOWzhzz7OrRqOEvP+qFxdcIAkwJN2jEkOWai5ImCr5OLI+3qOwH/Bochlfi9ALR
alfhg2HcgYu4XaC0csSO+ImlJ6lMQ7O4LXn5rqav3Crwm+t8OvGYNev0/Xaz49x6eH8olSIRUjeV
NrxdMXiHjVFASwLyGGo7WGoOekAF8+SuQkUo+pe7w/KYJdYOyJaIyij3hxonFhCbb/stny6HK+6m
+RCRRqu/n66qzOJ200fHkEWoih3lAh4HY2N8jWZEztGWcqGsTlxJTWLG+s8UcMCoHwAGqBYcURhA
LMlUeDOT5fJO1VADx9ENga5I7w93Lrmgq+Kp4vaC/wc4Wkz8VNA1qiGNTbc8GijfDYFkEQXO4+Jz
CRnReh067jlRlrvum4eh8j3Kl/Z9xmSA/efFz9ZVLZ6dLpF9TEzUwObzU7nR81Xgu+LbWyxzGmLE
HMaYdO68JQnUcY2UpN1811jom3AIKRpj7wwYDhBUbaBOiDNjKzH0uNkQmm/tQkxQbLgmQEq1UgyP
LSLFfjcL1zRzaVl/NhW2W5LDT0/em33YGTwMPavNw+DRz6DhVFb+ZvrviSvhLT5UYmHYT7yMrWRa
qMQauPpBrPaXjt7dSsdcweGmo83riqcwR1WHAfWk6IONWNCvV/Qofnp/l8U0Zsa626plMAX/XyoP
j7gs9dmyGPi4foIQzFRPKLmap9OsHqQiPX9U2J04HiiIx2PyAQ/kj/MJVNHVGa7pziEKtqSv/yLJ
sKWW/mYH28zfYiUr3GcbSJiDkJHkdMQy5y34NJGRMkQbjdAt51AXCDFifO3Tl8KkwQW8TW6fWq5v
D04v3LrZ/h+QV8UquC26WL7hIhlMw7fh9zqqAKOa+CovEtdQuhBkmkZIdbJV9DfZnlWtf1Civ4E6
sTPvpfmn+IetQ6hR91LJTtOws8ix2eYng6muejBdyB7BB2dDpf7QEkL7Rbocejm2mnIYAqZ0J73J
a20AfGFcLfAa6JcR4MgKzotDwy5rvBGPu1m0Tufy8FN5Yd4KUNYZ9ZgeZ4+/hPvwrVQ4+pfUQPqG
sjZA6a4+oXd68wl+spM2yyRhHE6JLAnef0wnFIEbHm5Syyts+UMV5blSBzqc7Z5OgRb1IARih5fS
grUTUt+iPo5Q8ZeO83alk/XhiLuzy1lRxm546q0FQwas0DUQuSujtoso+sDqFJmzSAB5N5ASOEtT
oWdxOeu6g1yNnW1UEDxqp+rcSt+bejTAeIgM6EI4itBcBUylQ1x6LK5X/SAJSLQN+QsEwdBIwQUX
3NkmEfEllq0yz6gOkmXvEZbmyT5gv3T511LWEvKd/yBmQlhsL5IEufolSSFtocKNqjfhqtQ/QPCT
mNSFChrtSVAST+yTyNL4tA99uNyHy9J70wmw5JMt0LLR4wxwbJpBY+v9aK5qdHiXL6Fy1W0xQiIS
BEZ3nn7wETWthB9oft4qMR+OEpV+f2JR2wv0zrwKnaOe9VIv9IInBuL6PzF13QpGi0Hi60s+zTh0
uz6mPg5qV/8H5I/LrOSkAbVqYH0yR0RmIlO2nCl79PzZxh8yWecJucWl2881g9cP4S2PuoF4s2T5
k9UEODKUenH/Ksl+r3iufzLxeuCUJorDauOnAqxrIDqDnNdlgwxss1fex2uoQEUIIAnn8KnwIR76
05V24MRliD+BqI2OlKkxZS+dqyKgmvLNd0iPzKCOZJroIr59lxj5jVo3izACR6hVpwh+iMxpOwJc
i8QgO8kGmyV2I9R/hJKd/qLr0v+0nkQC3bMzoFpRHzRxVKsVbUt997ABmGvzrev/CBO7WRBrMbsK
8RTO/1H7ViERpxkG0j1Wg1RDsJz+21NYk7NW3kysT0bvfBFhSL1Sg7ICEHpFRQo8NuzSpJj5omsN
ifCo5V3DEsTzP6eBt7egnEL8H7fmBQqJJWv26978GvY8u1Y9YwJw3GbYFugYJYPou6LYPZK9rXcF
+kVXY1SlGz+Wb+hx5HzLeJKKNAqEYV+FXEKDShYT1mbppgD0NkhkxUYPwWPifpIqoV1jGYSA2O62
JGWD7Rf2GRArtnWXtk3Yi4uB4cKmMaGRBPyzwkxnxA9BeSXBOsj0blmHAb1Dp2rQ4OW5mZFb6pi6
4p0IoqhjWYsqFKElhZTBXE3fN6u1/GO3xkYH13Mbm3mitWXBCdnFBS2XiMiz8Oolea23eAyr4VKh
CWniN8F0kYr0YSYjyLkWUuscixIFb8of8et26gs65IhrRS2z4Hbni02tDCqJGAeGrsUlDmvnjHjn
k9UmkB8VFHy5gsjcK1hMQT6Lp5eeAF47qMROFb9OdQpfSS75T2gG8B3pZSXdUmlTbAcPVy2wX1KJ
PX8j8ZyeE/AU/k+GsEZ81rVr26HhNx7vBUoctyfo3D5RTFdAEAFU/PDz1eglNTPyKmxm0sZq8IN3
Blj5jidRX9RpjwMcsgrqlMRgSZhRPqQJc0xePIaF4nm1mLinGYAjjUWaPk8bpp+b9UlS94Wrx4Ss
ecq2a6gmJtSC4a/snTVoiMmagjcOvl7+Dk8P00YFChPuqFdgSf0AZVqpMkWUGwNQvyWVx5bZUUMF
mT9I8hVitYIcObX3WnkxgTr9gcdHD5+fHjucHXFHmvClr7jkqVjZDJ4yjOGR1RnJO8dnlh5+0fEC
IJJTgYhVjgemwzdxaNbDHxRC6DVmKwoPB4lvedOr+QrWVQdKXWrKNLPL3enzUV2Nl7ySkwnigLtK
l8muw4ItXAcsS/25hTaD0NggSpTmKBSzypdnhhec/E4NF2mE5u2d6NWlmCBAe9ZBSVL5A9zAiiMM
K1hDO/Nkr4MA/QxO9yWQQz3vFaqUVZI+uxHGnOCFg9MYNPLDU3UXnHquU2RFOA6hL+z+YtfoPwW4
Hg7+tPZaM7x+7+drhG/udi7v/VX0xKkUCLyRs5JElDWI7GjHrzdKA4C531jHsNgxb7f4yivvWUHs
WAePCvmhhflBrAZjxFQdm0d3NzAuq2TzFVkCVbO/vxa0kxX6QTZP5OnoGV87wj02cSa5tPhFX/DO
dKDCaflJ2EyYFZBqN6aZtoBQzLEI/jv5njSSduGhCNL+8ZSENzG+X13PfPBCuVtp31iw23d6FKYS
Gr6HT3jPWjDM5/5vbVVrL5w4oFL06bdI0E754xa5CiSBuZY4HFYc7MXjbb+3QFLKnTUFyquFCJts
pXr/VVGyziNsZnx+r3gvp/QoA0iXVPhSjUDexBU4A9SuAJgbIhEJPBZhgs+wPBIppxH+9/aL+bzG
r+lZosElmvb6tPexmDuLgo4XbNOPgSqdBZVShAk1B7UkZIsUaAvrBygFcgQmg9+XBH5DOdIb0NTk
BntH0d5HCdLAvIM52ZdFs3xluc8heYucBH+H4mhfD1X5moiNowUU4bO7R22gW6d727PToLBngNjP
ZXfOtUOc7rgcdqlYQiKcGsD8gVQ0yFHnctgGdXk31lJ2AGsRluWB9u63/tt31p5jaKqa5w1WE1F0
l4jCbPbP6UPHOSptEa6qTknWj76WShGV7ZCqgsYDfttpkJKXNiuLseOaHVxu2sp/WIUseRJS9MIl
cA/smaXvPTB9smmyY/TTuZxHC0faq4aFGMr59vJpX1e6Pvq9ZQNn2KvPWkKw2425VYwUcysFBk/n
YL59p7l4rCVwDVKKwV8hF9U1YvjYxakMP6emN50/kozY0uHNyteJd8fyl/ba18rtCr0xMX7cAar/
Ft2UgAAg9DoYiFrk5vZ7O0oBBK5YtOJ73JC4rvIf346OQ3l5S+fdFlSDM+m0Rg40mMQV5H7eY/r9
+EU71AesUirZLPBwzF/PemFAhH3HKbEZObRRmEkv7dHYfeDcatgVpYpozZ5rVSYr5SQGJgiUAvqE
Tl7g3U27vP8gHCISNkOGiNB69XJdNXJGuLB2+X0qTqZ3zOEMuvQ5pAQeHVy7bYUa5rdLmZ0YLeYh
vChJyHwGBTYGx1xAoOaIhvA3C8ILLa1B/MOjT/QwbRZ/6NtpWpkADsxs2jCKyUioHB/Uy2QE680f
Syg73GsgJ2t4XIPNKyrYbk+4ZZ0K54dMRCCLfiRcvREsGRcTU5Czokki7ITBhAuz64vByJWNGIrG
dePA6kTbt7NmjJbjCIubyPUEOPbwMYaKbDoEFzJgXBf9m69nS0dTK+SXol+tDdqh7H9N2FXzE9/L
Dq0+2orQT9K2JG+WXnkDNAtFQmJL6JRnOeMDXX/E96hziVLtyYHF1jrsogt6RlBQ774DZWeGRZ3b
7zYnoKOf6mfFqFG282fhKiqShGp33uSjKG4Iv1qRF+rNDbqnjpq10+KRRg1R5Cm4HIsBPAv92Oxk
EhYr+nlZjO7k1gqBpsG2+nasqWfoGJ9Cqsk40qY2/7Ve5Ttse4ebPogks0Oo0u0rq7+71IoHKSRQ
aXjNlNbiRAKuUkuJntvHRJyTw+SEBos79/pNBnWcwNZlPZ4iAT+1uGY2fpBmLlY79+DB22NtVo7z
DisoCYFmDn5nTvzW6Qi7/6zWk1E/gNME4sAaRMFpvLZWRbvxyKjnSfE4+dI5oipjwXJ9tSs39LJN
cRJjrMWAA7YdeUoWyzjIuMG6e0ffDEeahwUHK90R44MG+zmgUixtZOTPDqcG7jvkrQ+IL612Pelz
RCle4jJH5R1UVWniFdEvqB5VExonv0z+PRkBFesZoPeq0wUWfpT/X8d7l/6XXDxrL5orseJLhGNb
DLVwoQOEvY1m/9yi8qB/2QmThYUGD1AHd1EtBzBTlhXuHgEoJuK1fyvPmjztKBRqmmUKZQdLRzKx
6hEA2JxUkSpZua82hyR7EA/dCNTP5NMZGUODbjm7IalKdx0sc7YtAO+w+ovpjx9DezQGYVs08Ajp
JJFQR862BTmSX9WWIPUm9XrEXKMTwat/h0x5uX42UAo6f9SE97M/gK3u8IcW0EbsROaEKkN/5OQE
plunf8dHr4xFnxJj/rRPbc5Pj4cT2UJ8omTDBQD+cvCAoqUvu1DnQb8uAIkiCAsaFul3WN+aal6F
WyVFPE1nggU2uZ26YFpB1WQoGn/W5LHwp3huy9nDbkNwwQ4ZvY/XW6zKSoaG08VvE8Hmvyaphs4s
lAQsjLr10oowXgLjakO+c8kMub1L2Bm0TorKCyljiFYSLw+axRLj4AR3kXB27Z+TeeI2KQ+FzhOW
tTdsnkFiwix5YJtfqOJEoUxD01Xx8UyPwbYbeC+bbkYN79UgdnNiEDh5VjQWN46id8+ZZRu+dbrs
MZVrIck2TrMotbEc0PiKHmTxac9ctz+XG+nPSuEj/ZHU9fb8wLGeNZ9LQNoyt7mAKl4yUs8CuUD/
BVv8tMXfBmspMM2KD2qwOXlVi1W6JlpNxBiHV3ssoit5rthL2QBiFTXqIo5ySTb7PHhGdF8MpIZn
vtRXLp9mepvJTLUVTtZgO67V9QUHspO8N7pNw2W6hoxH/oxmYz2oVzrPF3KbpDqJtY4WK06YNoVI
hvPjf4wUGOK0SW5xMuAbikCbNREQ84Ssd4TT/C58RnDnuwaFD6DHOj3wOVH3fGjafaOpQ/aFF7NV
qheJ0k+zeLHiuHwfccq911g36mb/+leBR84ejuKXBH8p7WM18F2oMG4znFDiGeD1ZU2ZJ+qQ3J7g
mHqoj0oG5yX/mTdK5MnnxVYojxjXKuhshHjNLNMs9ykm6V0qV9tsTdc14w2qCusitzYkxBi5XjQ4
TJqufm4FZzmx1gBjeQA+QDPrZyS29PsibNSt1XS2vepCKJIGuajYXydjFtyJFTFoJn4Hvh09mW+O
oyE4aKHsvMVXys4hMgqi47qwL37dw0wsi5PidlisnaQrGs29gzl9FjpUFp5wUy+hJ0vwSYPetB35
GYgUXU+WTVtgP2MIR94olvnfkmQogAky1NsOIqvcrcXy6/G+WF0YszcRX8z5LBa1A1Q0TwZAi7GR
Zbf5jhSdPXdqTjI52vFSw4WBmOWsU5AjNcz/IxONAzeni8EMHB86p6xWg/564OjgjRQymjyERyc0
WpjhHd50qMAUID6nHWMq2TRA3Lp84Yyp+k4d39Em7dJiyRzJQx7SrRRiVZGRvpKmKFRu8b89yPia
wKegv2yIQ9t/mN+AMiINuE7aFTlBnrOqCNV4CLS6nIA0VeUdfL+yUV0zU5BByIisaGrwLpjIXAwL
tWEn+Jbh2EzQ5GJKhQL1iRiiDBj4AXyro36QWiNDdrK4FYhaN9yvypLUH/Uguzil75t1AhnYECVF
A3v0T9L+7xLIBvdwk00mlrxEzv+XiNI629zwFEFCozPjSIb9eDXQSXHwli1vPYGt6S1N7x1+gXuA
HFS2FfxlaNT9jn/BGYa+Yv8SQKo7GMPRr8xmSuaD2SlhktuT7lewIQFVe66NSRZSX4albLHFV6lm
Rw30Fv05vclDct6t92Y4Oa5m3KF8e+4JqrYecFwVz9I5ceqsr867piEgjAYXYnKy8Qn/8bxlHEXU
vAJAAFbtzeZOpvWgllBugjdeeh3B3ws1o8xcQjhl9ABK7pMcGLk1JKOHS5Jgu2CA2dhSOrgazgnD
yKsaNhNgxitE9oHKSFZAJLndl9gWNUNlF4XbAtB9raWcobRtkL9HC3vSNbSwH89zVZExO8OiAaUB
qC6CosCO15JdeYZfBZ4pw3Rsa/vZgdmLUiLqYnsbr7zMRUxBeRbTk0JfL4dbwIVqa7SteU//Qhcx
CDE95eoSeGsnrEgHC/fTYMUsmCHbX0S6h59PFYjqxF2pFhasuzhywZsx/TbhH+NSR4UbwY/qZ+X0
EQaKL2oD8ATv3QaTuBDiqJdnKgpaYBQQxcdmry31GcvkcxPm9WKfP11Ms04OrnzG87X12B+c/MhJ
SJv5RwseK+npw+hjzMFa1YWln0HVLiscJYydRg69097zKz/i/54O1ZlSOAbdGuLSaU99BS0r6tSo
g/nYE+MJC3FIsqo7GVS9Bmdtt62oJ4uvaHkvv0ZK59GUqU0zd9byEvuUtvNbrRAcg3N9J2su8WhD
SNmL3ZdyqvHmLjUSU4rmV48f7Oax5PqkujKtbX1m4wsi+D/U5rX9Fgkasoaiqhl2+Zmg1BXruYLS
C7/a1VmrFcDe6H73X9llWYh9fbcmgHWpf1xx1ikDmJb+352U5cPoz9kV8HoMnP/UpDHFDDEfJHJk
d5xU4hfxvJXpI9Pj0m7IUo9epjCX+8xmqvRqQ+sicXiYfRC//62n/gNzGFd15mjyMTn+yzJCGWN2
TxIzj2FT87yUaFTOzk5JIWB+XmA1v4ZpGM6EVOgCBeN3f1+T5ABJHKaHMc7ocp7se1XzMpWIa3H6
6zSgTiXkN/hcpGhBiqgftCDzCyHd8JGLwDG13oY05npVhIuJvTJrdEDzk2iv5ivmSZMdRFTFX/Ma
pIURelN/HLIBFRYnAPTmzy+Djsiypnq8zKs5SPFDFxaO2I7qXypbVD7PJACL6pSLpUCgth4rpjkb
vvk0P4AIuZlFDY+jTrduBAk1/RwYWtKRSAM3JigsZRw1QTOKLl2r+SBFye3MvKhSi5UzaNe4/D1h
IaEsUI/aTXofkL2AndLlaBqbTqtDhWVviKB9GnY1K3nB1ZUVT2j3X3etcq43SJ2gFOy+fnaWKBrF
FqeX0Cmq+umXq0/bArcy2SM8lEydgN+0eEW49sSulPF+uZQD4s/p+E3IeEavJDig/yKvhkGZ6xQb
o7IRWH4Vmf/zr0yjW1m9pMO11ZpgjRmt3eBu8KcQWRKAEBJgNqw5wmv4Qhshpoi3vnck039e/iqY
0eaQbF0qj/Zb0QeKU5Gkj4MPiq0fANdm2K/qVHEw4z/DROT1otOQwi+CNhQuAlC8lSEV0rc5Ukzd
pXnBEbi52CgJ14QaG3N3sBXkY2cpuKuPqxada1yRHKpL2Z4f6nCvveaA2TtueKUl8bVIIrmboe7O
bXdUB9Evfzs60+79CuY7QEJBArca8vdUOKFRkczWHNoO21ianpEUb2h4XwUXMq9gWSUbRU6OCcmh
KtcSXTEKwyIVbq8ILlrw5anT8dyLq6f0njGQ0WVkSMWKZ4qcOn4pEVhTTOWVPM6sMRfZpasn4sdR
c1j1EMxeOT1UBCoI+g1JPS92jqq2UkmykzFhLdes1C88+Lt081z9anWJBV32YkQVjmUUYAMUkj+u
wkpMeucmZKkwnmUiDyD2l42IZTQPEan9wK4lW3R0unCKM0T0obuuwMkZ+22F0CArbdiPgIxWw4S9
TezweziBpAC/r09ndF/tyL8iD9mT4vcBDdY1KCMb3tqPJQYluV8uKL1GnOcBAB1IlR3yYxAsi2b2
tXUAjpabUuwomxr3CyfQh7jVkXNr2takEFtw6m+0G9mjPrX5E36OT/+4tbsB4edgWpb37Pbhapop
B0AOnbYPr9lWcyXMWnFgXk6SccA/G1FA83jVp80ax/A2ftOxngkvCkE3+mS130siD0IO0Uamm10m
tMcbtrFRX9ZNuMsTkz25o1S9R+NeNwu9GLA6LO7lsFp4R5y+EzXInzstrtuvEYhSCKAHUV2rgYSc
kdAdIq/jOmEAgQVbzX6zmJeh8FqKggSnHcTL+jLGSpyYMVt9w0f1OwmoQxxkTyysejLt/pJ43cQQ
cCYH9iZyAcOQrUn4myvnAnlUdyxDBA7mW27PebkCmil9zaY1w5hqgfgn8QuVsHJBU7PDdlVUDQOI
2N+JY0gyfVNzsFpnyp9Wfp3POZYRhc2Ph5XMV58uWBifjODwjJGcqnbnE9khzamnOHqSgAQozBfD
Ef+0yIbeA6Gc1aJkYVEGrOa2JZUzeqOVE/H4HdAv9dWRjN1NUsI6EerRFwNlEwB1DQQthfwqp7dE
JgMxdbRjSpKcA/T/M7cjqSheGtSjpyuD2Ec3ufwOv6/s22utlrX+qEmHnVRCGfcct/PKMtZ09ZHM
VLV/kxrAuUqymp0EsIZCruP3TDq63dISYBdJsOW6Ksbb51s2j5c5JZliCdeiGRgcAzYWMCqUA+bg
StztCrZ1HTaV3Qgtmzhj/MjiZE8lwt/ad9rFZpANisvIqmRKDfglceVdT3bkUy9PcWzpzFy1HHta
JYT2rsOUvexSABVdX3M1pUtEjRGKkqwzmjNpMPPZbjck/vo2xzlkSiEP8yjbB6Ne0GOgDVN4a9HF
fRwxUqW2vS1/s57Gy8Imr3tX2oN5jHVbFlXZ3UvMXrgR5uCpNyn0RiVEpV0iApe7DCOlMUF7uDGx
5AR1lAhASaxeuJAhMgmczKmV9xmf+EkuYO8VNEUr47atONQgqdoEE3441oTBCBmnH171Ihfpq6yV
5phl76+bOL/nQxwnzBv+ofzwBE5NxiGpIbQocW4UIC90+3y6kYLA1RhNiATRboVailn8g/rcrs84
Z6lXcFM9x27s+/+4PU4i+Ry4qgt6NcKdWJKoCv1SzdP4AO4powBlaR63w4g0qPT05Z7tFR8ZhjgK
EjoXfSDDRVAm9g3pxLvIRYSFoRWfp2enpWoqOnjt9igHJo5/ZObFZYQDql3xLcjqSnzr9Xiq4B1F
Z7mzOEdigKsU5NsLxG7KmoXsScR1lRtPDFYInE09lHkNwo5LB6fGBC3WoRKIdgK0c5YqirWpyCBF
r8DA1ABm0NbzgvAk4Dpl4pwGVQY+wM8VNQFdJwco07D5FRDLpYXC3wxnkVD1xhQGJpDlqOujMbTq
DOpSAKHNi07IX5euAbeR6p6aOUer/mwiKcnIU/Q5dAqIE7FphOXUlxDXEnAXqcUnQWjg5wFtitdN
PnF0YxO8SDrNu2rboSR1FYWszQwhJmSH+mkL+7i5JA5Eufea+gXozlGgdHOcLMJss8clvjvIP2nM
tPcr36Dkwk4VP6vgu8hN3lI+ngvPd9KcCxvbEGiyNsZnbHL/BRJNFIqbWx3M4zniqaDstQltmXqa
3r9z5VCVTdp/HtAqoykY6jnsEmnIlnxO+Kw/5yDtY6ssRZ5FIbIoCivD7Joal3em1CdGQhxaOcGn
iqgtcppanZGZO6LntCsJyTjk5WEyzO65cahdcA+SZwAeQPl86x82XbSRmVrPexNwdv2i7JQTdF/0
UOAB8ZKE0ikV47gW1sF/7dI53GfuyPM3nUCxZbjyPK/vSq8BbN0MjcxrrkT+Qn0enyJnlcRtaVrP
q/X6xC+rjhI5RtZ08WgCClabuGkeepnAJXEgob3Cb8sPcdpzBIpBsEjzHtzjwzuQPTUDIyhlHmuU
ur9f2PDCx3g9N5xtqsre2gZO8Mtvo34DvppXAV6OV09piA1Fs0w9CnOpMZW61T2xKtgq43uXrqIJ
GyaMyzdhnC3h25YlgFoTdjUU2WfiPxEYNe/b5cTCksJfyOKb/FMcDY3R+0Jj+n1VA8n/ZGxs9l+i
eqBunaBw8+GlyTiXESF+FQVrnZfbH/Ayo8FqYiPCWxHCKzsCnYlI4+wNogvpbW0oCLyVpg7iyjgy
bdasRX5ycQaq/GLsre0nczEjN2BtqmZZuG/hNoopQ0p1JTRizkVA8e163ok79By3J6IyaLiGuRo8
wllD2lv2Qx9JI0+ZGMMxuEFUNJx/vc40VKNGoPCJAM+UP1dxLcZiQLPPGxVjihrX/FCvkAiNZmBL
Fa8xIeq97ERvQ57PvMquBHXALgeQfUL2IajusGV/FBTYn3wYzSZfqxdKo4TLi+I6mlBiXFrain+P
eG7hK5gEgpTLF8g48ayUQr3qBsuxGtH9dYW5lmg0YxqtoL5HSq6TLRzMUbBU22/wUzXPFk8JQ9Gp
KMdkSavyyUc+XG2BlBKopD9DAblvEVmLldcI8Um6RRd1bWaF9xXMAGmB6yU6v6Q8sDhdG3aMCN+4
zirQk8k29ZC1rLYn1UxieQokO0KzQI372zszu0KFF4twKsGZ27lxahVs27uPGH8IhHrhvDnnnsEZ
sDNo48aQ8AixxY7n+axlZEvrfCxnOa+fZtSg36xrtlpF+Gy/cCn1S9KlXCjxKQtEgLEzmie5rDZl
LJ42PUg1IrZrMkN/lLC8d6gcUw86j4sLQGoOuvOEDTIDz4/VeVdrF4jU9de988EPx1lTrrJQaOix
/ti01ovU3ih63V0sh8ynF/+GIL6NBk7/tERewn8LnafX5Y3zXIONMBtUKaNqsrlDF5kcVKwExUcn
Ia1/1BSj4idrxFYl7+Rc0hBu2VEul+8rGpd1Q9Y5VEaqQDJUVBUXrUM656LTzb9uQwk6Oad/owMc
sYRh3IRfmI6YSIDEgE3iXVz6B1BpffqZJAK5TknD7aKuV00ZC4KlsPyQ5LjxvmxFvqTojyJ3+5+t
Bz5eTCY1MPnu+EnsnUF5Y97MICCueESlmzfuIUsW9LHc33uqzumWOrbWtiJWb+AkC5Cm0t/ZjAoe
H74JUP6g68a5AN1YtBzSsRilkxq6J0WsHbs0tZyvqyn63Gs3JY+ufm+1vU5RZFRRlWqdM8Vs3Ph6
bPLzq6C1r4NWEIju/TGK1aLMgkGLiZA1XJCnecwr7/6whUNSti+o4Mg/zDrBi0B9tDGCBqnUIRZ5
gwPtu4V7PaR33gBUf8SWGwDgtNt340r0KqKqJ3LcE+7106PMYmzy1bQDVDkSC8Z4zJ+OOO/lEctd
J1LyhVMoKiderBAMPPKTHBDqyWiqpZ4ziuDsQWyrx9Og2gPsa0o9zziO1wIWoBXaSClI2oa079mm
6aiNbm/xHCBUP2rqd1XLB6hB9BXXq2IuB6H2T6pkP99shNJRNK/JgM4Kb/O3hMTDswmn56KBp0XE
Aj8n5Y2vEcs2y4rx6bIj7SziDjxcWStEbiZvffvfbCEpzUB/QSxB26B9hf7R0LMv94SAgp7Z0EEt
pM5BCSH5e3Fo58quU2qsGvRxuZgE2TUXhHC+GG8Vwcqf1379ru2FsfOfqNIEOPGv/07o08yYnQRh
sRJKJxUTMxUHv/kSGI/1I50A86xtmhbHK2qMaSDnr55UMIf3GE6GZ/hH4Wk96Q9arwwbtCtRfCRE
vJuS+NMKgYtk1yE57AtgV3rStXzy5AeqAqagoEYR8lDucVz6u71USJQluXWq/M1hxmdg7/wB9ESA
uy9FKO9qacwzu21UbTxWOsZHuFLZvlhqpu9uQvpnkYb+5KVPtmkZwSfdfW/kRMRTIyQXdVJ9R2dd
Ak1YACPB+MvxZbWl3B3KB9Zq2klOs4lXfDjyn8BN/S305Q3jjJPDCMuj/KYAWJrwsXZXdhBRlDDR
9+4pUNFvonkvxj5UZZCOO/KOk2qp93PozY/VRPGrs8ZP6+XIOqFs2zYGvu32GCcfKzdlz4XLkaXC
1EzIUzssBRL3JMIAsSbaTJHRVuoBc14KHlEw58E4QmDGLbEslUBbGhxjNw7Mw9p+YAJ24ALKbOm2
9TajL06RvoveO5lHBCC71EzXnPIHVUDxEsQX1a5OL3+DeG6Ecc8O9B3tDWXTBqKjgoy1j6r5w6Bt
zuL8bQRMki7NTgcDNN48IFUS4RlS3VlTzCMfQWnhXTypv6HEfZH6fNXZoMFN0+zHV8Q+OoxpMOgm
Do7w4EGImDycW1PETctGKwucrwrqIApjqv3oHWiDMrQRtDhp9H9vLZ16ly+7dwYGA6K1sr04WWFD
uf1OCkBmYlFj9izwyWZwddeuO+AUNjjvBoXq8ZBC3TZiRJrNWnTQ4r78tE518f84zbmy/1sRK0Z6
xrfdz0JNA734yVJzHD8eJuFqohM7nrCmscVIDb2up3WPDsE7xa7r7e39HnWi/9QZiqLOSDuX1g07
LEaAQefPUExvVjwMOox1fbUaePzcWXbFPE/ukBjUBnj+Q5p5XNAcFTLl8/p/FADYFyhwT47ZYNRQ
yhj+GRSkhZsbC363i4694xsv15HPo4Vu5yFu0HddZVlyOXkQlEwV7+sKUIO6VmtA7aDiJgWx/wg7
QMTWenKr5USJITbvByJKVeLVdJVUM3QO++qGHQRhsJr78FT9PAFagxfA3lR/nTnABvMTPXEfyvVe
2yqu887vABxmBt85+INxcrAl/jyHXFf4N3Kxrqvr0/NbFgmxe3KfyiwE0v5GEzEv0WAta65eyHuJ
pANBNQ3YLDWXI1lfv1Kvaix5JfErE8VXiBsKEkYW6QO7iQ75zeQffKFXFxkQY430jZrOHe4hK9d3
WgC+tAtjegJIfoL1JtppDBZM/EoWazhWK4sqxHXJ+a+qZiZsLTNe+ywPYS7mLkgeia1ESo4YnAib
eNP7fgGgTjxwnXy/Q7w9riL0tKgkCjHUitiaDcLO8XffyXWWOqvq/sSGYYg8jK6mTK0Q/rB8b/vW
tBqM0TxABiyPNHOgwa8TXEd0E6jjFmYEkVqQWM4bWeXGzIC/3r9r5HHaap5VA+RoNZENJwTCLbiQ
xYPh7WkNtUVGNn1ufJgtPF4B5GGuxKxU8LX7eDN4dOC8gbMHVIAkIJrfhJB9+M3Kw5e5yvDXyM0n
+PFbOmaM7HnjDuGkmKMCixkOI0V2tWtfr4u9ERgCrmV/cU5W4VErhMrgoDusCSlvc0FoCp09dTOj
IAO3vAGERt2Xf6g9JtLejs9AKsf+o/cW8jEyqmc04HhS7P9ScHhqhKsNEEsDcHKQycPf9+OzkB46
M/45D3O2Qj/0gouQmwVO2hv5evNSDOG7Np4fN+xLPKSYtgfGU+KQyz/xfGCIx5ayGlW/9l2BAKj6
dR6cPltx0vGyRJYl7/s34DwFydeTUrPJfVy7qUUdQFWZsxvHMssKBA4vf7aE+OTlYKfBGmjr/Zi0
nfjn4FJHd3TxW+/z1t5o8ZOrBNzBMbwIgtYxEV1sfwOjqSDCnNK3odHMUM9KSBlRrEEs7VEnqIw1
KMB3I7ODl3cv3NJTpDi9dwo70fZIM8sj13bZ6jnSGbyCorrUi9w/jxeHwmNYihZs5xLD8dP7k4Lt
RxyH8/jkf1erCsGdab/x2x/zmYQnMv5zc8Y9P59bUq8HdTU4DZnRtsaCFNo5h0VzrNUBAZxNHvw0
qPAwn4mBAiOqLUdx2Wi+EITmdbezi3pOnHhZHowMhSHaA3atQt/XyC429liC7cs1F46YJ91z1fhT
l57d6tgJoSC5zcuAQPqo9Qvoxe9nedTxCE0QVlS/QcNvMQ8wknW29NJSepFw0ysuBdQKulrIzcYX
ok04fw6F/IWRmJ2uL0VCz4ENdLxxhbgbe0hAF5NVzVz+8PwlZv8vlaZVTBKKRxvrXT1jESqTz1du
d/XpfVlXOr5GdxRk9ZmPcEa/sm3tlMMjW+AaUPcBNM/b1IsNNMR87HBxlsbdf9PJwYfaTxgl2INE
I5pGLBZ0OgLxWgJKnFuWlXxjbNYIGnmrafxlkhY/7+U5WsjplWJn8B1es//dL9SYLLsi0dyxqQqY
8BY/w57JqEFQgXFAI/pmKaidvN2zaM1qwn253CqsXh4VyQU6krl9vMX4ytCwVjWy2DjK2acnntwh
jGa1YktPDnwtRwgNUpO7ay9VNAtgpFnFXIPrviJje4dZJVzbyD8skgqaOpCv9T6LD0OY3ZnMcSKm
QVnE3ooOCDRMxilVfQ4EC/hta0ylO0GWzRMayZRloiqeY7hMl7CuAvzbt8/LNsOGP29Fgh8XnvT5
TMncZZPUAbkwvO94Ht02CMQxUTemARJT/YxIY49Glf2CPAvRW8wQ8dzW7ib2skcs5oEKddytv8oD
IQfFPZoDDiOmKPRiKcn8HqYFdQt+Qtcmc/MjLW8E+a9Eq8us58uOTvEnGN5o+HalLkvFAlYDkscj
fLonvOHRYZ+ncdKfG1uCcFyJ+Qm0oFHBbSWzYCwr8EoTMJT90robUdz1gzBe3r+oJcnke97yzbgk
saW+FizZwhrDeuAjo3KdCdxskmT6rkodInj+CSnafywPj1WIkcbhlpwbH9RLsHnDjR5S02tzi66l
vQ9SC6plJ+LIM8LRXCu0aWs/0SQYPRCvl6EEDAQhzsZ0uNPIC3R8stzdBhzYXftVFZnawRf4uwrG
XNTGAh9a1JFYtxTNu7fA1uyBJukDqrLBhaGHHCs6mgBwsVvue57v1CjqHfNbe1nT84WIVVKvmm3k
VMXQWdFtQ9Yeo1F/JOOOv5mA6zUaRJn2s2LOsPqZGxdMQAaJYK+2f+J3oV/4V2SxBk1z6s6KZnVE
faeHSb2/POU9H1FglTFcSP3QHxTh1X5wBWeM/NoLjnOnvm9kZdtS0kTPG9lOxwmrnf0Xc77VIVeL
MSRrn85b4Ut87YuxoH6jDVZhmsdFZPS8GoMV3Zd/s5dfyFQSVmLwKlGpRAb81KAnJNKCzePkjYSY
Ev/QtsSMZgtjHw82SV6gksiDVWm7oSTvG+G2nv2btG95/0SrtRCLGDwv00nkewczduzjTqLt2C/5
DX91ZAYWI7P7MYlXi64A+Qeb7v0/qfulWxw61irua1aiL2HXt/gVJm4R+YKyFYYe7erUfzOSBZxx
m/s9GlCIcJmQ43kwqK6CKtxdoDCSxNg6kvCiuHXVOlt0+xk1NQdMTSc5Wotp6VVdwYKU2vuw/sNU
ruLDPb4o2PXj6zd5X7WiZuBhfiCjz4fVPFZHlvxBdd614F7mm1P7HZy8rFOnSj78cAF+x1wBWQBy
/iuQXchPtkJoMFP7ibLwMMWejUsmhTCZAeQJYe5nCn5GEeEVvhMASEj1TmlfGqTssdBh5/xmpp+i
hn0RL8jbUdGtaS3O+pVIeg0EdFdYDmXeqUUGkl7BzAiMDOS+sDFMsYH17LvmzApyShJcf3DIbBo7
6M5AEAQd1T1yx6mqEY2ffqU5rz506mZn11XkeCLIyW757iLZY+g/1bH8iOR2bsTww2sJPVVIW5Os
RzvlLw5X3UVH8bfcissIkWy+Xq8CTsLeUjAXHqzUiyc4fkFKGgNp5SmAlCz/38HHgSIUmnZjZoqR
QrFw6g9Upv8abx8SMJXeEB7JxhhWndShkQ39S0TUrCAbap+xwjgk4cn/7Ew3tNzaw7GR6AgcLdLe
weVbybVmr8vJOWZRK+oyeaAfB08gDZhyfcRggW0O70yLhJVU8G0JaDviZC+cOPQ+EaOt5/AR7PRa
VPgG71jsJuOxlign/fI6jX7uYZpJcEECkIA+dN6+y6040tbDbwW1Z8t5Jg8rjwF1M23hAdijFZkK
5GubrYoHZC3HwQJS1ZLatc4M/9LDMs+7FXmNYlER0eYuZkMoMXrEcvI+Aga2kEBBdmqGwbkVKsNc
rm8CW2Tjq9HWyJLyCvXq1ITJDKt92KtrC3+3jPCTJsXvjBYZNgDSVzg8Ov0q4/J/+h3bLJI4fcy2
Lt3pnFVVZ2+wn6ePSRXB5Pg0diRLDivCesLdNbxsvLbLCaBK6JEvccHxfwsgCKijltg3u7DZ1jhi
3+/RCHluZ/TwXxuDnO13aiHL8KrjVuBaF1/mDrYSLY9x/7AnOZyyy9IwhHv683BvfUDHdVCquzjP
ean/K3DTpCoZvBl4NGrJBCWVZGPY+5vLL99wcA7ibpj2IVmcuz6adcZQ+stCOxIdHCmQiuroO+k9
i+pVVeeNBSdSgBpCE2KI5J+vDGSVp049JI+B8HeJ5LVwxHrOomGXE8UNBEi4VZnsx7aoTfaN5lDJ
lJG9ETx9vpw8Js4IK0z6LHA02ZvQLzpmcPA0MjRqIUqQNHAtX8G4i/aACi451RSA1XVI+g2o0WVu
LPj6fyQoIU9cs900tX1LfBBkKaQYnLhLhkgOMovdj5dJ+fAdf0x4hrFWcWKQj7VJPClqZgnHmU80
qp2QfZcY4SEte7xDG954eSl/XKqg52U9KDXXJR9E57ADj/kv0iNJ7FHooLnq1+wjBw0mcf7yNg9u
Tw+9ITpzZl0JGw+5hYIahB5KXxuGlkCFOaqbXQ8xJxM3/6a60qLSRFs6hTrOZOEqhAESm43o2lYu
vX9SQtjw6MQm65daDXiTiHGpbNtn1sBrwjG8CN+RM+VIc7VSLWbA5kptm9FcyJ8e8woMV5W8nufK
zFYJ06o5xMUBNus27VhFrPS+eD5CA8ydAgLR8FEU9MpQSNr4UHsghG311WqRVDmVgeyDjZLzNaiE
YaC+Zl7njQLvfnjsYwM2SluOdB9xmz2FeBcDQ3z7BUkdEoA1cGNrebJ4BeydUiJptjt9JMOasmZY
za1brpks8j3JYc4ScY4C+VV7jLdOaiPpKfxXmj60c7Nz+gYKpHArufOULgXUK3qWk+VgxREZ4qfZ
qkn0srP7oCVHYccbprszvbpHuVdu2ohmNOXVIjS1bZwnOywDVHUWbxexNfCAglNoADcQxgcJdJNL
muj7xsov6V7RDg0BWc4PH3XIMX2fbVpdr9+tmQ1mT+0uMdysUcAMTcQKTzl4f8tFamCVnOeY3Qzh
aYj/n7GwnxpKj8Ztu9Mir/us9SgfpKv3D6AaAlHW34xpiu2gNCQCZ5jILFW+S3lI+bzJbV/v/DSe
q1yOAyvttfUZL9PNzsfUZofr7bcNFRDFXjfJKOmZY9n3sfpZVQWPPDmk+CysXtnYsNBATdIt+fSR
ioweprIUkFs8UiI4jymqJgC0FBppiKeIruWdbiHRhU0GWsetRfSGCVNTvUTBMWgwvB2KXu9HwO/1
zK9HkHeULAFM9xdMmOXeiL5UrHKy+Jr7oW2JGbRm43yoNUomfphr4+LBjryRq8bDIXF/EEQehS5U
taNQORqLsajAGRtxSzMDipTaBuJDXZ2FsCzLK8xzbqtO5FP+eHYSbLk5Npkt+tQO9WJBT6aH0eK2
Ah/veRg9mymopBwqwUCv3GnLzI8Hq7TXvmF8/RGKmRkfPkbv4OWp+R5ahPY5srAtyyZAw/CfbrCc
EXMkxXBP9Fwv2flhekI8IBvMXnhXBZMtkvR1yvyuVQr103J0Sm/y6tEU6CTl+toe//HA7J7hYpJ+
1lgUj5ktxu3hjXWL0MaDyjTYn4gjF0TJ7D4VHar18O/XVcS/IuSZiqgx0uRRrlPU8RyNapUNK5qx
sGRYLUUXsGZG6AtrtHWByq/CYZih0/QM47bR3skSdQbLxkwCMTpT3TdZ1GvH2F2xZU4q3vRTJFST
G717nW6Ayv42w58sw2Ayu9ohr/xO5tPnaRPsOGlm7KMOyapVU9RtzsFza/u53kwx9ljfe8HQwHTV
+ebs5KN96oBDiYOR1LbTxfFkgR/IeHWZ1/dr50V8TaPvjzi3xbHVcM1pEJsRgdMt950OrtM4j/19
tdQ6YWUBIhWHxioqy4OMAl5nmysRFuxybkcX6SLi4fNq2EybbYPlel7E0drn2ui9FXgN70WlcSiR
GqgkR3bLn8uWoOPeTjiUEgeMHFOZzqReevsT8CWBQ39JODcCFw70H0zILR/lplBGDMY6m23uRmDy
T5kSOSJc8Ph170kcxRuoFxGe/ihN9l9tMqFD/ygpQ8LJRVDQNUAWrJRD3LvOtlpEvl+QRXFPipAl
2QhN1zOEgV/n7dfacGW9O//D0AxO6EjTqqoZm2LvhLzq2wm+OIZIRCjQ19d4FpU5N66e2CHeY85+
Ga0w8S8zgBYtryQCJhH4mpQALJQLe1LhpsZqrUXLwDTGgVP1PTUOMDKpx/UKHJC53I2/IlMZqjlL
wtxMnbElwKP05LuQk4NfeEBrWFue3TwV8w4oO0RUz25jL81P/4CdDKDktEely6Cm5rD4icIwSFFs
NwpGk+8BuAU5NEUQNIagWB1UqEbY6s92avttglIkLPeKNuMRo6LoaG+G84Vozj7QHGGIA9M/5Kav
EU5ZNO8MgMUuqFgAHWaxNkGiIqYbHDSjzLyYHY5JidEo9d3+fcT1rHl49nBL4CsqhyRSJWwkvvjP
tNQ557Uu8V9lIugTUl+1BMGff7z1MFgfA87mimHASCd31Uo5KV0BukykL8lt3HUu0F7Es3UJhhNX
TBgDK9uQ4hQCMU406Z/8tMefXhIU6oPykXMOlwFdFEaJtQnDo/hgsw0gd3V8pntSZj95uol4LIc2
MMTr1SmFUN1yk2n2pjRCX4/V/j+O84Mz3beIy5uv+JX08PO3Zjl/SRISJ5HQW3UyJjzwfPiwZ0iF
Nc64HaYbR8cHnM1AIsD+2O1GWNHoTvPi6uyhUTKh26aMEFcxFbZfrhxBLIAp3IepO4OJKWEOxpFv
XR2dyyWGYnOL90rsR4bWf55mjZocX5VuwPV+UgGgGMGcsklvoMLGzrlX0/fZ2en75osbpIGj+ONp
DvAdbdb2F5BSuWaXP03EjVxHhPGpNCU/RHj+SWn3AFXcz3IgrJ3DgTWZPFD7K6KTNV9bil3Lz68A
wzQ3rJICNJgNR8SNlDDmXJCQdoKa1J9zCO2u9lMFUwGT7e3Qv8y3KclZTkvadHuKvgmmjn7ZdoDN
kzko9Jcajo5Ew82P+PJhC64FFWfRi4h4mmG6KFqgqeUzxEBCasyEclYUacGqn5FS5c6ZlIaSSZTz
raqa4nv//Xar0FE/n5bpDKZ8RVBqhCcJaQjLfvQJ36eytsfBNoo/bYBnZjkbf7SOY0fKtA5TIDVw
JG9ZTHrdxH/0j1K4DVEWB9arSFbWFd6M0SveeWwjx/UQhUFqPVgP2VDTw8+99pPrAn5PE41dA6F1
sZy3xNXWdJma5OkFSvIhdZrsVNF+s9tD+RghQKEWR8Sb6MuGRU8vEGRd435k5vk7Hd1KUgTAtj6m
pxsnD2qOrptfceITPUFhdEZNDsMU+mcV4TzLLEF+2Vi424bAoDiZ6p9YRWD3Kmav/QcUilyKkHGf
sleiyPgowTYFYyJzdxfaKvj7ZKPUMQfBXlHA0HNZwAYpxXO9gnKNDO/Aa03UTPlUiw2BT1GE1CvS
jMpyQ1L6kkNiaN/SP0pdzvY9uCXpXSxIaDT1PCnkcpeOiqvLYw+b8RdetVkp3YvftWsRt3H0NGMU
Z3OejX+hsHSCDYKXrjSawLIzz6ije4riXHMBK8vOInLxM4yMAN4+QEIdC/Dj+PDtyY9zfsGhZqsl
rGqnSjXtDuxx9BuWbnfSb1N+IVVGyVKWPbNA6zLbnCD3hnv2d2cwgXeQZsQ8koAJM6wVBDrQ2wmC
gY527+WzjCFLJqyjJjEPJMQDNnFDTzQmRhqKRv7kNc0cqYzqJeS/bu2L3S2xBPZmsM+yzDhbiDLN
aYiZfv+YP5StyBPnBqb4+QvRur7UrX6waaVZMwd1seOqVN1JvjkJHEiEZ7dY8nr1iPIDodAOEWNm
qRMOra0nfX847TwNN2mPJVb3q6kWWTOK3wtQnfsJoI8Tsn+es9jl5C4t0HjkPuQqvMrpIU/Ljdn0
bNhx5cijdB9nCmMiY1waAE1Jp708I4mOzkoe0oe5RGdFEuvB9i3nISaWCbkat8daKETGoxVEfw91
eAMPdMCC0GsZ3kE1+TvqXVyhUpXo83Cb1TAxA5frxkGidGMvJrgTDe1K5p357o2LeNURePgwf+W5
IUwxH66jaoh1/pURCcOBKyjrfW3EY7xc44/Hj5nFGhgp5vruOMtvO6X///rGbtnPe4r7/thG0xrz
sT3UAHEDGRtP5Xp323JJOtbZDKtEiXx+2eow3uwfHBLqC+xxwUl20le0OSa5IHlrUp9GJYziZ7BZ
1M4cc+xCf3hJKwICzWeSNNorDuBT1EJgsRgkDqvyhSLe/xh7CkNYN5zzydWKDApQ/otDai236Ren
v06hl3sGYL8/hRFRwxvxPVOPEFqQDZfdkQI3hrJPP5NkeoBVIc5yE0jJV3f+/sVK7SQ9ccOKW6zd
CjQyaoZv/zhPhYAK1tWjqjY3rXqwkROb4wFhf5alTIlDiCfkJVS14kKB2N7S+SXY6jljh9zW/fPZ
ac1kMMjCSfMPQsnnnnBLauxcAcArXgTihFlCDQDSierKzC6if4HXGqGkwFsM6SGhDz5fR//jEfjX
mbhFiSWfhJ2PrLuKk4vWjHuYbkADjEfy6P//50ljue6huPtluMUK3+I4etdm2eQwwAJ10LfJJhIv
DIf/qwtc+tu2PsnYnCIWxUsCfMmRKtQOJWtDAo7EuVGyqcs2xXu0cBB/XGnV0wGF7hNzymOpH4Bd
rXlJIBYQ36pRjGZX2vk2xBt/78/EKkfwSsy95zR5gZCu1yAMmUJGcefdGI/DmbUPxn89gws5qoKP
cwfBfSouVF1p/z3Y7Yf6ew6WmWIxZOOPjMnHkQdB+MLQ9gpKWfARdXQuuTbZsIHXUe3o3Bw/mWsT
/5HsYrIgBm41m+xoKqAP1yDiimmfQWfn7hAmXLtv8588h/rB366nsKuD4L7p5DN4T8NwyoM+7IUq
95mivl4472su/yxqNe1DNwhz/lrGC/gi+0kdK2jfhrxH7kZGBo45q9V/pSepvvrEFss/ErmgKMAn
kodYioPA9/S/KlQSLsmyCc6SgpDuOHM5Whj2J2NvEySOoOfSrzJMfMpZHBd1k5erjygUh1IuKJqs
el+eM3vootk2FPo7WpEa5l+ZBPfV3zcAjDZbb4ZTSttG5eKcbVXi9NXNCUhvYWOBId98tsjw/3sh
AGASFXEtXWO2BDIXSyLkXiqcVA108Mhfyc3wanrSVTQr2H0NPIYssDEED0Hvx3R/MinFs8x8dIao
weVPPDqLdyp6d2QtbYcZtlUPaNfe6IdrWSP/Laip3MQBWd19HJDnzij5+bEo7JoLMPJWTGjOlDA1
bmpsnmZOjymOXiFvz0NCFbvSYMgLAehXEY00QwvKMPXeD3WgHpFaFDJS0z79LPGYUILKRWY/ZB5T
5vgjKtVCBQbhwYDbTIX8xAMdmnnhtFT3JU/C8YQuEYhK+RrlZpD+08mq14d4CMfUCkWwDHUGv2Di
kKW/V1O+BjkbflfFe5hEE6tGiKvk5WdIDFONlMHSj6ldm5MCsKM4jsm3iKsxGYX0zegn7r3vaJI8
rFhTdxHXnHnHQ5LK8JtNaJ6uNvgavwlxzaz0w72yG9n59Gp4CtUQj7ljGd+kx4xmTuhy1avQxxUl
S7xcfxBfpueX6+QfN2MNGwjtge8vLPmkp66M+cTpoWJvPlSDqICaEC8THKiwRzyPOJ+Et/jjMZVC
/7Fn72/v24AZNGje8sNXdizCMD5EHXGR/2/yHm1oz/fdJp8+5QwCI1H2Xki8B5+DpMpbBhSdBsWO
n0YkZSVTUMw33SlX60xBS/nyicyVkUYd9P8FTfZuq9NjMJ3NXE9Q9354QCXkYqqXae5OU8ZEU+pZ
KKcLrxsLgu5bwHl6zxs3+oAEun2Ay1DKUTSOb0TAdtU14Hv/Kb84o1wyjL7tlGtvy0Bncz8/6G+A
MQDOIw4JRdiomBbgIXPvgpi6xXxuGY8i+rLtjXjJAt07ljsEGfggQ1ZRA5JuZHUPt8e/T7lWt5Jc
W1qdzIH2uuIRbJvzns0RAWBn7Mc6cA87vP+YRCLE6E8IN3eyqUagLGyHsZ80084wVUi+JKfbME3s
KsigPc/9uHGebL7bJ42soIt5lNByMl768dfJcf+k6A7eX1p8+TqbeMIks4JO52zFTUBXJUL5zpFU
vik/A9Q/J4cSESAh0fC3GQQQFxeENGUCPq7Q3eWgq6grNCeLL0x0mu1hHRw/HoR1qB571DhVlNfB
Ud9rkn7xtY54yVAlDPa/I6As2emJINbDnbDTb7e5LzVvpAef9A0Aj1wsVoABR9sss4R7mjhvozJZ
HJpphbFDfiOlPAeNEdWCd2KWmykF8xsq8DhuogD5AcqxS/fi6wiB0lBaGR0KnoA/oajyno8a2ZZ4
cB0fW8Wirh7o/lCHVDGaWbFcc109Yz+HUo9AmwvM766FbmDNYbWvSyVZ+j1lwsjzvON0m9TKixbP
V0uOBI16/Dad93zAYGfbOBgGPcrFgKoFSOKIwdKra/mw+ZDNK0Vj7uwRTYJaJm/PyHsblQV8WMO/
LGbJWqDhGBbhG2Cy+xu+N3R4C8n5yn1uftLPIU+CMlRzcwfjYghLn1aop4PJDgHWpRPFqcuXxBCg
GMcWl5A89TNuiKSWE2OQM5kbqPwkrDKB3LO7HK++gFEKz0Gqui3wBFl7ZtllaFUbZUYkyHIr9nj0
F514fw9CE0Raej+iAB/WSd4bimeXidVgOg0vOruWZywgW9ZAk9Lm2ACXO2Zkbek7SywSNTKa212o
WRtxC75+qQcrWiDizGfzN0XTs0d5LmHvx/e58rYYNQFgKsbI5Tmdox8XfGzGZWt5VyVCdVuo+nOM
UscgdiVRcjvl6dpGckwd9FtvJXGRKqrgauHlm5HVJkL6n4xElImr15g9A2fKck072fgKi12/XS2p
50qx8eXSJxJZA90EQFFRPvn9GM14QZOWAQT6zDKCImnYGc2J8PQPvbDZ+c9jNanCxqO2RjPJHz7n
L0o3kFwQhdJgMPrwXKU/SDbMr79//0x8XSlpoPgKGvPsQg4uG6mA2GbQ6JKpjzUZx1ub9DSH2Mbz
rh+YrqDUnza48p6HW+GceXP4hoyQW9V7B7tYumC4O8FRh0Kv7CAkOnwZVc2uaVBjQLaaQOOxLw7P
2NCkjzZ4NTbKtD08brHCE6WR9PLNG5oFcIt4g3+hPBI0hGykAEuaChN60Eeedk+jzks6HpGUecxz
oxDj3Yd6Lm1kSATd1UW9TRZNAqs4hQ1zYxUib8RUfUtZT2ZQiBdsbvg6+ucc3u5zyErlhLdHQNDv
2ZmmX0H1ojXiMvB30p7QskpGXBJP1rHsyI4jP9IiX8r6ShMB51DaBvK+kAQ07FpyJc6Grs82OxdZ
Qk0496BM6omyQQJBxb3+BQkP28yOgrCIws6mNYIf0f3eFoWx3+djXhuaUN/RE8JABf3cYmFrZ+fU
25FLvEfvLZ2YrVOLLQ8YRJSiz34yG3LrvqpZlyPSTmYxikUAeaVYRBrY7VZEMh1cviAhCF8ZvOf0
O/0TDSpYH6QIqtO/+g3jE7bIGvImRmGllodNowhNj68WPDCdBawwK8sJrTUydHbA2IwiCtEkBycX
zkrWpoqylhkTFcZqzJBjZXKyBFJoZSI0eYqGUcIG2W7a5vgQkoSJyripq2Di5S8JVVKT4YX7cvCs
eVOy5Rjo+TD7pZuViJ2R+VTKyyuRUcZt7nvNWvV4rfBX/5iQ5qIv2eKXrsRmNQA2P94m6ihwdYNX
YwjHR4XwsQ11twlgqEg0y890q+1byn5QDTa18J9gfNeaSgxvYkygdgSjfjot4mWR0nGPaE8oL6rA
0WphSVNj4mUZ3UMJyo4UfN31ZrnqlXF5Ppu7fnc9tb2NJ82Q9aRW7OF3kQ4awgXyR/xdn6cVwXDD
LB5C9KZfJXHfrXOLMqtB/Lk575IbtX7Y4gs+ttDrVJFp++nfTAoKAPHBXfPfKj4Xt+uFgVvW2wm4
G+rU2ZspBE0Kyp8rEKIOHxgMIQ44qC45P9v4ou+qi5qmr3Mgp4EAzCFKGuDI0ql2STUvxphTAGxX
sFTGhCDZ/tCq42y0JBZNTX32aXyy7Z/GOZl/FDezqxrlP8dhitrTwt25TrRxFQMrAlfXuZUQWDKH
s5pU4dx6CScH4kMf1CsQmFAsHsWI9A7SS9i3NMQtk1FWRXfQdSSiYx9cAgokSOBVxTKQff/l6nEg
Y2Fs0ux1DtVWv/YeU7iGCtebcHD7xWrG3wOE+D5dQ5ffpY4kly/wb97YUCg0Xz3z1yf6nQy55ZPA
k+ieF+QANE2p8iknXQsQCvA2sKFA9qKndtGFbK1uJNuVkJINxI/IM+NNhPv3wANss2LIujr5Rf6d
Wky9BOmQ0fz3H5t6nF16Kda6BOx1vV5QfXcp8jKGKa3YQNh4k2zIGgC8IlOQUUo6TnhoQHr9HT7b
MtG63E349zQOIYxxUB7H5d3nNjuRnBygSXTlzy2QI8G/SzZClOiVrN6WZvFb/jufGZo7xt8/Jce8
XWAsPVevf+rYwP379qas0JTuEK806pjvk4/daqn+HAAzKs8YGCpld8ja55cdokx8m8H+/CYX+82G
keKLBnWXvXsDpQitDmeGxpt2lNGqFfAgqqa5E/vWnBYTeHSKllVJ+JnsV+lwbRrXcVUVpKLAgXVS
4qmvS6vtlm0fYbLaPIwBwCo2QirN4ikZcdmy8vhhm++C9p80/9p5npxw5pRdyRgWFgl1QGp0vZyr
UY9sNLavBUCLlPpA40tOiIkcqQFyk8Q1ozTjbtWQHGMOPFTVlWjGRgmfpWCAtv9bwwydjaz0dhS9
3PCrUMVoSG7IGWN2p8JdoF8QB9rbaAIIacOFiI6H3bE7F2LyvAbDK23pISYmeXEI7BHwtPL9VN8H
Gkb4wbw+zGEVIvws32qMQLiB3iEeG3ob1oYA+mGtv6093DOtiWeN4MsEeyeOu63Qnno5q+UD/Ozh
mLABy1Uv0a1pfz6qAFFXQtCjscp/80lZmouMbtP6Hsc4fMqtjAoxZlpccfIeDEoo+TKuelt5d6gC
OqMKr2Yv7ee3ipTG8NeJyWuzIwxvFifCm4OVdQU0hiDFdi6wu7nIACWC3y8ZRBHqUWIYg6gYpMCq
bqwWwAtKYfVyy4TdQaX5aTD1GPXmNdIQ2QJz7JQjuzZc0BrLKpAGP2wKwG+1/6dAl5kBz2+AWVKt
vALq05qtSa+WpKg5+fxDahACG4vDW68VLXklQaAlHHEWZSGXBsMyOgpFXa5B27B3RviznTKUqF3X
igbHExbcp8JNY89x/W++Jw83gawe6YbknQmtW1US38uwaGYrjtaQMiuKBFau+zzRaz4m5dZnyk2Q
ttFK+/DyNp0MCyaDPrOR/AdX7XnT2rfjefhA5Tg6kkQ1CyxMLytZ4mbqheVlE+Y20jNHK3AV1fnG
hIrw4nLhPTOAQk2sO1W7cajxkEGlIX7emYSRdCZyghWRP1FJH4sc2G082AvWa6OiegEX8tUzWple
SAX7UTv7zKsGp/SScovavF+iBOj16mpJ7/8P+A3Utx6WZFjnCzNx0+B5SIZxsFic4EpjTrbG61uN
VAHK7AmufVBKZgteUgATQle/weCfGdK5FDgunF3BK7glHsFgNVl6N+SmUzvNAQ13aP/zUXvL2gGE
4atvB+7gi9mrONmgcXEee/a08BHEVMgcTt0AX1Hc9wpuvPQlr/lof1ETee1yX03esvKiY0ZiE2u2
czsB0l2TTrlxDZ5tdWismU3Y2ix+zKh6Wrh7WqPe6m18bHFERw/yRcZPa+eBh51pvqFxHKT6IDM+
5fkjdmz28VVxH8K/a94h1WsvRIHYxT53bgrjTjQk1u/FTC0+nuBTHIXqpQqsCNM19RZhQfrO0ksj
Be9f8E9HtbzsxPg3y29hS+hFhommhZXpY1d+/2/ibPWgL1k3uWTS+GdoNFKXcv+Ipo5Tb/3kKtvd
QXbHHRY3zPqiibgx1JmkHnP/3cL4ov+HbcZSa1p+XnCMTk3J3VFPQcqaH5g70Oj8eFMA3uP45thL
tW+rVT6LgA3xKG6t4F4FnSs49Rr8SGhltl6wL+nSTYqtECgf0160iq5OUl5YkVGL0MRGe8obK1tR
KKUTREwlsMHK3H6hQ6pKoyPJr/X2w8CFeho0GC1gKeUtdQ6uPiLJDiNEDLU5E68E3VT0oJns79sG
Zg20vyn09c5DsFz+QWckRsUh205lJ+YgnP/IN6BWZHfFFmL9n6jOxEqskRXzYePTh4JZ9zrV3ECO
IBzGHzVAU0cyCiCVA1JyTynY7DlVr5Wnb2/pvdjy7CzOwTb4gxW3m9fiHA7DfH2KnCQy+j+7sTq3
iIv5rVZgH4nkZTGsdIoTHkEFXvulH7MZQyLN9G/lTpALIFSB4vHG6Sv5yuUp7BrLZbxxQVrD5zHa
shFKCF9F0mBDpuzKtFVhaPwQ7cvUJ2RBFcI1tRhdOpcgwcI1eS+93RG9XUrQd+JLq8GLpdnYzC5W
4kP4Z6lBLSeyr46QUWzJ8pqgWhuFie8VtnOuFB13ADTUE0Ew8aA8FjzaBAWnyqJXfwkj3X/22b4n
QcutoSqMDFDyIrmex0a6qfjrFe7mzhoO+jRiwwa20Zx+gS00WKpv3d/a/chpiSl8mNomf/7Vxoew
1fFr/Q7O8xClPYSqc62i7WHjphkhdk5KTlrUmIpgU96+EYf/c9cCKw/iM0aOhrgT7h10MLAFTlqQ
hV/FRjlXVtGNHCfdiTnJ0zbpwixX6zCp3jo7o62+PJUbtiyYgAl2oWYaspHhZpjBOsEkutR/W/op
DczPdvr6YfFqa7Vh3EwdPWSIJE4nN6R8MmHC498OUrHJOpqBXA26nIQUJOEZ4ERxnx2qo8+cJC5J
cWiS6MtmbAU/3VzRXMXig1H1RycKwD/VO3SrqjHGlLTMEte5wNgYMwETymKxJnK5qQXgAc3Qm+Ow
KeFYbl4Tgxpd4jUOg1cjLqBwWFPe2204SrYk1bTjbI5TukLpYTVCCZhdFVm+jIXqYmZvbZW2mEh5
EN5Xn199fxGCtzG/6XcG0oOAVgGzosCe9jpfjaeaep5Azv5gONmy5sC3l4o1DcaN41IMA2IIaUGX
WNu9ua0gEqVSp1C3qH04ck0Uyw0RaulQDCDIMqosXs/dStStr5aj4kZhVd8UODMmKV4mbPwJ81/T
9NdcaBP6M6V6Lf/ljGXyXFjwwE5S7xoEAu/MC8I4MPGwDVMbh13gHeJtQcxYCz2xUMLGLLu6b9p1
Lt/CDyRrxZxxgcj8I4gQr9mYeHBczO6T04V3qKQQ+DCyHIUSNmp4HI1U1YFWkg6JT7ygUkQv0tvq
WE5ps9HEL3so0tKzuYnfl1eOyC0MiOkb7ZWFPEtK+p2JmZgnvvtewWWU5NjycxmWOfXzBXmdfUFw
vwMYtwq+2rinh5Wj8Wr/NjvaKrt5yM98DA1VNdSg1TdDf1PadL19zcUe5XpC8gYOYcdNfJnaRAp7
UZJWIvB+I8rPeJ5IHZ0In904SQfOrJjfCnB4YG8FzcNHo46NQ5TfiSsL4n1HAcl19mtuUz3Uc59N
xWOqZmzrLPimfX4Ob6XdYVob7xBZSJprvSf1o4LQ+WMtnmLGL8HA+gg5Py4QuEWjNsE4dksaLXaf
t0j8+GjlXDnKdj1NNyrchx+TnaePiWjC0bsYj5ebL2pPvCrSTOK1zVz7BG3hw0bBCRrb4nhq3v0S
gjWTA3xdhXp90uD7m/GAZ28AnSsnktn6MUWLPDcjyMkbcAjhPg0ocTx/VjBTmcUZlj4mddStZc/f
FOJBesOAvTRbudgKClWwrPGLaDyYugSIEqgYQ0UX5XZMyze0ul5jkxNUOuNBBYHLrvxeU1riS9kz
1hRNbvVDqDNVepW+Nz2NN5u4Z5wC8OQL2t/rDBpnxhCAlWwcbJJyoyNmoduw5aZKE3qEdFqmL2JF
ALdbDuwKXhudp27vLYqcWUxy8xstZ+UyyDNyn5VKo6JCfTHahpdD3dB/A/C5z+zJYwV80IhJgvnc
tj/2AjsEUyEeHxvsRzDrQsxF9+fK2wI++4ZAb5h8MnWXDnQ0Q4UGLeNZOGhhES+Pep8ztIXXp8YX
zOIPDYl2w8mPqdQVZ/bZWwZl0od/1hnOq/zYxgx4LXXqPbg0mxI4gUhIcIra0zYuKWKGzzf2RNAo
a8nVaaRzT9YyS4fvT5ChBatvKc1YzAQGujfa8y/yfctrQ8eqRonj1u2v9tsk47WQ+DzZEOIlmTYz
cs2W72H05rL5sOTA5pHRCQ5zlVnCSJgpSNAEZ1vF5W/QlWNtq6Qmz4H776M1ecNd7VqmIdiYsEIw
nhyEM2XDGbdn+k7ufKjOCLuSm8FT1/GMCB5YRwmTwkX68ibJvHC+jbjeoEHg4lqprFkoD5hla8EA
y4dE9pEzuC284/QZpln8c6/Z5b67lVvFKe1USFm1HNp+z5aVp7ZDLNGEzXnTGy7Fp8DfteGejX1C
tiHW7m78pzrk4WBO5ov7zBRHGZuQ8PZw2PJlto1JLlMSwQRSf4S/bf7J5aa0HUe221QuHietqIS5
0TbMYXjq6gJNImZBTQ9lXZsadZ2jeQpIe1YUgso62x+K1EIqFpSZnq5svqvUhmdASxGMAQMVm1Jt
PhWHh9aggzU9DkcBwLe/sxJlXEhau7b2tC5Q2hI0Ql3kZ/asrwf+AmzmGOXxSSnRObge95RsnC8Z
DUQhnCGKBkAVSxxOkKw+SOGvHAIEPaNQM/72AWc4RjA2tGPnXIoYaa+GuU3XO+pd+egNWRRKu5Rd
rGmQoE9ycSmjp+9TWBh6W89/CrXMX3+ngzI3h1qblxbZh4sJfKoFDjc3rdJkew1wZiBrpJ55m/C+
tqGG7MtsCxXUmtoa4L5gKPRpTOiu2NAIQUBaWjoAUIBCG2Ka1Tp7RdT9g8EDxT5aSjGvQFZlnyaB
4d+1/1s1b3kDgWvtQ7rxYzEYGcugwgv6xYkn60yfkyZSxK00AG4p4UznNMbmeswhJpVHYlRfuYuE
i3ASwhZn4LUL4mbN6o7VL+Xq2wcJFntB6chuE3vR5EqIcsUhm/k7z+tfpO/+M+9OhOn6XZMR16vj
4E68b2Y1+RwkqzcwaIjyTqmjRT/wqjc8rM8DlZRJ5IeTBuPSB8kTufW1PnG6OWOIOM5V2YUmw4jJ
wE0vPhgSXZYgCo6FSvNQIbNPZuAW1+3QAbpa8SGKPbOCkVyT0AIB8XCHjJwjPf0jV2F7b28FyoKh
ceZO1g8cR4/zqKL1GAcWR5HACa6fVpOvnFXGMRGkHZOVaTuYwH3m2+R+zT52+cyIaE+W3M3jBhXh
C04SpQj9Je0dQZ1mw310yuloxIvCDFxNx3nfpCEM03Dm5d26Am9eKlVt8b2Mx0CO34HgAN0/AMKd
gM0vz6ue2j5pvCS90jhVdew0a0M3tj09sAOKVFh2cK3ekG3igOueEtTSkGKoB4Rd1XQ+Yr9BCkr0
UTaC9c1vXPFKqXHixUpxCjZ+8B4wMGeHGL4eTaD/LGoNSQ7VFDYkPOHZ5HbcXVwmrfhrlLMNSUyP
vqI1f9VipOzxG1mS147rl0FBvJA4WpX9oKSuAPy/pf2nxSuFoKwtmfKWwWTkBIJp9kdfAVJ+8SSC
0GDjUAAtB7c7EaPO3bdPHTH6YvN4QpcRHiHaeaHOCO5vVTg35ma4I0BUR/F5lYWgqbuVOGelFxQX
pNb+vT7vI0rfQNLA6zUIpm6FDu9M7OBRkT7lP0Mnx3YSKbbyBHvb7HGeWApk5VeiCnpnF3Tg2QM+
QgHnd6sM1qsr84TRrohoMdcYN7PrKGOx0a5lARCqlMBbQJZ80BkH4Ds1RCEN0yghNpIdjACFUE/g
uSHL+hCMvSRwPY0mZQq78qZtGsczrcdCPZHWUgQz48aekDgWAeuQpmlHLFv9C3Nzt37HO6l5fRv9
DchsXCi3A9II7IybgjzyK3LNYNW8z4eN5K575DDft+9Lw8jGG/zXW9lKlLzTOuEi+wM1MQq8MFbS
zarz5CA/asJhWZkL6xaRy/+iv8hYF5eGs4cQ7q2FTsCBsXEqcdXLbL612ud4Y5Qv8wBjcaw/2OIX
W93+MXgraN4h/DIgAt3d8TgR6RGqpLXbSgxVY+OjShwm3D/Qfjw6LFHGXklLHlenmHIk54oWncF7
+pNSQHgrhK5+y0lg5AU0v9tMyIBNR24PGIGQhLRltk46aP16O8ZfjB+c+Mo5asGrRAFldhUX1Pnb
PkRiqmSh0c78fjoAHKQzFUbhDHba0UmldUsGdxr5TtVA6XwgyAQ0QkOmnZsdbcEXeoAFkdL+b/yH
+gZVXgJ/grshIR7V0zpW5+oCT12iRaFF41l3y513XgmT8iKM05Ul11y1gz8PZG//E6Hlxoxhyt86
rD3TDVeX5lZX/zPX0b+hY9ghhK8SVeoE0pvRTQuzNkW9Facpa0vK41kZ3WiacOcZXzFCD1CkrMoF
54iPfi+7oTk1Wu+Z4fKguGXviEAoaBUQcbsHYW8DsJ5ddKvUMAAysNP0MQe/RBPs7Bmrqt49lfhK
lwCV0JCW7OIFzMOzWLVxjmnWEP5wpaex+zPnduarsnRVSRbmYkM+nyFXut0AUXNFcsDpFxjGPcIn
tidu4JxOFfwPVvDotNoliqAwcUN+/j+l6PLhkmpYs2MjP9eP7fxu20q8G2Z9omDiWcuJ/XDXZlJN
3JN68jOrV21YlNgXdlqql5/LOiklW91uLwzvkCTv3xjyxUl1i/7//ch260XICuOHrVk/+FSGCUh9
qil5p+lCKj9GAISY6iKRIOpp5lf2YM2mj2Vb0yk7Y0KM1Q0jTdv3vgFO4nc8NSzWhp9pDb1CqtG2
0m3VvVdkX9CTAt3OV96CahgtMBapxPxYkWCDyGgYBLhL5m8whWa67jFvwlP20m9cCkfzIMtzmZZi
hALI85ONdATsX5Wkv8/lGT+vYKZQ+IqItGDpz9GwhBg9xwH01LymyL3K4jZo2YwBV2qFGEfUwhOm
S9uu9jNzsXM62FkuQo+v8lOhRbmCza5FLuaBRe3efuAo3LNYLI5R1Xj42ldkPZEpofjxqqSSeZgM
g+BFI54Dmh5kI+IrhYxEXVhFElgJNOJSRf3UiJtjz4BNMiG8pOEfwUg+rGEKHcdOR0NZSBtQ9Io+
AW/xIBo6VGrfYzYI7rk95c9dMLT7uowOVL3utth+SJVB0teSegQarpzkp3JkmKwRShIMjCukFyLU
5rQvX17D95mkhWA78EGKtzOfI/ozu/LUzLR5uaNdSyMNq1gz3Ywv5dkGgUTgZFUMhiOm8pqy7swf
tesrhDejtUFN3Rv1Blfx3CspxhI/LFHZhPp+v5FhgLN2i1C5PuSSbk2Sx1pAMdUXvM3YeZLw/mfh
1EamjoO/g+NjkGw3I6yEXMshPb+sEzctXzrBmiFj9iyj3NhP6w8rJD/39Si8FcE4GauORZtyAEXe
6m3iVOnUNQFb8uIZwfPQYVS7SuuWp46CqkbUehQvZ4cef2Vrdri/8bRB4YmX+5QP3oLa6CG1Ltel
7ugs0i3OiUYl5FKIjm6W0YPxa7CyBR/pzoUd3xeDDG41hr4Eo2YHSpytGQPXinHDmFsH6hMH+0xV
bq3GaAgT7VHuLFH4mXgGCPB8tAbnt2xWMUM6VFzpy5D73MGTWkU9pT5B4MRicSiHH33n2cuEaDl0
LIJzNR9gkoqTeodejZIHfj+IHBUFVJqVqyDO5p7he3c7khwe8/F/9T2YWWjol+yKvmXWtOrKXCJm
AIUzFB90e7JkqtQ5fR4hTOloBHxKhGzAiFWfSR7ELj6RmDoSMU/FT+2eYwsNrT2jQ6p20Vdr6HOj
smiLc+hQtQ1CHDQ9mn1+QkbHR6pFYfd00woIN+Xj0Znsyw1H1zSc0EnEW9WvYNWDT/S4aciADq52
QmdbYaD4XqLj+L/QAF1c95wph45BjaSafbeR49NTDKOuP3Lt5jdg9zPR0xEI/d+zsi8lGscTwTG2
wVdsUgHub4T2191rTzU/HuLbFCzQe4/pzM55V9+amOxIbv5zpqccmbhaVO/ra3w/yrIsYvstZkq7
7pejLTrl+wZfYZKkhxW+xiXnEmNky4IW+Dgwz9gt8hfqIMk1ANEpiAS6pFov7KEeZMTX6JhFsvYl
zLlkSxM3Tly43a9Fo0TJXujQToQpcLhBh9zdR6Do+nbS5ZJCU/8eWIJURhqqfJ+8SCW1WHw7+VWE
dwCCe5jtW9h/XVA3y+h6g6UJysWhamfoelKxFnQKNqhMQlfO77XkNuLAbdM0vBwuVT6zbb48VsUq
l4t17AcrvFBa9anXnD5otZhmj03MnYzZEzokLfPQyfLclhya4I3G90l/gx0C2h3FMOJwwRz1Y2h6
/CFivOjRRxLdOWVvaU7I56h3Yz22GKHoTmTWOfzLWoijq79/jdsdFbDO5EP9/h9ZvH8z+HOWdPbO
EBcgJytpiOgTNvbHLvfObBvYlNHvasa5TlzJjwwCR1bFWj8gZhvdveMirJ72dH40dcxAdlyDZsIt
aLThxXHcPJtQsiLnh6P6YHwFz0P1J+nZOVEW7XDurCa5u/IW+qeMHyHxEZ0HC6QHzhNsYhq/teFZ
Jmkaj+I7/zXwG654fDLQ0MzWuVOcj4/qgEu1MJ8thx/0zVz5JZ7NdT/EcpPdgZVbO7zEO0p6hjEn
ZmVOiT7810+jYREpqwym1ZemgjA0c25nVtWZWhf93vb4MmInqE2uzIiezgc5UjITHFlWHZYkh7JY
Ynp+oMVyMz4hSkjsntlUPoLLPegkwJcRPo6X6pRwsBD+1B74ZUObIWOtaS+uvRdrVrXH6xTFLgwL
BPkkQJv7KQ3uxrjln8eeS4vM6s4/cS3FMWMfiZB+Mcrc5KQ/7X4iIC/EwVAbPsVEC1h8Vgi7Tkzl
8dP8H68ISdG0/EUXw1z5YXmGQTmNNNonur53tzAV7oraB3Y9wXX0B1ASkARD220Y0eFf0SAc1oU6
n/OJfL8jtv0sTErfmM7zuNywoMazjlSPncWNMsYv5g7C/d6ugxOBRs2eDjIu3nJpxPJzY9tNHOSv
Jk+wE73jtVNk7a7g8qSqhtqaYkP1nLLb1jP+PD+/3AK6//07+CJxx5SHtqizdESB3WZeVidI7XpJ
FFlVOrd7Carn6n+cHC1BwEDNN8Q8w4Il2/WY9qgm+/VIpBf9OCNwJjq3e0gT5uDljDK+OWAtFswD
6zAmJm/gJs14iSEGWaUA7icZ+SFs038MsoQDjgeO0HQ2dr5JAKYTtHBDAaBi/tCtRyt2ZWP5X1vW
APB7h6npxeePo2apw3i4d4Txlslqbei5F9f1sifztc/sto/QWJcbGOLcHBh4d6L5YW3nUyoSKF6+
JBDClXS+o5+IlKAn14Rcnnwz31HYEm3RQ9iEkukSQmhVkBq/2yxf/WRBX4i3eYazZUUFIEknWBzZ
oEpwhntrEHdRrIPZA0KAl6EI3h7PwzpRocXeKdDFx7jQqI6ArEgt5dv0XHnfm9hqtY6kwVLRRNJy
mXV2zM+h3vnWMXBtdueb/WyIO5vigSXVDBIJkvqzbuyAeYgRxclrGKC7FuFHn2ZM9SiSpbXeIx/0
UrbEyZqQKH1LQxxlewz5Yx9vH4Ga2WPTpyCyuK9Of8Ktn3+BfUz1S9lUVnVsPHZpPJTL6G7SBDQj
MiUASYn391NUnlafCoqoc5KWbN1e/Ju2SVMcz72NCmOrCRa551fmfhVnZCYCXc7Ou3UIiZ6++zIM
tDRpZitV7GMERb5LYCIDz/e2ZVglcOULXpiNyZe7wlDgksamH9SlfOdTSnTx5eA3+VT6DKsfUWR2
LpjEthACo3gHj53qny5ktCNJgCjR39FfpfuSPEpdeD38zauRQJcoR+0/gbPda3aNEltrtqeZRKJ5
8OWCi6gGbII45qwS+XHXw/aFT8Ybyj75euEJb2TkosEuyDCdE3tKq473dylyh981d7MDiWDAX/zI
1Hjtgy8QP4YMmHSHCzakvivhl02M2fhEmiReF2jfnNQJwjMhkqwKzCXdjDQIZmPJxrnT8as9TIff
X6q9pg+ApmKXi0nevVQeM8/rOulMPrNl/KY212AEBVGeSUxxWa9kkqrn23dpApqOmg+QCLGsoRXI
Yzt7Cn772VakazxLBKYioX9H9b/zeJPgUC7tClShC/c9uP9NyoSXicz2cdvy0o1hLnfK0eOm9NH2
wtGXC4n14gbQNdptYbDC2AEhKnBpn3axi4ibf1AwnGt18F43xNNJf8WJDfa9Scl5FfEvVU6VaKyv
0EvBw4LxsU+pU8Azcelf41I7atWvv+PKXLPGU16eYBUX59oLOGIwv7H1NzkJ2yaP+oeXN93wX+Es
9secgfRLCfnnY8OlOHweDK+R05FczCO7uXkv03lL/xw3gzRtLpPtNezkBdZwni282D+8DJtTb4m7
qOjd+S1xyzNAQe/ElDG4VWypAYQv6IfPXOaMR2xco/FSVMRv1RChYyvVKh/wQMyvTyfXSeWLhzhf
igl3hqq04v+/eXOEhQLzCCvKjU/wE8K5z8yqs1cQxAhYKxJmBTbLcuLbKZ3ETVxyyl3KqaLr/Qqc
apRkiQ796WzCCezkS60n+j7vzHtaQ52fb9561ZrGk8JhmcMJLbPo8xoc5i0NvhJtB+EdaR00ct4s
aRe0O11r71cWOahoT6oho+FoPgYmT4Zr6eyO4I96kQcjlVTAxGqGKMh9hP7dqLQly7/EmPSPcsxf
1upCQPooIa9fP7nXOqhq3b/YMo5/w85XUSoRFuSXO8PCu0CRJWu1a+03d/Kg9pWyh6wdLQ5B6p0S
PNSCj30qvqxO3JgRLbGHVwypGUeNGtWg1GEl3CWXSNxEqIBYua6qKq7NL/OGJyKvFb7CVdcCa0f+
qEav7Cm2SRr/9IxuX8JU/YAnC8aptWVN45wM+gE3CcLJSGkxAmonE33I8QNWZbqNEhU+43o/4U8H
7kf+rT2A4Ownk1V5yovovehFYugR5+ZlPg5+Ks8tGudfYDUobUPcKMGJiKKwk9CAoP6f7ZSdLUO9
Y1v33wRFZBQ0VsnbybNLJ8XBwjoMDBTTGfpWp/jw2FAZoMERPmO35B0XOpDsl9VtxdF9qJ1GHgTP
OVXb/hFKEJm/ffUI7NyjeGaKTTIyGhojbhyH13Enns7q4ktkh+1vb/QuP2CNBSfGoW/cylV1xxRJ
xdd46Lw2HyDpUhzmOoZCRRuAMzE2EBJkijWBGFFt2ZuMrTh6if3CA0JAyxdMMGG5CETrowu70wci
7BuJegHSPP1XX9mZzkd9JBDPX+kZ7G0TYDg8C40KIWiD2Brp2Yw6nK7Ah/sO2dJhpiYvEnsqZdQN
DatXtmosTypyRA9yJu6+E+bM+4+tz7bfdpXSggpFLLfO0StDhYYhju06qlW6ONp3idqqUVuH/iTH
J0YkjluihW952toeRTjr9bwG2vh1Ja7HKisAIJmvF2V4pD6XJxMVt+3tGZWBPoIgG1CVoD+xOz4F
KGk4lmCvzzAOfrWgW6DyjvP7tXa0ojRe7VxSOHEHpEIzQkQNz/4bj+lV7Vo09BCsCyn6cNR5Y7p2
X+uZAoHJjxB83Do8bpoioa2bPDABg0LhIapo8lDMh4UnAaqn016klqa27fjjA4+fysWWRXAhdj51
tYhfj9S7hjEcVF58Wm6kfbUlURWD1l/uaEH8ZK7Bv/+62IsZUeBY4oj58I+AMWU8IpSwdcHsVY4Z
6v6oS9YdeHa0qdrIGdKzcZ/bR9pn6XXiDlGcqKkMVaTbGf/dYD3r5vv6Dw7U2Zt73wWgUNfUedJN
5twtZo+Ur80pvEl8BsGGCuEyOcc2KGaVP0z/XSehI+SoRZZfz+aPQSV3IMYeR1+2H4DgE3GswJs2
NtfdNl+YRdofvbYq3LsTpTyqjGCEQ8AaJD3CD5U5CHuep5LhwPWaAUnHMReVLWoAlNZQQp6gT8Nc
RlvUzgTv8E9mr82n2vck4pRqozfz0ICmG8vleNy76MNuYP4+dh4FjXx/QzbOXORsKrbiwQrP0DN9
RfzUvd1dnkYXpB9a3klL/1goJMxykioB6ykkVlbl8EfzSYMS0T0uiyFIwmDyS7jCUKLePu9V4pAw
8pKx+Gf4QFTPIaWVFysdofdVeMG2Jh3+aYzq/J0wtKZ5ExJ5+ejFQ0b/blxA9Wy1G1ut47QQhqkp
1nBXXBuIwo9lXS/9b1GHGdj1rhUDeuqWOdGVrYiSFiozjnwaYSf8GN7MkkZmetQsuP77/4gC+zDK
iFR1QNNiNN2df5IdbAtla0YbyDgiWgQzMArSMUuEwafFOPvSy0iyFN9eIvgeewdC7PXWxKliis+5
pJsfJrxcMliEXLzjpEX5Rtw/gyq28DzvFIdOdU3xrJFeOuyk5b5kWxpNm6OS+0zVhgUWLu0KL7Ud
LnBRDYivANoQpwziRrKimrL/0O4HxPAdtHPAqtK8KSwgNfhkRFgXfKtVWSppgJ+jz2fq3jHVsLO5
kgzu7bWnPcs7Ph62A9GC8f6X7/IQ02RpQNKhReskX5SQG4yieqQE0BgcWnn4PpX8Uf7VeBclp/w5
Fm4EyWDTQqGTAeDNi0AVZOoD6AheYk4fTfJllvHdxCgem6weVCsliuFOCCB3rHy6djAfaKDDSriw
o8ej/R+lEbxbnAmlj1C6Y+LhozGaqRA+VFmLB5FYRyUSGzOMWfvMm9DPZCm4TT/VcVgE20DmzLIe
oRvpKM6ke2SD+Xm9LK3Qcou8VBG+02s51d8RQqENsSFYcQQ7LlumR2vw5mZk42JzSmq9KypRCDxK
IQpcDHktPHxZDQAK47wu706gAEl8U/H1FDPchSQX5LA0VvZRPb94FAzdqDuk4osFbDkfYf0o8nNr
IdLXJKb7mdGwaOD6Ikn+/NHdkP8qoTfevQ6mmNrbvRE5DiA0XjtpJ/7LYeMYSww9mhswFdQVF3Pf
sSyAXJdswfTzT/crqJK1x0RHewQEbXXC3e+/PGO8psnObm+MDOtQ6XOn2yjSDeKUklK4lQPeO9O2
XDTOAMyQIi0+Zc48NSbJLy3Gyw92tQLLBSTULj4LRvgyCGoSDNlFnvwEyoa+KeAKI/d6leAYoObX
P9t5RTmcl11Hl/XPOjxOT9lCHexp4R3hIJZFXYK3f+atgNWOi/nBmF6E38CXqfGc54Oq+jH2hs3p
BtDmDMBj+zAQFtLtTluN7aqiO+aepvsvcWm9F8dTKcKaFst8VvcF8mBqDtGRwQ0C+FatkY8IBG97
bHwSv0s1P3M18kLmsZ882vWeEYWAMy4WMts1lsMw9bMjl8qY0J3HnGZZYTG2vDqRZunDGwkcznO7
m2z0KJKGfnmj1YT/O9oLNxgLUpJljt9/Of4xS2GbcYhSmNbeqr7lR2roczsYSm7mqL9qsnYTfOgJ
PyirKywtGExpus7ap7YLp4sM2KqPs9tKEh4p7uBluq0422Yo1h7a7loItSzw6JWZitHv/T3mqN44
YczIVn1Tq7BQdbJ8XpWwU6+txknQZ7LiXAfSiOrCyI4SJ+dKXDbVJY3e1J4J5prm5hZDWPr7dx1l
+gWcjZauRJMUZIhViPa8yteSnrp5QmM5rvsesi7PX2rWxIunuReXFoYrchampL4NifIJOzbm+pc3
TyOLlYyVW/ZI5CWOjuonG9hsstOB8A5eVFeFLAr1I6ETBSeGnXGWa7uS0uIyXWRRTy5v0V3ZdOEQ
2jolFxGpsFwWKohQKg0IZjyuwnudM9gIX8U6Y2flfnHuN0iD3V0EpmudpDBf0h1XQXLqkeQHoceR
DBlG2Nj58e/gFEGOvzNdOj4PhtwmIQhq9PCZ5F7KNCBfHjlc+MgdbFycVt42il7BKqti11pe5gxk
DEwq39XpN6QhUcqadVrZAI0pgXk/9QgjCUvvUXLq8+SabOMVWJJ4WW+IcoB6fqi0sgQAZKFoMB8J
AB6bGc6cTi1j5kOjGmFArV2HZuf3YmDJSYzn8bdOcJMbwshJXPDznu03peNFSI8YE9D+XgX2apN4
HflfGJbkj8F/ypG0ZrK+RLOyBXYtrXRG8MOMBBGA9+vaYdzPIplJS3zR8nZL+R1j/LXFKocNJ55P
taDQY9DChao2I69Do9MakHaZOcV1PN7YTIMPBFOrOpN9bWWURksoQ8juTGJLk4Vs8vTXVhFbRseF
VOaTLcXmbKc8Kcsqwfwf3/3oXa0nHh+Y4deAX2ftjtB70fxknxIzp9v46s4waQ2xaqjjfmFdVEtw
RzHC0Lm3diFVTplbDJWluBJx7ngDErVL+clIFcvlmzyWhozaa96oJtJABk2XFtbO6OIAALiJR7rM
y2oKPIyAlhyb1cOsqU+fnOBWk/zZklZfRHAuq7CCvdrQh94M88ZTr85BQ5kT3MdUmai/IUDrG+fs
i3oWVEhJuUUZ8mFdWexR6xEhJEfKUXr7qk4UcqiiUn0asymnDO3rhRGcF6uV+WOELAIN7pCmpOJf
3ZBdO7exMB+n4Gq8bPtW2SXwXDbceB0QY4vi62cesg3a4t+p6bMbw4y7/cgGD41DSNb5VndcSpAy
3xmdFh/O1RzxBnYxvzKDILAQQMHfB2VQTwpBKW3noV/X+yO5GXPiRUe3QeMI3uHt2xSjQvHAGFK3
pcz2ZwZDXShXFtfJPIBPVqXSlofDRI9lSyn9Iv88yA4BCFKs0gkqtO+sBo+v+3rm8tx/25jWXtV+
I31DtBAoc1a6IGNif1/xQLniwfOy+R7gSRCMhmgeQOZj9fX1usIvOVnV/CPqEUX86CMoFX4xTt/y
OFnRBlV0+w55T9DN7SF7U4O7Pc12prruI1nXhu8H6smvAr4OmaoVpn1qM+azs6UAX500BPnYEDU7
hNotMX1ho+G6h1GWmIOHklU54Q43g9oVBBWHfaeBqrCGsMCTvKFk+bN13KfZuIt9tolfvagrD9n2
91P26SHNZmva248/nSsmwJw4rFCJQah+rGnWJFHGRubAuTh5Jz1j2P8Z/6IxP0xNDpYgKwwMjWM0
FrUsfRBfJ5Oz4C1tXzh8KfFy/c5bwjnN3yC+EHwszvusfrUFuWOtV5gYNqoL1fQHtC2EzNnHjzP3
rdy3G+eu8Ru0/SBsFnomzVUm9Qnj63M6ti815G69/Vr8f1nPsYI9XpZT5ELzwaYPxHXeZ8WeYmv6
qVHXNIxIt3zGmQwMFMt8G5O57TuDLzmxKXAQcIJp4u58CnNZ0XRIwJ8Zzz/6ku0NaTeEffNl4MJz
E3+j9cwcoFQSkHbFBY7BJIJZ2cPwE6JGhY7W/Dx6PZKQg1FGoubYCWbu1Cow92G8hoGLTYD61ks+
CaTCdix9fhqbYWZ5uFMmf8ivhPq5w8G2GC0RU0PnOUKrw0Yarp/LK4Bv2MtXVLNS6syPlH4goSeN
aUWzLTtxvfF6RBalzP36FLi3NT09s8TWc0fNFrOE0IlWmMs2FzzGu7Piz8b4X1Q4UAskb2WvzMYg
L/1AcJDtsB8NB+zl7IwKy8YQ4YDO3nyRKGXadmgZMiSTTbuuZ5bQNBMR4qpEy8VgfTsReZLJbS0s
tfvyZQKAYp5TlGe/k+lJ8uMulURzfPs6NF02ptb559Do8ChLT+jDfYIFdap7aVxUfEcYQxGp/sfK
q7Kklza2ZBzODg5vNYM/gyoKVUgbhSniifJTjtFYQDpoqclfbWW+mxdpfeppX4kkxCB2+eoFZliv
kGGwipwm2QjE1lJx619pTVQlDaZodfBrZTJGyzPa7iGWfizSGB5WC0nOHwsDYhtptnkc5R7s8gok
9Hmieg4dJbsPvuAg4AHGjNlxwfPjRDu3/EydZdFSq/aZ2JJfMpJYfkrY9+eKf+INnna6dfRBaLqp
sAu37MUvgW6QlqJoOhxAsePMOvWyvEWPrb1qXFUbIyTYizM+eQJGrbyrcbiS5KxOrth0oir2/mCr
wUfWMiqg2quJz8ZAqJ1rUdBGsOqJtC11glLCitRw1FVY8LuBtjPVQlvLEO3Dir26tB4xIK/TnZGb
DUXxpsb0AI/C3twRoh58skUaWzHVeAHlC4YVb1dBVcxlhiSiVkLd7Rm7AMkVaY6eLS+ni2gPh6Cz
bBMbvSH1J2nZ+qP1WC5L/K2vp/mR7/9qjdDcolcSdenCV+5sB+P8kgJKMBYx5kD5V2G1PF2T2Ivi
aa+DJBsoLu8906mTOpH7qjeg/CZCkim0+JiuhYjvb+SswUIlqNN8TxjaQkfyvpvWAR48ICuxXvwD
GECpZV1mRrqA+MLqJXQSK97B4GEzsrSuHH3/2pgDsox2U95TAtuhinozzz3rVA3lttN8RQtl+4sV
bpgEEg/zkWRDzQLHnZ3N/916pZPeXlFzU6UwAufK2T/7n6NJgYmJ2Ln6I4w5EVFxd+pb85CJMNaH
mp2MvpVQHC4+LhccNBqbn2XfVyBaWsy1CD6gFQ/EdtxzOSwatbfEWWxRG0lkuALRWHDmTeBgHZm6
J+j4/Y+XErb3DmoRVwi1Cnq4hElAD20sC+nl7S1sogVKDEG86lfU+RH6vCzIvXrETQL04JFFOzDa
vLB/TS21Ywn47FTB81anZZT3Eu1K/5A1efutC4Gbv6YLXlxrFK/040eo+0JxkP4TeA5OjD46G3RH
m0E7No/UcUItBosS/NEMk4qjSZgM8zbLxtHY8QSetgtTPn+RXaNkcwdq+x5JWDGX69E7UH12n9SW
rvZq7s1xrK92H92Ra2qKkCO+09/2BXAlLblyYaTxXsfNwvWewtYXzAp2hdn7pxUFKKvLtTzV5PI2
QQs/UOI1+QT4x1f9jhufUVu/I54jhgTRSUs5XsdaB4DDNJuSweMlePpqzf4ByWAL6nDu+4tBrArk
+o8Y2RVgRmpsifrS4W1unGXJc6UTI8KBNGQ95+leW17xX2zL18LjFraGYXgDexG9aspqDgFpX/Pa
CkdZcg7hsOKvBgOOwMcOjjZR2I6shIKSAZKkCX3k4qup7jb0WbH1TrtncSUEpf7eJeFQ0Fhz9TeP
l0+WrNGQlOGSQX4TolNRp/F/8pmHCRia/zTkOhMD95bjFp+I9gtkoMO28LVsYw5L+sXdpBulmdY6
qvcublWuL/b5aodshsAVOhCjD8T5bQ/GmZmRZpRYf6N9xs0EOJMKsQmi6d6+tKzGkUXliODiKD2b
SbdW6f4gBPU6Redd+Rg3YFmmD7fV1ACEsXkI1nvWDfO/8FtqjTqru0FuBC8y6TYCj7yMHKCCV7YT
KESQuxZFRhGRi6n+DCHlz668DdsBwr8Dlon/dHCHPUCNzV2yz5/E3+drrHqxNn+2DEkEW+kgdoYz
FhSd0JKyrjoTKjHMtyviZeW3Dao+nVf/AznHDSW7zIQUM4eFbFtCluWG7nJpx1LagY4vSvdnseRe
IjpjH8ShFzCJA0Q0mJoUA5U1BvH26vCyoq3SvqtvvmsGhnfLWDRaHbDQgS6Zw7FxNaRli2Of7VSm
Eim3K9iHZm4BwDkEFM0oliggFVqxMk24kbMxEXt6a3sDLlzDRVuqkzaEB1nFJZltDU62vYNATDLe
4kiC/oqtwPsLJI7JQ0VEiHRx0IRnXnqZ+VYtL+JSCEjtFJ9al9XXOCJX2xAMCzTgsysZHBNdwHGZ
u10WaYAHaFeuNpA/axyewB5pB8c4gtiAjT7xT0QHL2jZrAl4z7EapPJ6N6UBDhj1McIftBvjKvDK
1cHm91jJofy9JYzS+mSYSiLBtWT8aqTYiw0IAa88PBTzPEavOkvd8P0w/t4vLi6GdqKfLcJtM2Me
9lAurRiwGPXx+Kky6GYlN9eYnNt+Fr+us82LHlI+/03Ezi1DKIQr6Z/6n5+kRCq8K0tGg2ai7kxc
WL/z9oPbcN4d9yyUG5hdSfWMHigIh6VlB9fn3vWb/rcrcgmtESb+4kkrwAx1rCTD0706LGyveafB
J6uwYXlgPgAc+7d7mkbiEVm0WwDyZQL7oL85itZlGfrtXnlr04sj+z9lO23JRFp+/GmrSge9t5uf
2+Ght8iw/IcyuXyXhst38hsTtS7pu6PnXKc6ehYhoqYGFFFeEJTyAT7ivAYDVMeMXQxZ6qCQL8qH
qzzW1Lls+UlMk6PIfQvbt2QefNv1EaZzAe30ZNsTri/F18a6rXnONv+ZLs7VKSMCp3ThIBy9qH6D
3kDg7CwYmNdNcXryG+jfrBZSbzHeqW4efKagFocjE86HuItOoV4+7TQszDOAbxkMRsnS4Lz0B5oI
ZttCgxJKTm/Y4Wa72VO+U+kAT/LF1CceBeIdrGNCikuvjv/L54XXxgBkifHS7ksQ1HkLMdWS+cbm
rVvw9lsIhDlSdQ5d/h9XT55NbJoJc6gcv3aqWYXJfbUZuU8gv/qTik/yIk6IIT4ZdZWUp6nrzplO
9c3R4YskJ/ep4uZlA/l8GCG1HeK1z5dxS0ckFGzTE3H/uMXIi60Ho6fOu52MrDsO2buA/B/9l2QO
ZpndXEJ2nILoKVzzXSALdrhpvWqlmAgv5iX+8Bdg+FCAQ0Q1UykQqgQ+2dKfYe0fAIll+/96iG2w
HZj+m2w7IqD9nPmBHB0jDWLHBG3Aw4hLpruTBQqEVSsyPVJ2ui7AmP8YzdrpD+Xn9xcZhvl/BCkp
kw6TqsxnW5EGp/iMbpdKvBt9wylEpR3peq4WmjATq/lzbmaXGAxWc5mKo27rAXB8QWzCghvKEcoi
InU95a9oj2Rx2kMyqow0lxy1HGKwrqXJjbzZwZmtm2Z7KUkEn2MBoW6aHQneRkRHcjfAbsUmEOOw
0mWsSLQGlTtH5C84U65nNxIPzbLsjWcHHM6/fy30t5b14Iucg8m4XNJQEM8Tzl6jhuPxmd62Vmda
IQWY7xTTpgXJwurZFkbOzlBx6dd3U4Qb0+mrJlE8mMg7iFjmA6GixQeREAIiOSpAlnvBRVKftQdq
zUcvaA9oETQC3YInCM61UBm9OEocEVooC92ErMmo1JOB0Uu94dz/yGHJQCMYvspbfHsqx53MT+/V
GZVFo/Us4AJiDIeNfJHMsubopTm0enErMOlawedtHtbGX/1P7SDwNgJe0UnXorc4Dael7c+kh+Uv
gnve3ouzhrccsOS02ggtpKeI3kgrGyLimXyqkrGdq3L8j6qGDZGuHhk9GUMilOQ7r7fq0Lcj0JIG
3/izoU1fz1t8BU4WMkGYtNAkVtXlaqjNcEwlhfut+Pkj2aHQm5PgSiqaXogImBydJicfEzkzthFZ
5pSZe/kVfhnNO+djukJQTKw/JBfqXVf3Q9SLY2VvqgkdvRD+4Khq4srlNiAZeDL4azchhVlPx1Al
hMR0YF8EZCdQ/jDrYGA27WaNj+C+sOUMVWKyZZO+cPld4pOCXq0o7CQyTCAphwLta5SER3I5qzAf
njGPjlh/Y9BMrGI+gIrhHs9RpVa1Ee/HFZw/r52mvKDkQKmMYUUPas0Y8NX0o58HBN41oQZxSESa
N0Rc1eSvS7xnxzcs8oLGMrCLhRLLR7VM1YlY5BzL4KMKihgMytk+w8vNUHtqK0vShFstFCw+3v8v
lSQBTsT+Xgxsws6rBtX4937CrXEecR/p5ZgVNz+mahEcTeh4ZaKOW7tiZSymh0IwE10rYiGvhq0y
x68BLXesIdrEnC82YD1frn4QB8+n/SWvWYVZGkrJeklo+IZb3d8V3W8m2F5L/marUn0R058RT0lV
xxHsvtZq7Nd/QJxW83NszIAZqr1cET9dz56RLatVZiaqLuIEDc06SE6cOk8Fg+ocujdj8OO2UVsO
7ZGDOKYJvy3OM46mTvU02XMT1DKNFzInM1ObmEGoRp6ibj7BpBP8gdEsGNulQ6UhbmtjhrLGINQx
wBlla2i4/EzdiywtjCgtO0WFZCT/z/CdAcIrfxp9RI3vL4g2VVBAACu9CACQx61m5+LpMEsJdHxI
Y/giG/O8rxWtHzxD4ytgDF15OcwnzMlXgU5F3I3kqx8zAlkxiXv5XRC/3I3aM1mzmYuGg27stPdH
pDbsObPjLUjq0Y17eZjPKXrjyqJp+Z44DiqSdCY8QXNvlL5qA1+ME7CN8D1tlAiK31N3mSiVzo8G
FQJmi672pW92DPzjX2DD+27cZ/wwVAvCS775jEFTHVUcVhn2TtJcd804pULmw1abo/SNT6KQdnpu
3HdGj5UhBkgRgUgYfdSIiiCJWX5fU+AvnoCVCAAgUuBSHIVeE5fLcGsN/lISq4AexVQkH3AxBqXP
tDJLpTUFMd9i8BF3T1TUL86YNOTxmBuKfcCUzVYWdm8+Qa8+nRaZXjiaAH0QRT2Dhss/zuzZ2oSt
KXvgTSu0/Zwue+N6Yxl/9AVLeenTmgGsKZzRMLskP6gCV7hnaafNnQych71n0E5ucPeK1WiN2cl2
01YkvORKkL/IbiHwaJTZ4Q1+NaVRhZnm2Cu6zCbcQyIsp3/wSD0V0VEUt/EMoOfjeaNsU13fttx7
cNeFvvgzxRvCQMgw0BeyN51ZXqgYoVozed7ML+vU8ujzdQO9OCQReC+Icw35+getE40/hOcf7mCc
yy4mAUJTBKlYnnFQeDhI2Ghc9AbuHnGMSeXzf9WUy8YZ5pu8vzVI5qJC+d8mq3mw7YV6Mq83ip/i
aa96+6IdqaJ/6XToxCazToQv4SnRQYXwrZqDypx4KgzWwF8WzPiSDlLU+PPB74LBqH67pA60xURi
0XbX7vm8bvZCXuFTjunwQ0NkFp9vZ5GeOVN/p0WmSHJ0aGooQGNA6B7qJ4bwLJID1YpY1DE7AYXF
qadC0ofBIYczhOsj3A6rtMrR2zhtVuLCf/v5tu1JWCakH6hI8TAVhNkvPfWlfY+PZVrgR1dm8Qel
tXMmdNexUksA4B27DmY8+95V0jLLW/7eS8j0vpwUfpaRlnv6+WzI4quhh+hAj3lBuu2EUyEgYDLC
kHZ1u14Si5mqXY+f80o/JuuSEYkMW4FQ93XLxqP7X5Hj08Tkuy2GfaOAnkYK4adjXn/SFYP/QJS7
cVFWRGQxe6l9kxXAVJpeUUgB/wAvQx6vGLATd2PvWqyBc1Mw9WsuEJGad93gL0b+Yik8sqjTWNMV
dWi7lx9Jqy64rvRs1w8qGo2C4rpQ9uwHjARNmohl+F9m8w8MNJ13PQMlYFWPP+5NBk9kyybbf/lh
iOgWalbOcIjNyuq7AiWKoNg+VW6PUrd7ExMj/G5gjefjzHcqOIQD6RwiWHbNSL+vjJAenxxLGLR9
U/k8O2TO+RQG1YQMgT4EZdDg+TaLwcUYL06EYEVHRVhcUS39YOqS1PqYM4d7W+drKQnwx7410V0Z
T67jIST/m+VIxl6QYEYwY2B6qpINSS1DuOWQHsiC+hqNKxxJGEdqKh9K/jaBupqryX495VTMWHOW
b5M8hong5p4YyPfflEaBvJFsrje8PsGHxDL7MtwolhJySWp9dG723XVMwgHuRPOh521xoneg3x9K
Ru5CHte3BkW2SJ9bzYs/f0CvGjqr/uVplFFra9va9MHuOHg7tSyiyDOKIdCHaDUYUWbj6+cnJpJl
zPJ4ozEL2e/HVSGeLLvGNMpURZsHHv4NOrhIgRLMCP2RwlIuylhOdjfyE/B5sFjXEsi7bP/Ah0j7
4Z2GkBf4QPx4Gm3CIYuGCn+iJEHBuw3XFPV+CcZ2x1/vpGVKVXLuflncAoblk3fJTNO++V/uccDx
MdAW8iM3gXs2KZCS5Y4BZPmMSCPA5e2Rl8JcYo7w8BLCeNj5pCgNFYZPbIS0F5LAJkWYcMKdRU76
Kxiqx65Pw3uhB3V52JGz42aFYQk5f0HTRxvW86KQL5hSwEs0iiprtvibr2mYhCnnZG7w9/6DteFs
xJBOz/wu+5dtqt7I4xguBKIPd8WcuNBxa+U5PrGLkqYzCr40feKS7IV1uSAqtmEbUBoX0m1AKDuP
6fbGaopLrkau6iHqwsetECk8mhjPvnRiC3h7eTr8VkDa3/TGpoZN+E2AKdvQiWtmXzKPgQLRg3Kz
VcAkkncAyXqBca2pLNKTT+zA5XzkdiQEi8CxLTj1CEKR2uaSSpA1FThjftWbtv4vubT3EPN6PwNf
yrcotqyGos6wxnJwaK0qtwXPTyBXWSlFze/d3T2O1op9FSr1Ls1P06MnGG442k6Vyjq+02k5KR7U
nEQ/KDJ0ecOOTK/eZmkkWo7tl50aJ1FvXQuRcRDxKQN6EKKPg4rOKKZFQV35CuvIfciVR02P8a9q
wwROKWzayz+P1/DIG9bz1QBsUT5LeE42u2p5BCAv/RPNLnY7QoUIr58Z/rTeAiW5i5RKQ86vtTey
8suf+RegYrmd1+67gDlEblJjzyfy+vGDSi0rxtxC83KI0Kwcx49eXaglam+4ZvMMaRj9dxRP4oHY
T3bdUCTPUSDM+80yMirFmu0IqHGNQ4W6GNYsp/RsQp9hKHDkwVpN1JS1JRV8trDwbNt0rxwDXo4v
KLSyNDvtaVAZ4Svzed6BcDng3HSU3Akd2U7lkbWYkHBDx3CljvUGgdTpUjbw7teoI5Kg7W34IyH/
Q04KaTig0g70PZda6lL0nuI4j5wM8bdjr+L+eVNainLhB6f1twMY6O8RxP8NOaJ93f5NXbXOm0hq
g/sq+JOGEpMX7iVlhwwJxfjrpepNrdb/CGlx7ZCR4sWAetdLKiKPbsFfDPeLvFr8NgZg8dJstvJF
vSwqKXAsLoPbVV8xn0/w2gbzO9EUJFD7BdPFaFTI3Y4BvowPkE56lGDdeXk3AZurQvHnQJ4C0P+o
/SVGxyYS0GAzNPDQoBObtMofUCxZqXbBg38ORbUzHwJ2OLf+uaKX5orGNz+edcjA7goD0Umwqqhf
9kEnAfDSwwWg/EkBZwMEvA8Itk3lBEtsgcS8pg/XAmks0L9/S02B2f5yOSap7DamC28fbqU7STPn
GXK4+dhHHrkOxhod4tCp/tjiQKbKdcNwQHCWzIjv/2K5Xys420Cud3tuc+hjui0qDRzoYU19qTDa
SB0owK+dkH+vg4CKO9InT9SJOp5yGtZOw6Xmq6Ay6yvnGws173bhQyNRN6/2lsd5YkvBODTT2CE+
8SZu+lqL0hs9NXtribg7V6vz2k/5edtp2exmD/ufrxVuzyAxeSzGPTrg0MyyL1bBfMHz03ZW4ibz
Mz4Pmj98ik5/07fVhD8gglH8t0C7lq6KYxEP+UiX8ARaxgrK5GbbTHO6owlSEE/trljdEbocm0Bp
U97Hc42AHelixBxUyRjJo7cj1cclRkkyr4LbsG47+/VoWuukZjqlGPl3FLHUdHryvkE+MaGvjGmG
72t02y3GhWSW020eIyzHokU+oVMLfIFXVNhhjiwY+4eKlaqIHBxVlMh+7eoIPnrdgPV+VriIuyEe
sDS06j6pPU7J4XTMPGf0U8esAtL9/pXIDvsX8TajueVT7Fhnbe0NMdIg6/TUvvCAWRX3PJWfu3Qe
QrMRwPnQ9pL2DgtpmSlDH+gTLnFR+N3SB9Jg+pFraZVWrq9KYW/YAf55EacpxFDotSnm047zC6J8
tLA1LRovUYI+bMz7qhU2QLM4WuqCBan541i6DmNFGN1+YQWt+uMXKoO/WIJqPIIP3xlxrPnCP0Za
werv3luHaZS51ZvOVUYSY/vuaSWWppSCzIfvxl5my6/+JFtUnn6P5D5XYqipiNK5p10N1acFIubL
H1IlLbutucZaFwUYg/k+wRQHPKZVc69+/349ddh/YzvhA1UisEX6uFleTTKKT+IdItSH0TW1RjST
4m93MfGhgp5idD8XX3I7v7eZ27MDr7gl5v+Lx2qpJH74CpP8mkz3UMDWrsVn3hGxtXdqXEf9sc6r
zZTPwS/y43rwAxc+s8goUt6qcW2ZCHgThngwenwdPgySNk9RDh9g2mXnp1UePeFAYO9rcvKX+hX1
e9tJTx7E4xb1jr97PCQ6vL9bh4cAOxjAt9EUzQwp1CrPg9QRHCKnLRUFc4I7zcQa/DpzA8HWcZKa
XEAf85Q/wEy7gEaBlZg32mhEZt1kP7v0ZtBMgg/KpcWTakoFKUJOYE+8LjIB+ES8lEPNra3kn/+b
S55VFnJ4oDYSKwC8j230Mco2ahyHwnCaXUCjMZNRhAHlctsn9Frx5XJ232L/vFNi7cP8NMsH56G1
+fS0v2NhE6yTqQGFjeJi1aYdctN467tzv6iohjEWcYQeifgRKmTY3UBQsdyK+qJMXI4VwxNnhk0T
Q/i8fQXwmCgskSi6zSSC617lFNafdUJEzJ0XLEu294yP238XP9obrMr3UHyeBsZRtF7dLkEI6ncr
VjiDWkIj+66XtK/vAln0R2EN0hb9pHEtnuC6RUB5s+LXHrkKfPG6fH0WEemufi5QKWYC+k5xQry+
SelruD6S0i0+g5/6rmKSB3RUPe7sOYF48YolDPCK7MgkXGzpNsyXvNgAanCykmfYlxgUzBVFtAdq
NuFpILtZxgl2bbuSbn4l22oZ0xDpPJBwn2Sy3EkB6bEp4Wj7RTky7pV2b5H+we0vXEQCxEbP/YEr
EKLeYhcwmWSXvi3cVk/q9QLLUfYGVlypvymnVNpOQeqBUHRi0xYbzPaCpSDfJtP1cCUEdbfwLten
3buWnxhlMOVh3vchUjs5Zh4oev2vdibggFDmhAl+V4QqffbwGVIb9+D9HrRgg1lHHTVU81u5rcB6
0zOSAkZM14NAebxf2Hd0N8NfAg4BDr6vCabA2UchC+It4hVX8/PBeyG+xlXgXVkt2gEyHCq2FMJv
akjrrZ2ojf9uNmrkDiOxUhqdNkT7LgiFe40yNFdG/E0xCrTLxOmfdZ3Ez4yW4sD09xIwxMd46u7T
tcmk27A54DnkQWS5+qIkwf1ynboL4gcNGaIaRyyyVyeLGsUFowGHar7Ycf+6Vj3b3HhFXYYsIpaB
WxSbCEufQgZ6zGUDBD2UONmroPXfTS1Tr2YqpuToCA/pyJ0gwz3LPY4MYWmDeEopJq9Bx5YqMG5R
4bnTa4hnYACZEhSKAof4ogVyAvu4g63vFdkDcbk+jMqeu/QR4/YEb02IdiWK2Md6xEyQ2ifPnxnV
BOAnWfYknytRkWl3N7oIYuRxFWTnpJq1XPCO1ummw5G6bJ19vUWOVhTLsmQZ1fX5+rVNbF49/lnG
HDTYS+aTI7/mycX2nEtSr2oYxioXcjPd2vVDZ4H6SY8JBn4A8AXbLRA2Yqkl43Qhc8k7x4MWsTCM
CH5m5aN+LbMDpZ6q11ePvNQrg+q5KlcjzJ5Kl0Fb3sxtE1gcP/8Hp9cCn4NZXsQTkT8j/Lms414y
TlTxIrd6H0I0DTkfIkg+aYHlvxlkyc9q66mi3O8tNCAXyZtRHKYJiocMBTEc/oCDwqfClFNI8yqU
ylc1SUiTfMK9XUoUpvYk5uyuN8kBGlCkK2Pz1f4PGf7wKWo4w0czyxf0330+AczJNFZlF57X0rBl
5Td/JSaGjvFboSWxNZr4myRqso9cX0Q766LgFLvkNCLNAl7IYhhbX9HxwFNRAY6D+FF3RqWRQ5L2
8qWiTNk/auzSITLe9Vp13+eZ+CSLe7cOmRvj+Rwg7eOxBtXw1N6vmQsCc0r9PIdjW5VPlWbpi5Lh
DkvfS39lrMAqK5ZBEAMr20+KusrW11rHNIoSlqoIW7NbFJ/PXyYW1qL70rW/SyMccfjKevZzDYhf
mG3XLpgK7wRUIJ4v7IDpNSV4MYgI8JXPaJdxfswrdewf6yJMz0jsfx7vd622YtXOYEEMOI0wC3Fd
DS3Hbjs2sLQ8/dhyBlftPDcVITWFYL0Fx8u6YUEcw5tJ3KQaIK8eJMGGcw/t6aB8tW89IpsycVvh
9LEMXcLyPS/84JgAAIdh1PAHFsarwjd+OBvzQM2T+sV6ylWfOqutH7PIrRFaJaxqe0p+UzVrHOM0
7brNiFEfC/NJniNwcDp3c2rDZeOG0B+h7mMz+HDGOm0RGjZjvXGyCF72tperlQn0VZRujH0AFTTG
N7bTullIacTeceXJolSgZew+B1v4tgPJGpcfsKYuRJ7Qn0A0Cf6Ms95xCpzem43v7FmE02BCBer3
iwyD+hJFsJBOte0b9zWiC+R2h1d7xbfT5Olb/+NlY0BzAdK7+7pZSB6HhPqMwHV+Tz3I2e9lKmKQ
VXFMyTppLlIG+4Bq/EXWjsOY97NsTS+yjc+wdnZhZas0WEyxAIaW8SI9JnoSX7Nxa5vSjwA2Ccig
Tsv2IAlGFIR2E92GqAHe+IQPzdmmzyEuTSQHyRggJlIcK0JU2+0qCJ8zN1Dxf8hiFZXy/FzWLuWm
0IuM/OqHE9sGkcrLuKMoEuVJ1ZaYngGqO2o7HvFwaCHbn8RsINdKsCK8P37h6o/TqA4QzEYcjMgx
8lQqiG8AutyRCvYAjJbDv4UKj7Znx6CtuOE16sOpWhal3MepY9h/N/zc5Swwlu3wYnEdYgBuP6ko
uo/Gp3imNBRafCzceXOzYjo/+avjsdGYQJJh1CzPscHtpPuzIj8qGiy2NVA8mu+mPsccb8TL8gZ8
GSIe0UdPtdCbj8OViQ5hKtQbdqBZnCoA90FOVxf+LezWvxQHElJMXJAXd9Lf4c44ghW5FcvdZY1v
evkbIxjKNEIRB39z2PI9KKamY5ZfjdJlsbsNTDTjNzyST6TyoKwpapKeYj1qO8xTkDZ81CPxzwJ8
d27IRJX/iV/V5OAD3z3Lo3zWEmJs3gn752UJ1z7CjQiLq3U52XLO1WEXH1f27+Ot2ZEs7iRZEFtB
yivDHxp+demxBZAMfxZ+QlffNmYlgNr+ZuT2Y5tQyld78v8+FOupSf7KZ3QRz0t3CaG36XwPYI+x
veLfgWQVr6cOEqTFMP7TfaKQ0r47OOXzR8DRCbMXRCv9nQhULRwh5ny9exBV8b4FgFakjw4T3t6t
6lsvfPhPmOolMicfYn+0vnhtFPZOidvhsOwDhAvWgKdIiP315IlKc2UB91HHKfaSBmIkDz4dkGnn
exa8HpzwDA2d8pJN7KtR5ulIOq+bwW4V94a7vnFF8U2Kd5FSSK4FdU5VrqZ01eka4o076ZpfaP6b
OxISVAj932Giq3/IAHRLery5WKleVCoUJQIg3MBBH+DNPScP0eNrftPCZ33S3Nj9+OtgMeKy3aRu
hphmJvLFW7A3A8+aqYEMCihAfvSkMeAbagZCeiz4OMUD25aMY0RX2mnqEK6MnuSUeqj5i+NfNq2x
wukSeFpFgc+NYdxgwEZyLmNvbVGJF8Vv6U8m17E5kBOY+PCUqI1S68MOBY3aIOpOq/pYTa8vrN68
qHUHqnli68/ueluZvqWaY4PEZ8RgyEdnv9fGKr1TIwC53rcB2gsdUMw8OaI1413TpSX3b1YUPbKX
wMRFjFI6u9qH1By0s5syK1zWr3x9eLimqH/bgvw5mlA+Q6BSePiHfLPwJ/jjnDESFEBuhrzeKny5
/PRakaVg8bJcDeYIF3iWqMIEDubKFrYLQjBSYZjHLy8h3Fdm4SS+OPEHqEvceCemxJ2JHHxcjx3m
jpqoHVi2PWQLy8H5TJpx5S9Y7BrbUyInXYm+b/qij09CYOezo+aa4502Z0aQ8596jnxNBv1+zD25
9Dq46neHk5ffL/Qpuf6KjplJM8enXKuEAW9ia+fPTA+/JEdxkyyWPT0Vt/D6hBSjUflMxCOlfDbu
LJJ1t9oSHTayV+9LMLMkOSiKrBA9g8XP009OWbAYweRuvA+f0E4APFEluzrLhih2jaDwc0pGh72M
1gJMUVJomw9EFF8S9hTkd3CwDEM4lGJaBgeIs2pH38RfAHMlaCm8uigjs5SOrUiqef7xLprd5QzA
XEHFiOicueui4Wdxs614H/PaaxOmRGhjmvPF86/YXtJf5fLChYlWOzSWKDyp7P5ss6qOOR5M1ugG
tn3jxdiaA/WXO8Yj4lefcDxNSCxkfSPUItxnWyNg8de7QPkiDmzvei5aF3trjVPi+pZ6OAYrDzeK
D+0bTBUN12i+qiMLIL6I3E7UyYsWJJkYuJ1ksI9bBxlVZUeaCH5Wt65hpVJl0JoiCm8uLTtZcNJ3
MStK2/RONS6fvomhjas8SRnrLin9d8NvGMSceRFeAHb5h3SNKpD6l5GkTtppIUerNINyJsOhDeTn
SsYqUX0FIp+TMzTgUhiO1UWNoeGNExmSG8wDQiix4NuoL/AuFmpdd9A65qwT+t2IIl7sFZnL6FxA
rkMp3fX3niCF5LPvb8qn3l4tg70oPXuc5cy1SaNTExxmUEWPfKkDQ2xSxgjDvou6Oo0eiNCt880a
56ln+f28x3OS2ojbZEtmvdagprdbhFZYHuZiGJ3bS74yRDBRhZ8BAVohZN/9OcaZHLdNsofD5P1m
6O6imQQUkDvkp2765ZGuh9XTZgv2hrTdEVg0Rj/YqLTxpMPExudiOxrNIXFAoCrQdQxDuLYF+16z
P3aBFRWpwAW7f9btKyB0WwBw4eltjNzqg/hmTootQjz5O/N4FIkHbv5RTum/ZtWzoyKs82CBO+3X
XXHd6nE8yl/YLvwozqlcI/CxpPmda+IcRTCcotGGR2SPcP3e4btszoR4EiqcR1o7G9xc0sRz6h6t
bRqe90x9AOk/+eN74YtLwf7lLe8PzIY5FeecgY6F2SApNd52siVRifs8LvWADdoxDdO2NYIeWgIV
eV8pFrfYX3Z5lN46erH/bAcM1kEaVg+E8Y8O/G8PU11am2YpaoipyNq7GV+p64WHtZJKZ0f8kVqR
JYk0u7Ga3gQ8Y+fxbbZ4ZBR9Sc/5wrHWqAGMQ24fR+TTaYc9IJ34TD+jo9f2KbxqHPOKal0gzKZM
AZhXcxh4ZlqFWrmqO5T3nD8Cqi0w00yzQ70uMQ57O2hrfZ7px7dM+/ZdpNnzIdvijrTsbvuLMqO5
oOr0gaoA97xkJYqaw66eEcnxd76piX0b9Re/v/OaVqEVpK/UJzwAAHIkDJ0Vz62s9YPd+oLdGHaL
RhUm2+VH54TBb4x0ErefeK/ncYpf4PpuyueVrIk9syIAAMG2DvFx3u6hoolguhl5RGDUV0VXkeF2
zQX7l59ufSGAifzjTtS06qoDyFEHsqC8GyIGc4RflU5/JMTkwL8qL/dzuYdc5WpeX2G3s3UKvEYL
w1y8Q7+f9y2akdFOD/u8UQFhpqG+RjvWdBV3kpM+mlzrdM/xAwszd8nIa7waIIYCXFaHb8Uxm+4Q
yPxxwim4jOFptPHSQLZDeYGcPSrboKHysf31aW51qkvLmjGsH5+7C4rz2pw0rYKRZpIiKnDt2ckD
MRxgDer7x1J3+CEUI173/DjpC46I9qxpRkVZ8J/PHtR/ftU6WI0EB4c0GNLLlO9iB4hnM5cpGWfQ
t4romQP5yNjvD3LgZmvlZ/K01oyGVtB99xJY38R5AhbrWlgzSrEM2KsMHnP6E48sPSLchCaABL72
jEUlQqTpYMhjs3ewhmg2KPbAYH8pYIt7EaV78rs0foQ2tc5dPlINGeXYVuDkganxdxrm5onJFy/t
qyb/LvvQyfGCaQqgKwe/yO1p8ms8/35umah0K7uoBzyuJMWjsn5MHC+CQmiXhUvwDRdHOMuizCoL
Ha5xb5HgnIGPmgqL2qfN3zpK8cK9nCtg5JnC8std3gy5DJyJhrbYMmVBcm4iUR654SLuQL006VVR
7H6kEJsF4Neuy9880ZDL9Zk/TilixHb21v1hyDAIJnN/dQ0wlQWbyMos887ubTV0wHEuGT9mZxkZ
qgBlynPNgEjjys3Gi2HKI3D18erEG93eo2Ymwi2S8j3ayXcqyUkLDALneV2bQ4cxF0Kpk7Bl0gQq
qt8luRZcZKeURBG/d5z0o0dtO7i1nCQnE5kJT11n8zwMkB1im32RmwOv6ZYjRqy8au24GKhLRFB/
Sa6Z5IzO/ydv9vIT/jDh6gnbQ1M//X7z4FAdM7ZHvolOE6uTMvRF8pbiMu683RWnNYRTITMCMOu+
EE9B+kfqM/9pGDryi45ISf+vJiTkbcK3T5lsn28oiP11NP1nU90hc4Px7nRYDqTaOts2nFObtjNm
MWE7PSxw8YB09O0VAASHGe3qnwvY8fTTb4a9aVuo2XHpLo/29CqnHm7HEzUcjH/+ZI2oc4L0Tczi
SY375I3rFSagYpiCmoz07vdco+hDLAyksqg8TvqtSDFC1QJ8pvNztKQj9Cu1SdEvJ2HZ2j4XJqBJ
z7BT3b55PD02gcjOV9kO/Nquo0crkTAf2IRZMY4SXINQKebE3cMMqjrRmVKBqJigs69rbB02uHvY
dT8tJ5Ro6QAdDx+c7i1IsrqW4cJnlu9y9/AkuxcOCrMZhwmxjBA+rb8n3WXnFtsucrff9eKIx/lV
77ArCAUc83vxRHobrWB4H6oUnlDlpmYBj/PQ8+R5Vrr4yRgssvKDawPGKmdIx+dQGYgSGakbL3it
l/pjx5xEplKPzF4tSlAo9kVeLeg/dR+T39tF01Uyha1cEl2ER1zZ6AMsJZFCdVRnBQ5I2umyAP0J
+5MtHWmIz0A5UF46CRGF/Rc04mS4zhH08PGSKxKF+Ai9Syj5KraXOvG/GE35cZDhpOrsUSKSVJwq
vVOvW9mDR53rEFy7yUuCx+mlpupa8VKnBHuHzxZQDyh2JV1yL/Lj1o3ThoHQ3vspCWg7rDYYg3vp
dUNuP2kVAFybxI8o+RyZXWykcuTV0zub55Y1w+OpWFXUXREjfiRWjqo+UHdfiY6Bv2P9rVZRz5RL
EB/mxVvY9MYeWH7YYB5VDeJ8AXzsUwIZkIl2xXV+2IFMd8Z1lg39D2vHerqXC7zc9MvcRsGMj34R
ZUN+TzeBXTGRArnh+MmazYLB493SM84TMdjrgdlpIX7bdWYMnPTfB5i15PUqMZBxxUJeiKknrFF/
vbMWpX5WWEodXD6fk4iZNrhhzRlV6H0YdRpkG3JtaOJNry9bPZfGXsalV51xPQhBq2rffTAXKYzx
R/5jeAa84t58zOHNsSNzGVJHr3+Z3fHcpcdcxAgILMPvslXc1Ily4slahy0FhWViQoY9CFN+FuRk
YYCBDOicmfOAn74UCgIC/4Li26DWfyjOkGf9lzA0h/QC7N4FSg11EN+ZMfQRJrOmeAgTyeBTgYrh
KqXOOsEU5XkfSM0rCUPPjQeqQieI7xzSVr3Vu/UJyWuDEM8bWE+ReFM63rDniTAi8FCmwG+Ajr7T
xnltWogiMSwBdxNCfhJju/vbCgmr4pKMFncQOS+QZbkJgRHOhiiR4+KWywc/fd9yakGt+bAT0Jz0
tmWrFWtU9bdggTpqKRfdnicTk/3rnj33EEHEiPMdWvHCZlLcFNLxmBI2MFBgfShTCuuvKlq7MoWa
+h0URhzEzRYPQjqp5ZFcWR8Kq9WHSe6qmAvqadF/EnYfJx2EM+WxZPmkOBzwjL4sBNfoOwF5g2bx
ndnq8/fapnusesl3yxlTTZPc84kUdsM0lLqMSF0agNI7x/dwZUomAhzmJCe4MnWyZHiwI21PaYcG
8UG3HAgiceRH/XAo4LMjrtUUYlVW9LLoQBAMvYAjcGjyXBfmIR2eWDVtAtj3kw9Vb9IT/sSRl19E
LQBiG3tZt2ykPLVe9qEFn+enbv9d9h/5tKuW6YPvLWxUAWqH7SoWEayeTtJ1RQM30kB1dq4rpNnp
XfQYzKqS/h6QC9YTbb+Puowa52CksbHOlj14Hci52kYQmLQpAKWmZKfmTjftc3Zce6KSZd9JWCRX
9BNJ15r0t3CVlOLle5iLzc/4L11yOEoPeoy9Q4siyiWqasBeKu/5stIOQjv1arj1ig2JmzY6Q8JU
nzDoVXE0UzEiDtM3rHjO0uUHpdDqMIbGyzadSr2zYp/DjO5+DouneysOECLa29s4Tg+0n2k+A3Lc
cqRSGT2EOxdh7oXAgopl2Zi5TXR5h2kOK9B3r3NXbqYZ3ZuBX/FqoPfTD3+fxBVwlI60m08YKS6f
JZjz/5cxIR16tuWcar1Q3sw6XjKCiWAWMglmM6DeXCP7C2oeVn48BiTggkDHs3AeVVxR/VQbhJc3
ztOxmhosauYpBQE6kHb1oCNLVqh76pSB714aCZ+fPi3iwt8CzqENwxf7mGqfy52fg5NN69mxo7A4
5AOieiuoqSCwwA89B3YR3m0iUCeQnHn26RN8dX1mCgep7nn/icDZOhYF7R4jOtMAeP57aUy+gez+
nzovKNy6FeM3JD2PYmmhP+S5MfwrPGI+dvSDoOuV/xKrmjUSWzQiIH4ybtaifzzwHofuwUDuYLPS
HRRtwksaA7H9ewNJQylI9M7uael5tUntet3dJQUUM7V9O4eaAo0SpMY5u/dQRHhBTQFULmMajaVS
gD0eO43ujQ4N4BGbx/HEFJLu0nzqg2I1mLdkj8fFqFKXGzQHsUPIPRQh9ZaYHNjNCXZfhtSbacKT
Sys0lHKMpKckDfmkrZwyP4F0dbNFlWGCSeBL3m0hZoQo1u5RzsEq+7NcAyBIi6Uc4oPgVqDGrbZF
BFaDLcMtyGJDqgjUYlnAxR63XH4aypjJQTzsOuknwWZ4smtfqEt8sx+N7AMevZ7KEQMizkQZYBAR
G6M7RBJ9e1OXWE/CUbSqLdtmuui3nC7uvkbH0pa1d7BEZusqxIwjHPwoFHORK0jxUN9IJWvpNnRV
FyhBWZCbgT7BHAwjnR+3FTJlbKYmrg6UOP+E5m5NCRmxIFFmIn7DkrmH1AEC+Y3IjnAGjtEK13Hb
avhg1LNN3wNtL7IFAomSB6AlwvRUAdFDsZZZAeGtPMECZ3lhQTXSzHu0E3A60xsiD11j+9LThLNK
X+5v7yqTM3eae49gKPhqVVg5T96zzxv5fgel9sFjBHobDEMX+qvp6fvVqCB/BdGVT827ovnoGrDt
ySliByrS/++rrc2SimHrfl4WtkFMwmkGZihEUoX9+c5fnoQ8TArP7XE1ptmCjGvyyYw+5LQ+Duak
n1p7rjbvT81mHZ0xS0bTgSk6VgFFPdicHfXT6cfvNRMsPBL2d2+EkIjuNmIUd0IBvwI27/M6jHVh
pZgmDkyJXUyQa0rPwXN0uivRU0sjZX6EouNnMygxRvbM7seux86qroz66S8fKD1tJfOCGnSUv4bC
kNDasjb2UOAUobg5gmlpuqeNM6VU/LlCzEOApIn/jbuIsR/oh0TZnK4WXHj2qUkQDiYmjsoal4B0
GqOb3LPF10HP0Np7u2gYKJyXN9EXtnbwRuCBlozxMIZwhIdX9f8bDt1jzr/LJqXqzuaeyNit+9q7
vf1BcgCudJA/tC82k2RNUzGsfmuiXOJK1971ZajYR04T7bTApp+fNriIIpoURlYwBAq8/BgnmbCX
0K5GPmbEL3rOzNKNBtNvmNtT6xmboH14kAKd5SeSXYyFpKLgtY3gV8ZVS64Ao7nQKmfleJ4y9N2h
t+9O1aU7PDxhBeLH8D3TMQsQreFiK+FRmLKztwNIFtIBAz2GVcwcZKP/NRlVUN2Mj7B2Y1PFEu9Z
yVJcDgDZDZjimG4+UWsuYjhmM1J4vYRm2mQF4r5IrfNbEnb1UG6SIqMOzBtbc/cKb+Vgg9iGWa1z
ufn+yntznKlBel6abvqSvvXm0aFeARUNnfcfsVhvwvSmL/uFHuXuIjRNW0tepnGUci6yFTM49155
PftMcuhg4tp9/T+ii1jLNr9OOkz4204Nx4cITsdnmTTyhZOcwZ2nG29wSv4oT0E2rr4Wnma7WVjf
vE76ni8N4ZXgl0fcPj/Udtb/+3oOhP/OaNeFOXZnUCwwuSf5+tWAxiU3syGJeUrF2p4WnWI7KR/B
nvwhmCi8O1oH9j3ecFxuE/fFPw6Vg992pY/1lYBn9YXEbyn46Jy+MerHnf20UPQ205Hb/ZjBBNNT
PKaKh9O33EmykSyZQUp+ZLdSK/1oMMgmF2fBw2Xhn0UDHeGbIygS5ZnHA43qCyhMmSv9dfgybCgu
+Kfiiha6EF9GCAWpxR1QBqOjt3wRlbY+F6PAV0I69v/wCJSEH22w77IyqknPJUQXPWeuRcH/LMWF
L5tNWU87bQ9SCUq1eRHSgXMm3mcXzGzuznYL+tUl/vmTfJL/nFiMIe1slBWxZlJ8RF/bhO/yLG+0
hwYgl3DRD0l+7GJXeajn7c1oDSFefT07YrJdq/GG5ct5K+77qV9bf6cZfPQInonEQ09+Ddl6c7uj
485ziFjbn6oX2qyAgYLEla2VtiFn42XZ2olb+6depJ3SUNoufjCBcRk4YvPvgp35qXK4DM56FQHe
89kUWSLBRuOXfGyx1Ptd6zd1ywwMlaYj3RWetE8jK4Ch+uSFnyGtDJszcm6U9TRk8W9K9ulU1yyE
G6SpQXW7BeBCRw/6oUAgEn5OYY7MWGT37Fkx8OiOAYtBU8wq28LEiCol6tI5Y6kKfTW0Y6o3+U3e
FigCWoKeKOei4ZQfZ5Ukax/UE3htTNU6XWgnxAESm3pkgC6XZnTZ552Q6SHT+8FRlCnZwJJBGn1n
YMgjM4uIz7C/xDsd1RWiQJE5QiEhOK3nQbag/qVr1g7gzzeepvLTyrfjpPohaucIvu1Msxnus5sN
4W8mEugUvFH1R2zyTLHLAA6TJq0M/zj8YLxv5TLqAgPX1VPLyx8SzmDLTqpSQBpTcne03t5U5oiD
QHVT7ztIcyV6IaR9FADmBjngrk5X1IWyJtiN7jmpsmQZWK0hCDwiLoTSjxaXedXirn13bDsaqIPS
384oe7Nq5zFUj9+65GnTARoUY1KvdFO4NJthMb8Hxr057LBtnRsc4ZaHJLspPSlAhygY2De2uU9/
0JXYLVoPSIt898RJB9jJgSbvJ5vyZly/R1ZlEj/FcE/0p6wmNefeYT0qmMOFOOYKppPiKJ6YvUwj
hUBBT5UrS2zorITew+UA5cXk05tr1iQ51ebp8StfRjbYVj3dg1tEXKVb/1Sq78CdDt1GAAn9Q/bc
H46O/mRgv8bvAnvzLiTJcXUfUGrATW/vLLwD20HyCd84/7prcAMrWFWJ80J44HU+QiE8/br2b+Z2
ScEZGBG0o58aMVE18Fhu5lXCcWl1aVW2bzYPsBYgbxoPC54ApWeFQRIdaPsWlUIdLdQYog6S/jwX
ycDZtZn9RHDEhDSqLGfxx709E07rvGNJ5HYbsiVq/47D5NlgiqQ5jfEYOpwvjzmFLPoRb71C7W1W
M7GXRh/aIp92jQP5XtJ0C5Ak/qNJfI2nbOJ5AaA821ORcosbD7mM9SUHWAfxP7PBssJUoM590ffX
HJkGxtF+758Fnux/w+y2hFceY/ifqxUJxmvL3xGNk/aTzTTnzyR9dN1gO1dYtzKiFfg/nR3CJ29L
FR6ixaiIf6psLvY885669ARZqPa7+u/7e4ppy7kEzIEwMUGcpT5YZuQ+/4BIM5NohtFV8eftZmFa
ao3zLDfW6qOzmV6wXP3T91EuZNWPXBobFXAYmmV/QvVG3HhO/t+NOp1yIkMtrt85+Y+40BJdn41x
7Yf7Q1UFW4p1vNLUPdNFJXdVEaOzdIaiQRCDh/AbbxnBx5MlWzGwsjht1H1rGO9EiaIVo229QtZr
unmT0YrY4CtGtD9VAfumV7tWSpWslHfHUGcZ+74doVDqrKALNywf09kwAgiNyu3Op/QjKgU3Ar6c
HJwvGY9kShfwKBTHt6YwYFexd/dQSj15oFICttcqZa1+aNH0bVYOk3cs+8g4Afc6DhPH3+IuLS/f
u7xMBHM1NTQqezKeEPk1fEUZqf9qYV9g+sTBnIK1YQctYV54xPrbChWH+L5iNOPKIFZG8UtE26n9
CPomxmFSuC2g4/HoVeRuHWRV9HJ0aKHb77284p+AKr0oE9/Xu9H+tl+qhDFHWlXEhbUJcv55DBhD
gJMHU4aTXRTSuYLmhjq9PDPLT7EOP5WrNMx2d0a69BflN5UwA2ofknJ24wQOFrQ3jlMPzRqDt1zS
/EmEoX1U/0g3+uc3sUIgF0VNVHt6ryNcS+zDTIpF5URwZYlcK1+aB0CNyTEo9uQ3NaodOcZnNFc/
TVbCQMV5L08VCUKOHlaa9yWZbiSf0ZubQhbUXMDVMMYXRNg0UUtQ9rs3xVDHOhwh9zjwwOm1fXi1
S8me/SVABgz6B6cAC4RDSz9YZCkip9orp8g64fdiA9UO5pHXG0ZNgwo7as5BjbyIaiOoKCoDJZ6D
1M/OjmspeadOV/2Jz09mdxdydZ3yuLadPOYQE9CfJ8vi0ycDYM4BdxA6Dx/rhb3xH0tMJ9RPgpHA
So6ZdWVMrjwRf0Gpc+UNZmsW5sHDKcPiiHmZQ/P8OXWBBAMWvA/zG6KYWaBRt4jxteoS+mjVMWWs
Rs7z9ZGBxGD4WedsieG/Og0rWqKOLfqd+phjawJj5OubT3XGRdiswjJELTyUR34PiCOd6grBtEF4
qZ+APrv0HB5Dy3+pRLwpJ8dR5Pd8QSNTE7y0WM3rldBOOc5bjcjWx1PH7Cb4nQ9L3YPlzq1L3JfR
RXyDvnjbKCtGp6mTSFsYHd+RsOuwLBFWpmAmqIcCUYObezqgswhXe4iVqqvgHT+Yc5JRAr50ddWA
4JAeKmPZGF2pe9e8vGo20mmO3VVeskWof9Rjt8x1y96WeLqEBHFPauVQNGcBBqlDYi6bghWBtRcu
W6196kDME6bDGCYfd0B6LxSLxz6oWUz8WKufFShQ+ItScGSrJIjJ7vdZ/cD4dalCNh4Q5z3k2R+e
vPdDFh8qkfzY6WOoS+WaV8OqqpMnvaQ1tOQANaTHql9FihE6/7jMVFW4SMlNNh0ZE4ajQPeuT3X2
ZmMCHWDN7+ZHJWK/OEtm+65myb4ov5GcNdx1UGaAln2wERhFruP86N4tT2cYfw2V/k8FcqK2IBM8
f0db8v4GSbdO1t7v7Rxfm1UNO6X/SSLNCGD0zzpw4aYuPl1nzBjMZ42TESdjira+65cdN5tf2kLV
iTF5o4p9DPNcrOLu8aynEI0fm+w1SmAAGrkkxD3iTM97/uJUJjxTqrAjk7tqelbh53v5eoIOhubo
odEmUrAn6BwepstGs3RbJQqi19KwvcY4b4WPcIKSdLKcG42mLXQuieKvuB6DqGw8ILt0fV+Bv+yL
syFfGhVUkGekuSXZdlKzzwOnJrYnI1SvqDTUQ7Li+XZFIur76XOZs+67QmoSFtbJbsg/uSzmM4BH
En6Ulnn/9p2u/VVHBfCJmB5SDL4ubwpsV/aDHdGHVQGi0mXvA0fjp8lUVCdoFsvyZpkL+LWtYzHp
KJEASvMAwp7ItVuWj+uetZ3xcLOm6N6omgZ8bHoQe1lmZHosMD8ts9DlV5yX8rdjHMN6yBnBAXOc
IXj3gLN6HFqWBiOZ6iofsr0vCxOoVdBNxIjQ5C8ftWUT5gTism/y9pIiaTJ0KbKc3ZvzwEreVRiS
NcmvZ7wc5yvYuI6Rt9+43yvZTF0RgT6hdB/nwkBpBVs8XhD2wySS6JbpDMAKI6CPA1Lx8sdnmXNn
p6Lcez9ecV/vpmGdF9XmSa3tRCZPfczEVnko3CnJpZVsOwc980Qc9lrH3c25BxxCn8QRgU8EPnup
6Afn4AbydjaEv02m+BtZLZlAn7X1o6oggG2U0W5+O0r+toY87ZLKxUs/cyK7QLIydSYYx69Pa/58
ltVNUbAFr8cTnBiTx2UU9EIeG8dWh3QNlARSxioPVSkmPHFsBye6mL35dNbkKk9Dczj6+8agyrTa
GFAhh4y+yH+4PiRYeIozlKxWH8t8s5+2Lc6nyX1GAwVVegNetbfLScA6omYf+ixrYHpQMBtp3Ypo
Hsi3feGMsXazwDKOoSSJ/T6GcjMNjzGxo4KUL6gD86C600yEWrdGHOr5WpmWBNk5WSUe1w41dTxo
scgs9exCOkVozRsGRTwcdKHP96zpJJ2Cf+xr8DOrqD2+kHpTwHblBFCTFBPXMwUReiyCRqwz1qlj
oxSpky0f/OTSWlpCnLK38Vk042UHqY8a7fvnkIAz2cmnXVxiT0doIjrO2SBjGmr41oL15CO+90Xl
xugpEhYDRjPOx3JTFLqtdNbVR2K0luD2Daa6XyNYtN1mX8kxY2IGnZ28kQ2i5yhTA/aQ4ymgtDzG
N8bSxkQFqMUWCVCYI0QNJzPbbvFMz6cEKlHzng5aXQBxpJ5TEqUoDgn53n0wqzQFuttk0qP4ILQ9
+bjq9O83znQDuKOrkEsMhbJBrRJ9pTABd5tAKQZ9Ncx6lz9lt63/Ha+YP/+igRTU2SUk5IiJ7Nh4
0pIagaacnxOnQO7y0NTc3FLOr8AdIEvXtTrJMVN2nV86R2VSjgkTJQixOJoKaTDlKsBSqVic8Pgb
pcR+6+fA7HPT3u9cMCHilXOAe3FYKa6dhaaqWDiShD4I/18LeJfoe0U663kQ7/4/J06WRi1RZ1Lv
Crvy2t9b3ZtfrsWNjOZK72P48+6Ev+CzBaVy9RL7o/MHc0MbQzJ9SiRDx9zhzj7gsBueh/4AlIxH
kPgH0os+U9wICQf0SJud8K2HUM14dzqYD4skB9z/Cub4KGTJGM2vSDfySvzJeqsTQ6pl7oB5AcST
dPJ8nppeSPX3CC4i4Kl44lngGpMM6brcsMoGrbawDMkuO51iVb9WvxtyrHEmtKYYtILqJx3JXrDT
E9F8dPLgrHXjNZ7wLdeLGibsY5hT99k7NzZRCpgq4/uZOtxNwjyzxirf/bfVk2pTmlrvBuMvSZtS
KOM0KnBxI20Qm6oeiYKGEWLTMlx3pdY1fyX9bNHdwDS7z2EpouI2ehjQuUqGJ9bN+ClP//4LahsN
Vv5ocZZNMikl1ezy2ADpITo4iN5IQI9KXUW5d397sX4Mt+yMHR8cwHMEzQR7lRNSNi7PIZUMKhJf
Gbe8XQfsMgMkFGbtLkbCWlOzsm5Cv0Y1FT2dq8kuMI5ThIp27G+w+WXL1nN+wry+0V2l0/wZDqBj
dyTPxOsZebpzA/LS0pdJnhYxvxhlUdDq+cdS109mxmTsZVCDO4dYAF9fqL2iWgTIysorqoCbfK2s
7ZuqyVvDXsMhCm5eaXnzLNgdIfzk+JiGUHgK1YGnViB6jWTCFgIxbya3B9+N3gE9D6U24RJ0HReg
De2wSFVc04tOCYeWITRWAUAQEENw4CnPfpNefeTESZZAToyEsfTPUHjgH0jKKXCw09gYNrAgOzrk
tADNthfluufoB+/YtK1ljdGED1K+VnBGml9NHrdUH+RmOyvMS/eLm1je9UdzbgAlxT9tMpqmMk2g
MPnNbhvrNrkn2GzI4vG4Afbamnw9OQcZXCRPU2CY9jDKPRHzh6NLrkS7AOUPurjhWYFis8Ajrq4l
wbF12X1bVqiG3ey8JjBVmocr08NPsKHMxaxOJLEDoh0RxuEFqk9DjY7/8G2eqMPdwGA34ZYCfznk
OEaGxGt14IJjMfI4HpOJiPro+z2Dnm8wqdeogH+INdNgawgfgMZCIyD0y5/qycdlkJGfxRwOXvbP
tKea+dA/rZ9LNWfNTzGQnEIAaaJ/+rycnEGRxDgFG0vmHqfjJ+UB/0TwzxfpthhNPLdaJpFM4CBh
xyyMxYNjwhp7M2Q4pinj2hGE8XXLXk9X0kLI2LaXaSWQVSbcy83Hv0FZvvMsrtjoD4NNLUquPiLn
5L9I+0bzy3Lo2MMXbXVASivVaUXVScbyQ96p/0X53C63orDvcmtKgLu8+X8GSN75knqPANxhESRv
7BmnHcmPgYQmZf6A3yGXGb9rMEucjNLNJPN+cjdot4TO8A8Z9WDh0Hb5MKgioIVi1k4oQqnJV/mH
8As6oj5hWmgAD6uXoMqCZMePnN4bCnvoiso1VuvB1y+STo2fxrIPbPUNnrQ2zPOFMZO3yqm/fB6U
IbWzViU61gPfIMYDw2JLZPFhXoigzcPkawn17oXEYhMl2s8Nanjj6rgLHHB4uQEZdelxcrrVnmZH
iWGVc0anYq1fwjcqIuyCKq/9XcmaViCLg7mEcXLWIj2MlYPVECi1c7xDb08/0GQhyKe/qdYiKS/V
3Vo0UcW2lVTw2UXlvgUo5U/QbJEOXTWj8UCmoBnmHv3BLthOKP+LOjaJq+qE1p/sCeIWjirY858y
TR2Tn4k5PPsHplyvRWFl6fQZTMu9cPQRNrDF8o0wzjSm/VEI3Fu+WaQkmod6VvifJdiTBjcOLjdA
Ob0bjG3dPL5+HH3FWtrYZyjuxIbNauNTm3c7fpE1S4jvHL9nlH7uWgTuUcmi/s9oBxS+teUUOZsJ
v/awtJsBEQoeZnQU9wMAGHxnhsX/PMg0Yhn99DrGtSoo/gLbxr7wG41Y5NdOeJphND07oEABcjbp
plK3bIm5NOulHa2bdkTk/XPUwheZyz6nH3YGY2n49RdLgOpAMlRH6+zqWOcELNlQqVhhMdVWGFeQ
0IM0/J3xG8Nvt/bEv5mqEDeILTsB7qiMbP0r9Uy9EswMdC/VLqqhv1HNmnFdqjL1RgSpZOWCT/cr
qQ9dIOIHubsr0R9Uj3U569teI/BfyVpH1biM526nC3Al0Vgok62IQa+BrY8lPojy8XhkvLeNc0Ou
6fJykiTESx5Vp6Mb1DkWDacgherfKq/v8DKT+9/R4d3jhTrEh4ERzg7QLWOCKLFbUvj0VZQg/Up9
G0PVVbW3oKPjE1CxJHeqXlKGnQHDgtuuSYBpwwPmO2jStiMYT+o9U0VofFlmbLpOzlti51+SfoFk
BBSXbfoQFVjzt2yPEIq4KOB0U6UHZOHevqLBLS9tcS5AlKs9/Zw6DVpSUZXa7YQ9Bvpdr0so94wI
t4YgNfMApjwWOeCw4kpRvk0BkoikppCBAyvKDBuFrW738Xh7FzYAcHisWdkDueKAXIRV/4CO9YPE
QlwENy7mcNegnRs3UwAT2no57TKrLdgXf1nRFJfh6F0rqhlVfe4Xn0uffw1Mdym7Y9V5AZwtkiIp
ay9US/P9rA8+xe+opjt5yEC4CGbdLbHJCuyB7kUQTzkYPRkzkk9ji7/qYf3bseIFDuqiJbR8XlYj
zXjfcL4RtSW59uqYXTXJm0E+EwIEmCekL35e7pjtab1rDIvgB/97c/ZOzIt2DxX8YjJRyDnWwR5n
PdDdfQnAGH+fhxYOVzmAGc0miMQrfAi4JJ3sqQVsJbjPoAZcYE1orrJCyysLMULEokQYyKLdxhsd
xovorg8xSroEOX2FadTjAIs5gzMRsB5XSGhdoil8lSy6rXs1pW89SoeZcmB0OG0SunlxRxh0yNZt
Tk52Vi93GB/5IckOkyeI6L1dFO559dk81VUoF9eIGXxj0U+kEPbcJrvChbAlXLzq0jGIEQ4gv9vv
3fqfay9OxgLneZ4FrxCdW+dz+iy/84ANrEi6HhErOF7BT97uhrVCNkoYRQKrDuznU5nQjG0zmwjY
YSbqBgIsY5ugLiM3//i8KzHeojnXt+/qzw9HGIwCIr+sxpynwbLfPZejI88eREmIeR25ZrgRWLvY
17ydigZypf/deZEmRpiR27Hqd0rIz0O5dZYghNOb0h6ySZDRwcf6v4tiVpD15XeZmk8/AA+WnJfY
bMNG+kQGbhE6+tNOL+Y73YyBHhPtTh17ldg6CWGeNvOoOY+J/mvhwA43N2+8YdonFhEw7LOU4NVb
d+cHm2N/nL9qWKzw9cw3dhWB9JK0v9bFjxSj1S6Rfa4Ji5cJsAm87QFpOmjjxbH/CQD/sx+ebPhC
WKafy9f3vkjOBJFcM6CNUKH0n3Iw2sckYks/MxaAzpLnyayraKIetdmNhAbJu/BZ2AdT15FiIMGO
Abb3BBDeqRHmlAfNZZDsTMQbJMEsdm7TIix5bgSuv+zzN2foLLg5ZmZhoQpMVxI3WdlPs909lBKJ
ewiKUtMMjr+DxmEgpyybkqn2PO5DlkhRw64H7xuX292MkkHGVuOeQqTupkuVR/X94H2/ntTlHL2B
FZleDZDopFMAlYvDsvltTszSaskwPQpVz7pwlvh60wcNKUMXkne3QuJVg73XatXhcXKjdl2LG+Fn
DT0lO7efIbn4lRU6X3Z6GvDYKogy43Nd8rc1ccsXY1Wm3UfsxYrNy3/NKxi8lSQzbD8OSl52r12H
dr2DQFbFbtBpkKb+l5TjGCcLwMAQt0jXJV3D/fsoyujsAJnxJkoGwf8Zqpq89JhUIPM1QuSfmZYF
WgjFM4T8JK+cNi1jQBYyLpM+wpS5KBovmQ4dOyplYndWEtyZyerbgscfxJ/EtUlWusloDP/tW1m3
/ZLXxEAq0J9zc6BVUY3ipYbJXoczdp6Vyw3unIF050jtRbV48nie879T6uCAoNqeh9bP3mM5X08w
0srgxRBYO86BfYAxsg4oFNVzzvnonlKCLZxlQimyrs8LtAtvvaN7Ayhex+8k+7dQVjIaUb8MR3Zy
vwqIfWb/srGpGLX8+VduSv4c+aXzSk1QwdKNDSx4CciONCN1oBAtE4nbqaDXKTJtlj1f6YDb9P7p
TrnAVysw0U2BkPEmzGMwOEj4SGGcHHEx/EU+BxwehhQ4AhzBPJdPMrDAGRMR3H/5hAQ+Qwc+7G0e
xQuLhYfXOWVOMt+duCzN3myyIvOf+YmgydhnH57XsaKgIjnRcf2IHjPnzelmgKEA5yClvPRqNAOb
Pyrbf+jyiS7PsCTAq6Ywn5F3S85fmEO/97fFYIbeuqSviwjS4263SkYDlK79KqGEXj1YCcAPgqRE
TRxj59N7Cubf/fsfKeWIXuuH9EWCfA/QsNSaaPydDtTgNnKn1luZUSTgxn0jv7DD7xKwFnBb3u49
2iYP5iT2o453bnjII5l8FZhBzN4apKTaUfssseCcbSjLEfstgoWXNF/iS6Lb8iC732UipEu8EYxB
6xTL6P34Y/NmHr2VtD5ZX9Fphe4DZ5bGDiElHWRl8oOuCtBJ88PsGdFeqH0x4Yh1NObQiUVaO8Ju
YXS/dwGkj5Hkx1QeybGIiq9FbQ2v8ehpBN50malUb+slQ+ebYxXUt+0B+x4dETlXbUf/S7tVppG8
QkqnuxUmRxKfT7OwGyawhelsbisDWxpv9ZHxtwRXv7Frfo+HFvUvB0yV0Ra9sWk0uTe43t0EjCRC
LoqvK1YF3MCfgxLwT471UvtrSnZecnzbnSPsEqyck2ycFw3JqY4w1y0WSF+G/6BbXCfecw8DNSlw
9PCvw0/hbrbfr29d9+WcZ00V/EfTViUDOEBvPIg3l2KAebN09O07GVq8cGwD0MxZi0rl0jqgiYkJ
SQGy+Fg7ZiUPRnuNAH6LGx+Q48KWqzyi3t3rM5r4bOFjMGPS8jO5sm6uHczL/sMS5OzoHsvJD8/t
Hn26oW/1QD+Xr3efU0n0j1AZQ8mMhawcR9eHbRx46dhgtvwxFvch36m+1DtPDctdTsc/jnlJuIQU
0rmQgzPSEo6d069k7+b0Ge5OWgBJFXkJlHrU/GROAXO/Cnjgqo6AOgu0BSdFZSwRrFmoivXKb0Zo
RJYdtfy4n7xQBUHlSnwmYPtbBVrsp29jOV/r9GYmNuHYnlBmD0lpqN5b3Lg80HkyQQmwx4GZ25rc
zK9REGYCg+xp2l6z6f6BXcF07vM2RhDdAr/TlrGHLAIYxcC5Do6AAr6QzmN7K54KNVA+vDGhTItk
5O3EXZ56iF1JuPEk1v56YnChzUNtpegol8Z/fGZ7mFmvRqggXPQahIzsLK46LHNCaDCCzyZ/8hWm
ZpVkJDYdJmjWQRHOhSMTbXgN/Wi/W1tyTwNP0+L2snWGx2VDSvszChB7/c9LouRRsUjum4hms5VJ
PudPMVn5nmMUN1RsYMZ1qWEQaQuIlHDX8/E9AwKHK84alFGQC2CGhTtd/o+OAm/Zm22iOAcLqqDB
XtdCYyIr6p1qkGdmavxE3naSkRA+CelSfvfpQQUnLKtb+MUEVz/yj4SUPaQ8uqzMiLrCdGbUVT1r
Qaat5B3BIqKRyOYipjrHvxuIyxpR3f/p0mP3vtNxS4iu8rZWT4WrCGtxMrJbBG0IUJ4oW3FCvDsW
WLJ/3DpDJybYewfm/CVSGLRENLplXCKDl2/qSM9lG12MUQc0DZ9iec9NZUJXQhwvBc4Dd8HenQ6C
o6g077Mo3/b+tttR0V4erysm0dcCyM3rZYNLxmE9ayup6egDPnpTeWLtsNuoKkSJpwbmybZTfJ58
0ynSVlEB71o4crXq9oz5aVzr54s+c5xyUbjNjqWXIP2CY+kSg0ERNh77PxTGx5rj5f+8gD0XR0j8
4+tl1exylZH05r78dA4JT3CF/NrbikJxuPo9wCNr+p3stNrCHiI+3sv0lL3JCUSVNZ10SJrfgJb5
IQLrXircsoiFSP/3fi2YllQQhtt11DDUlafTz8tYwRbBEDXZ1Bp0MdmpmbiotIXSvn7sq8HsqG1m
i6SLY0ZI+BLwcqzQ/rLZLDaRcDLf4ADIVL+Ke0KdVuoi1oziHe8RSG5IEn4VONFDJoHM1Uc7iTB6
q7A1J5AFGqwWdrIqg863FgCYKId7Jr0h6Tk1jvE8Iogue20Eb6leTlHCFBTbDoDJwL20M5KFDZ8t
Q/9ElUJLdeQ9/D6fS6h0hSyrZp1XqhiMx7rPwqdi9BJxazsFgXKzqQ3Url47QGwKsPbxRWDg/0xZ
aBFqXaEDcD45Gx7odecTY4Ae2O4VjcZM0xbbYPAE2TKqOFgiKl7A3IhQ69f09FEIPQ3rLiapXA2t
+VNnPdDhAavQxT5Og9wagK5yafh4YMlk3AZEBPCM0qeQLm89ff6gUgtY59ceHQgEdoXL1/gJaggx
crx6pLZZ06n9NYwFJzjOhYKIbpT9TfBd3v7ysQZY0YAdsIs6FBgBRL1r1tZU/7UAyguDn94VTcBR
4xpUMBz6ctK7GEtEISm3wsljumfRuvAx5x5Yl3nFYtkUCReN0Rq/OuvepHBP+ZinvmtRApx9890O
sTwhr5NLxOHKapC17S0J5/nRnFvtFWPS1DPVg0VNeWHnaYpVBukAvO40ISJ442YYwnrGS9cxc+xB
KQDnAwX4kR/SFOcxicayUSyz/U53x8jEjUuxvNHLdhUEczlvHsIKeQNmzeiSncMVP53e5Bweh0SB
E7snPHDBoL7FNjrOuy2aFKKvFOF87/pMaV5It+78/7sLTYr7RVCCJZKbwMOLO33UfTeN2/GlSW6i
p9WVXGzmn/jrkNRtM2sXHV6aV7HyVOz/9gYnQ9MpimotskGN7J/JHtfzq2xwmeW5T4Myg2xTbF1f
LCK2X62REzHc75hRx318blsTWwL2dJ9KLKY9V7VfdsfxqVQ3FJrRm4VxmIJ2kXpWAECo7E7BIhc2
SlhAprgq55/TmACH6ys9YIcqyHPZvirOcOwptF0lgYRgx7q9lw8PXJoF1qyy3oy9CRB725WOFTbA
j2zyUA8NuL2GpJg/6zajVVaXt29wircPuZhNpBVjAWomjRtdbxjWQxivj4+kIABIlMRU5zV16sx0
j4S5C1+yC2pf6I+Hv0TQNo9dH+yrln//8vRVjERmitjEBDNyQCoDVOZTaSJbW/q+7cT3h4XJmvBg
Q6P0W+vxr+SaeAzr1rwOk4q0dvZdH1gzG6xB0UloYozwNM3UTBY1tn1EGApMOS8h4XPMPoOifjCA
PGYHvdtPxJJ4YkOvdUM7JFPojc8M8JSuy5bBY8Si6syu6/qerCgoM5KTy1OZdBdkY9qzkS7SsbpO
DvgiBuy3NmwEb1LX0/NlNbea/2AEfp+LyMFp5GtVte/n734C3bMDgwn2sDv6y7psKVujEIfrPXe+
DW93pRXT2vnh4BjyL0jNO6phu8ZaKIExIHqZMWuh34UcB8R5/Pq63yuN+6DNCF8pCOBONbdkkJso
G1b0fOcGq64IJ0wXVSUXr4lxI/j2UMnIU34tjg1RTEaqHvT9vRT2553V5c1Udd/T3J+lnPxXyGQP
SISsA8QrvW+AIyjKOkUpn0JdCeiGE3Z4f2Pmmw6zzpNKoGL7/VSG69xz0n2EMftyy8zdEQ+boZE4
YRGZz4M7Y6eToE7ViLNrnFtHVvHp85vWyF54+RH/eSgnboeYPYCkcHObS4B4PmjB4SHeWKceKBmQ
c3CpP9BGsN7tjHW7lX9XK41eb0+4ApmPaF572yMRI/WxhuSRNIGH3WvVTJ61++neDobbW0XpPnKu
y8UBP5eOwPJs8MreNF88o0/PA3+kpCxNxxaeNqCrZ1oYdgH5dOum279eBE71k45d1fOXBZPxOT9q
5VwE1bQva/6av+MRIhr6DaCNh2fLXWgI+HGwWGpL+pSRq+o0P4ZvzO2nrfR2fph3CVfVauTzXPCO
lgaJMZbGsvebG0fTmKSgQG8V90VYLx0jVdaKgg9DkuXg9IzUj1NZR52Oi38l57k8TGWyzfmbxJXV
ppvLpn/TyvZZqSWIHbj3QQBHnafzG0s+7fka/vFbydI2ExZ7CrD1EbCCfDVIQkG+7idj9uPLLrkm
tvx28ANxdJFZvhu94UOWtX575hs+OEwtkpn8rUSH6vnC11Ys2p8+OOeltUOn0WdCampTMoOdS7/O
DIer6WFsWWLrb80+DlgzJ/rvb5+Iep6UF/+LQtnRFHsjGrZxG3VenHtihG3UbUEGD8Xar2R6cBAm
rYdL5KNn2cxLhrA9eODb+JnodoLIUgAnK/ssH4YgXA7kdxDP1StfjbNXTy2w1yCvqpdQVSTubrtB
2lRHRi4udCT7YiIqRAXkmHuITbcbfAYoUtEzFMmHsJbKx8dD2gE8dBu9tpaDuuTeyvkyyTiQjJ6S
PsXJO+uIi8gYRMWuo/UahSUiow+bs8IfPBj9tBMIHcwCZ2OYsyBpL/84fOTgzeegPChIUS18uOIP
OQi4kMjg3Ozb5xvx34R04Ot4YHdRpoAuzUjk++G31EOdV3SrJJb2NQXsQJlru1ktJdPQJfs+myDs
IP3lvT3LTJEbsfQhIPl9WO4CTyLcCGL+X1fT4kcAyiW3nCWLlT7lS+7zcTE8XTIC09vEoJCN2L7u
VMQLrmmP5wnUVXMI4Ly2mkwW/8l50hidWdWFAijtXlqPtQOISTbddg2QURe1CGVlU4lvBf8e2WU0
s9DV/PNYonAGvyRGGTCi4oqujQda075iKK2ZmLCIszgJ6nOMPqraFO9rkyhi2SQwzigYoBMPAwVm
levUqHNgJAXk/l3zZXoixgK3FZBXFobnM9upmHYNl9MPUS82fpXzSNbfUTHNtsNpjUQG83GDLjDZ
NMpNoyTMnCYylqqOadmzN8WANFOPx7aUS5mlESO9q3fyxoM1Cs9lWrgBAPiegypERK9h2ciqlAtT
5Tn4bQtY9Lg96NmATkbULJD1AUQeGCxKWTJPfUpc8dG0W8Nqhi7eWgNICmwJCygUNPH/IWTdlOtg
173DzP/HaQIC5wUY5tD3znTNHC5zp69bLqnub+P7ugy771hTM04SEVjOA/imPoZuptF8WSQsMYfX
7PA8iaUwlz7XoNe2X9VoK6JdMdngoZKr7ndPubJVjEuMNiyP+eVl+K0qQRs2XiOCdX6/JAwu1JJq
RQZKwNlPsj1xY81C7lpV8OuPhsncQruS4qCEZxc5kzkl4+joLg+o8u5Kc0MPhVpM3qM5zuhDGiP5
7xbuMHvjW7/YVaC9JsdKmGbHAMn2sH6fvi2VuyZC+qgT/UHApjcIwJ31Rzx39z4YfvV0pmUUKlFq
V04+/6LK25OrsO6/E9CD2a4ODf0XdkcSSPEnMVfPnyunKxFdz6ZZB0wk66Sr3wKZ8WNtAFd7p04g
XgyPNa5Vyld+3YzBxLf7QmczW+hsLY4rDc7r5QfGbc7soHqAVIK0sUMXjs3hAabE0pTYN/keL3W+
3sBCPbZk+/04hdD3AOluhZ3a6rO5xr6btuVsDZIvKIimAm3aNMf8TCvNH3BabTNmL74XJYNuHE4E
uzdHjvRXKRpXAhvMIUv3RJdc7RH8z1c8yaVoLTYuhGFQ8rydGWeZA2KvgUPeXZipvy5yUuCu2vHI
HCDQvhDY1USo+sIsj7gT7tjmP78vyHr54jyimqD9HFD1sU4P/80ay7TfBh8vNKV5iX1vCy3wHB2E
ANvS2h8ZffoiosAyR6ZXLjXW0L9SK+LlMeNW2/IQ36vELFNrJqZmze/f8WwF7cJ3NFYXrASWENLI
t8BpaQ1926SZTWEkX0UrRHMJT6iOhTUI2dJKNvf03l5O+u5YkLdhMTQVPKMSkDWLrPfw5mrffeTY
XqUN9s1iOcTg/S2QcAsZwDBLjzH6hfeJY+Fm2qJwE8ZfxWUUhPe/42ruDu2poELPCC1m64KymLlG
NmrTg0WVQiLnLcIQaV+RfdVm7fv8puAy9rk0KhTYZ9wfjHVSj0O/+JPRZjerwrOSMrhNm3RB6VwI
gTt3UFsnAxZZioYHGqLbYNH3IvGshftt/qidCI6Fp95PPQGcjUOg9o29RLUNEfHab27r9JcgLA5C
hM15ATdUetjySXKOUp0/gRYYSNJvZE04Vj6p9IHw5aKnalWj1JnpfrKlcQtdVlwQKAIqUHYvJnO/
oZbLlI9A4/KgN+6kYX/8bwiR57X2CjvaadL3U5C2ybu3MzAsq89BgcH5GZFUnJzrC2mMOEb/wvpb
ouU5avnt0z6v/n1eRnPoRaklYF/CL46U36l9p3D9s+tjdnhJ2DNQRCLXoIBh5f3RaIlzb6Tyouk3
jHiOPdGz5eUylhplS62leQie7R1aa2cBzVnHTTi3KRLzN6ysjnLeKt4IsnAPx9zpx6TSJpPmEZlb
qDQP6DZVfrpYQUIMU9OqprCA5C6Fiy7tbKcipkT7951BxJvZYHACfqQ8vUQ3RQ+IDc9DQGia27+a
SS+KRojEchqpyw9VtduD2yU23wPKfqcff8eB2K77uSLt1mTAxoGIo25mqJ8+dQOrHiKPDECT/+bq
nHBRN2TT38VG2Cm2zUX1Lg5oCj529pkLPnHgITs7/A5+/jFVhoVKEOD2JWuQq6jA2jWxaH1MixBH
Ugn57qDmhTwfZd7AXtGrC9SvF6qsniPNTKJPmsUnTQMZ6K2jPkx5XnScTT3DKN3QiZmyW6+i8YUG
fac0dTRpkI/7o9yi8xeojTqGT1PEhEKVfLYEWJJhaeQIoblhq8EBr2Ho415mpCZ48MF2083hKoQ+
jxvX8ljeUOPCntxLwfhW3sPUCTVDFnc8Lt9NeqfosGHloUkJMw+nHJ5JhmgKBEemny5N54GN5UsL
uRNxbLciDBWb6dDClhAsJ8GeWK68hMUxm1U1e3LAovhRtJ0UMeHxXi1fSnrHMAiUrn+9OznE3lyn
0atI59EWaP7Q9JzbdNalmSYODj6N9ozRLJ9baswRUfpzM2tKniEO1Yc+SqWr2yQjKsNGbYbo5YTy
w12ddUVNF5r9IReRAKTAtvFCHVrsnMywuFvZep9o4vuRKiUGZ9kY/xgUUbsWTUzoG3wGGT5d+E2g
jQSXSkR5VoMkaXBfaF2jttlNbem6f04+g9coj20fnzHVn1YYxRXRom36imBCxmROxcqJC0Rxoa/D
3aqxWY0Fi8nGBKuQzHd1m52KNUnk53tNN/wleR3LQE59oNhyzOv7eyUnxwPMpsz5Psob0Ei/jA8x
hGpzGKzbvl9i3eONCKDi9eHULAAgjtd0zTzoXFEdg+DuSxbNSXKwxy1uw6G6UbLmO+e69YsOH5mG
VpZ58sH7dr8q1j5tgPoznKXvHs66cIFYflRLuwv0Qxec3I8IGsWMII0o7U/c9QMTtqOAFJChDO7Q
JHID6LR2G13fWwJ+PGdlRcrMigPmy7vnnz01LfV3GT7ocEel6PwouEr/BtY/QYqfKfrTMx9+3hNK
x2/uX/T2/auz/lPwA3IzUvLQN43R0DwbtVbxFE8LOHRl040qK2uWMaPFTDh2/oEA3y1R8WHFMIso
6RcPHH4aZ9RRnhkREyQkmeVewm9MnEaKJnE65Y1qsQN5GYT60Mw6JAbXU2IAW/x/LOLCDvhON10p
3wpleLreg2R563lcR7aNHI3TyhX7wVXpbKEYUy4eqDjT6xJfA1Ln3SJswga4qVfcBaUX5IsXap0Y
GSb2L1v6nKGHNSpCyzQZA5PeWzvpqCEjuwXTsUHRGFw+d0OEatRHcTQ9VUPBBPVWBeq8MmP4HUGc
AaAaeYItklUcLO3ase06GKWkaVVspu85V5LpTtRC+KuObDATS60z+xj3GydetZjqWRKoXxSwwgxG
z7IAjBLn4nDZzvBStGG6k8PlwGwnQ/aKCgk8doBNQq5XUb6a8p7b6hL7nU8gq4BoIMhLLZdH2O6O
V4POMErW0d8ujhV2qozzhmtcwtX7r5BB95WDByJ1HU9MHkjzK+KYLXpT+ISYNSXPdvRF6aWcYyQu
Xkq8GMYbuolfIXGeS+AaEf27QCKFrCu7OqoUnoXMbKR3D3621jRhi7YdMqDJ9Pz4a1L24vrtQ6z+
YGXx5u2+mcruAUNN+IE9wf49i/hbqBJouTe54D7IKUuElKuwORoRHvdxoV9dG2d2JsjiiJl9sKNe
Z1aTWKT1jHeJcPm5OslYImy1d5M/toH7bg2vmzOHtESNHFEUw+sRvVHIXNMQv58c1/ig94cG8yih
sUYPddFXdY3+DnYVRWdg0v4U1UM54ThHBzIkbsjxZix/NILr4BoNCdO6Xjp1NvKKxoY7LvaQutcF
Ude+H+9gsCSOEMAqWp58yEgUIhewkO2YJdjgaQxKfIzfHiSrUAzMLLVIWQg3Qkmor2jyq/29yWY6
RVX1H/yVs5F1erraTzVBv3wLH+cmuxqiNt5I7n+vr5WI6etefWQ7uFrpyYgMfxRXH5Vd1C3JApr7
v75eONi1MoUejzImD4hx1S1wdf35HcUUQmqKnD5OeFWhCkYRUVDlDQjnd/bMQsBFbb6xNBVM659z
JUiUUzgyFduSAX862BaQWFJ2aQ4/L/9YTJnhRMa7vRgUYr00G5RMxuAU6vfkAtW/MiDQgxmBwqqp
L6BDOOEj+VPZ10f4Bwgdl/sQKPNTz1+WwdcDS3O+XZPj/0bTx4G5oSmWtHgFhDDnkeKYZy3zL/4Y
J0ROzWVlz16F7Prs9iJy7cL3M947RC+0+8n0ZVBuTiU+vwHaOhkkUZCCnyqOS9jVgIJo353XOX5q
89tPYDXrjSVFbW/M3QG0Eaqv1g7/6SJu/NhsfFShEqyokFhrvblhn4ruU/NQsfdqv5JCrw2BLeFh
tILrbGsZJgHEuBg1yJAilu0Bra8mdBISZTOG/DuXUOWm8hg2f1J/W6qQn7Eq5D8KpWh9Fiurjktr
syjuYWuyS4/Sg8N6ff1bIl2U85iNFH0OhigDxcCGkVWGQmf07j/79F9vUrvinZLGPvS9cJtMLwyJ
kEW9m6rA7I/9tXUqleDcmsj6j9UhwyaqDuaoIjiicwsxGi6JMN/Y2dUZJz7/PuiTQd2HNTXhgHO5
qEpLJ9upsoYAX9ciU+epLOUwOO/P6JCIWtBaqqII+HJjnqs8l3LLmfp0vNcIVdas3bJ7dJczkv3b
wG4q01WGUGNHrUo+JEYWwfECramJcEeW1aey/UFzSu7aDi2w2nu4rlzw6hz009DjuLvOmXzYj/x1
nrK4cRrVlFQoAs6VIZhVNF8CnxHhS4xj5xVU0mA5bfRZWfqr07E7OqF7phzFHOZjEKtugG+fSaLE
UiTKUpHesWvro/RTFrTpKCEeeFEbkrYgcpPB0Z1SdFZIGFcLCErmmKONHfK8T3odIQeQjKojVAIq
LngUJiWYBG9CtOXyWN00Wh9ctfJRgJe4X9888jwBDSRHVenZw0MXpRZWEdqeTEa/6VwPBebpZ0T6
HNT0SEJe/kTUDTCDWDU3FCIoqoOTvcpR6M8C3EWpXcHZ8DyxuWuEwZSCw1xRTi0DL8VlIc3tYyN4
MrdSNwnHfSX8qefczaE+pD64uUtrQkH4dC1t3An8mmvcd0D4X/tJnSGgqWv+rVL0BHePPS4yXC9Z
s3Yk6LIAutxAD5TXVmpjuwgCexppiwTBJ2xpUYH0GZMRYkDP80mz409u/aeesl8YYcoQjUYwz9Oa
5HtWrW3L0bXVIVRWwVcMuqokt7EbbRUDw052q54tEuPgjcorrBHdTg6aIcnSJnGp4au4b5baHK0e
mz9aGkUsqAJO2FtZzxDrulNRK6K6oXg6X0QvjZ9V4JxYGfIapteJ9FDdqlFO8jyNc9OkkjI1gBL4
PvcbUIHCutW79PELtoPoOLaj6RBQI87xVV+Mh7Y9AsqomM+Cmtlnp8gVbzrnKc++AAHNGOyEtHj6
NvWPsx/5Fmfm3mD7LqDuouPZ2s/LA50C/aWlJqfY2uY5J2K05M6wScGFNM/g3FGaP7SGxCAZtdNZ
4g3L5heDNtehy+VAA6adIo8QtLf/AiM1DEqKqNNqXHtoy2pCBM1BYFCoto54HJCCC0HmeQ3zDGcR
azCtXoVpVxnKOvvYWVGlRzbkePc7hehAoyYTMpG+G5rLY6cOH59w4aflIH4Eue4jrpvm2ToP0eYm
D2Cz68S3J2X9ZEW4UgW1KnnvAkfmKtlbctYrdmeaMhD2pmLV98MWYxlnWtXvVoNnfS5an0lmLMVq
lRx7Irzo4M1ud0XqPgwoYlWX05DBRMj8Kg7WQ9I6BxVZOS6KA1eGf/EyJwiR0g5qkzRQ6f5Mr/CA
lWUIcFdssyEac4aYEr/+g8ZRHs06rXZDb17+LETenjKKYfZtigmex87qhILmx/k4t5PtaGXw1qdT
MpavL/f3ndZMw4gm8gklP5Lq1uWsy7F30DnSSxv+Xb3fCSI7rz0B3mjd+JaD+ZZ6VP/X+qbeF03J
8yh8WBgjJ8kF5jn7id4YEJKuy8lsbTI3OxoyEgshV1/TI54vBSNO7E7cwTXiDAvu6yfFDekEna1B
MLVSkZzCwFR61EbYXTE5ed4pzCqq6jjPK/9Eex5lI5p3jhKL/lqC45UCwaP1GdNGd69WL4ee4UQA
6Otxc3QdzcILbDoabmpuPzS2Sv57FgYAXzJdoaa7AKoQ4Wz7ugjLAtb/ZyIRtQvPUf8WzV8KwStN
YRs6odcHxMOMWwDuh3+Ttpgo9iQ5VOBfQb0zdkKpNih3rd0nyKFmDyzPKN8Ff+Zhjm4pFZiOia4s
K0SluGUFOjaUFH/oGB+t8EZbFP2cF7lJNe7g7FS6V9kMjVIKSS9u5Y7t0S3hatlMQJgER9MLPeBa
2WYmUeSCJg6GLpFNG13PVbqJs8YXeWu/OR3E4bE1vRnGLpLM8IAx8TKH7/FtX9yr79UuhQNUv0lk
DcZXTsq4gIpWOzbQkutp7ZiOOIV9VG0mLLA4zpdw9B6aY66jVpJ6FhyDkxvcZ6+aJlmeCibiuG8w
KRiLwfiVEb9SMxUwgO4TrtWVebQ1ANx+mEFM7oPgjonB5v8lrG7Nxw5DHldDSJNcIW1RPTiSnPaS
bbSxBcJWDCD6TnhiwsLpyHA67X36LaNQCzY4nengngdnuvvuDtvqaRVtWQpzyYtWyyFFZpS/gxCd
9JI/uDHvtYbJgnzTvY3Qd5SHkXtvGfot84qMDn8tuCyePC//1EyOe7T7l32YrNk4tdegOWUDWCWw
Z/ei/1NxtYkN5xq6sTGy8XClko9EdgCNuW0b//zMfjcNQcAghRtCKVmhtYB19d091t5G8+1Na8J/
5L6qjXp1GMOQUNPQaOWl2nujONc/ANhdaFBWJWCUNdYHDgJZl1AI7f7OUFtcu2JtZvznvI/zlGZK
3AvyujtLi6T6XTYzKtBtOY1EHap9yqytJNkhMNM01U9ErIL9lcmStRCnHAx+Pb1IoE7cY4rd5kYG
3IbneChW0xnuNzdLDAxIASjZsJJOT390nORquIrl9rVs/7jOzQmrfkKIcjUelwe4fv4SWoNyxx0m
3Oh9iX5dl++hBL/ig7PmCoySFzCB0lVm8vRaW/oTUCqQ1fudBduzqwXjym+T+QfuerfJxpL0JN68
LHFrT9Ak9wTprb+tov8Ku3Qpor0WmLkQ+NYDkkAPFO0NMJrrj80g/qwPKi1o+7bRlaA+xIKawqgt
EbUyljyxVfZGfx5huKNU9NeYHlTHs7hRDHU7gEy3LyoMDdZ/KNC9gUbD5fJ5d3n/P0dMtl9IC5XB
6JVzZcnO6DP3Rppn2Wgt4l4gF980HGTTvNQ5iahWqwNq5mAZkpjibazjU3N5i50MsZEXMMjgUg+u
enLIevtbGzhrZQcHu2I9Gq3LOOInk/wRkFcf6cFGgFsgg4cnfePR+fwXUpFMbyuKLXneOfPUR1s5
HDwm3eEMh7a5COZTdb+L6OPvbgX6XLUXT0vphZxRa/ruTxzjnwDFLtqWIertNh9w7sScLh8Rcbjd
EGcsPXEgOK4Qah2dbp/Dpav/eiuxc24qavJkKijXKVlGMkgiGFvknfrEBwQrxiKG5ncAshBgJu91
LS6dV6tUjkxjP3HUMloJCmq86CTXnViFl4WGH4hAg88uymByC5xuSxSkQov8baEZhCMGPiMjsEgH
JGNuYXFRpuAL0XaG4m9aFz7KpYgP35V8uZf2nj6U3dfVK+A40deHIkHLOpFJ6BJrxwvP9KRY9oHJ
gXqJd5/bMQ3jsYlQvFvbTOi9tB+iE9s5NFTSIHb6+71OdWt4Vpp+q23Xr0ovH01E5dRUR+oTmfUf
ekB9EYyPJzDHI++NSwJoZxXhT6eyHAEwNHzwh6peXVfXNWlEgkkm7qOxSsy0eLKwdqMLSyA2I731
TNOmAtfzDHLPEFdfPvBnG0fUSn5RjSKxabfV9mSsOGpeX/ke+U+G+34AshigflBGkCZJNwwFg3X4
vjLEkLDqqY7/uuIrvv/A9d+2NtZni7vwAeVKkjCmEupVMQiWwub3tGw0sBzM7Fl6GMgRUevxbP3p
ZAB3XZQOO47JffibdEFx/Zt1PTPpVBx7Wj7+/QLuRSATl7fS3c4wx+94rMp6KydR8ZCzg3HFuQ3f
GXaV4xXaUeycPZ9Sikr55qVQIGVUP6MAvAq1sWTm+c2FeOZfTM0XDSG9wDUBZRBjTJLKLOClssBl
pbVG5kFNh6k4/tBZYnw7UyKXZzlYNHUN6ZeUhyV4aRUbTqvaj44eo9JiLcxLrDsDgyQacWE72aXu
8JNQIrShn+JHbl7hsF0QLVquR2e9I94t+Eg6UHiwfKiPgR+un0Ejn4/IPlnUfU2P9/sPmzZstb6/
4v0LqX1j/02YQGDfS95piIa+vS9uJKylHMm9aeQXFjzP3vEGpyfqfKiKuat9kiwpdr/JJ8aPPA/j
YMYz9yzG9dMvSrZ065xwD2sPZ/dGLxM1jKPTu1VAfjTwWKH/yqwbq4L3MlclQA6SqO/d28VKvH2d
eGVJoKxf0+M4scOZoXD0STeaWhzk4Ulc4coPZCbMfWV4nUJ3B4q6Bam6x//QJvCvI3U4lJqbdgCo
X2pRh73Z65wkmqeAQIIR219bxjgwxgrIGluX3jAPw72Lth7iX/Z0cs0KBz941DioJRiwTf0IGaqY
bL/tHNHi//3Bt+hOoBlT4MrPTupnwq7ZZahGm9UlCtBekkNfyBZGFgWj231oVO8Sqx7aYNfriHnl
LdB8CpTUrXk+ZUZuRfiytgGXREF54KTYJxrRPC4pgG/N3bC/oMWfcWS+G6TLuY8k2XDY1sNMxMkR
U0F06OCORUCNAaCOPm3L4o8EQkeGgWPSqwNSGcHNghNdN1G9gdS7CPPDu8W8lXfKkNTXBwYxunDC
4V9uIlRX/AfIMWu1P0imxJTrjY+tm1LICFRw/jyd8iESIcYATzvft1ISta6xBp9zaDz0W51b6Mfn
RVbuDj/06QRs8SSK3ux46IAbNZgt6m1zk4wXvQG3mfwr4J+3004Dmlb38Fz57adue0M5XPxzvrrY
jxEMlNfXtcr/svR8j5xDkHu7TL6T99GDP0JheACVG8G2whGVfQbJDlGsnvJrQlpMtFHRr9VumdBm
J7X7peWtD+GAZDp8hcHqdSt/xsOy7XulT9CsMfooDmeLIxUm1/HhWprtc3D7b51tXBCQHwoobE2g
YPqMouQY7AAGCtZznvnufYfe0mlxYDqxX6qr0m7/4wEh0FJ9W/BsqjXY7XQBoH1Kr3Wt6GXQmTzJ
SX964QoxaOp6IS6jk4MCYPruVlDEY3NwisNY6y0Us+ocwxuL+2Xj9ku0g2qP0L/Q3C+uPRYv9Jus
hJr9P10p4MILzleKpjqqvt5hFPS6L+skI70aOEfyEKJuxLNV15XP7vPDqHeyWZu8jUQIY0w5utnT
3EqTPGFfgqFQD8S0rl6fKA89IWg487HKIFjDJHv+WuxbIkRNMhjtZgb4FfzjgPmmZIPQygM+SkAg
h+f5EDJDDu2tqdW+Omzmccbg9pdaLm0cZG2rPwksG2tHh1lW2n/euNzyeGOWSBJR0o6bDIXa71i6
5A9jTqW4J7ackZh0oFfTe/8CnfRY5WskMHRnSWruAi5XWF46r4hY6Aet/6qbagFaFtm3WAstXUGU
F0u0yolXgUN8jqYo7p/I1rQNsiN+L17lKauimyKnMlL0/BQmz78GJBY6YmXxftSw/r4P+aHQEWpP
u9Pmc/BIXSknJmEvzg6mFVv7EYrQfeQbpvfaLwcapqtlERXM/4ls009cdgTYfHR9wJ1y+xBMAhPk
cSwdGI38zQbFK2uyy+sXLR8yAdf/dmji/zdt4Uw/ZoFzqMhTz6pp90BFU78oQBVofxrtqqH78tXg
BBXIcfnMf4FwFGQec6XT5GaaUCVH3GspV2iZNqBxorvDXuPDapokKYQPauCmDJdP9FFim/Ez5qhZ
trhB3gWYneLLbMN1PnM4BKcyaScjYeIWxajWRlR1iQhvS8bjGgex669gkb+cdhLpNnGyYyITPOQ0
hHnC7uwR1iNHphezp9AbeJR5t5drYcka5884KBJDX4qn/Olv5ygQsx1/edUSC6GJ1Hxkrt9rmA7L
hJjHUQzUMsrY8NMjDhVHPgMOJ7+9u4JNtBrhRm7ZhWrYLsJSyJs8G3O0xQhlE1iJNZpEUWkSl47J
ZhFFxaapIPRFoR2tfApFs2+LMaLu5irhUeKpZ92MIui6tZuzzhlK8R0DShaDNn26vh9ezKOEEjdc
tzqKcdPL62++SzfhXdAAxDw6BxQ2PoaeFirU5nsyFTuLoAbFkodaZ9BGobAnwEc9FIZ68P5cbOXb
Y/krTzmyzukOEmSeouiMDA7KKLjSK3jol7JMvlkEa/tsZmgzbsZtAzslYMYO/23QveoUO3gagBQJ
7Yu0FgV3xE5GQr1GidKc99LMzSISapoL6F5B62Is1S0nM42Keankln4FjOYMT7UlhlMCpnZmEoTc
DEbSlUjUDbMa0wOPlwmApL+xWMBq436hcT8a+RLiaB0wGPmQBB9TqtVbV7njZ/qybgxa6zFN4zjT
DRJRwP5/+7J052lIXf6XgprgbKsoI+WuY3AZujO6KZu2nHwwYzZ9uLgvud5hTYc0neps7A3KKSfh
cP9EWsxrfwe29wtWzEIxmrdE92LDNIgk7tAOlRv4UcgdDgd48kv68Ez4736eugXwt81y+52zhGJk
BggdMyVZ3pS+hmk0jhMxjzwMa6G+SEsZzBWVJoG0n+2pls0o28K1AhcxTZpzgKlenQKEdEyDydXh
9OreuVrEfI8sZU1LBYFgDr59YkGAUEQjXNMrKGHlvM//jLp5ayukz/jS33ELAKs8w0OcLmMG4XDl
HywQEqGIlOgorXLc5m5fVoHxxfhcyf17B/fUJUW3GZRfOWcW0tIPuDaHJTIVyF1jhdGMnCKiZj5y
W8cE7GyLOlnMyx43loiZhivUNVcINdkXLTrA/K/0G83JIPOzVAO45n3jej+FN55+XXFb67PAnDD2
SYA6gU7lz39qE/Y17UtPutVscTYJ5cy0rszAhqUdfq2Tmq3mf4ohnzw4cruft+ydU5L7kVQ8kTgy
jOwBQEMOsFZo5wQWykRXtY1hTmp1zPQVQci1KiC+kSG+IvBTo1C8no4lqCWBze5hOjkPX43ZpaFy
ILKuLpPVHh0raYX1aaLheQ6xvTzJ7O1DjiJbRFFBAiUxpnKYRupk0MOys5XWwtinm8Gc/7i9GYvB
GsvoNqJMjIKOWKNV39nn+MGB/77XGtbu+Vm+SyBJPmiKNH5J9wdh1SWgGxcPzyc7adEP8Lp+9x2H
h92epY7/eeQMUfvZmcm1LwTU/QIqxeV88y6G0c/5kEioPtpGqaHqPBWqSPVThdDrK5KMADD1ubDk
wG851UgeIpSGniJQOQ0xoUn6X/p5me0Ex6pArpI5S/e7O2Gxe/9Yz1OR3Jh8ojwkINt8nM+/o0DU
9R/LD+/BH/usoX5/eCwfWjkUolfeou6VBzV/6LdaB6W+7y+kgHwsI1Fzy4BK+nSdB9E8UACLSPFq
wQKAN9XsAigR/q3BL48GZLEpakRbe/oGVZeZVyhPRiFoOy6Y36Km96tZs8LuMsopXAtA2o3TJ+PL
sLzEr1wUqywsLKJGfPFCpKwvfsCe8KdxygkwK3VP8ssndHAScTJQnpRngADRUpIF+t8D9rseUlAj
ecRc70GZviu3OfbyWofKd572J/NjZyOP1u9nTZ85lCtYML/Ob86CpWhvScq1QxYKqaHLNY+COy1/
yUfXVzyHyjbT5ElJYhk5ZcowSS9Jd8/++jpkWtnKkGd/SD/apI3BGNrWIbZrkNMSXBMOVmOskUZz
mtHZ9ztuzed/oF/Zt4xireaQL+zD7PJvYEUkqIfuOs0DzmoZn0OuACIjgA0S8TD3chPRu/6eFFnA
bZDxSemdXO2r0CJnl/C97ORqKXF4okgMr75BwKEKl44hYUZHBxTiEM5cSc5cU5WWrj7asQTwJoiQ
DZbKwaSLy9yoxfJItQLfVcXu+/MzPS1V/pcQuLAsPCt3cctS8r7BGtEJUV+LcPF7CHngBkpwBSVX
k5bTDFeainSpmIon9ASVdMqA3U1X34MNalRcmxJJ7YcgTzu0B1fCQv/bP8D9sUFUaO20BwufZkbw
vzVjLWntjrkr0D84xi5TQOnBak38QC8UNmT5MUaXN9jclepVaYyHGmJU75RkVOr0LQwwC0J7T78y
f4LSK5VZ4Fx49x6bOScP6ZGpgGrG0eYnAdE+FdAFoueX4/2U9/HvyZWg2e9jTqrgU2i5kDfmF4eh
PkJj9v2pTxChx2HJ86QRA27nFYoFi8fEmbwBfq5AJcpaSdeTFB4ccCNqom24Z4AYwk3eXjfBumIa
AnBCUd7S9032lfnPOSuWEHJSEvuq7sPZSI5WNq55mk2eI6zRvVXhbJILkc8I43ArAADwsn50biwj
sAsxuXprJujeOG/d8WnRFhZySzfh+5ct/kOb0cFtk/hxp4k4vO3zTDzqA3LocXwcjeMNqOAfc/wD
9SiC2jDmV97AmX5WHDUhEgmt0PRTy2swtobN3k1VkFZmmqxLfyTu3e623LMGGAz5od6c/lFtZVkx
PssBdV1OOlWU95+YtqHlPX+16NUjjAN3NO9KChyN0zTXYIcCBJe0I3dwiUFq57/nfpmjhQXpnwCq
77d97rPCzyZm9UJx40qp60OjnPOwVXf4mjXTZ1RGFmwwRHycBjroFrRUpUaiO1E1/Ym5DvPkXhbo
ujRTdzE6mM7Kq9GNaypZM/SFWqZt+App0EqEkIm0heb2XsOH7IOHU+WBURT6lxG67eT9N8vjx+v/
cvBMA0xco8j/Y8HB15q8lFOZTzLiJwCmtK2td24mwSkBHXkgv0pUM8jbjB0spb2/bWo00iu25pFx
inPYsDh6sAWlsQ0wGsEp3zvio5FRbX/7gm5wkrXUfQt6fbsySR++UJOoy2bZr4ODFDR/4GdlBo6/
6baAIt42bna5U8hFusJc1k77rcD77ZLW6pGqfNQ2O5r8uemz3f4riMXRgpgAakXueaJeW8rA2NuG
Ra36JQf1EWyfBWrBIEfXDvHcLGvA+wr/5+Hk2PZ/Pko7iAFYRTHsAoTlV6zVTNd25rhbNs5xyPor
FY2RcX49gj7HnTHYeDX8mAEl3J5rsELJGg8KqIazhwM5l7QatAGBr54RTJAt09/fzYVO+uLixWXW
UgzFgqfOJhWWBvcv+gpBTBjUEhVuDX9mCTCDZEtdzSm9g7kP/fmfhQries1hD2+oxHRHJ4sPjogn
qlizaetl8annzarZpUqnrUQRb3sRXoFNyRbv2yq8dQfIrWmq7TgrPbOjgoEC4AKYnovUVEXeF5NQ
OUxJMzavtTJdZRJp+n6vddVmpdYkIfRJmpOJzV2mvfVvv2E9OXPpXbOcGMsxw1nuXNziLIqX64/H
t/W+DlqUoUXtCI4VOJ1Nnivmfi/p69qfvJVnC03B8lNLkrThXZrdgiCzxsQ9Nf4R3FAg9xlZCLVC
N94Obm5QzPVGvfOLwiGYEom6bf2rF2Dg7zrSAG6Yi54sbxlngAnNzdCDiXldcjRzvjm7k9cijRcP
x9+iPuSw9dj801M7rtsKJYjJlCzL/X7I0etSpzimCGCNdJxWQxxOYqc9iqnKp7kdUr3VBYvOjRXP
INqdPjfod24voP4fKeq93sUMHcc7/X7vsJeQ4W3fEJPevMMHxnc1F9czp842Em2niZgJvutnPWVq
C+YKhNexvnniLBG5vKSEDZDMGXxPmiidru+0wUXPxRDbJhxlxdX/BETzIwRd0VgZByY8ECdIMAuY
0nnOFEgmLXsK3F+7avIXT40yWpUXV29Bp3fzA0KT2SyYAsxa433IXttuhRGZAsQ//iC2hI4V5NGF
WlG0MiichF7ELpvTIdbQPmAOql5Rxa8KY54Lxcmz0LCtWnIvwhgEMQpIAQfYxb4j/DftuhjOZxU9
J8JSBYYfQf0PO+YiJWfNZXd3zkCRLfP7dpdZjQaXQdCQIfYTi0hxU2Yuy5y2h804Mro1VlwqN4g8
3ziUJqeULasP9Rh7qQd30PXTQTkQmoTWRM4tifvhHsrrZioXrwHIdLgLJ1TDZsWrwVqAlMAiVU6x
sXgPEm8tPJuai2AIi7y57VT33FmxoyKd2VRDfia+mJ5NvP3jbeZ1pQ8A0BlnpQCRMDrj/LQeHJhW
OU9HkgzTUx24MLm/yFWvuF+gA07L2eD2V1RNfZoMUB2gzJFhoBjY6TYzFvX/Ccs6xIUz/u7gvtH9
TEO1Es3jieBEBvQWK9iObS3tYGTSLfMTTgV85O+KIaurBFtfH52Q21dZzpZvJmap3LKbsMajCBVE
rP8Cs9Vc9Bzfd0yrqhox/44zOvYKprLNRhGhAwzSHtSfRz+fXzJjvqbgbaMKna7cPKdJMndMEgo+
wMKclxT6lrkiWe9b2lHcjBasRcuCBXo2H5ZvwjcGI4ElIj5ZzMppuyVIqBz7WpeCJX41ywmxw/Aj
e8vsv+wjjM33Y9lOsUbGhOUwAY0OQJoLS07BrS7O1Zig0pq2gM194X1OKqPVNh2yxtVPdostszl2
/L0l8YT6GhOwENDKuD4lBNZWXjKfqbruu5KQsyir2mNPO7tiirior7bRcyqO6vVUjRtRAV8TIs4m
tluypRIvASKmV7hiQv+nNl18GcubCvmycxNYAqNDzLj/29JIENhT+8mpEvXbUAACie+tHtPzISQc
uAAYcLsIqQEazk/cic1jNzn7Xop2VUEM8VYIMuuCadYcK2Uy3zyAJ/s9XHSOfr+3X2IN/7lyc0lz
AQEiWMwPc/VXQsFtDpSTTxOmXG9FjIWFdT5ICVMyZ+qVFB2QSg60tlZZpalnzgk+cYdZkClaWls2
WeyFkZzAyLuT/7DNo2wle8Dfy0v0zNDWJas4VJ5q9BEb+jH469EsQn5KZ5bNyZkwuhGDrsAav7d+
azNB3oYGV4K+ntIkbicGD3O2ZJ/5fJMn1o2D9lE3q0DB3oNBIXQMvWcBXGxJ+sRno4F6nfmDDwFa
vI9jgRIf56a3qIhubs32asTUsPvhuKFotbCuFAFVbZ4gzLIQpWUZdrmaT4VkoVGfOau+3CI4CAr/
VZFSUzS+S5R+FIgbyp7XrprDmQ2VgMBAn651aW20r0Xd4kfKkgIJ75xbmIQxkd0+A9yDl6WwfRfk
zqZNgiuzhePFtXyVs0KDOfLKFgx+W6EDT/HcESY/8lp+nDU/8hjnMa02rQjoAydymJuWAGsfARyz
1DHKSwabVilCYkfmCwDryqyUom2yPA8RMPOedq0mZLI4sX4c9vnu4x+1XMBKG57GOU57qtMU92ZK
ZBO+lWNufEkQv4xxdpYvGb5tDL3z5JxAnvx6IN9zUBReO6FztxPs4qAnzs4tUDbrd+Z161HUkJF1
BLmOntpqeW40wd7dKcsP6gUZQQPUsyciOy0aG7yxOqPuR1AXXlkCEHtCnGon3rcFvu1/G368GS0c
xq10imx2RLu4gT88IM0+Q4ghuxT2N93aP7ISayCqL4tBfN0bl6hg9Qyd3TIAsGv52UcktpTTmwQv
mR09phS+iI+CMeCccjnXI2QyyCxbHMe6+JGsihEFfiC8a7xFOARM5UM8rGKA3JG381rU+Lz3eAgK
cwJ5ATX9t+enxSrQMcj0lVu/etieOKwU0sNg9LsndUQWGu/9QF7M5Cw8D7WtWnK6QR8yrHnBTNTS
JQmaMx1ITNFJwg5cEh6bt6Y6gzKWOBx8SmL9kaL3vuuRIekCUlIxhrFJa0BkqhpcHMtn1IYaFzoy
CAWbwV7MJzvOV42ESBzqfjU6B0Xkl+OO01dlFr2wP2igFWzCTBFeqvhqlZzsz4RkFvfHOdPhUQ3X
BPFbR0U1Vwry7O4LxqB/+xZTFSyX84DNMN+HolpPJR1aYvl9bOkaPU4D9AV+0fdi0bMJygnY/5WU
u55poCuw7s9Zhwun+Bhrfnt97LwhWT1Fjmr4BGfFOPYpMDesudhLUAUiMoE6qgr5m71fLe3yMNv3
Nm4P074Giwtjc2fORW0TXYCqyze1FujtBTOVLo5ci8Pzo+KO4pNpPXU3jXQGtJZYUqYuprL/tobd
Ycl9Oz1Cf87bBWdFmri3kcZV7zU5EQ4gy6Mkgln4+6fRRI0+r+uWSU41RjQfFX/hnF/iVZofIV2E
9MG+v07ZjtESfzcvM5VFWu3EtmkGFhai6SbQEj1MrfJ+4HCQz78yjZRRwZ/74as2YAUtGIH6200w
VS83t9lL5VuZA4d6eSHfjiVFkPcyji2wm1zvwqdQHuZeFWzU4tm1qIsaHdqu9dzg5xTbjremO5Cd
eGeYuu60a/zP61yxdNz0pzvikbcnzn6Sw6aRMFrXRwOwRPNvfUsmWyZjBb2aSteakAjeWPvXhzEs
rybwQ5sH48naw6SgLjQbud2gq7Dms5BpZwL63CTu676qdRP0NWvWm1uJV+ApT8Fg58XKHlT/M0Pl
y7jzmuCh4eD0rc6GFC98JQNrlMba/HYpkRjl11iwO3AV/lkW4CpfL1UsMhfzwBWH81XLro5irBMn
ArmgLyjdXVOzNOobihCZZHm2vgEaYXFBOCMLzF2gRAlAoemg5e4D9Ed2JhNPjKF93mlhhhNjJhI/
cc04AsOf10lZ1L+BpYbmx39vicwyEsVv5f2XbDPpOafa/RapUnFBE6gd0mIPiV3IWYBrLAezKeo4
LFenKrhnRllhYH8lkUPX24YkFUcWcO18xpXd4XBcgsYvmlMx6CFp5W5nE5janmdGDXs1ZZglZAdM
8nK3+t05FIR5udH++OprrLZd1ruz/kzYAxHZsSGX/MWbs0JtP/onGKYHyqGr/GnQvtqAJALKXw+N
PBNE+GVYXMaJMkarp6Ihbds4s3/owVtII23GvXBG6WK6rVdTD9w7f+9wA0EPuXMktsKbiiR+jpT6
8tHP50emExXzjWuGVvFR4aKNN8iXNGIBZugvrsGXERemRq5+/ig74AdxjWPd5vtyZZTWnU5HKnad
ouOcT/FWMJKAigpiDA/mNfFd4ZVGL/8ZtilB748ATUvu24/S8kXp8KdpPwD0GuYgerPX9Ofh/PnI
JlPSMK/Qk6K2Oo1Jd5uK2ADXCXeX3PMhFMI4vigzGgnBkwIwLZJqYHZtLFNmO5j7XR3PRBql8vz4
k7YAjt/qzPsb1/0lTOSu3QoeRIYQOitROcg2L+zKV1S3YQs49/D1jgxbmY4S1HlwywaepE0HU2ca
swRe5mFLJhAdxE/uDLB+f3BYGcbagnweiZ9GkKaExQvdCUOqEz7e4fzZdHkGuhQfuBeH73frjFqY
G9TSplfTsfvZyPKZ/itUvPdlvPUgJBEjOgYpmSmtLrfeprGcaLbb776fLi5BnwQohIe6ICM6NiBl
QSH0E0hvm15ejKXsirlWogD1dS81nrzSUIQjUUI4Dno0M+YQ1HKV9xfMk+EMPaREtf/wG248+Aqx
ZusFfub9lv7sZG+wI6m1oKIhBJ9/FOXzPrOYABg++M50Kxs9+vMnoj1SpXVWyQbB/tbFNpq0b2PK
z2uXBg6TFX84Bu/rxBdghQrJyuMAvGAElTaNXQSV4otNfYnDEFS+Xtculj7dNYD+ptKAHBo/5+9W
sm0uNgjeEHlkZ1Y+sejcXqYQEDQDlFSxM60TOQ8pDy/7+3tBXHDDMiU9FctoRYAd+fJmX/3qSJk/
PkSac58t0mnhQgXTcQ5fGKHf6AYr0WKnRZWxzUXQVmLSVXyJbdFB6cduVDdPPIk6MPd+K70d9QoP
Y5lmViwhvJa3kjcw/NPgItKWKarIYQuyhX0sHHXeQens7SJbfOGACtvMmzHcAyPCwYkEvExuzmHS
yiLVw8gxYpX9Gim9islmuu273bQK7aozE5b2Kx17s/7VZ7TSNcAJgIrKT/Awq7X560/cvgz4jRkg
XorN5UqKoO7fHKJPezFjRJg+tcPuVfWOifKsFHPy8roG8v5bL8lsXYnYQ8M6wAMzeN6f8FDDVKls
/zyiWlgYVS9ko3IyACB4NIZfn3Eoffc876u6fbDWYAJTfNJQjAno5lid5mhvnoc2VeYJ+TR7DgAx
+dHgpk10vAvsjM1WTdda3lLTv6mbYnHYKVgIqCqljj148TixbT9/wYJ6/7QgnvQHfqlUJ3UVcHnx
gHbwDZS8JZPYRbmNkX5Mx0XGNesN5PhAxmeQzcruqyCb/knRoi1i/5GSZdcVRJ19qX1J4ru+FpN3
xMk4kBnnXddzJwsKddNMD8sx47KpGp6aABUhqAr3nzfDpLTOWiBXN/bKooDDNz3gWwDzlNsh2um3
cBHoDy41i2BMNQH4JQ+eMVOvRWJFGgsy4me6q5ofdtNukNbHUP3kxRERKFsQk0AMyiWnPTANARDV
WMyqo8MGl95BVIfdeTQiuB8QAKmWLVLx+hN0ccj8fTiT0LimKwnA1mRPrtV0i/TcRVNr1EB3+SQV
ek6lrBPF17DHCWiLDjco59jaQzb2J+Vyt+i9nGc0HCmUrdzGb+kBwvksEInnJqHJvgDK2l9Qt7h0
CKkLHLQai7aOxEY+DSYKlthBe+F6/VPL3UO6AQLqWxstp92K8SkiKdbvzbafDrIvRgbbQE+CK/ga
OQ8bsBz2jQRZi5h5Ek/b5kN36HgKYKI7bMN7e0QBIMzdnH+f6M7M5vM9LxfL7WpmxoSg65fABua7
tKli7Q1PqT438QwF+u3qUJujiOxXb/h98gc2VrLoqJyzz+7oGG1w7KhgOUEgL+mejCDoGFzv0Ym1
4WWKgFcxrlINMuAxyprpI4zzDUEaEAdlAdonGUCm3aF8JGgIGIa+MEw3ELh1EDlqZRJzyg8FIx0B
XqdZokcUy3D2Ha3cSqqImM/PPtLEMFtDQ2QyBGr+6SmpSa2lhVY4WOozfD0NVYpRZoYo43hlsGc7
tHuLf8lQDp0NNKWNkD0isrX0ZltnhvedmZBqVh/pCMdkfnPJIpWG3JySy1TUiNj7i6oKv/idY6DD
a3C8098VJCffvd2b69z0GjBvLwRLSfqmrhrIEfMoMyTmNw6smrjxhxgP8c09DXBx0dab+cbV8cAM
UN6EmyUiKPBi4Vi8qsAAJ63kO10JNIRxFf44opjtwF/qQbb8XodbQFxlOXzjEwEtaf31iWVjxuLw
O8maKG6kADV5gO2hy6wUdruEgZ1j4uiLwoeN2dgrusCyFwg6q9gnnnWetydK5YyGxxLPauY5nEDH
hehPiIO1TSCu0P/6MIiyCRjgXaVOF8d3Pyi20Rn+GfXwVBYhzDrtywvXuu8e70a+vyZ0kYHAZ2E+
FmXlwLjssp3m1cm5UArw08BltKEG+vZEgx8gUzADCrUyQfn3qSQ9NwJWf3O6IyId7iQAKTOoNvlz
iRQNmSlmLpKGIlVtqHI8E37W+7rAnedrdys9N6Qv22/sriSgGw2NQEexnKqtb44etUT2CbvFQHpz
FgE18t5Tke5duiLtI6f/hC7gW1oDIzMuWRgIm2BkO+oIyVWloaWq5Uo9orVk/y9ZctHEogq4Ahj/
iNg0q49PLyty5JMT5shEVceBXhcfhjEJSXfxMy+1bRTMP2UM3+CnV3LEczEXQ0nYVH/HRiUMsmOU
W8c5r1fYwyIXMOidiS23nuD9sP0yIPpCk2FX+RutdPPjzY1oJ+r6j9m8MFMIA6BQw2AjSB/pPbUD
TqCfPeg64RcajVVOBqb/RdulVocUzVAJC098751lLmbMKpj4tdxY52c/pvm1Q1v/mz+HBJCTWaQ3
clL6EjHRYrWtc4S91hnEeGsrOexT228DuX9vD732cCUlVnCSfhH+jamOOjcdGP6h2dksS35T1bAj
dvddbKP1ekgdiGdQHcjvQIqHDpm/FagkKIcvMMgQ/+p0P38UTAn1kRZSXItOYDbX3dr+2L4Y12Yf
166ygvCC+BjYUBtTyS0JEHqECzdiyGmhAbnKGuL9UKTmJFsh/9mUi9SDy3QBOxVQIPMTmR770TUR
vGOFrC8Mw5+hGp8aKDPmIJV80uK68n4lz77SqXTVkvLUf/SXGsGUo1bRV2iDf8XGkF/FYmjYSF6z
/T8dLkMJzr8znGi3taqoYqOiRkOeoSGsOzHkqKXt8AqsuxrG7VCub6cm0hV/xjXsXBNPCSGKm55k
lJPrKFJNXovyLSwrXLQCpeWpGBzRPV+8ysPdpbtRoiSx54enJE82VxKJ22fZJ+dOnmRx5bfmzk/X
QeTZzvHBoIv87Upl6jA+3ofMn3uiJ3hLpNL5S/PVrWucNSzpm/BcqPW3V42DpeXb7InlWQKX5IDw
0GZTNIkUCFQewDuRGM7ykZyKiBKC8LjaW4SwCxyUjbwJq9dUyQmLfe49axqeZZ2wYB0YHrq4DZEN
8wPi6RxSVmTtknsZTwA+de2Cm6EGySLFinfwCsbLp1xub9KGWxoBFBl5VhJg+mMZqtDOuT36nc3i
P17mKDX/u+EXVL2APa9sra6mVABX9kXYlj2Dwf6Wwy3raAJprvq73AmzHpMbwubEo551hwC2WdTI
GoR2PpXGvOT73MqK8ZQ1ayotCncBeq0P8ZSjuXX0TteFal6iueBes4Iz0b6iuBL3SA5RRJzDwpzz
6g+kpCkBVrAzfXx8CL68xicgstLky8yaL/4b2whbBqp+Agq7fP5JaYZgJ2Uu82wJ0nw2uS0TOuQf
Q7zVI3AOrwDySvweMl23t9c8xnXlvVtR2RYhNPs51UfqUNZe8RAYDwFQwnWqIP21Ytjr9ocIqud8
YXyKsBibP5N/5yr0whGGvglX0zQ42camwdReqY+SS/an1bFTQ9CkTdNDtEATZq8YSaUMvZkH0DVh
Wsmew02mPrrRZRWi/zwlQgUVRwyMu/A3Ya7SoYhV+gVgPBTNSOr6pwP2sKLIycXt+MT5w1sKk7ph
pBbSW2kyDUOCvObeo3iAGR4wmOxnhK80dpzt9yIEYZKpRwg6FKWi9CnYu0MrcJzJay9rN4UE0vMu
yVPDIu2ZwZjyJrl2AuR87ogqyf/qLDJlegAMzhe4KZtJ5rX5F/XyxByQ56OKbtJvAOUUxJD6UpfI
Oo1Be6xaxQZFfQ5VMHFmCRUl4pSqMRdrM6l4h6wxsodN5i69Y3idHYeen0v1wh8dYy6DhetEZdA/
q6Ib09f8LgNJQjRX0sSNZMPir+840XdiDTfebkFkseQlu3CpXJZYPz02JOJzhM1sVFfw+eYRg4u0
0VUCnpXJuOl2tAueSeQp0krHANJ0apdT2Nj3bicYKKm3FtiEurYD+eK4Upc/sOheWg1kWIeaGn58
uZzAWA8ThnY4UIUGkxSF7rmRYzsfMOCqnexKuk0Wjz7YHKxY3G9l9ykkvHHIezibfexgBO/oAT/G
HgmwSpd0MjmikS0p9vJgy+doqj+sZ22lyxD+rpRklI8Gbap8O5WTAcJQluJcpHgEKLiENYyvZNlA
DuV7HUaYT99MwfjSj9nEtMo2NriAjywg5aQ9c6ltYHASasU2gnQ0FxDxHQdRuCuDhr5k3sumqQ1z
fZRtK79m0XpQnyMfC3M1xnl2ch1BPliD3SDX6/XEZLWSr6ME9xSsTEN9LbA/xF1vcZxrRlSgkGsQ
6wfb9UKxLstvZwlONj/JLMMMy4+cEb0/xy0MiY290wsrsldLj6Gk4zYysWV6Eg1CKYmyEhAQ/Wql
c99ySVogWYTONQ5C/BypkPd8SbWIwh493GiWvsHRdCWaQSu+kPwu/pHATfcXIKKh9iEcEE8kKu6h
FrP4MZ2h8YJ8lRhBD7mNur4CLz8u1ut0bitGrbfzS2g+Z6MPOGw91oxEHiDVGpFGLWg+1xHjvvAA
HS5QrYJcz1rt+hj5H0EQJ4b2gErJoFLMydiBJk1p+eqVsjhCnCNgrybp1C+dgD7csYQKncag/dSD
1h5PuWsmBFFq3jBsb/mO+/fzqAeM5graEGD43UqvjEz1MPdY1O4zgCNxxPPqdkeTTnRcye7S4IJH
Ozuc7dO433H0dW7eDusswPFHJm+mC9tL//K0Qo/ZBPdGJN67lLW9qfr9Z4y9u12e2aneAkDMYQit
mUKB/HJfQwsx/ntj2ty85R2GayPmuMeZqYbHG9Op3tj7+AW0xn/vT97I+1SEg8NCx8M7xsRBtwOJ
FlysQr3gIiSVd54UsREuUrQScYrTPMJRd5VPOdNbU8dJRAfUr2+6ihpUo4gP/wSWYNWfuvHiZbYA
maqdVeWr7ucujo2p/uITEJ+4Bij3Ggs+u439M2bvqNa+8y0+HgB/wwcT2MkOJVb2AhoAKRCHufQH
uwbdVRd76yLWAVL5qDz83OOGN9lhDrqE/Lmc9CpiE5XrReTzGcMWPouiog4QejxitQVyaL04Ge2D
e1KpZ8KpKWWnOtc1+UqOSgJle1GkqB1/j2iQ891ivQjv3YVhdVff2jj3t9MIrG6JAmjgWtZ5+T01
R4JmmyQnjIS2+wP7TOLtkwSoVlVXWDtlXf9IZqybteMk8I+rzC7w5g5L6kZ6hMdOW31yqTP57TFF
rnjMqrY11rDB0rU97IhIW+Us6kkfyZh2LKxq2Fi6ASDn4wRc92BLnBfuEvMYAS0yPUhQeOchUuoa
1Hu9LrLiiH/7odjrFoVoD0fRqFbkGo8GI2s1F9x1LK8NOcjkaJ/RFvp4V7bb4jRYilUGzJ4zEdkr
UVjTm1QH7VZdtuDw/gy87Ch9NK4UlSKd+ysGSrUOwcP75u+yWL/NoK2j8adyOfutLBcXfmuGPyDj
uOxHZ4zPJ/5QlxeVEtv9pUUgsMjxPdYv6+HRJczJ0hojC1Fp0lMzRYIjv5EFMrDFTzTD1Bf6XfIZ
dFxP31oBRR/oNix/3o5NFhqe0b3MzWL+lmUot9Rnha6X0upnx/MB9bu1PVi21Eo9n43YRSxv1Dc5
Rp5lYcryGZR6m3Il/44XGOwAmJsT4grmZB2vu3kYpSPHQzh9uUC8ftN3peOSWowpsJjUCouLuHBt
ZOE4CZfeHWl+0tGnriBK2hbNEwSARkfVnQbGrpai2/1TAqaCvU6g/SMzvvHtNW3TKhP2wmIUDXL4
WTAOhFlP6rp9l1+wCer/gY4Yzz/k/s42TzkanNyxtqP/7WpKU9OUoJZXMw+phvCnFVfzKpirZlv2
jc1Z1tYjMZwzzbmQPEjEYHTt0m3FEpli25IXHdvILMdGDDXB9E6uWD5DyPqjV4Tuf6kwkSeC7rXR
IjD6WircXvJnZ8XNX9iFpRNdCYOpKSSOqFKqzFGB8LOHpY/b4OjTBGKY8gSPif7Xxko4rM+ZWsUe
YoKrzMqiTp4rw/0rYolSubWSty4ik1SMi1P3FsFdUnhGLTZbhkabPrC1HmTIcxXc0apHg5H2jWTg
tZGQwArOy1j91QS7PJDWH3RskSnUuiJxjZ36In6ZEKVp0rdWHzlmJPbFHhqjwTtKdPszoqJDmYDY
LJvEuY9fPoebIATyxhqaEzveExWDS3aU+ctqyBcBtndHvR1jBTqajoeUvLpipqWX7csK1s8X5OPS
Yl+nYkZNCnNE2W5u9gKTWyAvjMQ8xTTZd8/gLoTIV0id+pPAf4aOup0v/6F9TxweTGaVYRRpjQte
KZ4LyfOFj9MPLSmIH7qjL+8KEnW78SM+U8V4OQ3uuKl1SLJLe+3UuFW4ZLJ5U4afKkh3ocP1wLk1
eBTn0pOTf0yOlHd5R+f4KxJOz9Ax/6R2rRfShgvc/AcU3L/L8zxfUJ8pUl2YVUkd4uZaoZGpBFuN
GujdBMuMY8C67DP1ZdL4X8T+/IJcq3D1L16kat7XhIfFsRM1gtl/snRg61UFPYfJSRqTGu9u58UA
k7mxzFgpckW3NOHx2vzIZcxw4+prhjKuTqRA/eLe5gHsoPoWO+70QYq94tFtp8mFCo/Ueh8zpCsg
LvTQloaQYXlom7y7prXg5oZeJbHZTx133RyjncNx4f5Dvpfhn1yrLnoQiHVPhBF5H/SJvJTfxL6n
tW+TN4dl8hB71EFP49OUCP0TwP3thnhqa9yFlNAq4jZfVR6z3gm+XM/m0YEGSbc5QLCyrmxR/jhC
CdlCQuVoLlhQqaE57ruc2i855A2NC3C/iC6OKN9t7OM/De3H3/qaJ7x4gVQUhcLLIC1yJLN79P8C
EAUGOBXYBZp4/9VE75UrPnAxX7+Bs20vRKcZ+fP7MZzh0Ku2uAil9QfWshxCLopQBrDUMnFhEUw3
AA9y20IGJZS3c7dAksD32sAxBTTdMYkHfZj4vmGYUE69LDrPrLMK7w289MsAYqSiATMbOeQVXwa8
XZdKX65VTYUXYdZmGrPHZM2kKSQCWCiUsCy1hK9nHVFML3G1iYrImagbYw+q6Ur5tjFCPJgGdLP6
C4ZGNFmYdLDKyNNaT4Tw5eDrkD1JC5JZHT5tW7Cc22OqnC0hLoBgVblsIDxAbe8WqUXzE8nPO+nK
ioqmJo2DBV6D7/hNyEoibdIG7uPm7RmRBkxOhHrpjxLYoR8BPbcQPzUtWRiZFUaCtq1FdrdQfhZd
es9rRiuPwrVqD4mApBj8i59pqWO9cy+4e01pLM+9F5EovZ6daMi10LcyNMzZVcxm/4bWMVHY9Xx1
Ep09BraUo0Eowy5dWYvhrgpeD8x8/i8+l7otHUqSRmEXuwxbHflKtYJli3phfYYRIl0BoYNLIXg3
D301urrtllwoPtFW38W1ArqcRv0YqzzKdurUCOiJj24O6s48dhRHtpequnw65/2EmQzQ1RdpO0wX
oInPyOFh5nEF7ZNK7pHyl2IKXnxj9O9NCjUD00PskTZFWm7UWbFnM0KSdjGEBWtz9m6Tm+S40WAt
vLXVkMQR9Q0ocM4nbvI0TFsmt1pTgomOenN7dj7Wvlulpgq9IlEn5JB9KFnxCJXCJ1E0OEuKf1nc
oh3khk2Vr5zL3p54Kl35m7bK4da74wi3XsgsG/uoK1K4/X3nyYuHnosgBxPElyILPc1qNWB/TiVa
EVtkLIYhcGjrnJ+mU2OrBU8KeNCJXYoF0YvfajZW1/dxiETi97KGTVGfrzBLOrjIx+l5rK/ssfnC
DgasCIusmXjvD1wpyzTAeOIph0o1hMvhEJSlz+A9YOYAgMDhhO0FVgw1Dhr29NG9JKssE1Gd5Zjg
WwCn044riXLbESU4q0H1Th2OXeP9OYkLTMFed0MRX4djLkkHsWmWcAmXN15ch7d5w2kC2wm2aRU4
/Y4iRt2WpxavQhaYTkeyLKdY15VwTQ0xs+GFpmHJYPRwmItcBLB4qeFrj6sQzxx3rx8B3lRc/JwD
hvy3+t3oUhN1nDtoMs/bYnXoQ+WmiZCDt943G0m+tWWceRqdG/45Ge5V0RtHMDsjeAKm2SUgyQ5+
8nEAjjhdR4ANC8g5IW68yXjdl67wucwnJzlAX8SUQdnv9RYbPw5PgbDI9eUGKug0m9uGqu2uS+XZ
Lc2M5y1/VDgKPPxGYHayInJD29+kd7eA4g9znQw6H8vqK7s767r8LiKy8jhAYG2B0zRD4JKEhKLb
a7SDIVPu/1WJPIXvKd1eSImnpejLLMdSeSYh2nbTJtGD90B5R4HYFIhViJZuEXwtlP+/ta+fN/XS
6AIbTQW9V6JIRVkw/T62FvBuPCvGvlMWaZZmr3xwBawWHd6/Bx5ot03l+I0e0AMAIzXc7fvxdhhy
ad9balReoXvNY8aajw71otx8YuieLAcXNOcEB9l+ouZWaLDh2utp95RI7pEZQ34GpQKpuUEmxpZ6
Bzg5NBAWXBjxeMjBl2XomPQV13rsOoOHSEieteMcs8npllipIE2CY+e3sLsZaqf2qgUi25tXhjZN
u7cIBhhCr8+bJ09pBsV4vB2xjjBT3Z/T16r3mKRRERge8ruq4IhoMdoBNjrkK6LV4idjVs1WBtwp
U9KpYNr5j3GojxDfrCfHKQ8tM+xB820QB4oT/UiOUS5Mmek4flO3OeQCRpe3c2DVO/GmHeNmjd6t
eEO5+EJZZC7tzb67tbGrEIupn4wNOGCBDlylRHbmxDWpUsRnaseLBJgl/QoGU1FSwLDx0PzgsHpI
E3Vi2k51hRzfrblgUVEL93kP41XF2enG3eGEdxUpiWPgOhh/FuB4tnAcOtym1UvjqeZkQGLMi07s
JSjGmhtl6/iEBP7xhP6CSmSjSMT5HGff3DaDvXhK2WkGpzQO9ehWYdC6Jub1eM9JeJ5goVZMsayq
y28fdLM65ChuA+He38awEDyrPOv9t87ursC+e187ARKqTyAzR6mTlv/J6vvK9f3D7JxNCGqZBgNK
09+O1NPK6HLrtPe+WiSeKtozErKZF/BqEg+fogngIyoBrWEEOfhnUgBvXM8EDCdvo7C0Xx5z1Q4h
lLg3hFemoyk+dpEGAd6DWUtayoAENL6DiTlBxu3hk89QJaliKe+7y3ktd/S/BHA4sNqJoQSuWZk3
s4xRnG/+alqroBFDCeEQ4ZbLlr1U6nmDiZmVKscD54SgxybWF0JJzoDvf2Xb1k/br+gH5gDH3ywq
AyeCe/6eYuM9WRAA0IoCVmVvOwjPbajo9m1mUKhh+g6aW7+M/f/xzwEcW/EuhO200TvOAwb4Y9l5
SzvDz/HDTglyyWQZ0YwwaeTWhSMPRYxePS3tDCzUeTg+PIg73VqDn3+y3smTRLWd87+HHJetf3yJ
lC9m8QFVJ2X73/PT/ltXZdhQRUbaMaepMWlc6hl2DI2HCkPTVKOJrE6xjkf09LcCtZ90dK43uFze
jA7JRtwsYNj9YkoJkQbMBMm92/Oc6iTYOAABcRShl/qTd8lxJ4pckDqYcM1OYQtMarDp5eOtzs+H
3ipEsbb60ghR6qG9wVZXHFzfmBq5TDmQJxc+EP1csmfNQCr36jMY5iKPEmXvJViCxSUjeK2MpW99
hPzAQgfDEC1cXcUVbescNYdVm/PAL8gmKI+wU9WSzbWo9j2y5tPyIFYeLWTGrq/3zUJwVxFdizwW
D/MLejENhFD1FEs/Z3Pj5eH75kcIPq+8ZgSeP915m2OyEzNhN3eT+KcqtM/SikIf8gxUCN+7p34M
Dr6K9HeM/gsVkGxS17noWCtaNkuD8aY2uHyxafKfeHW0AT3GtVWA0IpyAKxr62bgm5lLLItZpqLA
tcYEYdYJiD1u2rB8OFGD/V2uTDjEi9YTNsKuqNfSo3AlHxhWJmfrnuS4F02+9/yRfNnOylHkzBUH
zQobAB8YTViYcXdAWt7uw39apCUkKJN89bNgaMZwHxIgGGKAiW4vMnvk2E7LjgkAyNjuFqUDCQ6P
z/Z+ORqwq784Lx3vAOG2yzwjJJHIO4k260Q93PiqKQ6G8CyRHudGgVClcrPolrday82sfA6SHiAw
M4c37zzCFGXDqM5WfV88CSEsEILQQBLGnDCYSpldVwJEIxzNU2OxegYmQN1V5OJhSOekdOXpKjUr
ixpJ6KRVdnqbDEjA/Q2qSJIRrD3pGEThioRnPqcQ+Eoswb+h2/LE36xG0gAEakCNsDKwojMXNWXD
OE6mqgLLPw60q6YMKkZPGWefstQ2n+3fVxoINafj2DxPQkQ1Iz2EhKIF2ePg3ZvDeaacYGc54SU8
ACQGRzYw+9ZLFYo//hCUm8sgRYZJlPX4dhqT70Zhm9UE7Iqtm0AbMjsZhFlgeQjwmV/ZDd5qvCtT
VTCGgsRLKHSMb171471hm/4TLmWH7kAcxcf+bhoP1xjWslzlyyzXIYuVcWnG6OULnG6aeOfQVJ2S
REF1PIjsax/sVYMelqDPxANfyyL6YUAhHVjq4mGt9mwzzqwXgWnJXHq2fQSy6kSBNYq10imDbPwW
hHsIxE1FJF7looWl8q45nNBZ2D70FPur5ja7vHwby4DLBPKmUV7LdZmzEYV2KxKJ0sAyqlZ8hxIT
lZ3cD4LfOn5qtljbUbCupi8kw5SBzyPXDj73aQXqLyrgj34S+FB2KgRUR3b3Zci9AK2RS1ke3dE6
JY8va/ZQJ8YDrMvxJPBYJvjniPPNif++M6HLoWtuZaNoVej5eofIbB9p/Hh6WkFjNq5/P2eOemJH
Y4px4mAQlmkkC7cnmgqnq5HoHOmkp2b5IOnbpMFUBWeifm2lM8U9Va2IhP06QmX+ik5myTBx2Vv6
YpBUfTsnenzEihUPpplMdthH+kj1okzt8PubRTlsEtjEMwSX63rtZv4Echnx87GEEMg4c94GZ1BH
wSJ2unhs444jn+ZxuF5xPvvApoG4vgjgfL09w4V5AaDZrHwz9mqmRP+GWofD+VqrmCj+vLZvsN1W
NSbYjEPc/pnEa72cufwjNnDuk0oLQh5eYmbeChHKem4Y5P1CCVrXNSfFcIjpdyP2AvVB6ND4Cr+W
Dsvu+7kyq7P+MNlkjBK0abK/6uSP1L2Po8dQ4iitkYxBsevEiRlcmI4d7Xtl9g4eogkNmu1EYGh7
j8++igcxSmsrJYbjNjGs986mn5GOorQzfYVuq0Xu7gOAamsSx9nCWREEAKzGMnUb6rCHvqTFkPXc
SX0vuZBBHZOi+w8/zgLL6V30EC3a+ZIGOg6j1rCuBoeksFlQ3Opyh7hO+7MqFtYynMo1HCwF9cpB
eBP69RuE2PcqeztbpjtBHE0YLQrG9d+cwfm53MDHFoFsLk3BTBTYNlzyjF8PKB3qJ0Q0JqiNulUv
GwJ+uKmTHUjOjjfMs7OG2xNtkA2MKBvEri+0VJi8/7vy9p+B9KQdm6xYjSMdJuvuMOIw/UPvEe9E
qJeUiWnlVx69P4e1iW2cnBDlp2tulV82fuuaRvTWoXFvi2J2o23jhnVbpWZQ/jk0t7VZ7bMugPNf
4coREUHNA6IFlpmE83zZwA89ZTDLplDtajqGF7RqFtFN4icvbCe+So46+UuSrthDGRD4OaoAGRhX
Pd9fS1FgLa1Ymrr1Rb4jrSK5XrDOWz7TRWnm7bFlOdRkJPd/hNKcxE4vtsoj2G78K4BlNuGorA0M
5pqnZbCzUKAzDlnZ2GVJEJmoFKZb0yY2maMtoqwcqKhYSTrVMyQ6M2Tg5mgV9EQ9gKqB2lSQ2LgL
OEQa59ITY2NeQka8idJrgA8NvJDN8Qt2RUHw1lfemUqQ01RSU6O1r5MeotF2GAtTr390tQzYj4wu
PIiAeeP4S6Av2hNdS3kO1SAxp8aQvYktbCCn3/PYEjswNv27D5nRFJEfZi83ulaCXulRXZj5utpF
iyBjqgSSyrFcQ4QbB+bve8X9N9KkUZV7iLTVIxPDhtpvw2Frkbqcfy8Zw1/6Im/k54b/sYRsQF3W
kUKKMR9yyV3djkzjbuEFYMd4iSA8zzjD3CSvedDqa3aVNyfBZ3bQMVtAUdGXMPKS3HIrTSzLqfTI
GYrzu8EG7iTuADpOdvmogd0AcJvK58Z/jTUnPwXLNE1wd6VsvnkKoEtzE30dRLnMxiD0JbMO9sVa
L0jMF+59aWoOroBj67bWfgIrU9JwQY5y/dpXdGTs3W8b+mbcrFLR/zkfO/+DOSEaECMf6BM6FkM+
dk+mJBvCZF5pHZf/EubmGvoXhQiAzBVaWGzWGG8HIbIM9tlG5jlmU2dizvt5csQ8SM4AAe62PTrp
7wfNOIY5c2b/1jU8KSBdI7vTscu2LSt++l0mJve6mZ0CAFXnqthNysssIjSPIrDb8tNPn8DLxQtw
+B4DyuObEv8rl++Wxo5vUq9frsvW9IgbwGuOCnLcOucG4X3f0erPPJTWRVND4kftusMXYsKkch5x
fmDBUTCwM9BjSfRnFFyNN54H6G24A+/YtWtAiavS+Tj+DXs38dcyPcDRjcQPAvUEacFjACiAymgk
/aK6Pgm3H67dTPXMoQvM4pQfG8mdaOTGyvJF6/89obwzZaRkcKQwy6sEdug41G51NIYm4aS2b4lH
jEqYQx8Di2EkuEnDLUp54J+2MjTJwZWqy0KIFZ4Cqnn/drWjijObYSF3g3/iBSO9hWv3VgCBgiUx
pi5nS8zpcJ8x9Wsah9uENeay7V5S4a+A4uJ+0+AcLRGE0f8RDETbpUzXluE8LFYzMlRxWPk45oZ5
MooPadrDjePaIWf/jrkmPgi4qVYlVAavM8dTQ81AKIlVaecy7mKr+NZw2bd8sUx9P4BXLjFqkym2
vWhxsIJoEwr6Ba9/M0WNFxeOt0uTSVy6fjVp84AQ3btrmWlQvxeXTKlMB+4J0E94pBcE5eP2mxZl
RoDXDBLl+XBQI2hgaWIQe3qRuFVzCGpwhPPFSrGKtpp1ZGUgCIjhgtmcZ+H6MhsOa4Qdka7cxOHh
4Tnn0Iusb9Re6ZQw2IqVN8YJZxUD46cYlyInQk1p4kLdej/vbwD4sSkL1+xR/YkB+c6GcPy2NUio
D24XTpr9j0+uQ4SZ0HeIOx9sY/o5JljmmO54ywB3DSs4KckEcwqE0+kFK+r92LQzDwq3WkKhL61D
c1l549sq/DlR46T/P8JcSdhD+OB0tfIyHk8P/SCzbzzSvsJhX4+ganckGi9oZ9N4QZOTrF0g7bTk
cmqThLWUbxTR8nNC0M2KS8MG165pL/RnP9BcsG9r5xsfFU5E2laMdedTeeCdyh7yEvSMYJqOwH/H
b8JH2goUMqXylYpHMiVsFcQbltvXTnbUJ2O94Ib0TQr/DRcl2N9GwPb9+lWgweGiu2tAP6Uw8Oau
HsEHktfOYhPKb5lj4jCJnfBJmUyBIJ4vFfZeBbIe9Um+eJdmPQP9X7k9BY2APdmLHrXyOJqD9qmV
+RuFhc6KWF9rSvLcwbksfg8MuaPaGlsrWSHWL2mgnFuJwkM4T8rpQBJTX4vtHtFEaVkycpi5MCib
h++uN7fH9WOhELJtcg0P3qJNX8+SdpLdydYl8VfJCzFgOk1lq7/T1SrM4BF3Rsc5Ai1cu8jVFxyn
ELCTPviP5K9qphxkB6eyy9/C4kRVN8/jsYyz8N9wxfJmIduEUeefK2F1ZPiC2ch7K3EahEX8hGVP
z7MFbACaOwtYvTMAFB8ENszygzz7R3I//5B7KhqdqF8a32/+k2uuDkthAc2erd7tHOTFeIx8/W0m
9esqwNC25n3kexhS/SOhoxibPERY0FyoE6cjvc19373NEHviWLWnOfShqKnfA3CDK+k85c2ZCwUA
0g2o70l+s2sJfpW8u7faZxQS6EmQz7dIaEvXl+/aY8mr0ZYpH15XAtnwXCTWW/bxbQIy/EIsOV1p
ug4vcERUBsTLuwm6aEvP/gi8C7ddbU9K39e6cAu7NlmbXEC90A2QxsjJrRAt+vwaizgDv3Qnu7OU
lHFZPDUjrE15em27SRjgJVMSmSOVwMXzdNc9OusuEZcZGEALQXFAgHVXvcLFJ78Nn8oHAKuiy44H
9h82VJnyTf+mNs9/C7Di0bO3VHKtB6yGAPNM/LLTGMvbhr2tO6AwTT1Jdoyff7wFL3cL5A4Bq4Kb
svABaz32PCoDJY5k5RRGjmcnbeOWXNXlCz16YIScyQdnrzvLTCtevFvgMHHVjvPFGB283m9+eSMN
oD3r9liltqn+Tu3egZ6ZLN7O9S06xtXMwdlCf3X96in93YCgkRvvRtmss3bSyfzC/1+UVoB569F/
0vfZc9W3g/AJRdRIJYkKbOcWZ/FPNo6GuXonp0Rjw5vV4ZekigzleLb9GOkKwKK8MnHh8V4g3Z7Z
6XQQkUdTAbYK/MOsoyp4gi288vJRB1uZ6GR9t3E420JPd62FEpIKp8Hv0N4MnXzXjnKfbFR3K4Xb
4niNKTY+nyt83wveKoBw47QhSN+fg9R9KH2QkJFHk1Al5hEFUpEj3V4+AejSBCJ6h23Od7f+vH2/
CDe/cgJ2KlCoLGxAhvtgIpV5S5JOhth0bvwB8YB57B6BZmOR56KanXxpPTyXygCkEAiOCxIGOE8y
hiWb+6CNkgbFs2h8P5fIJRjQWiJ7s62PFjzpOSxYbOqVItqDzRZs0t5hAYrJz9mMz2ITzh+G4BSt
MaXHZm3SScMgHP04qMv+1roR9KD4VCXEfXP3Ug98SblAodW/vWPoWkdWXKmy1YeSnjY74NIxSmrZ
MGPKouQt5o9okmWtnxoneK7mNroRc98MydCBFZTm1YanTCqoklRJ/gJd0Yc37aKTTcyBLtN7T8Ew
EU7BO4y1+wgN6v0qAMhwO49bcjshmKTQCrB9r6h7+foQ0pVgQwobHWE9lbneMjrw6LAv6n8F+j86
Ywin91OyzIQYmpeWu/F3qXAtq3WHcfON+8flPhK0JRD19a8b06WuIFXHDNcHtnC9HdlfmQ/vnFF3
HyLWtzB1e4htacqThDEGrRrdWCh6+UZ/q8Y+rX7PS9e2yBQ86HMMJ26fT88dhRGWuMb8Mo5RYD7c
Icj0dNbmxVEIY04DWJk6d/ZNqfPbjvHKhea3dTnkS05XGV7mcqFSx/kxg6RWbqATBcs46m/dVVql
zMpKZXVTpgsz2tZBLZ58s1xmybPvkUMxOg3VzuDr7jH4y34j74lJGkBiFzHFbMlxtyg6TcdCXAN3
CaVVI9JbPOjsII9kABFgC4pZFrBUKfWt6IrG3h4UZ0uZORTvC+LDJExfhMGHImtdulyNxuVZpwL6
oQlT1J/VaZPk63kj4YTh5mrGh9TGTk56dGxvhFEOW6PoeqwPh7qKp7LMM4J3ZZMScWKfg0eqsvEf
+4l3+H4icawdpE9N72sRp2qILfZCXF5fIORIdkSgQ96YtGVpkUjDDtHQAd0W4U2kIQZEnQSpH39P
brgsOE65RtrTxeFKLk/1pxXRpV96q1DrMPUCr/Egb9s/12BpWEMOrndUki6Xj0Pndm+gd3/X8/p0
PtVoZQt+E167AkDIEn3lzXWGue/JZjI3lHbawqHE43lmjxGdRgcND8qRoT/2UPgoXKqMViZQj7Sk
UmGTP153OcsyStVdC6nf5BdKQVZ6kQ2KH1KRLjPnnWRDUVQmMSQ/B443n/Tl89XIGDSFVyfcBgrC
aXZ8537LNyAUTnRC4yyjaNWp82JhRUoQF0z+a6w7j/8OTAIeZycWvW6oIXnEUUE38ErXHfdoIeVg
X8cDFblXwgdFXrx+1bw4JLQ0yD9R4aLvRdH8M5SGW1brakmVaj1BeP8/KgPaBwEEG11ZfH10cgK+
lfZspSHSiWbJDx4My7ZVOm4AOdTO1dF7Vuo5w097uEvCT2k76Vv8Frn4xIKjJLibnwhXPEio+1K8
M9I1pK36FutKO8eikke3o9jA5Ttv3VWPNkR6UX/ZXsFlfoXvqa+ZKMeo5J7els3bdTxJ8Ao4RB12
KhWKb9Kcs28SoaihKwJ3rjr4/fd8LJKEB2H9rb199SxazKQCWmCRh7TIqTIuv7B10ZY+V1fPcN24
yVjFqykL32HxIppbGYMLbZRFgqUTH2axbusV4gSw0cgLTgI+K+OL0f6n9tbtc1E4uKwiCO7fw8Zv
uFV3A5DwquIaofyxoXZ9Qb1idnT8u5esP5ot1Oqpka6i4bRpFG4orIXGZBlPQif4fLsdW6bAV0/a
HBz11ImWXoWpFhjH+8wStZzGS1mzujVotKISbnMnNR+p3R7hFLlExZ9ZIlCrYVkPUM5hSqyuiLEa
xfXpjsu+p256zo2oIehn5mhYex6jk/9/6QPb5zFX0sy/vrfoIKIj0ZSVj3DLaOx8kdX59QfrXg9p
FBk7BFt6eg7vx0BzcLxkbuOl2kBb24mGbs0w3/jMC0/VOl8m7i5TlbX546CW+wFsWzeA4tYN69D8
daJWLO0qgBYeTFLPq4Ipiob9U0XT73+h3VLG/sqKQW8rF2KjtnnB2e2mNxCdvc22YJKpZnNiYnTm
MdsyK6uNiSqoQomaYm1KBY+GzKkLZguDZXsaXVg5Nri71TPLa03jdO1Fi1xbxZBNAV68F+xRZahu
ePsKP4gx6ObISR1y+KwcXhHW5GcqX1HjPseKwvm89XcKdJ8Yr0+RhuRikeqaEYmZmGiW04Sy7gjq
QJAc49paSpxbmAcRBLVAwvdUW+Yz8t94giHY5hwguLwLEIOoMj7/0+nyNkhoUJZTArW8FCwXupSk
m05empuYetqyU7Zui/qcZG0nptJ7mvvLtLg8yxs5MeqJ6ufw7PG1MFaiyM5/A6urvkPIU8joylxN
x3gX6wYu5jCVvF5ZaMIfsayfN2JSa2H6z+9tapxsPdwHCQVFimNqAtcTaqsCCbMSTnhMRD8EpFsp
RRZjm0hDzrb1Pb0p4JrAmYIR73sEqq9CKWLeXov77dONzlRx+1biFmoHQ4vBSITuD5tVcHwiIzH1
+kuVpKxbBZrvJTiYrh71DLnedbH02hz8hHGQSV6b/jzLuGrbM8VOSe6bnFjU8cznYB24bOxUzDHf
fvy4Agg6Sx4ZgsWKxk/uw/aSBJeour3dZHtAJhfFrIPLqrwGK4Bo1p+YEMteCqICKPTExJhqHN5G
H5oKi1+1X3FjBk8AlrBBV8f/1v151VytDvu8Zbh5nWxx9sp5EMf0ApJc+DuZWOnxJLe7LHApg02t
J4J9U71uuZ1KudTCbDn99qCsG0tib7Rlvutb0UJdRHMR2rW0wEx9IZ9+XvJYnb6SFskn5208YgwZ
NRUNkOGof7E6X6kzGDt4+mSSqONXDkAQtBZFDS3SSHS+YOZwpbunQHs87p6rvJ6AVJFsa5irOs1I
AfkuS0jD1z10R5ajT0gxMabdw7GfGiNyPcNup7yhwsUkwzExuaf1JM0+dhRbdFu/YY8k793TTyfm
86sMUkbKqNlEpV05VCvnxfi6Dd7o1JH3xQnHnspKpCOfN6MhlvbEwB3E82a7A0CjShZgIRNqHnhy
Z9Ylgcjj1BqYDwXxWMaVx7dF0Kt+4gPLRflAIdFLamYLAiKQG9MKpVQRhFqWeIzDiCzvSBOV5tgx
kTFF9yPU4HfxdECHOASgD4fFfizliNyn/Fn74Y5YKVGWdtxY54kIbIMNoggK2Mx9tRy79lnAvFl2
IhSubUw4nVcFAkqKM8bJx6AvlPUreeycgcIIMm7fT+c2Ouw9mR89Ruvm2VuAkTrZivbqtcPi4x66
d8ZoT0tyTINiBdJ8eI6aJXZa8331NHWiToY5bpqMWe7CZ6rzEWBBjx64zZNX+68UDuxsduI2GNDL
iy4AMbTd3dH/QIhGgikJTxVBEcDaR4VLb1wKN4LyxH4TLJr+2wx2upkniGN4lh1DB6aQGJ3w5iGR
HFnMXGjQE1CUeMmpxCiajEOmJ+MDHrKBfIa0JHnYjiXk7IIjIbd3gUS+1pdO2W4zVqGirMoTlGIO
3pqmVkkm8U3jP3M3nXYuqt20hBN5If5Ni0J8CEBNebgLCPmYS7rGpsEx5QUOvy0h6gO90rJ9LdkE
0B3SwOC4/8B4IUJM+8FKdLGyZCPkeDmskzX9tohM9fivJrkE5mzplq25R95S/VeOomTVy5/zsNFM
bCAffjd8fU9Y8oFV1mcWg3s2I0QlcwANaENXOA/qpad+vwGjAKAtSIuDZbmQKR4Qm0hi+Mi/463n
gAFU2G46VrXy0nK4cJP+QptnCClETqiW/pHArmDmMOlPCgA1T3D4Yf+iNK2hle9KucT3jIftzdR7
iDnmCfbwXe+J508fhsfa+6xFA8VthfEHqXx6m4soizf5LCdLHFXsFVgkC3Y0IJaxoOwGtA+YJbCm
NqplSrxx05XrvFAhEISZlW9LMyJxaWEgW6ZWcayTIfAt213iiJoWSZsDvJ/HvDpeUvdNoCsPZZtB
eI/t56gy9XwKH2w0LLQXpJJf6wO0kUTSvHwiYwdNsh4lfR5e4jI13PDubmhqlxh/GRyXWyqljNEa
mfnTgGGZfr58H6TddekMl68Dp5Wu96KpwFU22VJoMBiPpkU6DbVMHxM4WvkmWNTmwvpG8Q3cjWld
B/m7KjmMMX/jzNPj/AtNldHeQhX3sLL4AZMZgSnOIc4v82D98sjrBm8j8ju+BQTOH6FpeEN0TTpl
EHnfAOZmbROVpRg62Se/WR+7RdF35tUcfYCZ3+QtevoExisWhxSEIG8+9Mg+cJ5cm4mV+vt1kREm
js+fPHthvcnfMEnv/HWuS2H3hyDX9+3Pjy4O64XxxAgrs8QlZEWZCH2UUlQBFNBdCxeXCUUQ3zU8
5ZLTobiK5NB1GYHPhaQ62vf5hCIgShCk2oWjnDnpNShclrVUtyxu7Bij93vPvtRMyWQSc1lyYwWB
EnQX9x6odXpDYvMrOYiPovhNZiDyJykBNXX8bx+Bo0W05qFQU28Z4yDTUUndbn5qP3eYZtRQc/em
Yyh8Hurp4Zc8+pdnlZsAQ70sY5n9+audZXEbkmRPA8wGoCXmwiwRBuCxFT/F8u+pE0JUhG9p2R+q
y6jMosDBxSOJ7ejrL7tTqDUjAE+nDAsJ/o1/RKN7IVL4r9mJ6md7lEs3n8I28nU+LcyCqvjaO5/B
iBYR9BsH2cI4cEhhTiqj2qXNxwMSU6R2GkRigpvPo/JG3TnBWOO77pPhaJMMUYjf2mvqMAXwkdhw
jnsKiYzmMF+43SFCZd1KQzTqPYQBUCUl2BvP9XXUA8gbI+eZKZHZpZkafZ5atjPe3f+wNmnfDys1
gnFgOA6UG3pHVC1l6D0fd9Ndcf1jPuUzs5fVe1C/i7uKxH+Iu8uK0FqB2sBcNr8yOkLifJwSx9s9
5rAaN+QIwpiqU+FMIiDPuoHc82uNHdltgspSjLK5UwlLdnEaapJEukoD8FMKNz810ypTGdfuOWiK
UtDJsYGMku6CnQVZcnTkg4rcEfeKqL4WctH0MZ/DW3+sji1s/GNKnyocFc0lufHK3T680nYBEmCj
PPqTcf6iIceGsFLTKOoNA75M/OkIo18pvDDDaiUIwfZtRlyy63HTGzfocDSbfk3FJ52rod1UJmW0
i+3KI298lKAWXHO6h1GYuiq9R6S91Y1AQ+jInxNrra50ouyluo05AobE+UayWj8VqlVjiTTltfjG
PtMCIO4ctjCW7zUPCBHWuC/uKieS8qAQhX0AFf2cuFtUINU5cHphAlXTBl40yIpOxhegevjpi+1C
PaRpTqUuljI1/y3RKN3rNsOTEY7606EHKbGv7Hfa/AZfQdioY7HimxdFWsg2hv+gZfe48vsr2x4z
XryVnFkqfMzAF9H/cvVHkGnMukCtArqxbU+PZWMf3G8In9vHi95iTHtwt3BAcRCE2aVXEDw53AE5
1KX6wwYl59Jq1eimbSK0wiFA7ZyaGOwrZlkSdWihHHSKxKSVPZ54oHWUFg8LdSP/uzN1+Jh76soM
FxXmRSQLloNbwUS2a7rW3gXMokEjybZD8JLtikuqaXgbeYciJ/3pcgwebUmekHL4JZGmxxzel6K6
GMLnrtjGG/dZ63E7oXlj9HC2OgZ/iKD/+VKdBqLqo8qVEe51O7vzEbzayi+jYLWhB1JxQvoceCeK
i8E+Rsfy0zeeFx+pPK9AcOkKBF1lqOK0wDIGObbb4bHKS8S6L0X40PevlvRR49o4Qjpq7ll0wdC5
tLeeHfpHK5L9I/FGKh24nVyBXhcNYtU2k6qmrPuKKH7Whd1gqOj2refz58tu4i0xEBQiDgEJ3ryF
PXs3F+7DrzNgksF2bc4TCpUUUKIUP43T+4dC9P8IXRGae8q26BmK1OFLnCeTBGkHwaRXT9gskNCn
BOJS5FPGR7iXYQlqJvAWrQLilE09IsvrrTrJMkCn2Hy9QD3FoEPUWab0yfmuLKRsQRQHQtdJOaPM
HF7DmUkqyZzWXnEi6bkmhLSloeAgpT9v4INpYUGcdvmQ1vc7nB6PUZnp34qkCx+esAIBRu7sTQPw
GJUP5ilnJEC5sp45moUpTSBoMAMw522aUOvhyvODEIDWI34GUhZi0TxofORFrCT3c7uawc8rhQBm
mKQ16c7D7vaGdvqdhKdtn4PS/Vb8/ZrxfBuasXcz9K+tMruZ8s2a7ftNoQYLod/f0N8jbyO1X82y
2514PUEWuzQVOtBDVXa08M4dhyPtkh1ZHgp9nqkW2aJdkYQIYOXGqVOVe5CnHM3alKRSMy7/cdgS
zhLdNc4n68dKj5y/REWR7S9oOzoTzuG3NmkeoCjMVonKD3l9coDCMJG2E4ShlZujLRJggUqbYflU
x7LVmoFvSRGoQnGvCCvghAv5i6xThNR/k04MGxShN5+pP+BKXy1q1Och0Jjtu9IvH0k3JT6Uyi5I
T2UWYStO0unFl508dGK1npBcM3UEgS9wZ24FKh4TMRae0sLuEXiPgEx27bhB2jfITHbtHLLreEuf
+Bn0mtAByQwYZ0XjS2WIA1kGmBLZPMNXwZdI+3qwgJ4Hkc30uETSMCAQLqdj0G6m2NL7Jz3tr7zB
JTGMfZY3D+6Wt/Tq54LosbKf57yKMl7bprIv04NBUb90ds12y9OSvxljJH0Mktrg9UwDukvbGqCU
JTuqS/TEetwoNJqCpbSvpVTe64HvSK79m+U9HLGp1DPjEscTLsulCxAGLz6ONPDfB8dXAD0OFAFw
zaSoEs7W5j/u9hNUI52x3oeijlR9AaNUFzMPJloJVf4fENarczdST4UXolpAxY9XZDhFLYo7e8pW
Ph1U4OHivum6o/yO4ZQDDyBdasGSVEG55X/VdJDlMIw1/njuyED3/GMSFckN67zW53OqiMP3cQB8
sGltqKg1GxFUGctGXxV86mX5NdWVppJUh3P3b6KSZ0H5DS9DyCmcZVJgNAWNIvRT2RyWVl4zS31t
WQpYs1dkSAkF4bSG1BcJluGFINKX6uLu3XkMBTSuo5MPhD5QiCLnAcrr05+qZeurq9vspqLYhPg9
haT9oLqJzFvKBSWlHVa7wOaeUwoadfTGiTvXaSa5ScU0kk7LQ/qWWQIDfIIGpzqZ+QwsuhfnUdQx
QYgwhyTL0qy+qcIAlT9najYAkCxw3Wza5HCANf+JNYpY8YLGhK0ZWJhCVDCo3W4V1K9CzxX/j/5g
/S27xtlQorJS0594SSvqhw9DSHIc3hL5bK1UEIrQYP6jL8wzQU6zAcOTTM2Dh9GcKBOwQiUESETY
vhj5ZpGY2WaivZusTIQzkvyO75vsEr2sSH/FK7+aRKzi0le6Ud4ngAkPY8i/FyHpSrsjkQL5WpKB
vIq43Ksh8xtlSfoRZE4sF4Kh8tJiG9h67HU29wBJLkRIJClVmy1gAROoMwFVH1hhhrYeeBQPVgqU
y55lyKKXJ1rRMiqZRWiahGzHGeFzSZMftuynDNqxHB+mkPc8yyiynpUJoq4pnyagRMYCYG3H7i8C
6aGZ+rYhJozMewBySWKTi3wQyj7heSbdh+67M/PcH9WcHczoqWeoI3jZP9BRvpw0t7YbVdJvRZv+
FE2tiG11JWhxfkJp6c9Tezu0UIgiF59xjH53iJQY8XvmhmVtkwr6LA0Ex2gZflGlac+YFFz7+QSj
LWUMKbDlsKaUpPJ9HeO8HbNHDkFhiW7a7xqoTDeRsdMat7K+zwxqyBK/SnjjxXIWyTZkQ8ZoPXjV
ea9v0HtznzsYOjrHMpzDiDtc+vmB/80EziPTRL/yDs23Pni8aX7Yuy16JWAlIref2LGxCCT8AKii
hIqvt7Z84NxM/qLI4a3IA05n3VQeoX3SLSm3f8HCoDKnAZel6PHo5k8UonIDtmXqhQGN24fpTnZb
Rp4FrPfGcWJOvrDFZBZJlrfn692wL4Um9vy8YAqngvhDnCCIa1ZeOQuM1VweQht99/GFhdzzKOVl
N1TigdFgtL5AxqNR867aUdWDaGIK/7IaxKwmP7GvpXGsbelXB/QZxusfoNJhkTSCr693vrCJtgWc
9kg+aDwxCDGKIJApxfA9v2eLyi5vqPwIu7ynvl2EYce7eUk211JB3pVWKECJAR5tfkrwBH/H/VHU
FtOXMNi+93gm3Cze7fftaxwG5UKNgGv/nRqEaKkiBWyHQkMIz3VYmEnP5c7Zj7UoeMF1dntpjP2y
Sv9Z/klYgIDn8Xr0lVLcCJIb69ro/XXSzg9n+/F7qDTjsqYqbK8Br1Nvvui40CLpold4lfgJeYHL
zOBTnCcHQ4Lv3ouynsG4+bqut8L6FmSJPjLjLr7MWRbeGsvn0rkATY/bVQe/NIsm2+46xmjHPR3s
Ggdv7TOPgee74AuR3Qp34kmF+Ms9v6RVm68J/6RQ/Dh1AzeioTnVhsVZhBfLfCOLDOs2xaz3vvwx
cqroBjUqwhVgnvvRfzcNHpYejMiDYBKFlM/FFPPgyyJm5dBxB7YwJohzJOH/gXKE/HLSk+XiIeKV
gepQaTJfa7UmgAihupOpQXWgvZHMsexD+H0vCuKaiGm5CKoQldBagsw9ND+6dUwTNaF+Txh9rto3
/dxCT7aYM4FdFwf4LjH8PWiH9O9fj5YO/7K7cf/x/axz+a1+p9Oyfi/AtlQbmiexaOteVePQnxq7
isXkvG3xQFJlhFv6SGc36lHEhG6ZRcR5RamrL92fRPXIVY7pL4XEGC95rahgJTZbn3w9VWqki3Tq
kDEbNBnM8++wUrnoaekeZiyzk/eIRrfLvjkeTwLEeMNqZZotL/v+MukVLqoIC++Nd1wYqj2FnGuI
CaGI7eVUZcGl9z2QxDw6/iJxL2kZ2hmqaw0z5kr6pD0IEJsfnjdjvx2Q7B8lNax7/i6DhGTl1bL/
XyQjaBbTJpBp4m9woB/rx41bdmaZOoELSFmGV/7gSrEQ93fQgy0AXJ7ViDbXYeVGmvlXZ4dkOkc7
Kb8YBVcVk4XHOp7Vap1KAwsDJcDgkQvCaWisbxwaRATCesYBnSSZBMj/y5jRek4ZB8j55GcmDEZO
KqyiGbdeDLNIQiuA82bN/lFb8Mrm3BRXJ385IIqPFWEa3yDVG2OPek8gVqiMkF8ZRQmFvh0ZNMn7
cOhXaE0sK5OJ2iwDmPEUIIhuhhFlTeQitWFjZ+XgDT/NpJBtlJWoaNkWdJSPPI71ULOkiqN2OWYT
G14445fkH1QTdRBE4KYzTg9NajCm0zC/OwTtG7m0W5S0u2KA/dDiO7RHex9vdmK6D6KXI5z/Y65L
glOSGm+mINTHY057LNM5vEnazqWl5/fVsMbaxMp8nMmGhn13RD6FyrrVNjmHO1kE7BYMvs/xVot8
mOf/BJwRkZ6Q60PAvIPhyzS8miH3WhN94AD5Jyzw5cpxSQno6DNDy36TMOzYNlhMnO0GodXSQioN
PrMYiaFcRs+TjY5+YX8KF/d1RudfSoXCb+9y/6GszRXtoU++Pd9JNgJZxQUYKofi//adT6IBmOcB
tE3QrklXUSA3Y952eyl8akXukfy3xHI4D5xOT9Xbbmhb7BvtFbvxdqRyw6qVstx9zrNP0jXPRnMY
THDcyvPq2ADykjQxaKzjXb8nvlB/IVi/hF0YoDLlGRYn2p7/IMLMV2sVNexkdTk/kSOCaIDOv8oJ
nzXLicRG54L1nbXIyPgJ6l8GBPLn9SW6M2Q7SUPYFtm4kF9+VpgKJ/A95iw4lOLdcu5InnOFPBPJ
FGFLoEauE5Sb/xIL7wMiv3jIsJ4aST+HM4d9bjZS6MwvZkqbTgLR1d7nLTGGsN6ynR8+vVDS/Eq7
9INEIN4ENNoba8gOZBJqc4ENjzGCkdDATkV8PHhPxFDpsYLjSI4dfJow3yZLAvT3GOotDW1jVJ5o
9C7v/U4YJSrMpkazGzrxEUwL+87uPDRLUXlRBImuGxUtuo6ABsLaJDpNG1Z/4J42LDTRnk9n+In1
w14xODvKAVc4kqHPPm+CA3QcqKITsUHaG1Spee28y1WleX4tJEkYNNUNtLMbQlN0HJDkSQ1vuyyG
WWGSkO2qvyaOePWRDf9W1NNlXP72SJ4y9auxogKjEfRwGVofbBQxL1CyUq3npwJoNxX4vtEi2RL2
tG8tXcxyJg2wc0FXQK8764B0llzMOlKCZpefh1M6adQsKKNIdLzmNwAqU72mh/SqFaPA4OExXixa
4sow8rBu3C0TaszZ6PywZl+QDL8JB5vTIHrcaSEb606qGIpf/Y0xR00aovuKdGYutZ44quXUZA7T
scELfOYU4/Tt+qeCcsBWRKkekT95ybN49luRGvqoRRIoQzEW+kUaIW1jkTKfaS/iSWWyoydzTNxj
MUnu3H1+32FEUajmfoX/rzaqiDQTr9xXBM1JfmG6Sx00i9v208gojlRXNC67enEWOKxtku3Cfxi+
Qe7bafQvUA5aupuh2NagM+8uABxgl8ZhS+z294Ckua94yWApYLMnFT+y8wjUq20eYTK9wENi3zes
wW1kIkd1SOJhtJBz/FO5YLBqlcVEJerywM28pTmBjETUUKoWoLTT2TCxfVT/BdaJmkUHLflb113K
VlIwXPO5J2maJkn5vJZ5R/nu/qoB39Kz9swKf5riJumdhJTQx4wEtDHpPDH6Ec535hzd3CPLXali
br76hIy3GryTF0wFGmDiNJPxva8QNepwMIyu4VdlPIwxqcKZz62VcDrOYEs3XNxXxbcjRarohFbg
p/N17l0UBMn/inz0AOnmJl5k+xhujaXW+JKbuwg5/avSYLXEgpcW716pBuYwEhDGMJWx+VWiRHBn
m/r2kKkc/2MyxRAEmfJEnnOQoWNYhG86Rg3CQsCsV7JCxmR+U2qSTeaPPbR5A5eduXQWbXQMfp+0
w1w2E5LTeWhhwuBnUqBNmCzoZXikRRhJgPo27x5lVFdyeFicUjwrw8LCiuM3Zc9a1ftZOwAXpT/m
jwsDxPeywzyZiTtdrrkTabOqT4GyHPN36Ril//+kQ1wSdW3nVGf80lA7dP1Mq7L4WJKypTD1qZiN
5t5ZhSnVSWe3dCrgGTh1kFXDbsUs5YApfV/v2wtUcj8IJnQ1eG1Y9yDjHlcMakdt8ZChxN9dCpNC
lRtjUWYonMMPP7yrBz7JOsBENzDqgS6dpvhSXJRKjp16H3AWZAezKMufYKs3bqdUhPIs00esm/Ie
knuStMl7iRx/YcpvjAbfA87TH9hr9Lq74A0XevDMaTVU1OM6h5joCiQ++YQASn+OKHW3qPPN+5Xd
kj4FEihYXJmPo/msUiBxjkfkpz73vzGn89mH0jFnns7dsM1FeQKXiSPwfBYlTKO5dQJx71XPPe5i
S3UbQl1F8e3i6nEGwTIjvlK2Afu1rzMmfnqD1wH3xFQFlpBvBEqfLuSUuQhnmMwT6dO23ZIV2tNV
US0xkLS9PX+iopEJgc6nrkx2SfmS7QvRiVWohfrRGD2R86qunkw3G3tz60gtLypILDyxWafjLw7B
cWuJIRSlBDRy5qjGzRhmVGkDMgd+jbIPng7sRkJhsvAvqqHm8j7vGc0QPRus278EnQO4CI+A3rDy
C/sYlaxPgWULr/ydeNBYByApKjHAIOg1c1wQrDnQagm8G2xfGSOHIsoM4FGzxqRxgLdg9hKvDloF
OIl2+rTqEdH+b4mWKhMzOYjWjLfF9pFKHEP+zojZV0zMx/bQ6J+kKE8qO5QXRzfK8Z/KpmeXcpT5
3xsPhLA7vlyvtLfTKz3+t/luMG9pw7uJsCMo8GtiySYgt1B12oxeVs82VN1yFNqwyIO4tTsQeFE6
6nUkgpd/gpq/dd7qQ/UONEh7yPAF80HdnalfaR9J/n1hnj4oNMAWi1sNMyePEH5N+/vnJhhxsreG
ksiWQhOALzq87aDLs4YCOVMUM4oW46/99YMfOfvaDBOiN+wDbgm/F3sdGE+qFYatwkbHY02xWObi
Q8xMK8Q8AKeoTLU8nmMZbmzGLmYY4U7Bm+RLOeLAyaV7G0qVOLOsy4/P4rBHhy0A2r1ZaoeP/P8N
puuxQn0FxRRubN2EAw+ZgJTkHON46ae2xxEGBh2lfeOajvoeDDQp7cy0Z0oP+H9nNJWIMshpcTFF
ocfeu+13l1aDPzBpv0daVVLw7MnJGT0GcYiQ2yQJfRRGbsF2b6ml0F6F6csJzcqzLWw/mIaHSP0o
r7YEhe4BMHSThyOfGI68cbZYrl3dJB945+4pavQFp0WVbxYNgfG42Z6Bd1gisVknwC3RrU+gFOJ+
8HWX8aKdhq12ZeNMLUcrtcTrdjqhV9bj5JWEnZNKEyFTK2UGl4psg3Oypz4DSHP5ldHTvv9o5E9/
GtTB0I2oBrscz7YTdjZv3sLGrjYOpgFi+4gBPLo2jvtas7YX31vt/4SL5Ot8nj80lUdwbwPvlxcb
RqZN4jqysE3kg/PFQHr3CWa+3TJeFRgJdAmgxFCk3/aRZOn6ctvvARnJoh95L8xl7AWFvAi+u4hz
Etq0Kr0ARbR6B4vrPzngtQOL0RKCS9KHky8fugQlpIf0J4SLN6n4ufhUx+7lLGx3qUwlGZZaNehU
sJCxyFn80aBqckksNoL94KQH576PSQ8jwhZIFIps0xBI6I/tnwk2v9lj9SqJe6MoiJGsgOSuiW8O
6thAW1xjSCw4PaDWsmPZIOmBgcYwpHeBzPMzFFeZjKyeRDYV/Ops/DTIQWgtQS3EG+/N7iRb+uIG
XZvmAskv22f7fyM7FERZBd/Xwt87jDAM4jSUaPc7BjQsfh/FeOtsn7jGWUMVRm3dkykPqlYgStuX
hxAnnVie5zKvYdKTGGLuLKkOX2EmtCeIyQNaIl5tZLTr+44vE+TdrarhICKnvPFre1plCWIQOv6I
gQpH5996D8y1Gb2xWUNyXjAZ5Xs18qp5JxCVPXqfaamKR6aNpbgRj7B6f96dlWz6kN9xgDQ0L8o4
Yb2ozGaa7MFM7IWgGxZ805211C7aQhbzurCPXgWE/6IXX5zrULYni4Xb70Y+gh+y8xby6u+p2efl
20t7N0QPFwbKNClxDl3fU4skMdvhn4ErwpCzvSHhoXlHBzURmd8A1b1AUL9YKRtsUjObOCBljP63
udmhKrPHuuBRKeFK4EYo+tEA8FgB5Mo1e32Pmg4UdY+DhqGetcfzB6zY/N+4Sbb6aTfqtSbRBLxE
qrnnyzzktx5HRCkSjhdgotAPaa23nQGCbaZXUoQTi0VwkU4ldLFKzfGt19RHS1Fru3CXUAhpsqnK
Y1dR66/mbkwHLn2Gh7upxyzqsii23iiepmJf42ULqHMfeuIb4/UGsaXALNh2ROxYc6qjMHUDCxl1
ajpZh55VX2F0/5NP2161/Q3xRiAS0s1K/PUyEZ+Ns0Kx1DnlLDVCBDC0H2yK1PfAOixKRztvIvwL
SBDu6zqMs6wmTBzsyklR3wMaCRt9k/gOR6KCAsGcYBYbvn8b76fiATFqoRL90GcrdWAkgECw4Q7J
ITxYqaYSnJVdbDASjyPIsSCir4FkJLDivhKGRA2MBILbHpv170z+9UgAlx5dqp/HwbFUJuVNKBTG
/iDJ4/OOtDBRudgbiQm9sXUk++7YRQBR/fn3+32o/eUxvUS6SP0tqxIaXBe5lBHz5j8ggdvexJ3j
ilebyxx/wTouSFtR4zsPSLX4+J4mDOHDi3POC6JRmI6cBm6atlGbk1vqjcVuruZOJzy8OZmNq+Km
H1e92C2AOsV6bUMWLppd/Ar83jy98FBBlW+2mRWFRuCk2qya1jiuThNZ5XxaJikONzjrYoTtVbix
EkR4emuO2oNdUCjOyv9Hph2MKr+Z9v6HAqPQ1VlE0/67D0w+jd6BGQEfVdSf6UUFg1psZigZKAUm
OniwgV71G0vXRaRER5kE90nLScqak/OAtdBAivHYdVCMuhdAvHi8ffut8l1SJcUAr6sznmY3PRw/
9GZmILJfeZeqIYOSDLn2MNVmiiqj7XaYV2zCBM4rz8uwtZ9CrD+ceKFu7Lq5tJ/NgcNGcnyH5zsB
N4P2tMVl0Dzh94W3NycH+CpAVuchj4ZQppvgobOb/0LNHVGomZVQelFlrvznezHZspHYzL4SizM9
5FR2gAHz5WcGfKGYoiNqTuXEfAzUGD5DNmiIDoVWZdPM8dzhdXbQZAxSsuZa7tx2XHjrnvj3X1iV
1/2C3wKY5sbqYKw21T0J4ZTMv4z5XguqUyo+fQn1MKN0YWNe6WSDaaOULac8OGYeQhxkKSJBv6+K
qtD3YzstsyDewjg9TWPU1Pjlw2yJWu76myy7zmbK+NIgEIjgohrfANjfng4FGRtD71j0IQSE04i6
DyUipEwFC6AWq7dcc3j7YsluTanjvYe4+uHczofV4E29ufsOmFPNNBQ7PQVZEwOOozcUgrJIbtpX
CIRjZVJ8Y5n/d0HCyJ0+ZGeS3YVWxmuhz5u2/xl874kJmvBKFsKyJ3SsIQgSI+9lnTl1BHUYSglB
acAk0lcfSRK4hPeNxdCmqJgmS6lF4iJwlUpsQ8cgElfHeWmjjOFbR1iy7fo/CvlpeFadnAtDfOmS
7Eig3fJyTuL6nCHtpqQquZzaH5D10HKIhp57dIDKF+nexkWA86QJzewHleFXM1hIGZbCES7eNcFg
Ndg9+SHtxKD2Xpd+wKnh+YKbpnXKflpDV2K6Wo/dMqdhb4DmB8wkCHLVz3CGBfS56q7KkZrAxElA
Vsc2tT45Bbvin2dexnPsQ2UHBrEIW9wqodYt6D/MqnPBJ2PcFuj1lsNrS+9+jv9uP6BhvJ34Y96h
01R0tsY7jgD1dO9QV9eAAlFmH0plZUQ2sdz8k3p5YRs6zKGVnjsCifI9jmibay5qLvpbHmYTDEnc
MUM1JMQdH2rc34b7QwkUxvJZCPiuleylV03H7pTEeL1vSR5EimGOf2ZHC93SlSxXy919tnBwmoOs
l4ZRzpV3PAS9uv7VNo6mGyuaIR87cV//CGRvTgTjtMFCBaYDCuE0gN5d3B5oJivP+HMqR3/NpYkY
CeBbNhAzOWEmDSVxwx1wmGjl3nx1qCwVlPs7w5SsZlvgXHxto1aqWC0fk/4JjemWeVtrcUsYpcwn
Eg2SFUL2AG3JE/JyRdx/QbOKBOA8TwdW0BiPP1De2QumkP2KllRy9n1DbtfHWc+DHsBaTlVwU+P1
Lkca70yoF9MV8VibHmX+OQ+BwyOGWvnEUGxgZzD9lZ2LlEUz876dAE+e8F4/SNKmy7L+Y/Q7TlsF
apQuir2l6FOxpLMe6iiPNZF2LgO2/K1yPfdnPjbWXAFwDi0WADNNXm2Lo9J/mWpaLkTOpRMUStiO
SamBeBCsFLhyLXs+UfNEYgly35zRmyepmd54TkSs/xPzuN4Frk2I40oz5precwi4GlNx4mrHQZqD
5IxqGH47xhctNL0LTQCrk84cxVPfNGEoJlZKtYIpTHX75s297C4tXBpnidRwty8BkMNVHvmH7mkp
1neIKowvtJWj7N6fcw+lGsz/n/s27MGzho706bdTR8LRUjclnIvJszFAFL+pYDIqB9WLYEp8WaHa
ynoPgmn4/PNbVCwqGQcANVDJMoVKuYhO+NhTchBsfeDiRp4TB06d/kMNGPDxTcMJwfThkEbdyi+R
oaBSD1RfOZ0wxVvhuH5W2imXnbuMqY5OuQK6pyL3YyCDbasdFylleSdQ6YhGZtt0Etn6i7Uo7DEE
TGYTRIWnsyJjilmIkl53Cx82ZCDJ/Eqkne75VqhsuE8AXNENDZTLimbRtzo75NduvEG40ZKYiHJu
4G6LZE113zbxGnZNpLbz0vaksqL8n5itWwdUBCoktAPC5PEs54k1UhVPpVfqtrdfoiXNSisMceGk
QS7rw46EM90F9Xcxaq5v6QE0MUrRqej36JQ351mn8rc1QobKq5vxU/1x24kDBUSV8BS54QW1+CJn
F28CvO9t20VZRr3ivPIBDHTmXkHGgajqIHo5sk98HblLokukPohL6py5Djj35E6xhLDWQWxaxrHs
5W628q0uKBzWmqkimIfvH2NwhuiUxl/NBXyWQZCmUrIPgz0YAE5DUuRwors0rf5rjvlw89gK1Sla
9HNKuZCj5VRZdkrcoLgtTSykaQtS1jq2fV2ZOjtTzaDaFaxsyxq21DsJ99HTdj3oadVNwQwx1NQZ
YtliKJPgK9ueeKL22jX0U5pwha6g2VHIv0VTrLiImcgOuPdYAk7XJ/+Gah0TQ2eX2/LvsMgnx4DI
AW5o5+iv6flzpjeY+/vFDoOzloaO/24ZqSll90DwArjTXUf/pVFUcTMjxkhgu4DejWlX7L1NZLYY
i8LuRr9bQBaYoJFuPriZmAcISK+jeARvKrxF+95bY9tdgzP7/uuSHSAr2B9q7n29mKW61clD3zXg
Z+iazWeJJ1JLTwFaHO5LrRZZQOgFP/caaPHHzZg1Ee5AfVmRUsl2YR96g7j6RgYk0OXUTeI//UwG
izRpVgbgj6Sg14KuY0viMrW+ZiWe8w1nohqjiCp1IkcpaCCo/NqE6XeWLqzw9LeqcVNgT4A+E47p
3S5Eej+Fy/PaKA77L68/NK7ekIYJxHf7+Bre2jysVoOhmKykK2akhYfslvJ3NZahGQFOZzqRu1rl
NlTdfiCD6nPcsv5VTsgOZDQ8pOHT18f2znvdWsh8ox3Vco+2E+c4q1acoPkqfLTmTbaB8QceyFgK
fIa8ci11n97d/LssuZGjjjDO+LhxYQsrrtrc/3aGaFrZaxdy8xqYpAS5OVM+Qo4S6RpII9U8B7Gk
cPBxvMS9vPw7DUqHpYo0vZ8UXWCzf3evjsfLad/2QU9KF6DEksLjNdeRb/8WGxA6iQY/It7rgS/r
4FFlQFmvCCP0k00DGA4emEDiv/2Tbhn+1Bd4Kc2QcubV3bwOuxpzybV9af7cZKco2AHpzKyJbXd6
WiX6YKliisJ1CFnbqydVXSdcEaN0eiZ0arPNe6xqthqX+OlP7bqPNlrr7RNf6NdZmtxB5ogRBTMk
TfQ7mMKVMTFeeBOfW4N/sBLkemXqKHRxT9s2m8vZJJIcUlpR5n+y+/5lG6YwqYK47lFQzMpSiiw8
VU/z1GyHRa0/QTCTwdqBJXn353rw+KPlnjEYc5CkjCIsKAlluvMl/bCT1XJ/S4nbeEnHXUG5ecV8
YXCLa2bLNi06ooj9nmxjB6184qr+7RggsFvsrQxA8NAOntG9LiamK1pkmu1/oX1QskWPneuizkby
IJ9fMalzZ8ABmpTaYKF6t+v/H8fg4RVkkQQY945PE4Sf/FXa0XB5+K0q+Url10JwTVgdkJ2MXhpk
jjca/qa4EPEOygZlBtQ9pRnG49dc0wTcXI1XVva4TFnN24DvqnnsjwoOUnU5JoVrryz85DecJQwK
sFElXV3uWDlsF4492m3EzGDYrZfRr2KiNWDDFef0HprH3CSeB+eILvMHOxiizm7NgrGbP01jAu+g
yiUlv2zr8JI1IM0QnsZYEds4PHrUsWUNAc/WuybANc/xn8w62dZG6PvhSbLl7TDBZ3gcbsNPpGJ0
gBN9O7icWwtmiTHrwsEuAx0UeFGQB6mG6wJPZaJJac7bRPmdVyVJLiudh3xmY4kSoXq67eSy2Lyk
/xq5I3vvWjwyPbNE2hrnqrRNnBcEORYttpvrUc0gUCf32liTKJPJw1CswkrhTs3WMmJGhFo0Bedh
hU4abP2SXNdB8SCo1XCphI7taavl+dyqvfksdi4ESoobeE0Z52wnRHcgVGpe8uLLhZbnVLyAU1nV
/nKV+RYveX2At2S8698la/FljK4lNyeFf7pGJf/oCLJeTYIcUZUmNX9ej24GuuKYmfWJDxm4r1K4
nVd6v/45rQMzSf0s3FU9gAP7WQA2MppWlGJpsVmZF+r1J8pFFWdFwYz6BqNNpsvaom4aWpqQ3Ezg
A/NT2gOrDjM+uySXAZSyzpVWKzg3gvSzMpSqVw3JwvPiBE7N2iei8QCBDlG0kPWp3MT6rCro3h8N
0/0sMcV3bj+3KS2nD9C5CiP9cupRmaJpbaPQ7qORlnMLZy6xvOHf2q4v/RMMICL12rVVdyxrgC6c
/jXbhdk5LbTpIYgxrr1akNSOJw2+PdrNAQfy23CPA7zc+9whGV8E4fJru41iWhXgHNdoCkQ8xzSf
ZHk1VC5CUOKPNjxRxvHCwH1WAFKPmpNCG8bbioqBLR7Mrfp3t+acbMSIUtF/CoToxN3hSopLL6lS
fmX0Q943k2PU3BtpBUCropvszOEmL1JmMi6xyNiu8bIQPN/wlKkdNmgrVVpCVMes1Alg+eRLp5y3
U9auI2HyQ7hcLwbU8eVS+3abAW+eXXhSH4PYznIISuKmtPMYgY+16kOO5LLjC84wKRIv2lLNpEml
h33WawvP6jNWAxHT99HnoI9UtL4P+kYDUzEgDVFSS8M1w4lSHMkzs5XTaMH73E6eWwNykqUJb8X6
yez9Srcdfgx2/YcyUvb58EnoDoCtCZily0/UMr8mcpRln1A1XaqjrsUWZFViW8B9NshGkQOUyicY
hMUC/mS2aHOLs/fqdcGSGgovzv/wq2k9MFqG3Ac3SyClIra7HjuO+0BawL/swm5YnNd/NahlYoFn
wSiwglliSyan2aQWlriCe+VfWw70uaSMR9M7qoSB842TIFX5gZRQ2RqxroX9wxwqD7i1QwjSev/d
S1U5UTZUKQD8GIxPrk3NoPhSte1vCSKOcias37QBs5+tBN61I0bGue3TQkd9+Iny8MS4c3erg1b4
PiR0nUNfVAJuVHeb1k8Jk+CJLNFs+8EK4koY8Q05wffjzXpgG7v+FjDiNoXPOQhkH5vFKg8pbpA4
fEaEkO0eaRbS5qedEVE0LPpQBQRDO23soR3GNLdQOLx595P1XHFaK2s2QPavPjmoG5LGjzAFcv9n
KoLSoba4W4YkE/xH7vfIrjByZJ6eom3jff9MK1iBnN84eHYnaoL7ERsyoiaDix7Kb/5DMA0Lq0j2
KcRESuQermjpM+cRr8tNVHZEUD0m9wV+DaK+fVgz3M8X33XlE2jl1XNA982xiIS/b78U4o7Q2QGc
bR3zhRDMQLtzU0Z86HNEqWDNwPJ0plD0aD8VvVbAS91aUPnQsuI7lceXEJLrLRjhyY9irT5fSmvG
/uEfwUM3k1YJHJTCpPVAF/39f2u/6IjQ6HYNp1f/TSyJAxakarV8xxgaZy5O08L6iaq3YlFnRC5I
Wa//bGhdNtMUf/jQcFuciYmY/Dy28X9j+MfoVxLZyG+M+TQmN7XacFmIGd+VX3mDpiBgMJWscEsv
ZW6s0bx5S6flVlT0bLcsLQisyeZKn1fZ0/ADHUVZgfTWhTn62WMJQMjg8ohKH8rxvR409OXSXqCg
kEp+ajymtmtq47mcu9/uMEAGQCg6tZyqvlH/JpAV4mybS9vC2C91amvoBASZKmJA1NSazoNo8KYk
HLaZnF7ywTlCCtSA4oAu0174CDckm6RgydRndOiE2+xl6PrXfDEuzI5juySOPwr582ahiryUQLPf
wY0xE7A5t5J3s3sIZoOnOlzZmAGns9EpkTe9weDO4XAszi9nVlps/fFyakTHaKeDUtexIs2iwTAn
82zAG6rXInlp5L9oyROnnc9toZ09Pltz2NiFE7zl7fhLyBF3Gyrw5fiCfucxI4BacN5JC1YCL+vU
Z7Ga7H2StsmvcBZy4b9HmnvCoV/9/WEq+ZITuaj2iT8+IZmLscJCg9bNVodp91LYe0hzElIgaJ+2
FyCqt2ecp5yOMuD9E6EsTtq7q4Q84ti1pITsWEx6utbEzuCwU2fvWH+gLknBHOAE7fvh/bF5vliB
+Zr3/V+OGbqqYBMAel8Wx+FpT1z/wA1C8peDFyOjhq++FLlonYa2GHnRRuKF/0Sj7snl2rOQvjOz
RXtU3VdG1RLYE2YYvZ2gV/5zQO4OiUEUwEIwLNhiKdyU2SV8tMaIXif+o/iYk1g+rE0fj7mYowty
ca3JHsHhWmLyNkXo9bEx8/g/zoE+3nvuT6hYiMbBGNqDHH4WUibSvaCEo+JQqVlCBXUx/Sdo+aov
R0tLhwtK3YZL0So1VasdAxA1dgVEYk2nhkvw6B2kLD/L7016oaXDg6zXKwAwNmvagRFwoqqV6+7X
FA0FfzRYi1czWvfHc/ZNY7QeIUltGNkadnSHb+lil0t/uE+N9/Kh17wmTE3ds/j6zROoWbjKSE/H
XSgEWWHeLlRbwoqi4UhuMby1amryJD2Mo96YoD9sthhre8I61fNnQIMTtoBxSM9XhaBZ4ACDMUEc
H4mNSi+TSyHM/9VRhqoVAffF3K5xwIzxMCSqr8pyTqfaAQ0D0VU+3uOp7iruhgsxNnSO1VbhAtDV
vtqeu5XxRd4zvYpOwYQCvzzH5BBM9e+yuwL1sHKHTyKlrwKbuemy3b1hEJGVN5obXeQzKNDyUnBa
99GsObKkWYWgFXfyqQ6ByEfsztaLAlcbGbbx4oQypmleDpXA08A1a80bPi3OIoQobO/Hm2xoGqmS
AwpXLF3EIQRuFlVHaojuOH9xJFA+hgUbDovJm2oiiicQ3Wz09RwGbwlSlUmMkwn3QT3KZux1PY5g
nBZYp0icsy4n/zRaSyUZiNlo4gTDcS1iPM3N+kuBf8FRJLiNz6NSeggKRJTjdVCn5jGOfE2OmkYO
6sO51Bxk1Z2/fTy7m0VX1locyBvgvi2muvQto2SjrDgQt3oISLzC/0eg7ZD9B9nWbqYvsRexmgLX
fZuvtrGoj78dKU95g820GURqzjtYVFzj/tkRNlu5m2MCeEssWl/P+Zp9vAxP6PiRZGikWCiKBS2a
0RFxQ5emD9sT0AU5Ki+KJxUE/4cVYoZ16RNc/oAoBTWeovWVGHkt34GLw/7WatEdgZaItQ7HIZ5Q
9ootCcNl9lfdkGFPBUA+ewQFLdwhy+qcBwWsKTqp+90L3oloywyU+gAOZJhnby0WDKcGbkctdVOK
38mEcXleT/yGPTEcSqfS5xCgss2m2DuNZv0sxCXLDxANBO5NRJwdVWRjGph8kCK/KQ9D7ArxD7a9
5IPy3OtsUUlxlw/NzERg/LRmAspA1PPybqDlAHBCfRnLJrGQyEXdhKIwqtyYLg3rFmdAZ7rPlYjX
roxf4mderUrg9iHKdofUmW4vrBEzv0EhmRwcW7e8DSLGvzPvu53ks8KoQyYRvNy5u3zpLNwfKt56
KYNq8XVQNcwaIar6NSKBvvrf2gvaehz92Mh9fbSbPkF+Ujh9z9RA2L9AURBysYJY0OfsLwiz97Al
PmrM4rkrGYsYTidDs7DcoyPXrg5L07EFl3a7QzCQ4EDbFAOU/uvPONxv8CNHaxrPSSFyTBTGetsn
CsWIAUQSRw9DnMjO5WMVzF8TZJuakHf6/9+9VTscE9JcViXoAN5u/WrHC6IteESAtkVheKOXDZYl
UcEBaaDTXTSFv0e05yspRb48uDWtJ1FWc1QPwwZVw20EWeaOOIT5QzQ5dKSLBEGRcZNHv//iNKPG
i6MUba+rDrAdy9Fjn4JQa7X5c1dJrDrF2+ZebyN+zqLXvLbzUZe7EiQMDTLj8u3qw70STrL3wm2a
43omIvZgBotqFDM3YE8majbf7NmSX7HP5B4b6gf3beArZjIrWOxWlOHqZ4iUonAbvUOcqzAVpkkt
wl7moIGzmkbGwYf/4o4DB6PkZhdRpyDIQGD7Xd4DCjlgJ9/LyaeP5LhkRUXF2SjaJmM0KzAXCw5q
1L3+vpAWMedZ3z50FZygv6D7qv2+YX+9DRoqamT7a1oA/4tkHFHPmbMwEZQxQ/uYpJZ1rKS9gCBk
WsBA6j/5QKLyGxqE+Amzobxtud6x6TABgSGCNzXMSXQRRCVdQzYu9oYMDKF2Dt1IRZGDkqz6L4+h
bIk/8Ts+tczhhcvEiwoI0iC+KnN6xqFU7eV+/KyxgrN3Ur+oogtG8isebZKbUzGp5fxbBjKHv8gw
+fFIK9aDGmRJ2fmo5+NGFFhXN4gLWW66hPWda62t6q/v2OHXxAE84JNir1LZjKf7cNW1v3qarryF
8NxhvYnZqftnWnpdfUZIRFerBCvv5Z40lA2ysre9ex2Zkz6AiqdT5491+CH9NBjyiyJhvVoyZ5p1
I/ymFB5Nu2Uf5qCjCTMPQHBOXWMigvRCiBolFHZxu0DW1+xk7lSBrS+8YmHdleI8p5Tt4B2Dehc3
W/Xff0ktf01kpulFBgSz6fooYkWaLijg/8a16PDJwvo4MgZ6aqNfIzOCpwfPHuY/Cpt+UMbmseKO
qW/aWSdiXlmXAbalFa7aCqPa2xbpAtIpYoqPxUtWC11lk3L0yiCQDXGLUfsyD8DcttzbnIuO/G9t
7PYiubm0mZQE+EuLlaoaB5IIOgCNHRjRDZnBIP4bAOgf36g14ajzKR1LUy320STQ/jZ5GWaFZSO9
iass2pXrEbbweEkq7NsEPyEtGMmvsNfcjtXjQVAQA1Nv/mbDWXgZn0GdwZfhWfxEfCAUEW5XJszs
LgE6TxfEcHdidmEe8iYeyOOGgE/OcXqOT7ZUvZnmcYd3uBcBr/u0MaL1F+BSTmlEAF/85JCx4X8I
4wZN30BWRIdaTXlMKpNARO+VydNiDOYkg1WiABSpdT+Qb4slKFWX9OX1UKp6NckbNBtpzQY73aOb
kI3oqa/TXPKdCkBS7gKlLAWkTTirSdelHx8MHUh2oHQJusaXaGQ1alup6sTj7q98N4A+jAERUOWj
i1BTGr7rk6ygOOeBH2GI5G+SJHBcknBUDiw/ppxF7KSYnM1y9I4raOJ3A9WdN97uDAp26Ztt25X0
X40/gmRGrqr3NmmDcWHVpxHxUOpJT1X06E4w2fMmWFgutFCnyOmka87e19wckbF3hBpis68eVzho
o85O8UQLN1aIrcQaWG/gO3vXag18oXaeLrv6JDx729zy9RZHKLziiVDjrWqf/zLXVCaFGmU1MM5H
73qxIUZmtvuR1cuFOLTmwJarPyS69YC0CnfKeKgzxIwKz1NgHD4M8oViy89dcR4lR1LEB8a0wPKX
8xbdTjfumWqejjsZrXt0/NarD+7A/j/fNFaokGWg9cr2DAIPQh3w754j5U5ItJOmKLajbNlV4Hsb
cG9xILiVOXWVKu7aCeZztgLbW7U0eV1FDnUoB12O3LusLnwtX3730b6Hc2VljO7I1n9vKVZ+T2VI
u0JjxpSyCNOCVaeuwVFlS8RehSPASQ5Qrm8E/Mdl4A4E2wbStxJw1HlNy4FAirbqm9P2tocDy1XG
2XPh/8PM+CQzrPpyYOnuOaqd5F1+vrn9teghiYmEuOMXjXIkHQOFmVSs7z0lb/L+ak7LL4GDkyj7
gIc2/VM/5yHrU2GsxUfOSmhGPhP2o7ozuZagq/safQzubOQ6MXAPBhyhz86u0hSB8u/QQEs3/rUc
CkaZfuHmP0ra+x9H++hvIR//t8j3eP7ZTZmL1RajQR7ROAOT/9AtzL+8zQuZm2uFjngz4qkz6dkf
oCsoKDgvqmrOMPHwQ6jb2/K2cNdIquUOS9R9xl1N/pa6opF/iZ0wnP3GMR0dLQpwO3QqdRsc/KSc
yLBe+IJY40UdLEyHnV7wcxbo1EQ2t+4p+vtziD8k5R5EwFLewJxXqH1z6k+vGjkBKyqrMXb4LVBP
Y7Dp5hYBr/vll6aoG4VepMBh8kQg51MDwPHCv1j7GXL9q2bx9EygItglcyb04U5Z4A7usUUcYINI
HjTQoICt7zipC8eGZ6e2F0BP1XYEnfaFF5QS7bpy1xGC9tVWokI3aYQlLJMhEdJ4ErJYAGLiuDk/
j0dOKK/0zBqlnP358yY0RHLs7n3bGyP2981SmzDBFapygjrsXT5RXAD7ARQDGEbzbTy9H01bNw5R
zHz0K8VEPiieHoudSBi14x9J0APr9LRSns4OHoaQHR4+zx7pOMBnfkRyftYOyXQFwfYB0vtkn6nV
5p0mCdq66JYpIi7esg6BCnloSx5JmvfV+fdqegI6aAujAwFDHDftjuwiyEqojn/r5Ze6nbIv8cR5
k3On6eiQNf19ADofBb2KRIUfrnuKju5sPueRInflpKBXuV9LjqN4erlGpZ4RRqFiWzqQ/yPv+Kgh
Pw+NDVHRTLcZodHpwkqCUJh0945R82denkMSKP1YD2jSWBv6kWpDAPHe/8bpQIeTHXGcO1quJ6jg
mbXYyYtwW3t23za2e1K9TAeh4PfB+AhK3Q03bD1NWo2oi5IZGYmvVfdYRriOkX7UvhU5cuHj9Uus
BFgDfBS/oKyQTHGW4X0Re6QSgtX/v2R9FwbQpm8kOFiiPh37BzhbuvRuLkHzW2+IPygNbnLVcINW
26rgAhyrIcKD1YjRpywpNEv1V8lEMcXkY2hkvP2EwB19mvdXPnwepRA0f6f7Mt0QlnJ3vSGgNWGU
47sqpf77y5uLqcBj5j4Jjz9leSmTbSMoWvVrBwY48QSlg8TZWmHisqBpqlDUiweYuuVM6V8Wf9BH
uF7V8K5JpQVbLuf4yReAP0aofxkDEXuRLDVbh7cScz0Aamxc9g3rMLIbO9YgmcRBJSqPTcxMT2+R
Q++9JUbwa9liEVMmslCjMtW64hpfQitRMwchfSqjk5X0IGB/gyX5S9qTNZOQ4kwGn2hkyxJ+XQO6
j1/qsbZ2W0KK3xARTAi9DdG4/NlHQxnPtG3lJnwfxrzv7Zfj3VJJBKsd3sX6r7P92kqVJwG0PnIO
N+de8qbWv4D+IiSi+DorsoWdnOLgwniLt+K8UBtmv/qiZWA1Mo/DIHPbS+BrlbuzJxQTfpuZoh/x
AEBjghgsj6shwgwMSzJzreikz2QzwnKAuyZ/piadVkgMXevBBcEGdzGI+woi9GIR+mdddAPsbjRY
+6zJkM8NRcVqsDYjpToIwMMqUeKnl3O1yvaycEcep9evfECTOIn44IibqqKHJtNKkjV+GXX4Xen0
ZKOo/LmVBDYdRY6SByx5oL+2HsY4PwX2oQU68hWtaik2k8EAQggWrLIDdmqFZE1M8H1vLj09rdjX
OaSwFAAObO5jcr2cqiUUP695Mc2yoJsZdYirIJszh0bhT8cbpNXUeq99PYAs0dzJYYv8uKVzO6m3
q6uBZ39MTdv5N2uxv4O8QtYntvaMkeOYs1K78roOK0BJNkKwiPrjmKywdIrTczvSLTpzJwCIVOa3
b1gplmrI2cbEUgu8f0437/Uh28f/N3ztlPC8FBAtoC4QAPBUVkhwGqayIRlccGb4h/8vjnCzhPdr
eMgxRI1VpuKlhZBakuTjRJBmfRImmlfgrPabPzAPsP/cehLeD88CnEZ13ZDbySmsB2QSWkpRax08
KVgDVaT7WTjc1DJeZ59cSnQW6f97Rb1dBBkrWDeWu9YaK10V8waXLJYaGnDXqAku/EXHLOpsuMHg
qlvxtcaKIgFNDnj9uMbQ6UNanc6vly7XzA4wnl8kj0LvJx8V5/jOAfq8Tev3V9T977pVFKwAsV94
lMoh6S18hfpHOYzNZ/Oj70X0qIk0ELyr4BOwbdgHM4/qXIp6pOvH7W+jYooeYp7s7j5u1cNbtrMI
dcqNUN9TrjcbL4joWaPRX2ObN2cHxt1UtNDrs+tlAI4HP3SBiX7zkck2Qh9GgZfbrSAS93rJbAAa
se4DqrfcpPnW3xCChnaHqabQ5uq90LLIrq2MEdQNmvU7XiTdz18VI/rXhhTHdvcmYg2waNLsSL/o
Lns08GIdh2SYmhJ9qrQkvwQKmEj+uc7O4Fwcb58ukVoDcjUVzfUfpEHqK6wV+YZAYZIfJB0XW3CM
KltvuK8jDSkc+zmdGcd77oueRfgjjqSY6igv+2fTFETTC8zb0iD7+qkr9u6U4ee53BolTgXBoXsn
8kFyHczyLnT/4ZU8JodNX655+lYN85APUGc3nOIL7c/ax+ylOy4VT2BGtsKGPOEvdbGOu15aRWqN
USE2oWwFap7cZVZzoa2UiZMZdXhk12qzPdGvlUWfOEcouXHg7ldLVb6H7PXLi2GssDu0Oe2FN2sD
Y90I1Uj0v16XEYVWOWk/7a1DBfDpRUYilgPMQ4XlPf3YAv+3V3UyyQVmewZY+p1AZq75kyheRK/r
9mNSfyhOaZU111oO7QO6o5HmbTSNUwOIZbHAUrbsihUUMLbAr+sMsnVtzY8gAzn4zKxLBLfijfrt
jbiZO9mW1N9KQGAJihpKeLqexjNQVnJs53LU5XewR48ppbg20JGq0LojD8UqGnRCY2sNjdzvcv06
T1stUirmLVlTBG8yMu2v7AGZxbsgEVpyrPYEyTuhZTdMRTN2xRosNT7XW9mX8Y3wKkNy3NUHAAjE
wplYb1jRF9YylE+rsifzj5VIicX2rb++Lo3lyFtfrUIsNcFxc9FeBf1pP/7vuAca/ExPjWSa4rKg
X7kyOXDJzT84KUiUryeIr984NSrZwsPMIg4QbnW4euLx0JCuxHnPlaexSBGejyREthYxACy3H5/V
hkuKlsfvyZpLDBvBL5XXsHHGJYMmSeH3zR3t1eBjb2KcmkH1jOyj3KvJfTj+S5+N7gsjAOdELFoy
+f6iO0F+8jHlrvaBykC4ljN/BQk7azlOrihKokPRGGE2VAY6QeD6G0F/DeD3Q66Bv04j19z+8RE5
kOh2bixN1SuSE5S0CB40fxN/opZsuS81TyfUAj/dZN/VH7CIt+W2s6NIXclb3e3mj1Kc4vmx4XEN
Hk+kKQk21eSYAXnF3spru/wI3a1YAidgdQSkpo4u/rUKn6gqiyhZpl/Z2ojNkLbDrzK7EodF4qXD
y6J00k4+95eePiJU+GvfTAujS7K8CI9C6ws2E6MxNGvbpM5Px4ybYBUdLpJCfqyV2RcvbYkjy/WE
BsD6U3pXBdMc6ynPrw0evVOEv8tFqRob9FJ57hWnIao33LAm60deEdxabGkQQ4m7HYIdhU2gqliU
3N1YVj4OOOh6QOgctAAd7aqz1E8czkX0giJ66Fnyri+dWcq7DnNXEFDJRhbV9dFHozTTCF/COPAL
q1HalbJxKzkaZFzJyW/WkCvQCQvN87bpuRJ000YjVq8yo8QVrLDuXWzDV9JdDEtCgNHTUM9kMGoz
3rG2cA3vuFecW88m5Wvy61hxOMmSwWsw5cAJtkA0XOj2NtbzhLwU4tIX0z972o4DFkQU0VOzaeTC
/0BowFXOG7L5ViD0wubSQs43kBghcYhcnMbi/9kF4SQDxtHkJFv6fiGXGSD/jF2vHBlE3+qH1aw4
n1mV0veenJIMhgi/GF7B1MURnsk3KKhyCfEBGfSw3OfVXeC1IAd2k77gQeQYtCn7TNiBxYtLDTGn
+0e3U3zTIMiADvF7axExg6ubl80S7KaNEsDtc3zcA/XZfYXe5xjbbSRc/da+X4MhC/XYITEHaXNP
gvSwMewcJpQiMYTL8JdevZpbHhY6tz+7ZHBtorM18ny/wQO/SW0+Xyf2PNUiOSVL3a6+H9jziaQX
nY0zr7hT+YxtMrNYteIPQr8jMuGcdjyTFOamPaJoR6KYIME2FeXAlEZMiwVDqwd0m67uQ4lbb+ua
SbQFdrDbDVmYHDAG0fjHEkvQZ54NqD3bjZXfH/1mF1u2L2/v6Sfv8AVQF4l9RVOA+45jgs0mVv8Y
cPsAz9rMmt2GxP2dY2CGw0KlVBsL0MlTJzk/xVQnSZOQw7FMx0Ix0O4c55eBLbqy9ySGNHhQuUq0
KQeilJ5Qq2RtGn3rbotVk3WEcWMbc8Zp3BoTBzu2qud1kH0gZtZ1ifuttHSmhfkRGpEvLPv/eTsP
v/sVLxModD1WGK8IyQHkBTD07KqMQHxBRUTQUUD9XnyFsnTMjb9kwxTmwz5paI3S7a0bJ/RprFKM
ACZYRRo8CTyeSJy5oiIAO49dZPVQmPmjPt/X/Jn52UpSrQOhc2Y4RjgAWprKbFJJMI7oemIncMxX
4G0Y2a0UKjAztkAgQacrmXp/6XR77adQhPem+0tihULwCZtyfRsKruAjDCdyxLI0pa8STsqUqxPp
8s1I1XuMil2TWERc4ZmNpa3c2rx//uz5t4gDVvo9fjRmo99ejv60q5d5wAHu4PSEiXyqR4mreFbS
xWsFcdvk7i1RezAZRNTd/XJA/u6Ju2TB8Yozbh29OeAIhASLpLHRJhus2xvdJtHhcv5GDrJv6aBR
TPA6xXN7vJii0L4cewxSoKqits3gvvDMwrQ7mNU9TSiSBrNHJcz8GNHIimdUhmuQJ33SMnvgGFdu
jB957bC71e0zNpnRIpjd5c5UqMh/ut6FKpNEfCFOyU0Gw9hV0XZNLClUWUezFYnF4iRYYYa7SfsB
pGWq7VshHsXSUBzJ1nNHVPwKbfUwjNwzWi/KVvGQZGmKt1YFOMOdcIjnQ1/T1BD6hsIlaJGNL12O
+8RakYbvjbr0nrDMxGPiKKk3ZfE0MrAXxHgqe+2jh94lD/v3WOWKSlVbYF3o7hreQ7Acw/WhXNR8
J9rLqBY1bQPsEd1fYtD3gthHtHTRHbq5klYaJRt0uMTSQguA6dQVIaU48+XCJ+Pclsh6bVyzx7xt
DS8TuzbOpT4Tmk2DersQ08yl53xq8CKZpts0i+HUIwnF4V5icJE01ZvCxWSyaLhXqOrcSSJflgSW
e4zoU4NMIrLUpGLvONswnq0gExVffMgxuYiwfyPOasdbXKiaU0YjRoAMM0tqKNq5WcBfs8ZsT95D
TILdZbvSlTLZ5RPO0d8wDaWM0bPevAmm2DWp1VaRpLEyB/pGh6XXRC6ZUkiJN1xfVGpNstNRTP1U
zJcjVaE5ayzHYTTJ7578yRiTSeLKcdsBD7eB8/T5YwQwyfvL+C1lbfGnmuE3Hc/dBykv5Qu0huw6
OiwsbSwHFKAVqBuBHy8YbR/0xjYXg39Y7+PxeJO0vqrADo7l0dEdm5YliUgGcahgYfb13k7sbl33
YJM4/YafEIK8rJLNSHllog+42dIdjRbWUG7aTdOyWH2FRAMNEX7X0rrnsGkB04NO1Sx4cAO4donK
fwk1YKIZ8GGmpA5LIrpBZBExZiLtZAWjMqnG6T2XwyuczdNRpl5ZqxY4F79h1juZx99WCJG7+llH
n7uvLrDxYbas4N6pSK/s711D6tFeK6KUrXLTfmRBZqPwx+BzcDcVDKvmwjY1sg/8oN2598lrbeHY
iGhSP8qTT1CycMm2R4gYvllstsPzvmdX01dEjp0a4d6egZ9zoMWh+ihMfrxw00VMKqpIn7E4vJ20
P/8YD9jWvGGTabKBjaION7+IQs3FjBw7OT0h8itkkPkUvGK/YpEHAs7rLhhHPAn82l3AWPGtzpgR
XEee92tgLNRyRV2SsOv/j9WuTkucKKBVwJBf1z+uHOaptR1vAJLMIZ4p0tAUOADCZywOsbZ9oIn/
TfTSRWc6BxPt0PA0afeBFVPmEjbWICZ7okZdiD7aywpoTFbvjKJejCureZjUPhJsUwJxAQb1YzO8
DAkDl3PdBwirtL5sAHj4BKTmX2lN40PB28TwbjkH/JzBWgWHyR91OR8wriFHnLxN2VRd+lScj4kI
OLJ30yno5aClNK3G/XQ9eLTtxd9bVaBj8r6Sqz5qhXedccsf/CeyoXRSCf/7UEfb3bSktAw/VDuA
X1foQyz1Vapx4dA19R7W2QJ+XFKVe+/WQleYWA6rwY7QdYZEncCbHkwJqbvZ3iozfOcbLGC7U1fD
8nmRRmpTWc+kXMpsy/7lqmicV1jmJ1pOmdSbMUZQ8y0ais1Vq3Ay3jFoZHcGbwHTXoqA9ry3bqS/
jO44lJVKEgJJjt0WZGYVjv9OFtLgmbDyRx8Yh/OLKC56ddfEsCOInvLiY/TooFikBdglHie0UGKt
t9qHmjzk/uvpy14I7TYQHJdDMf23rMDbTiZWQ+46tZncuYhO/sZgIkgA2nmm0QWfY5MfVAbxT0KG
HCvapisc/NzDH1ASNbBBsayVAzCK9mxkaBgWD/gwH6jk8H+zGN6SrL9ou8Ry1OJ3NhcBMW1PP5fN
UhY6pCvhXh7z2idfD5ve+zZU7NdBKHhsp4vd/GPqKnbOfi1l9IV944rpA8bGI1PR2tXr8c08nGIg
mM+zFoHFuRRsWjJnfq/jELZhOjHJVdDRR6k+vlrhkSRAEwTGOSUeqf4HK2zkfKLkLVlpYuZFt2hT
fIJF39UfWVywE8836FDVIbWOcgkwM8l/aRr5sUyQWhm5Yc0bxgw4/9wIISrp86s8XIss+g9Su+Qz
FDa9Ue4ts6VpI2UZQ7c2wzCtqMf1eA4cpT8sT7vfkifjwR5TYwKyJDGxRrYsMLgob9AArlAD5WRY
V9TTj6FURiKxcHB7JjIDMpPFAV4GYKpkKC/AwfexqBELtRWkd35HfB24l1fzlbHhtZTsUtcdhTRU
w3E+sq3iB+sDBLA0H4f6YuXdKmxsanE+KdAnG0pIhQo65jA2VxqgeGl4Eoom8ScC1E8NP970i5b6
GJQVDsqcw47YQAB9dppFACGrCWc8O7Ipy+GpWAdR8O/9SV9o1pujdxisIdaRn+GifI0o3fJpuUgC
QLYeYri8m3l1vtVUlOGl0DjmE9XM8tPP9Q32/bVi4CUnflWaZdheDuAf3POELAhlOnRF+l4opBAe
uJRB1b/sJO3qQJtHmf6hwWH7ImatpwnpYgmdj+FY7oUh5F9GZBlzrJqXjn40lrCGB+G4RLo7sojR
maea+9i1cric8rDRHIostyKsExThJTCW0vuDtaQOH3SKcsf6Bppca5Szi1Y7feXrDFky5QU4dl8N
WHX1jLRYs1pwhedDGBioxSw4JjaZx/B4s2AinnOS3KECRInnjrVU9vsGmsbz7FDHrDaa6Rmiv+RR
THkg+u1ZZgtAGRw9wJUP0EFfBaMIYv7F4VW1wInB4vdLSZF1xoz84wdEc+Ntp8s8Itte4h/Z49sW
T9ndYNgCsWtT1Q7cIXURVVusmCQnQd26zQMrmBum9EhMmwlDFcpsb5JEVB9hyQ9YtsdEsxwDs+tA
GYtcgK+k6rBu4uPOWABK0rXY7LHAuDGyHfWiXOzG+MuegEoUilkBTv1xzIsyow62M91HfLYV8n7y
bnn6xLZJwnjmm+My0Tl8z6O8Q3hxlpTdKReeWCNIebbYtz+erZ62XO7x5F0O1DX2xUdyo/A9Qftz
k7q0pE3i3tmaWtFk4/jmiNAfjo8sVr2eS2r+wkE8uOIgQepR5/UvCZzmppmKpzZ7Cu5QrZln/LJW
TxEvF+fC69rFzoZGYKIiesXQUfOXmqhE7XninfXes167TLtKcR/n01tP2CLrbL/ieDZ8AZonymZL
CRvzo1+pXjR/an6l0ZB95Thpw9PtTxQWOKHC1DsHMI2p9TgntpANs4O3jLF7dsZ0jZ5CLbr26iIa
2ADPMBKIbqBmgd2YZlpPwA3BCaL8Jya/rYnH1D30Q4vmogwPgIwYYpykyt7Vv4P0Yw0BVAmC0goC
TZ9QWpj87FY/D3nLEYZqalzyOAax9kC/ARVcAqMUPg0CCQOwfSCnRRBi4ZS7Sv/yqnOS5REvPIkz
LlapSct8Hqxd8bQeo0L0Q3MCshzgW88hNhsHz34Fc6yDBQ011WwnE40irzv8zaUZNqUd5bQEYpf1
/JIT6FSf824dPmDDsFswnGdlG64uP/zvEkO/TaBt7SyQk3SUADxHjqqXjniRvsnl983k2lQ+fBEg
dzl5mAcSr9RfLdUtJZKPrBWl461TA+sXuw4U1xySF4T22mtT0Vu9d1MuDdCjZ8jEEOg27shcyEFx
ohSdiptj9YysMapDD7amaIrUP0DGtNn3JVZKyOFCYL5g0GbNtz8yDBfpvWvWNiART3CpgPleWQ8S
oC6D3IHfPzAGjh4bg1ob4faqpGtd0oa7wgmHT/111sSxhj9lk0ENfEXuz0qR0X9bN4arzvyzY+YZ
lOaZUYiwkCwR2RT1J+KgcPY9zSH2mLdMfD2eFPU2t/AzPXoEFi7WKgEhtj/P7f5yqCyeZ6tClILx
xRu5BgH9SL3UEA4pDQ71sYZu9zok+QVKAHVPIai7FXv55AAvlbtW2hGqhx/+2mhW0lnngI12c3JB
K8+hSEXcgGu6GX8ZC5pFsK94xWBdjyUGFbUdQtAhIP1UF2PlHMYe0OGSzx1YT8MNtZKwFFbGa8ke
rGgnMxcguBaFwyutz52wM4+sDeH++dth4Rbk0UUdNOvhBxum8LeBdfbUMNfNN5sPGTU+g5ulsKAf
rUQdkPbKlU+QOn/A7UE49DOq276AeAfPw95CJ/h7cdFI3zHS6jKfwdmWsbgKsAJ1p1j1LcjsilTj
USUA3BgoRc7AJpM9KhkqzCglxHv8dcZLFI11gDPJlBq0wP3DrgmDOaDh8XuBVCkNflLq+pHJltpS
y9+BsIKEhwXwVF6+7rGLK6+8um6Lh9D8ziMwASW1cL6gpnN7qB6OZZSJIQhINqclPQpEgJKbef65
yjshPfKF6E7AOiYq+vIwosPJw+kC4Gxpd/Awgrn2RH6DDOVvlvc2n3Hzg0cEBplISx4L1fTe7+sG
EYJ/xf/tdg5wq3AdSuU7gadmNVI1Nzk9Aa0SoSy27QcojwydI8emnc4G2w+UeEN+I1sCl+qbsJxl
6GYizXfi1rDY+B3YQN2yim3OLIzFfifnJi+TzTv2W6Mp90SMzwak3phGVBv6QWx9WCLV5LEGGLw4
64OPZNiole17UWbP4p3pILSHFVIeQ1EalBEtm1gc12WrAnFN9hJrP7hKfgrO6lUsGXmlgJrAXXuc
LKMrouOwMIbNH2TmyPW49OVFwYSS3DM00LpUPitXqfztUk9r/BVky0yK+bEKGetz/p7cIPDHL0p2
KLR03KhWoiQbLzZKZn3oG5y/aYdc/P8J8dyxnljLo4+7cS6+DgiBCoRcI60WoChxGQtapnwEr7UW
fAOatcleI6/M5JSaezzNa/AfMOAxVVIN9/UK8cecKGYAiOOAMW6q2Pzw4iBX6WV31MmQ4Np6aT0p
2Cas//p+Su3TNYbMAel3HLGzmSNGOzXYvoZ9+BG1ZHq+GtUlYf8HbhtC2ZTkEKG7Y+LqG/jySe2c
ZFJOI/czkI9XLMikxrIUoOQTmp8vz6mZMz075dCB3hXtm4wfy+RH5dNF1tjNjY1olrDEkHVnXQN4
z71ZD1n2iK7k25d59MEvuwDI6RRBCFsD+kQuDLggeqmbczpHXD7tcbY6OFzFslN0Bl1xbGaD6mtP
QiUtWym+M3Z17uRsiftVIanoRSbTGuuTg3fQDIXB/RprHNTYPKS6QQ7eUKrCkqy01oRndtu65jpO
UjvnvSM2ZWH0GoCNFSVP4bwtUi0u3snWbO80ziJcGwAVuyLUM+kXoiTL2Y2UIKnTMzqSpVB5kir9
Hx62Kf/ruqkfh/HNRAJ0VKbXYPWd4Si2w1MQX2NJ7NV5R2OMeNSVHYumwWrilQP4iaiqmEeu2FUq
fwM1HNVpTM/uTJK47K+EJZrcut3LSD+1k0xZSSFhLZmng0pFmpdiiJ+6fGYnCBI9RDhtUbBa4Qxx
ni6bJ05+n+m94V074HQ2Xc7a4LCMQ2INwxU+RcZUfGjDLsw6htovfvJeA581bH+5d6JHzzMDKG44
Vm903nvzndhS4VgfINAy8/0A2R2TK2asRN92f6b26uqVIGSLgSaiPWEribIXxug0tEnziiZ2dbQ/
w2CD9Yo3b8K2bmFCfxe3Lf2CDihoFZt8RUcLKJLwOm77sjCTvwlTk+eTfeucfLRuMwI61BrF2+CN
9yIPjS9Hdu4XRyENkV8ClDDVqxAqfjdDaIrGU2sD0ZaEI4tzIGDdH/Uetnp15cxdaWmDL9CDbUct
8Pq+OQYZ0KSo/NtEgpjqRporn8MR496ZaQDPOfkn/F/rJI8x0qjB0EoNyurCaOF1Wt83LCAQSFQW
OcC9fFtoc2Ue09DV40x7TH+PVV6r0JfvXbQzoeETbbF/xkTrTqJTakoR+rWc7ILIq5eaLfayXE0F
H7zgpAWCKKyi2Xkpf8aHJYKTDdzcxNsbMjxx/I4CINN+aB9jlEYyQniVLdCjwMJ9r/wlVVvw2kEo
A6k13RNGCy90dB6OT3akQEgky7UksBINdMu3JdutL/x+85fXYbMvXQ7vKLekgRvaxFqHl/0orvxa
+2jerEGgWwxyjpCRDm4CGTrl2AI/tMkVB9FQ02X9GQG8vrOW3bM2bPI7cgR2imnKDXxAzD0bT632
ITTznjipxCceK/qLTRWZuwTd10sUHqf6nrD8DD9ziral8rtyr7CrbUiID49iFcXHUD/qBRyHZzxi
FXzmkWHNfDCI9EFefbd3cW+s/N2zOZepQe8v1RCPZ3a0+GjXraZ+uJTBxvD2WLMzWicAFkc8/Wbu
IwwbU5WBLl9yGtrR8Zwn2L/dZoiRtj5SUfVrNM7z+Ig7rP2nYF2OC1D8MPMVOuyIlySR76QSipOq
oRofVKv7IOnTTlMyKeRzsQDp1zQkqiFQnGEN8pomD6qbE9lPQRDJwwpotJZDua58qTwkpDtq7BGY
RBJoWaCyS/WdkR1yCd1xQpU30ljGYvUhcfqnwdvI2lGU3cH2u9P1d9tpm76KoGgC1CKWxNAwVACt
TlC2TiV7er8HY+SiNelf6i6h526Uf2BbC7GRjYawWg6vEBChX3pzfPtPdR5vEAnDPY1hyzGJQCda
zEa+FLjNJaHJsdxlNZp0XMT6oSiTTIheA2VFUQxjgNXU3ro47qgytFrfY9p5PKaCO7N0IEdtlpJX
dN1CI9hzQ6C5LWVTVRyZ8hdcdQ3rkUrsnD+aAt7fTI1nHIOpJT6aHzH+urOv/jHHTY8FCG2h4Vg0
HZp7vQ0snzdAp/FGc7CaH+yyWr2MwsH6zADcQvi2ZSjvQQroTzmCm9IGWxNtiqnsssxas6V2JEvu
TrqccZlpYjWfM9gYOZm1+1C2SppcmJk5GpugI33ZR7KIMsdUGCyeik3crVzjoTujYqSOlYy2X0nO
HyFWT44QtdykNQcGGC2U9fwbzkSc/TbQiqtb0kbEKPu506F8KgrOYiGAiKyQAKuCSYpSOdt7mAB5
v4GKcq89kv4ircvwmEkSMpKuvhQGS0JuPLVF7O6W0xdQrLNkQO61VWTkH/myX/UcE00A6szny+7F
/1kRUPf/uU08edjTgiE6xJ/6jJPgAmqNV9NDJKWkWgu3hFWV6TpL+BvFMoLPn3/MonbRxYquqICt
4zmQqisLEcihGstVgPMR216B7E4Zr2uVQK2Hc1wty0jKyN8SgKvT4W/7qfEEvkiNSGgEKF1gVg33
/eA0Shk2+Fgk6crrx2TDVV9nJViKpUYdbtEUU+XAKRe5ks9HZeK0AyCygeKOuR5Oz5KMyyS1uBxk
RBqMpShyXvcQo1IQ+uOmrI4HE2lCtk10bt//G+R5m3eTa+jXxkgLJO6/d3NdwkB/IB0GdzNjyfhN
XZbATXJZQyf8vbpFck35z42sK8sG4QS8LNUKkqDFV0sqkYmubtoSVwT94ez0XK3LMKMUEbcudVRC
/cqjpNSeWHgfLGWXpGOYjb4q0rIlyo9/szSKYZMgwyfDpemFmJq2swnGEQTC7vUoEB4d2RRbkW+w
5QoLLGYIVeBkDd5HDG+ameNMHzuBxK2QGzCZKAEoqJP0l8JjQVI8JUNplx9qCUattrC1dGn3ON40
QmaJhyd0VpUiWCV4qL39vCw5oxNRPL2gORdLjjZXEWp9B8HlBOLoksHT8oEx1pt9UFjeZmZBJAgo
IvPhc7xX/mQWF2l6PgIB5/y75sA54ShQm48VC6p2j87oSiwTnwQzSbJ83KlYHrmb+K2nzGambFZs
GlZuK6PNkhLepYqT+aKcd2oV6MkkbRHYKaWc4pGIISKyrdmhJC0/JsDpGiodf2OQnydOGzaTJXLN
SevYLmIo3ZuEZulTgWRNRUqs201VIN+FPxvIcdmXjW77xd3GMLQVOYBqNmqvPRRxuunRPdGnmMqM
W1lyE88vcILZkMj4C3eszVKGavf1lhFRTIfIcrAU0JNs5k3ZnHSia5RW7RQ2QDq5pxN6xB0h7lHP
O3+bPHRsw+Qbc8HKu7DOZH3fmEHcVGbopFyiZtkM4uvB0MId1iyiVW6/2XLPkHk2RArftck4IW14
QzRDTIymUf3RWbMUXdXTD9WlbFq4IbOE9fXL1yTvVTBvrg93jSXWrdSuCPJkKdWu2e41mFJj9HgU
JjN6vSrwsRRkNnVuFwhuqJwZkhA4yACJ8g0JoOmpN7CpappNQzCclq7cLjrHuRoWQNs/aeCnvIHa
iLIEWMuIDhQrVKTDkwE8VQunOMg/kgK/oJwkhH0X11Czjyivmtw+RGD+hb2MANc2vPbAXEXtFHDm
fNqcdWKDvJ5fvG3oBsJaadfIDyo1VxtGtW03AMfrGakqU2wthHOsdz01YiOl+agr/8pXqYFGZH6v
m1gxgF1TRNUBqakij4/xqrSGR8P6CVs8e5aqrh06sCIZPjOldZqmyeARCx/bez+jKk9xaPPRSM9C
1Xh5JEwYBxARX9Xo982Nv2EtUWdziBJhfJ+sytxmt89SwGkwWZauQOw5vOwH1Nd3hjRPH4V8JUO5
kWt6j/LEud8nlnA8HTaxy9mxiymKTT/Zg6O7HStPO9gYBDEcUETXcPCjYooTAXBS+lCzjKDxGiM7
zKuBgz7jDekesXuDSqPV1bevMcAgVJLJoFoy0ufwnSYInuhk1KSdD5rzbySXw5Cljmb4OiVkijRx
c9I0Q6SG9izj01rWk6IBzjAe3QqRUBjJXCl30gu13fQKL+zlkprvBu7lNy89uvi9wFcHITyhsNAm
sFB8qAHUB84D0tal+PQxwrW6PsD2VTeV9FDxCj2pkWnpKfVvSza7vDLLINvOyqrHuCKGRo9ZguOW
eojtc36gAGMyeAHl7YCAuo4HcrxByZgYVQGAVuOHzYXYoEjWeoz8zRt6TF4lrZ4UcMusLbIvRVg2
tWg55gptGFaByOJ4H8ADPI6LOrcqFZIf6ZEg9eWLXGeX63HOIEhSgAhyYt/30rwMjjQNx8Us9sy6
pnK9YrbdXYRfdPciSsrlXrj1mAEwlYiJ68h709k7LhtA/x+i5l+0EpkxmCrfCt6Y6nW7sI7BGyCR
UmcuGIFsMneAycg/s1W2aCGZs1tS25Y98ZaMMNNXjCS8pz31MAhCrT/cGkFLU9v9D0UF74JyCl8r
lucNEqmZtP7IpfZH+HKGsFM4TN0C8idc1qdet6OnUlojfAie7hrzgE/pWQ5hU7E/XfsgnLrvBcfJ
WDPRSpHNlvGGmrTE6OO2iMh64N27EL07cB5dQWX2dZbrOVskJrhB75OPDUuABVw61/6Esbic2y36
qxea/eNB8BWVweh6pZ8kqU6YA8vxLqt7xgzAYtxEnnbfobOKAjsznGMAs8b+nZ8G5Y5IUCVobK1K
hFo05+OY0i0/oB/XFLaIwmgaW10TbiMigMs6SCXHt7vqx5OWs2oCloPKDgHmG3aomTQkvNMypeGr
C7hHR+C1IrNnEAq6KNYFWLbf6sXahgr7FjDo4khnaCQKbnOtr32ruvEp2QSlzPIJzM6MX51bTOBz
MC9myh1XHjgC405djl1J3vv6kg5doeISnObUFCwkp6gmPsVcyYH+1ac7Ck8ZKAhwRYUgEuknJ9Bq
XqHZwDbMLh0lVfESVx24a+BFjLZr5pQjvzgouV6I2d6udBacDus998O913ExiaRUFTX33d9iD7Rl
GBudwUEXO4CtSCY0L9xEdyr2Lt3uK3yvqROJ6LsekybLHKPOgVui5nInpCPAmYgACZogSS23twMp
wiyLMvOO3CDrI+L2XKdANoGOQuOKBywxwA3yLoXj3lTCAoasjIEmmQXQ1eAOSEWgjjewKwZwohvI
ciY0VpSoBRQvpgPkMJWh+zFMydKR6ip59yr/ZMOyfriWGDw8t7cVkEGh1KLAyRJesOyIetaA6El9
2toiv5BSRhkfgxKqcdIEKVOrlRYXuvg5vDyIws0W1Ar7LUhIe480qGkkn0f6PVT3AxTR9mucT+ra
UmS/IHii7oyG2ImqcbC+xSEbDrX+hsFd7Rg16Im3jKcumAOz2WYADBbbBhjkBKByZ4B2JfQ5wAWT
YkWPJXWajyERZnJiNkg4qlHcv5dvbrNA+sMENNw3nrVteplfphLVxXRoBhfsh1Au5DvgydtrYNsW
38FzJifUrWDVn5K3rFv1dBM6DEQIWBX3lKxM02uKaME1Yh/SI/eIUwtAWDBJbB5qjCrULLObi8B6
3SRwvk/kwJiMXprL3gF90baaw5vOs2lnAnvTPamQnre1PPYoPHG+QsvJQJs7xtahW5bk5AL3FIgJ
f8PS+PoS/EQbDfbp9DYE0WT7PH6rZr4VSQFB87pkox3LRAzqreIomjkf0OzsWz7zUb8QxzhChLXF
jPtPp62toxEWWW01Bp1g2184D9U6cg8PWygvP4viXwfdhf7xoT3N3NGa6ySj6Y1wxguKXdSvOcIb
IHAIbkfKOoEiTrLBZxY7V3rx/ctqOzbz9F7F+ppG/GL6w2jw9iQ02OZb9NvrMCkLjeRURkbUGT5Z
8MUNeM5uUWPGmN0VShsSdDjLZKcxDrPjF0Eq9G3PzYUUeMsXOSbQIlGYt6js0iprJcwQWD9trQXL
nHyCIO3izFsNgnCQCYXeio/JFtmDvOLBWSTEDBIAZNruDbYJGKoZg8LwW+bGT+TEK2B1wVk3eNCh
cUJ3359hZsoJc4F7qnjEb9YnJza7Qox/aqGkK4nSOMubECU+EJupIxKZNihlsTRc/zR/j+tk9T23
EqGtrkSkIy94Qiv6XBSdQIMe61Qr3g5YTrVLuEbgatxMHU494rutwk2p/eG4HRx9CW5BFdk1YNlf
I2jSQ8f/2QklUu7DiJC0YRFA9d1hCjnbOpys3xLC/bACU92aCAsWs6a4Zva9kcO0IPntIiGGjpsI
qUNpB3dQ7U7nZkDthakHwmNuMso1rm3G9vBmINoJM2PhRQGNr1MW1/qTjo74NAMdtXxcn3qEJ8rX
P5Uz/BQIIXYHINLuA/VqGE6J5omyOSq9epZt+4IKIAXTQIfjBWJ4AwJXDuMsh4SJIXD3E6x1B/FQ
7HYvjI+kHyPfhnTzg4aS/XpsmZqW5SnHvFB8Jk/dJ2SYM1WE7/TKZmLY5jV41Oa1I+D9xmoXT00H
SBio36F1gsWw/oeDirzlucroyJwClMLpXyao5u1EWoReWSfCiyYLomJJ0G0lwkb7rycmQui72fwf
7PtGcx+U/i8Kv5srpkyN4CcSFLPLMMZ1368YP3KdFx2E0LfySsvbvIGfJP1FufG2o4kGEHL1emym
SFCbEP2huPIJDKUomncyzYGMWO2b4LmeGQnhhZXOKxS21Il2dVhwXc3Bcq3Dodg7R2q7Jfrss5W9
UXN2vRaVnLfBHp6piJlDjjrH+Gc2ojywWjT2lYn+XhV9DrQ5ejBRRT8snhWUygwDX11h5tR40Jak
/Z+xNTnx2pKDjs4/9n2ml/afmLkSxUnsSjzFQEhilIhzfgqDJ4Yndd2DX5mAGMz3ys8LIKsDqr0N
NWgyD2hpENuZw3u4vG7Xdoc1oKkTkub10k+LdH8N/CP8OvaPAbJ6QAfS2kvcjvw2hxRV4tjEwL+I
QckgdS+2PqkZghwcrs2vX7utkDblg3TzckuhvzwSjEtAwdLQFqLcN3f3vsiJGjEjB2LcDnZWl/Nd
M/bvst9bD377Wc8Pc8f/6Hfn/zkQhg4g409+YeKoBfDeTG/9tuiJovcRqCuCjn0lPbnVIjeVbKF7
dTaj1GXzBulqwnW6bH/KWe8kVHUexLtXjBzKwrkDSE2XfBUY3DwJitU0jB+rGPKBrEdtHI8BV0Of
Majeh7xGPZIOBDC7CpjbS4r9BssWr89tljrrImUSYc2SCBdwAEj5C7JgdUlQrqjDRTQDPAuzMCQm
Jb+UBmcQB2d7k+i8GgBWgUB8OHx9S26O5jhn96PNq00ALs8guk7fqP6oqmCH3F0GEfhZBD/wm4D7
Sslf5QnWtk7aO5KRVJtgMM+uHGb0QR+unnqkNev+hLJ8YEtdJxu73kSOFjolFv2JzuOj84MriPNU
vfLFCyCMQFQf1NOH8JviBSh9Up0rr16ECl37UgjIB/9yRmpI8R8TXdkyELzWktU+LW3CCJ3XQTKU
qG6AxtLhqUVPBAg8K4BjgQnj8aNFvt98IANN+yZvLUfEXmvI/zgvrGt7JSTftOQV6dVCQg8lYluj
AQtIC302x0sgKcIRT9elPTHfUJVHmIcnNFm/yu4Lp5PPHm57mcIvv9/mjJpBAiiN9FiYiksE7DC9
gJBNoQy9Pl939SVCFZDCTg3pg61bkVTQtKaMWgj+c5hUgdOY1S4Upd2vFf5CX5pmyYN3sxEw77pm
L2rHCifHAIR2OXVcaamHF/a0IjYmjsBOZBkspUa8kLDtmkY+EnxmjvfkP/FIlorb5YMUs7rjSj6K
H6/MHe4fGmZKBftQMT/h8alh9uFX1q7yZl4h58iFIsPwWnZU2VbYYyKading7QcnoqINvrL8VsrZ
uFSCrz+fMhss0rJg6MExai4j+/v3VzE4L3f02PasHb6ECI0l/nvThNJ0qWkSCoQjeE6svZ9dh5Ci
rCY+BVzfWbNKBC5s+nQ3EICHqzVuh7Mz7JgeK6BnXO3WOdWfznhqce2k7IV5rZQw43Nj4ej38sAS
KKhNRgt1DSJSQe0DaLBGhdRSEgSycy48tLVIf8ahUf876cyfGVDljaSnfCuA1UaWnkZq/odL+ygG
q7kRKEdD4Xgjmc0PNWDiePlUcYDr9b1slD270WTRj10D383AyWv2aeqKGs/5TOz9D3Yd2TAofrv7
wB7NgpXWsFKoaeBfGSKVyN7G/C5Cq4G2XuDv7+qfeRQpnVTxpknjZfKVLUxdypnRm7BJ8VObv4S3
hmH78qMBBwZNm1X+iXdYGGx5THCqZPTdAZXVNH+1j5xRGZ5MtU9qBJoiwf6posv+tE9eZIkaWylE
Fg1P1efuPkdgOAIZ6k50lV4REYoogKVBDpdW0J7dB+yhMUwJAk2HDZEtv5PqTKHAmVYEYOYXqxa3
6K112GddjAvrCLL7v5kqthfzOTyhXA/M94Y6xkim3zsK1zPE7yDWk42bpLn+7vbkrvmsXIGAYssw
m1mDBrvlFhcyG428bH+J9s/ejxfy96xKuXDXhPin0uGZDV2UfR2hzeBK4y/t9mSiSwXH3UNr90l0
V4JGUiROz6YjMMHKgYKtoHM3pomOdDMVIhuBKe8M31LSemEn8Ri+wo1GKlZCHKNQBGqafxjR8zrN
DajY12hkRKWN2FL2ay6OIq/dQUUON4qJdT8mLxBeYvjEyjr0+aG53rysMgP57gqXumrSvB7E91Hb
aJTZjSKt3GVhOOZNVVpJ7O9lwczdzDDyNHfBv1oeL9/aYTTu3tNR+jfqHCYOB6kPVjA6qJ9dwNT4
lEYF3nkNTa3wlFQcio42L+FnAO6mAvs9pDP/dYSf1Hhi2jO2Tt+aqHBz633eigUgk4EmBW+GKqpi
WKstdNlKl7c/xpMOy77aydIQ/vEZKVtSB/O4So5/JOgUijW4IA1ZtyJgBl2CyUrD1v+1TFyn42Q0
QmowoLd1tP9eX88Skjltoi4XN5sjJsC2TpbDd4D45Mtg34K0iHnaJfC2MlGgucUzFuT0B49t15DB
u798gEhYeiNFHHTdrfpQPEVclnOD3A3WNR7as5nU3LQOypDfPYl8jEq7YJaQL+J5Yvry28K5Gkx2
EiOQFfOtW9qorwQikeLhYcvTJ4dtSDJP5YoHsVficaPmrAfjE9b8kEe3wIxuuo6QY+9zYvQjHDjb
ABezv/TqaWEJzQCI7Wyn4pYi7eS7XmAqz57dnYeraEPTqgDT5dXGRu/S72AllhDy6lXpiDZhwaoD
zNtl4tIlJjjCeN1SyiKDpIYQ+2NgvWsCpsAQbk8XvTJxPpw4KW9zxXZoM24Tfd3lEBYIny0L+zhJ
JHHWaa7CP3PAbZgwgU6UfNKH7K0k0FuRTDHxRJcqoeHg3eXzwxp59hjCvNa7/Qbt2TERJqxtnG1C
hLcSah6cagry+8T1JeuPJrTDcD0sTDiLxi6ISBnWxxILNzEHRfHm0eYR60q1CokeWSxSdLgjwkBO
2GpNGSl0B1qTEBW5vzx1vazLo/zaCkcYVwQV8tPlb5qKH2rb9QUXtb4O4QIxBG5t71MUiFZmDori
iIzZ+gPP53yy6/FhjAlIu6X9Z8Unvp+is6uJpdsq/3mW1L3ur+rpip8i1lpHK38I22lheeG3qX9+
QKNFEZNdNvSZ1tzyacgq+ku6CK4yMz8EOL29kK9Du4376mVDotg3b5Gq61v7GHmXPU5DOuCabaAD
cHtEGgF9nGUJ0JndTlf2JwU2vDZrAS0V8JAm+PWKU1+MXY3Lr61bsx4gHLuJPUFrNFEIWIFMHnhR
1NwjumeEQVW5NDvWsd17l7iZWHEdsnR7C3ekCz6q5RfAO5ie+Lo0KUrJH0h87hBCGthh5A/lJ4ia
h5QXdyNQSMtPC2+IWieOYf4rq+lkRSo8E2zaw6Nt6KXR7s/S8WyDuRzj3FEXBRni3hbxHmkhQQZk
BqqGoALBHdaD1fsOhN3FIhSKxrnBhD1tpRMGGrh51xhW+D2PHjx/O6UC+1KcikycKgC74NyYtkLG
Rn9CPaNkes3Ebi3UliwtJeiEpEDSwfnqUDj39sE6MPuJ4NVmGjyyjfeAc26CpUbjoF4g/Vy8VD+5
jqbO2MSjGKDRlcQ2/DVMMoLmGFU7BcfOCZ00U3rC/DPkxXVUxAgh3nWVf/VCgo5wPP8G3dOTTqF/
/XnHwsQfEW07+UarNsIZd97333OE4VdWb3WaxTrdshkz0G5VK4ZT+0MdTmFDhlL2lNeGxRL72OS3
BYqyit4SHWLBZTGaWvaXSwdzyKHwNJjIlbhWS2DlabLq2B+oZhJgjJpuXOF+UkV2qltn15aVlJil
F954a+M9MKTu6JBn2M7YUVlSgP1W2imZmz4BjVMeJ6e1AR+Ipv5FSq2au42mNnW6qBUBOuHTyWwc
yMd64BXOi8mH3oWD2Dh3LMQ5+FnIoq8+VgL20DxzWUlcN+m6KXxPI5UCvewfdKL9ptAYdhKTK5Gu
0GYK5Z4G4jRirHlkBytytX2taI8phVksxF8P3+UepS9zsstlr7s/uCIB7qORa4zbkWB0NgEfnAuN
HC0nnKBSM+97qWcgDUlFsn2YPNonYu0c+OIyBdwBT2w5JFSSLcWDsnCb8Pzb+tBouRTWuBiNkJIq
d8LCbMHuV1ad1c8QYJ5PjVi2QETkbNaMoLq6E7On1T+RvqnLenvFNp6iuLc1FYLWM5Ndq24i4bQ2
kiBVqYgU8PJ6WMR+jHQqYaawW00XBzRQMJeTvxNfSQ8QtMaT4g4a0uMrT8gqsHSZZPyEmvfUuBpk
BaqkT7/xG8QBuLZ2UOdyAdkDdd+jWusnWG2yBtB+LRKP3k/mAbBbfW6Tyqew9sxgwKjAEc3f1ksu
4ybov8gMG1Yp2jbBEYC+Lpxz5s1SF604r17qiaHNf6ks6E4XowIGq0dELHwedZkjgHi/9hKdO1pX
VWBfyRysygVXuACwEgeTa3KCfIBETFFdqklz7EBPiQCX5XNntIxZKsSYz9EyknWJS0AEQEzGnGrf
rVfCC6KORJ8zEpAPmAVxwtk2lFBLfJCpmyGRDPinbT8BInRQT927GPHeVS5wgi5bnqdCCH8I9i3Q
iJS2B38deWAZzC6VPHFtili+us0P2TEmJ8pk7eK41Nh0gyJ20Vk4T76GBnqCS8q9AKgB5fNeLwFo
/o8a0BFDUAtlJjLN7EbRgcCfOkHzEQs+dy3/2ijOGc/ddQTyHxqsqgxwN9lImju9FfLFa5QUZobo
Rrvw0Qb3fyD80bUIoLTsap1l0CEDpnvSc7Lywd60vdcu3kLQDF9Hl2KL/FT0SNXRqjY9b/AYjwyo
ykEqNUkEIhlh96BDWdIVi8XbOcafsQlmxzK2FUq5Vh3NTlnCP3XbhLBxcL2/HhmK2ZUfM17J7o5S
0gS8Nru94fz0DYthZZ6x9C35dX/y3DtgwKGY8vePj+3Ic4EPzoG0sHdXgTLSk4+Q3wzWgoIyDksQ
DsGnXmzAgP2T7cHEsxiu5uf9KSIw7Pl3kHtJ+Tbxt33hQ/tz6jq+HiGKdc5UahCR9epLBh8+w77W
EtyLzBvya1zEKdISAhCLwYZLZ3rHhdLCkDgUHU2WDkm82c43v+FxE2taD4gjB+8Xb5JyPtP1FsG0
HYGyxH+gb4FtvXvVD8ZNNxc6EYBNvRuv5q33p7tqHBbkaVRirRlib3OzsqZMtVaKGyubP9+MXi+o
3v7VrLKmZ7iPy4dfaSe9e/DzvVWzXUGg/slhQGyhVuD9+lNuhlbL4HO7p0XO16DpDZAWpjtvUuOk
nqEF+2OV0V6PuvqADSn3E1m3kR2EB/dpWVQYCH3U8dX4PCYEh5ccqkH2oEy3AVDOdwLzps1SlXFX
ADyKszDxJWcFCB/uer4RaqdSAwInCr+sr2m8Hxr8aGgNAQUqdZI9YLYM4ptZsbrRkaV38+ONtHLJ
3NmnjWDxYgA6I0PIqwVIX/YStb2iKUnmkJ80GNwoYczB6CIBYIhIVxK68w/iWskxf9WeCLx0rxEe
E8rU4CLjbW96+rT2b8rm1u47JHgfyY9NMRW4hoqrHRyEjf+pD3a76r00vSM+lIAlI4KMq/EF7d9/
G5yeQqypyiK0iOJ9HqMBAZ3G8Sl9/nnAXGHC7EdOg7vtqjXkUcHOJrNbHPRwF6FLm111RfG7Mu8B
tzNw2Q68RT3aLFDOQHsGUNC/X+gjycXuz83PpWX1vhIvGgURmvQK6QMiCiDt2QkRNyPcuZejJXx9
/g4B4M5i2cZk6FZcyc6DQYXC08mAWOF1cwGpWAjkC79LaoF+l5O0yYPA77c7Drk/miQEOFdVhiEG
O4BMR7GzcPohMbB6qNlrp3r7m1cYsJfaNffX2soN51sF5GhbCdjibIeY+Xw7UIy8nmYp8ffGZD5T
646CH6Yg4GpgLnGqV8hZr5enhKI1BA1o96GDNIjLwnRQdX2nuMCETa8gq54cPamntKCkT3SgZJUN
4SufSlAIExfsL4HgwC6+gLhlCddqsw0sauXT/3W+FXfQ3w30FcsF/k3pn+wjgUGj0rqNYcst4L5R
WPbV7BbbbcdTnv4OTixRFmw9wBj5dY+CXlckZRW0dv0PpIVXWEB1Pxm5SMMdBSil39eh87ZcyzGU
TYsQwsxpA0qlUjpsPuerbx33X+k78MffM5zpH+X7lgLCjw3IohqI37ma4cq5ZkWjLoimi93aUPQM
q5WGpZoYQ5xx7yif7p7UoH70871U8Kpdtx1iF4xZpLNZd2YBUKWH53dhfqrYQ3yTvgCkqALOZmma
5/EJOGeRKm3y6/yRWOxd2ERoNIB9es5zFPJyQqnPTjpRWfw34G7uv182lXacSCCfp+fSGnLD0wnj
nBRx3WOjGWeMHnO9/5pZ7ixs+tecbbyuLHX7XLKrlBvHMuEpxXcgvx8trPR26cYwFQc3shotoCwb
LhlBjkZPWtkFguF2LZROZ+dwQ0tlje+ja+s3mWghq59teuPG4/I904PadEOfAtU4FK28/X2JZHrB
b41tobdSv1p3alyQvT0T8HPir6YsU9kv0kPRuTB+5o42sJt2oNc967NomtsWEcoQN35Lmsqo6iMP
j7XNfEewrmcuslOTUOVZ327NpPaWkm6GphPCutRwlq/YXpBhslnN6KONAf8Yc42fjDTZkXrHDoso
u4PCOJqKiqe/WxHL5IZA+4k+sCjkyR42yJmaDc2uNv5fnskMH8rXeBO4ufl4QpX2IqXBSH0KUl9f
2wXozFyeGAyVS4qfRU5pV31Vn3qosSNJpHlkA44mbRU92G5pXJwkxmbVON7q2kRJM601Ehoa0rnk
Cr1tAUnBeEr6xvx7otmkGNCqeL40IqesNz3vV1kFBJTbyDElL/YItlcP40/S1WSOYybmVDzy9B4I
quyRFdfA7hrG47NeXMKS1PnuUVXWIowhM8DwzGrYPkiVhEPucqcgzYHEcln1MaBUXxJ7dA/1Yoxc
rlLX8RyLLkOhvFciYpzLnLdDgEwGcfj55RnoYaEoIhgeCdlmM5yQnG86RXintjTyC3bhssqpAL7f
dbHvbWG1f6A9MkHSn9djKZTp89ZaHFYTaEr4flD62vSG9YdtHM4Wp2uA6CRPmmTnJpL6qA1dkNgw
91AbzEjWnVBaCj2FqXLCWQlK9iOZhpygDNWwQCpjJQCq9a5COiT1mAHtK5/byCVNsyNhhKX3NAzP
NGsQYVkIvR9vUnrcgvNt3azQo3TWxldmS+t4lysaSUCNgtO7WfZ9FCGO/g8g7+JaXC5Pu5luqfB8
Vy9n/4tIr7fWbMTZKWafgkaM3/caOQtpjxDrTnuw8CSa8PV82BEa/4SAu2bHkKjUl5Fchclf44i5
jkcbsCl0MtpLt3BREDEr07oPrsNjZGewdvToRJKE2cEs0cj3Ejryk2UrwdWpR1oaflB6YjFLSPfJ
jr5RImhB1/h88/mCF4ycj9FohFmCfsWU8WXLsMvw0CWz3LuIscugu+ykJC/PF9ivF4/QFpbytEqy
mnojWkDx1xFMn1wEapiMRBwRrW7PbIE6aZNBFUVVyKTI2MQoy5k+VJ1Dc5ZCs8iVFXm9m6DQqqq6
Qlr5WOFRxh1mkC+0dgGc1lbm7DwDV3ccbAgRyZ4No4xN62MqIaNLzGGCsGsWsO6+70ye0bh6OSFf
H39JwxsRCiUV2YGijbATb7YCzg80AYCtvINvmE0kw/a9GIL8DBTWmyBGJjcKARTnLIylKcnx9uae
aRE1a7pivOcG05gRH0hQ4Al/oH2dVhVgR1CG2BOtbRnlYtYqqgvIX1StAQrg1x24B1+EhSZ5GVBc
6yrBuGMRTEetILlU2e+VrmzzGmv1w9CrjI4PKfh/T3bFqrrfG1TIkEomQVKRXP+Xyy8ghv6/BTRN
/KpVWkPD54QzapRynTjl3u7TwMEh0MpBAJH+ibUR+1Ao/hiAXLjSGBEL/3y436LRCmHt/nZaDp87
eOeosiLF/zgrkpF8+sGTpvoTl3K22XscfIc1UlTtBJPfTx7XyJFvQssclPbli3q+whKFh2PTdwzj
8jAS3Y/O649FWftBGAFTzf+TOIYw5j3eR6VuAB5qsj261LY7EKO0grJg3xBxmtK4tmySEsvtKIQo
SFe5GfT5D+2y3MVlzx+oJU+Xv+rhIZsoyZ0DYL4Lo6/ZgRQKBUBvC28a+HpBWNLx6BinLxV8lgQD
qGcuxd0Qgq2Sy2aDtRAUuIRwEZHpR0GJa+U5khm7cC1Z/Nk31E2jdl/+JTRVav6+u2s0Zw13wOZo
DolYIyT7fJDKgrs1I4ar6okBhxwJl4/teJP+gNNtzq3gAwVYpDmnsvPDHZ7JFzl2gO+sh2+jpgCA
K/v0eWW2DNFMemoTwmGcGo5OqQLkPDJxGqU7mFyStpQib56GK5mctWFVp7PbxPWTSYTDmZAiPVH+
87S+CgXvUjTC/xoShY/zFzZQ/3jQSd8zb++o1NW0zPTEuzW7+khJkC9DTCFyzIM8fF4ObnoCWmTA
d1M9A7TNSefzpJXdDvLZEEC8sQODWrjU3QOZhUKYMMu88Ufq9XLmFMUGMqwwx7E4uksjHaYSbqKG
QLfSqg6Y/1wGxpb5XqGt+vryYJd1vkzyMesh0vqjpHuel+/HVL8g3qpMZ02Qja28ZxAoH2vmaAVn
oTSVN1GQJLHl6l5vy/6lnsd+xFL1EaCyF4yTa0JUir0FFiPdfPAJAw5wUmwgUTaOMv/5x3AnFlm/
Wh/WTrN63emGjcHwYYfABovPOdX3jBdh5KnQ54n8oLg65fjeO/zn+itdVaeBHx7i0sWXETrrjNi7
r4k9kR6+G0Mhia+y0TY+jpUz+Ebage+8Tn5evnRGtck573LVr2k0yJxp18MdB4lFwLdDVMZXqd15
emEQG7jwpUUZrqwaj3+zhLfhuB+Hd2PRbrIxDx6gVvWEJ/0Uu92RNwd/KyDWdUDbPfNkInMWrd+J
YjFTW3WhIMVEs08Hrii+R0OvKYOwo9gJhRBWx+3pQc1teDVpfGRBfEt8ywVTXhnKghFiUqDZH1mz
e4w5vy7y2GD4ERcpoR1sRrfRMCw7ATCbw4X/wTI+5MTL7JZmwkGT+lbtWuUJegNkOQWJELBgZ0dw
qcp4tR86rE8NccC97TwmFVp+RLizyMgHpJ5wX/G1xnc7DrNWuoRXERPbhBUJdmRnXwZYSjoA3VsT
Aq/2VypUSCO0QIBWHxXgoTVlqQKnckAY3QgJnM4ZM/LpsOVs7T3yuDJSixcCKMRH2T5eJQ+EV6Ao
vkmfRrobL8B7WfyJV/rnDXxzw1fK3GseqGxf8FsT86ufbDHCgzy/eyrbE3UE9PNzfIKwOrvqJHH1
vQ17xpIgAmXBUgYNkZ6X28HCekfkkHRidtWzfIaWzma3BX3+w2bD9DZ+iLnqPtj79FssPDOX0+8/
DT4dsSv6l+bbMpwFsyViFq4bchRs5w5wkG7sh7RHfL7PfKMSde6sG43EYK53QiqVh7KpI5r2Jgsn
Std1I5/vhx1mH9SXsnOii7E1T5xdFBMM9Ky/Nw/Y2LEXYy5d/AhgBaKwfjHM8O2lDxUwlifve2SY
yZAkhZRPgj2urcIbnzyekyMKyXAtvL/TZCfRZLQV/y0Yd7kjDHNE+Xpga6T7pSqmmZl14A8dAg5V
OvQBnDvQQPzCsy8WRSuic8w3jq54pIPPeY0BwHDGlmAeV5qOaDi1ZGLFGngT0CQPJ3WQp9SyIGnG
Y/FVcMSMPZIkWtMwaLJxPmKXn9bSImAcz0Xee4hDjciUkkHwB1qDVG0sJRiPoqYVllB7xitANdGw
EUh+9yfBm7ywHwtoSoQMBt7aAJcCdrdkUqeKxl7jCA8WnC8RpjOmGZ3bY2TKscAVrc26q80NZ6Ew
/DbSuqEStdh3r8a+lEl4+X8sheF9NXnNBsvnS6ob+4wTjSwnnLik0hH34trXJ6Uco19yN0j/e36X
nitQybvvIwRwAKYTKvMCa8Kh99YYdhRohNLdFkh+3hYidGjeewYIsjHGrFGAXTFquaY/QssKzt51
84UB3pmmkpMQvCD3p12eVcwvUu+/zWjt9P/jiHJ+Dd5xVkngtQelvpJww5lWFfVtMhVAIfcAO+be
ZmucbY48nEv4yBor8ik7fxwuHsSRCeqZiCWrOnFlOhRKrw/ku8gNN51QmxC2JDKowV34aQZ6xMQE
VKcLX9WQiNQ5KPxfpeBC5O4NZ659LSxyI2Su6uZt75g+whmHCc1VbY/G2Vf7b+K1mJTwSCIr5t1+
z417wgwJwwu6vSMcgPVg71KsVUF3d+8CEn5GgNFfWgoSijdXGnHl6x6ZBruF2WOe7PA5+INONUFq
8JVWWTRCTCWxunfWD2hxZQE3xtErM5+seKmuWxVan4oYzrIaKVjzx+284C2vg+2cQlk1xapOYdpH
D8KT6/pHxuJw5Ldb5PJjlLo06Jx+Kp7uqBhBD2b9mR2qRT2UFPkBCflnBEg4VKAuLiMl4m06KgCc
bEeRqKh4mA1nJG/JEOd7bVf6vR5eTrr84uxkPZeXSO+cTLQgW7uvfzeWuHSQZ7Py5cFpw82nWe9k
Re4FLzXlgY253eQWJ61KmQSIQ1ym5JV4WSYTnOEytulY1R1tsgpzDjqhGepy7PvccRYT6aMu1UNz
jW8boiTsQDTOOSx1xAUXBazHZh2Mmx7osHDzlHafgBrUY1imwkGH8BPdaSjaP9Kv0feacwsBimB0
TTgsq2ahq0sKFN1GyHccHHxBDrWTZW43egykgnsjlrKEf6ZyTUD88QUFtYc14C5PAsPdE1gx6dvI
gj2e2kNAqUeArnevGYXIetgn4XnkJAWHg5PQA99iqegGiuj1r5iYQv/txk663Pc3Ng4jQM3PHbU3
bT5Z0TL6yvHg69JKBWQIcNpqBVfXLSf0QkW1q497NlPbvEy/l+gf+XId9G635O3meoYKcnaAt7KQ
VP5mENAx7HOVJxk30Pgmsy+3hTqyx3zRVJTeKKCEDdMcnqkWaULbc7HtqQ1QBtNYosoqOc/lxrYC
2Lu/ZuzQQgJyZ5fAVuaGYyU8cB7kWgsIk1V+hiZVC6oqNB8w+36vJjEm/bX1SXhecVWNkSaTTzVr
uSj4tiuVHi7PpgxT8JHLsUme8yz7+E/S0nDQos+G6/vZ95EDaok22xIRBnJ7uIEGvuqIpZ3K+gOJ
cA4NUyF+e7dssHDW/1hS3WFdTbvrYeZV4gF/pBE2plwaflrvKbOjlIn62swhKrsk69NhbFW3xgZS
0g+cQW1n8CEn++DDwAi92BBMHZf7j8P9vlj4ViTc5Q0PUDhsUhSfEszpSQJ+eud/+eqnr4cIqg4o
MIk2JX/AJwC9xOgd+mt07ODFRlzVBEQ0RylXDIBraSj7WUFZpVP56LDtE8ObV61Re3CHOAOBhxoK
utk6ki7jTQmhzvYLLX/fmqBF957ln8zZ3qCjiZZEmtLqQdqo5LvbFgSb7tRkZ6eVBies7sMmaFO1
xv2aIs7YFq3qO9iFCsTlUcIp0dv+IFRtRzJm70RBG+sOf9fGdQgXzwwjDPOzIUm3a1GcLY9sRz7O
WReFMeKvGIE0c2TU2KudRIo1xkmjNjZrBEHmcKg1iZf3fDY7Eno7Z9m6PM1cd1d0jG0ttxLmruns
WlRK89Vj/xJdxzIZMxsWqZTsxjsejw/1lhGlWIcrW6ZBlQD6WhgIYUFt28SY7BAK43M6mUwP6Q6B
M9xEPF+YvllZGqgwSsuXVgvafuRV68Suq/wd2CK+j8Sd2OlR7ulWYn3AouAn1lYXtdYQoovtktR4
BwfnzzdZn65XUaAqTS3ixqtwfgRO3RmDqtLTWJ449tPVV4Rlsi2ifcOYCG0njNWy8OYVCBE4SIpX
1xs4RHqU9T3m1LtkicPGkyQ9JknvqnTV9qHNLGX4jelEDxrJXTgRWJxD69TvHZ9E7xtDgh04WgRp
ntMq+j//sF4KgFy01rOIEjUYSzWKkSfg39r4jXgzz+gbCaZL49XUzFRoXiXACaHiX/QwtP5COkDB
zS18hEtgrATkTI44TNrf2he53PyWJhl8U3CLKUoMLkeeNIClZzifiL2rEa9RmGH+x7dYAZ4zVuRr
NqRxljwNYmO8RCTQRth1cY8kNHoAfKk4l5GASO1kZPqahOpSux6vWZ1P+epVEqL9t+bGL9+OhZ0Y
ZNl3r7s6MW67PYR0tsWJwrWNmLwxjeqsQZkQt3DTMSNWqDKbYfBh5RDB8WadJLprA1JX3WYbXGns
xsihuzIP1kOmmx2Q8QJdv37mUKkSE7SZfZko9d880VNnZvKJFenTtsTvodAjolwXIOY21CERTIFb
MGoP0sK5j9p9P/2JDwD2FPuCzBUmd49rPq6YEixYQg0uziPj/mHSi85qnOk5gDqSktVsTV2h/rdV
PRJmNlBXHSSSbkov781QLYoZF069Kx3DSseT4Th0fzVDiWcHA0R4NxdT9YpZg/SYM4zy1mVCsD/f
E0vgzu+fyam+zvS0q9J5ev2gRAD/p3r/YTUEQq+VOfqgCzpdV5aQRMGtbBK1ibzQn7CyfqpfI4ve
lBx7TSzwXGmUd1kzvNgB3SvePEqbPQ3lVvAqowMjCk0Ycbu4fc+pV8fO4VOxrUDAgnLBFSBfH5OO
UL0L6CqKNlc2YVfK+f7cLGdWvhQvq3cnp1817FoElbL56xPTe1i/Ny9J3qQNrBcx94aAXVhH7K6k
HNimSJYWZdsH4JRIz71PbQJFYVDQkpXgpfT97CsmH68iJbLv3VGfJb9usBPz4zt3CFygW5OZ3DIB
Z2JirZMT7Gchw2VF1aM9J0mrAUQWv+Wsp4o8RwzMdEUByIYNYIu1o35XLqGPHd09RF8hP3VA3dtM
ILiG9Hwz2UmIiJm7msTYWC2IkB1jAXh4yQ5jgd4/FmN/yxVa4/wnYRuMiD1S5hCtQ3iJkGDulm+F
axefNLG3FJ82Td//WwqDiQ/43iPjP4CS6Wi+z5H89iIyybuTH9FKwLi0W8M2bTAOUK0Ep5uo1zke
Wo5TNRt0bDyzKVpXlYMvZXXULXgHAs0F7gtZjHBSdMD7261TkCV81TKJ42QH8HGaYfmdCr4oiTpX
sk5ixL1lo6HFZ620VOJktBNUEb+tvve05w2193aIpuuz4dkV6xJEXGmyj6SRkQilydGPxomT7M6z
BRfMoJrTiUFy35Y5OftV9wNuDZkjPwVOUfWjWyctRJ9iChY3F/AzdrObdpYkaWVTy3TEW1F42c1A
GwOzTcbUE6gw6TDTFa6QZwok5IxHB4Z9H/+LFHXi+nsBhQa5fdHGL2sZVl0VEA1Ln5NTzALWSwI2
g2r1OUCYFxHb9UoYthzBjYZp2Kmi1UON+GfLT5ad6Lnr0x5pKh30k8NpdWSsYJ+xs/UXuZ+jPHtI
4TRzngijANmBoPuQyrH5Y0eI4rj6+QEd8+jUE/Xri4A/OgfGM0VMAdY1PhR6GQDqeHX2/CcKBNfx
2FVIOyYIFcL6zmtCoHm/fdlWeWXg12eI0+dZ3FO1NtyvTLKILXAdchU9AJpgfmNMgFSvzQliefcc
JFqDHdvd0vl6Nb2Zd5RYJTcmA5AkM4SZwiC75IOUm5QfuQ9FHYv6bmgaElJw+nLbSlvAmluqIYAU
Hn+5XNVWhbI5iuvK4IvuUZQsRtHTPrkAT//o7v5I05W3GgSFfwA+SxNWJw+0XQLduWk68IFyKUWY
8TpwAMuk0bztCx3HBWYe5IJjSHGjBy0aj7T8fXS7pxde+KKqoNUOn0CSoepyXr3F/DwXjfq7CF9t
YoLzgOEL0ocaoMSD81Lmf9tfOugQldVfmcJvC5mMLF+bYJJ0SvHk2nDifxw0E8VUZoTBJbbCfLEQ
OdO6EnncyPdS2xOUr/vxZrtkNwka9SQx6pJ751ZqfcUZ2CGc2Y8UruoDIUgRyYxfvg5rcA9AxBWz
toQh6bFo8Z3ZTuxd8RCfqyAbHrrdMTnGkOfteXkVTO3FVFbHYZeXL9+/C/sSXG4CY4dOASGDZ01P
Q7zMhr7OC/8pIvrj0y/Ani5JbdNLSDqt3JvMIteIHAUg49raIMEXQZeyouxx9+ZysqvES5MO8NCZ
ZLM67xliTQa21v3GiU68dG2fFs3pnxz3bJ6UDj33z/+tmA+TMKjt8hlA/B0QFfuLOVI5vU8Q3UWr
eyK8QXmDQqlhNgaR49lwBLAhIytSGLztmYCVNuH4hnMQqfUmHAL2EcovKDg/73blCDgY1k04lkIr
I8WR7iTgOpnwEw3F3Ldi6o09+MsAE6NnZt8Q0iawIOhKzYuohpwp8U5fVjgHWhStrFGThJWkWVru
XCM+gU77gJk2RS5yXBY5ytyq5wu9L90ADrL5rFxC72okSqJWQO6cka6tRAQAM/Qw5+3OujEQNEbS
bc7bFpsGLie2Cw7Mr5IMDNfiWIOJ69d67jgKDLin7iHwbxld4Eaf+HBChPTUpl+Z+u7Kk8vHs7BT
2gK3j2RbXUDiPXWhTCg3EFCGYkFHKvsNSxMGg1b7VADzHRgWtEXSsOE2xX9KFy/H+Y3UL6xRnZCi
/jjzjfkFwFzBHMTUIrjf3ulpHzvRku6eR42W/IzAkBYfOWWZi2HlCzW3yaraQCCVmmAsb6jgQ3Tl
4Ygf23bdJgfi5EMoqW/umyWPqL9vV3tx7CHS6Y9BM8xb60BB2pvmmYIWNOrE0ZrdB3J/NXjF32iK
JyM0T/UdISyKmHq3Wgw2V2SQgKrZIUjyPG2r8nrMZhuiRkBXG0ZixavMhFIX2EUP+uhU+hPo03nO
m1C9jYS82OV/dMsQl/7PtdeF1YVxUkneLNAFQp23iQe/sijV3HJoBzrWsetF7H1+3Q73eUP86HyJ
r+xodZ5rKvkEp6AP3gms6weassDXxsAceOxQyhhl4HHOxsMnyi+pIPRoALcpPvQvn1DqmV+tnwqf
Chtl9wv4lMtmBa++VluBWeu9Pya2k2dUWTh4dREad2QLtEZq67f0EYuoV6k/twgWHur83apaClzD
vuBDIrTlZfRjiFs2Ae+enbHvYBB9f3IVc2EbspxsB4sydGIgFDPn4tO+T/vFzwMRsFLUwYvZQBxj
RETmbrvJ7pDknkEAUEtG+ZHZDzwqSC7lOQkWWAukqbrMqAEK3o2KloVlQms9j7FNUDYH0daZnqWv
STFAdQGcBZrzEcnV1Z4ukM5GBm0HrNw15mAXnYwzrVtoAyDOmQTMyzXNGhyC83WIsnmzbD0EqyQ8
jF0+AJWCoRvcAjIDaX7Phf+Dl1p6RZng7a5NJ2NiLs+EJiPWrVXSi39WZJsfqf1y/7jH8byIjsbI
vSYFdwYhOKZ04UpbPAbB9AEYKzr/svE3iqIh+QXbg5vNi2ckfpNp1iVF8bgTqjGWiaGUIeqUAqac
CstyK5w2NtAGC5m5sPwUzyq4GS9IJCEb2P6ABZ1EKgmfaQoLOjirEku8uDL6re8t3EVn8ffAzPsU
4Fhp9URUh8gGrwoCIQshemgSgcT84mz46rTVSVC93h0kNZEJPx3dbScN0mHbVWbGWKKlajSWlV/2
iL6n9Zryiv7/+1UvFBTdlR4dPftIijxmn0GkY7FqQ5LkcOvupEpOgKW9pNJ8nSaFF/CHnPG2zXaw
GmiAokOQ7HckWBYNWpoeEhaqUQCzYIHT+6w9B1Gyv1ETZekeEvbA/BZ4LAdM5Gy0OpuPs2N190P0
EzdcLy/8CqoIZYD0XuQI7rqu/mDCFC99yjelGis5VmJG/r3ZXD3ShNmKLKirW2zggepRHlsFSfTk
VxxwPi6Zuiuhj4cd/8zt4Qu/qbN+kvvkK19nRjJdRjMP13dV6NgzPQZ9GGNNUSQw2W71Gk7zHEqK
84G1MinJLUaWCXg8oPPwq3ao/wOVlKEQI4MzMrPukBWXJ/hy/2TUII3hO+L1Aql4aHSORCiwy8RU
0p2IBGKVAD+rArp46GtyiqTu51H3j7L0hNhw50FlI6lk9sMW5ISrVj6aIdq0/zNipI51634EPMMc
Jy1A3uvZyaN+MzB9JwSP4Jxk6g+ZXw4EM11pyY/7oSiGC2tCjdCo9IV1nbdyNdkBds3hjm1TMPE2
5JuhKcA1wUg5YvhMtizVAg+O0qgg8Q+Uc+r2MztP/cFuC3WjzLDYnKAiPkv4WHMeZSbJWFa2mtaH
asa5cEn9HAAoV35gGru14ztYATa6KmTU6Zmh6O8IgTViidchzQN/y2r2sZY+3Ib+wOyy1jyrpT/l
zGCD9ZKGUOKaWD3LFz/J6w/UqebMusxqRYCWCjH2IPXVvfLA3YII8UlqhqykfuP7PamEi/1IHCRy
qrixOUGr+jo7UJ7nR8m5+Q8ZGoShmJEljMH5Zp7PaL8qSmbYez461Zj6Lm1fxwMTytjItS0Xu0rb
QUdd8sS2GkpZfs+9Lnv33HPRDzVUt0B1JW3THIBM6zq+jKzOewmYBXiISd7/01XemsmNva64nS68
/KF/5A7xwTOc1tsFaA8TwFHwcQ3dIuIX/QUeR5I/yGq+oA/giMo2ywVgjsOSdnpAZ7VEjJP1d49k
NeAZ111jc3JBk880ZhsK9crlN/XpdQbttpfF4vfsmA6K/lkk0rMB4uN+ym95zf4qIsh/NpVOCFpO
YS9TGRRXSBB05haSQVJNOdhNxBjJK1AJhV3O4vxOszs+xKHkXZjlgHkXHiOs3029Hp4bCUfIzMfX
vIuEanPsk+QyVLslFJ7iiiMWipg4VL/pUwkClZb2q/dk1feqM4RrY9qw/ESSns/FTMvDoR/W0oXi
3qL/PA0/EZqjIhoNlRX+N4cFVIE5AIiZklGQnPRlWg+VCPesyJ22Y7QZ91qMTvo+EOI5CvCU51ym
UdFJXsDBnNbh2x7E4Nt2BpNp1xqRHnpj/ywWGDE8oxVbGVbLOCLQpaphjmqtmDtslzpyzpQP5tbR
2bfoiabnO+Hb48mcFe4NJPlo9IihdTOZPbZNuX/y3P1Q2qSt3IT+qAHLmOzU9hz9gGS7/JISchc7
TOZWXPHD6gI4JpxxpOz8uhNJ33REZKA8b0gjqOtQzTqpeMqP0pHzEJbJbVAxewsNGNNJACtXnJ2D
/ZWIrcSNWMGMwY0TsK5k04luQJQNf5vrjzo/QVJBLv2YEfJCWiq1f6SABt3YixV3P5ydENV1F9Pl
iWDE6EKUlc8eCYpbZ89iP3zayun8Ja1UDSk4RRx2tWmOxRM61omHLc33Vn+Jn8QGUeBenoQTvyev
tuR1JJq44qysVHFrawmX0lBwjs5IIEQ7x7P+HClwWZ/n9poJa5N+tgReTugpnEQhLQ7ocOi4pfjM
0IhBPtMUR3vWFzv86PitzCZv6vvhOU+MmEXbt0dfZSJGKBNkrSBUZDKUpsHdoG+c5JfS1bmc1lvz
h33uO56+SWUtpPXfGuFmldfNkA20BAJceYhdA82VsO8Fmy4LyrQkE6+kuE8Eyz1TTSt3r8vdNNMP
WcExvJDT+FG3JPtuCpV4js8N0KFw40Zui072CSPAkQ9BoxY0meb4k9yEMLY8KOTDGuakCc+WiHR2
2EyXdDjuF+sOaZbu1yu+sp9/7c73PqSoR2BANWbOqTvYAYR0OJe7A5s84ykMYqcCero44dNTgonj
l1LyMs1LClQ3nqazEMxw6VJtB03XUHtA0CDxlAJoLfHAqQaNTOuYq+bqmXhHIp/gq/w7IRqmhlN6
oF5XUqiy2HN6mN2Az6wusoiqQ6jcKoWYHjOfKvVxQq3XmcQ4gwyCdEeIqJJ0oy7rAl40gsG9sYQ4
jVul3HiUScORooKiY8wMRjF6EARYb91Jh7AjPfuoxFlWcITwlAucOpcbijYm/n6/Y2U4vf0IQR/6
m4nHfE8jSi7b1RGN9zrqbV8K7BL4y8uuQomV3JhgJ0hEpij/C7K3YWd7lnO9TxdRWB+ygpVDXUl1
6zCkiC1CUsvHGO22jJkreQomXIEza9Q6OzG7ChpKaE0vHq+2AVgdfrx88A7As0NUlMV1ccuiY6Jg
GOAzEJx1wKaN7o+bjoZh0u2b8S8ujPcg18CBbi4ZrZ1h0wOfKa310XOpgjYa4UnX/af53c2b/Ufp
99kka7lFjI4Clv0no76khol2Rn4r1snt9ja+9VqgWS4F+HogdWVvkalrIYEomy9uWoQwA4M+HvPY
8/m1kk/FaLBFh060IZ3BfmP43T66y/ahMhBrATUoXgz4hMNlfccQyT2jew7KAiwe3+Zlu6NVdza4
XoVuwQsShl1NwEDfpuJQO+PqutllZbr9JEPEWrlPeBX7kqbSPpqQ/7qPJbrNNvfrK4XtDJ6lVgNE
BmiFfXbK1C8shadssFVPqUzOcYDpmZSiQau2L8k3uqeGN4r5WooWCHFfMwoUHcgeajd6CX/O+OwE
DIfDtajxxpGAIVL8WRrbwwh9OPqDhs/GD0s5Op+HECvmyN4sQPPWZljyZwwP0ofZ69mHq4gSrDtj
vj8205VbYxG9edOQrYQNsQ637fpiw9yNOqOfzLBO/DpHAVb67B2E4WRQYfxsh+gM2PLpfIpdRLfd
GeYAlkOWibgPBdvs6rVU3o95Uq7C7MgMfkUtBJXXFmYNbzjlYQgvMfS9XkHqbcuzVJYJVlsiXGDg
Ek7vyZE0Qg4sADw9knGZk2Kj7+83eRAvbXER7olHcx3WoxOEDA95i7AvrV/yy5m+o/9+nNdpctcs
AJ752Vd9yPzSrt/1axb0JSEGpYS3L04xFOW/bqKs5iUvWQFEpzeNObQRBGy6ioB0Tq8Y5QF/QzRQ
13K7GFGUmYkdudmlLbkCBHK2T5Ibml/TnLui9l6fWCjXA5yUdYC2LKjQsDffdlDGxIy1MXxJy6y1
/QHgR0kKcNI7NMmOjmtIW+n98Pzq5QrJro2tOSeVFDLWEIFaVzJzyHtjGOolsR58yOkJlqwPEvH7
WrS6f25DZ9tLHdFuOxfUQEJ3csHq/CHy/b6vgXBHtwv8wWyxaTvXG4X0AmU7WBRBDEbLLvGXhksh
0pKHeNKQl3lQpbH58Bh04DHm3X0dLaY8OBNUF1qEwOr4wDjjfQk9imIAWDqR+++5DdvFF1Brj9P2
WjtYTl10AXBQEXXILgxj121szC5nuOyFLNysgGc5c9fYdbKTanEDFlQktu6lp2gLJ7gpl9vtlKfX
cp5XlnAzIQvd/d8ZZJ02UKN5FReDJahK/rX6pEJeQ0nfaqGaKZq0c5eVIcQt2Xih/VnLvPLLWPMy
oDFPaJ3uzIKqJNgwJzD1gfmAvhtYNHn59nAZYCKIb++iXY53hx2FiwoerRlXjMwDkP3UgDmwCgvl
7mP9VTkroXqJK78lb7ZUS7IJDiQr+mQ7jEzgpDy7BTwd1VGJvBOfWGADcWSTDJMDMl91N6OjFkgb
lViW0dQBPCZuArDSa9pdUwZNPAJzMp4TgjUiJ05naUO7UbDNVmUE42f+RtSVeToxi8Y3djBT6JkI
h5pYhIOxMVlI8O8VkqUwQxpXrYmP4XK42zaQuPFFMZC2dkDB5UX2Ta6KDhDYDYPgAgT5RUMW2x5B
HxQUJdysR7vaAAdzdEwQxDkoBwvFXWN+rp8jwCD5XW2rhe8fY70U55uUrOetWvKseoCYUp0fr6Yc
SU7GKYlytsFncmUdumvn+Laz7oxxKLIM1srUCorHo7BKvdn44ACuGx94y+EFPIhlcR+dwsgN/9tl
RqCC32adJyMOH+jaa/tkvXYP2Fm1kfrbjbAZPl+zebzkt0nf2NQkfc0LoRt6K6W6g6T0pGAF+7z0
uWQq5E1kl+QWWgYz4EWraktosMS6tHokSsbsqdQSabQC9ml4sGIsu9k/POXsyIutFt9dp7U5dwa6
LonG7+JFfPrq5C51fIvjWF8z1aYLTiugpCpmvcURrwe7B0M9YsRIVuJXx/9kyTKIfhn2Ewuqk7bi
2Le8Fe5YsceXjcDIzcuqhEwOSImcWfRuS/EqZueeDO036eBtBPr8YUEK2PSbpZJjnkCvTpSih3Jl
oQCuJTvm1b/stC90EjkfAmJ4F/b1fwxkFSqRF3gdSA+TeAJ9lay2iqR45OdLj71WsTjgzvce1pc5
Wu5wAVuzlyCZ0xhMI+fbheXe6pERP5yDmJbWFZUmkPXExbHqYh2ONmbBbSuQ/xFvhKfga01N2slp
PBSZdELwYX6eC+A+Bx3kadbqUeTWYsL1a8uHikG9rZJDh5uDb4cZtOQ5n6CbTdhaRsS7r+LHwnfF
W/wSdrpDXPXHEAKVgh+VcgikBVD5O9UhA6c+6tQkWXgUg4kDVfyZmIX6AmZigypTTWOYeYVtnPZN
QRo3EhCaJtom8VmHn7Q339cllCsRYbr5kCe1QgZF2YKzqzzJWxbYwZRF4awXnUvCnOGxPTJ1DWd/
H0z78dX03/ZQI26Avci9n7uqcs/gZjIhtpSrQQW2gS9J4YdPNtsMq4swnKeTEvtnFfaVBtyN94mN
AkRaL77vrAt05WVdsWSXbiCnYQaBb8WJKdwmeuYH5+FhrDqgzvkZkT+l4q2G1lNZP3kP8cx2h3xk
bqSD0fSkoUKvWNA9sp+i3aiGuv2Fn+944HPCR6Y7UCYmKlRbPV3th9p4sV1kaxFIXA7rAmfEa7VT
kHG2ZLDHh0W89l/2+RuKNp6y1000L310igGLPjyUKvxsEW/cghdg2g6pbexJEbWF+4By6sVAnS1n
hwiym1S3Mr1XgiTYjQ6ko3j/OxhkhGJ9adm6V9tel0zVLaYsglAcihdTZpeDFlt+4YDxg5fqeOur
0HQF97X643fige4qSlmbFKTG26lYpVdP3n9Z5dezezyzmW0vxZVQRFwqc4/+70c+B0fC6/bgi4ub
tO8UQlgbxE7yB0i5Rj76MkOwJxlHR+FNmkrcIduMlPRYh9gIQtm5t+uUCEzE1DjgR+R+1HvScdAi
nauZFg8P5Pei3Qth2fMYnpDtsTwoxlCTGlA/RBfopCoj3F2kFeO9L8c7PY0aUs3poGxvWXZEYjhK
18BlbYtuuwOciGMLSSkH75NWh6EynwsUpvSPGwIvC5IjnMCXfGvyWCGq1xgFQbVqbBzvTTYwS3Tu
80xw0CVUWfNFmEyZ+3krOBMYwmja9af7YCF0tbru5MeTuNKnXc8cr/lYV7SVpKlA5+0hoW9p2UVf
yNgluMHvyRBJT0QNjjUKvYS1N0M25Gbay67PJtSgZJOPgKQ8SgBjrqwElYAbnODlQHbDKsrhHoNw
gZ66rJ8Y0df6PST4ORPspra0UoVg/rXJYmJD46P6bDTTj5QrtjNW001Iihw1iIkV6ERyfpu5+eep
wNzJQb2D+e9bzpyd4V887NOILBLxcQSi7RH2VXsFzKVDqBtwXXRpyRJX9jgFHyTa1tz2G4cgd6ZR
IboL3n8lv9JKjzWReOMM5Ze2FJ8JDdI5VApNmNMVU/ypkknDhOJmr0wJEBbYufTfsSHdjbtgeLKW
78sYGLzHQcZCLpjihwatv3i4O/z5UqHEEyIRODZ6EedhnYyRDeMtEKuAm+3s/A13Z0sTp+gGxn+V
9SVdMjYyw/4Ko10BeY2VsdYwqjNWI7LMA/wyQ3g9R8GgPYEMoHc1qDLEOtfRqow8Su7GR1oyp4Zr
kVTf4WPMYGTeAHozkwKjC8BkGcn6w5CwcGOukSP41opzqGPm5vgPRH2R3ybd0yW6rRBzA0w8ERda
7G+ctPW7PCJ2e1G9B+4V7vUM96GKIaNBYgF77NAWproQbhq3LoK2ktpqM19rIupbUDKSFvMvSSNX
EOLUTSsQKTI9D5YDPbBP6KTXxAjTfQCcA//dH8vokKCC1zh8+lmL4j63uvpI0RMd1Lrt8hXe0FOQ
rP9u6zex7zpiGfJiz8P+vEorevS9pqPyx+pWCYRkNvOHyht+93KDX9qFZSsmlzAFNztNGmE/2skH
n76Xm/3oA96LhhpBnbQf58peRWt+Rpb/b1DolaSQK90YxGwhH1VBclW3r4pWTMgJWJqUd8c9+ebU
cXmSFY82VbCTlv0GZy/RXuAU0vGhy5hTJD98O7B+XPgxYf/V3XbQBNDmCdmiUFTBTaZsMXZfAeR/
6/5Zh80QP4VOdhDoC81yGx7aj6aUW78Ccpm3KAPkmK1y3zDixSWRl5M8CzW/fmZ9M1u0q+RaP6wc
+lB0yvxIuDHv92qA0CKs1FiKgJIDfk4e2nuZRvI9w6fAcj6AqYJPOhSP3TwlwiSUsxINb5YkZBOf
KcHAKVczL1Sd+Cu2HCRbihR18c8QbZ2Ccxk4sS27vo61Bqm7BRyFrU/skmoqkEGcr3EEdM/i6Qri
vcSBqliqXepoMto55chURm5wMhzXFQxmhMIKvRKMvvG/7eJjtJI5boIc1OFg27XcJtK41Q8jcMEA
LEMFy6nG6vRTRIwyfyMIfE8RqVGFTO9hZRQ5JZPI+sdq3HIx5RjtDt2NMGnachTYsdt7X6seA/bi
oxrgiq+XznfMilmhE26ffpSxwxGsCuzLjOzo3MZ1+X4vLLygQavC6AkEZi1I8keMB4LuD2W/IIn7
+DM4ZghC24a6vNfIemxBPR1HKIEFDk3CaMmqI90JSJyQ1Xof/oHtH3rj7zEP3BKCvzv2J+tF7l0/
TqTVtDVkWnX/tqRrmy3zCJZ3xeSugReCP1o/XweiBAC0AoPqaC/cMWNKKbJBCwgdZ7YqiSaRn+En
qW/aPKuqf0tFWkbVJme20p1SV7+DebjD9qiwKOQYtd2GcOYFu+k3ycmJoptkMt65YGeQMj5IrLa1
nilN8e2Ge9o6Z/nVP97aG4MV7pZs1Afx10pinLJOjpBCFAF39ZKdYHTyfbvBKs8wmMx1N8M1d5cP
xdu1+I/bOkk65rHifdGMvw6+RJIhRyT71IkFiq0N8MHWA9KoFmtd7NvdDuQqXkU4tFORc1o77Yyg
Wc1WBnUPL1L+u9zUJrXrLuCJFEi9ORlMYhl3VoEj8H80KLim/vX/yAcmFl65IbKrzs7rYr3DLQA3
D/wGZRXwV448xBGzdNW/1R7SKxnf7OaYnFJ2MZ3fLmoxoirhsfkQYfEtBLGIofvdipTlL4DiJE3+
YNrHrXuZ51iPs4c/irrfKAYP8xASurs4NznqaeGrzoR3EBBixQLb6SX0LUKfHO0bxwOBi/KGaREz
knKGUrDrCemAedvfKeFVFVRY13FCov+wmfeFQW7VOOYEiy85l/yvKIuecDPJvkTU9v/9AJomUSWV
kSugIJhYycVaJKHMbx1miPHTSGTVpYTrbuD4jpDWcqJq6G+mvVnQ9LWCiRhG9YPhvWIruyBlOuqu
izFksNGCGLLRor6gbBW0q4XJrcOVYU5br3PnPB8aIirzNg1xIoLgTZsHC+CqdTjXMwJ3JSODoIdV
QkUbZ4LJUF+kR8dYxQQGODzVshsr5hN7W6waaPObFhIfGjDNyLTeSzcI/31ZrHoeSFRUYWfN49Rk
R4L1U7GGy56kqS5w1bTcfIJeJu7ttu5sn7TkXQzEoeP1GhCIAYgMDSidpxv11AA81x35096wSxvf
5QonNGTPQOGul8MXCGsLhP/NtEl8z37A0OhrHhTFbwLGpJoGQBi+MuHbHYbbrQVSDkSyQPM8rqQ/
oasBjkXyBfdkzHfIMxBpgYoaPdPbh8Pr+StZxu7jecy9lvZn9jU8dw+KKhA00tHTSVvksYqod+3J
KgE9Dkq1mnJwby+Kpzi12SZgloO3J6JrnfTv1ilTmzmhkeyc1Pobbnwm1w+1BX5izXIrkQaY+c3y
VEMVpQfihVO5HISld0kmA9E/49aC40sugvTJocLcgb2v7p0si1LqSKg+zScBjUC26vMQ6hP48E5T
xwn2oCMxcbC/kMh0U4AVjEWURarBVD22MKx8TCCGtd8Z32+DePoY4OmY5Sf8mU237JuH9gCJyEkD
HNRTF2Y3SP2/q9mkbZi5eyY19zmluzPDuLH+D7mqk+0GTmGXH4M5K3JVQ6dTVD7XV6pcqkLS4HBb
UswxGjxJq8MDD4xwguUn1Thq2+2pDan+u/9PYPeAC4piLDiWhCWH2V849t6hS7lI8ZT4UEY07wtv
jrfDd3drhnsRYrPmKhhfeC6ZcsFP5T6Ra0fCZJ+gQq6vwFM8HZ+3D/jGmzly2lc068lV9HU82mjv
wwiyiSiBUTJK7bpyKD4qwbC05hO3DldjB6R5zQidwC6fbY/kCGvetgaDqAtQyxJ2LeWCu25L+N6P
sQokW/SCKT+7Zu/l4R+daBCD7A82q09bwhLxNN2n+zX2PDp5kC7tfeDBJHRDCjynjhSdONPIhjmm
KooTyxxGEGZxirOoiWpm+h/WlvJbx9zKTSHTuD4UMLGVGLZbFoRgh7h29kXGhuKCwQCWXwEy+Dj0
3JRGLvIxp/Pbe9fcCrTEU2uikxocnKyDi7EZ5etKXBxDTIOtyv27vHMCZru5zrAMJ1rfJwp6Sp43
ilLG/Zjn1UbF630zzrhnhI9s+B/8rXyufzp2zqGhQRZHhXAQR6GR8+3mEmKpcZfK4j9fRwZg2BoV
4GcQIvqWXXxRLVAfzE390MVHBh0zVRfhU1gKShBrUUYjPVb3cffFzBTIFFt8m21y/4phVt0say3F
VsG/QpnXTeZjsavwfX+Y8SwYZfNv++ARYQT4MOLIdQvCB7q8rt/BxyGEhz14T5/6QNrDV/Cxk3zN
lj1Qi85f3ygtmsxOW3dU5IGCQAmfEoksE5XZPL6Obja+hh77ZobgfZY6RsC1ALHaMGrvKdTMcySL
q4Wyo3HB90TCFV/XBcbZggj5hyUM0jAn6UbpSkNfFfwI9Sl3zTIk0mXS58u3cHlRhy1Eknt8w7KC
PLX054KHVmMOnVerN/A63Mt9PQm77PFzrka4vVM+Iwp3IvbldoB59QtqZpZSc524uS1WVCjnhNXI
mEn64Lnb0fskC2YbGEsDo14JbXWPXEmIkulOF9KuP60edEr7itUJWyV9ryyzDzfmagwilU4b4CMl
1JdoxMiUoelVk2jONDITSmtouPou3BBNccVb2DeXB09dJLj8MGfwZ/reLX1L8OOOzTkjdJMXiXCV
LpelC8tAeHKi2T8D9/wDtIR8H8U/D77kQ/PbEtw7YU1IB6XdMAaNM+zvpasfoMdlyWBMyIpnqI8C
EtE+hnD+qeU+6fxfBwQig6HS0A8mdLLBgudEnA96Qpxi21cqFr7PbOKqSj5qa0DoJdJ7qvulYDZ7
2wu8vrZZ0N2o+GBrrQNskpgC5eB5QM0VSEYNd3OE7oxXoXP2Ebq7vTX/eNIClITyuI5uvE89Blt5
zy60coJuNlHJ/y3Wta24AEiLxPUhQG/vTxktroqIcSTFU1edJdL9RSyztjgzUiref527h+gWWq+9
WuH66UF7dj8XiDsOE2ImePx5NBRKj3A3Lp0++b9v0gLUM4HimbpDGxWrpkJM8BghyrwQJZSJXYZC
uTIA6DhEhMF9V7Izt0tEfbKAHpa0O8cq7lQ4G8LKKWKosg2FWE4gyWmw/6+QKO+nQ9TS0PETFcBM
vXIakpVc7IIYxqe+5txjotpkoaC2DJK1d1+TcA7FPMvBOfel526vGhpkYnJomo2buoNLomORBfeB
qS3V4fsg/9cKH+//LSule9/bikvZwqQ0+icD6DGiWI4HSJOR28ksvAd2fg73lsAmSZ0MjTjqbd+h
1RDsJecaZNUS74IC0UpRtthPFlW9Q44VQOpmkXcrqsEyBZcEOWfdHlcP1l+Zbwaemv+oZl7pbRxd
M1KCj2mxHWHPjZkcoFxNFuhP1PdTxsmnt0lkdgbLgGjq6tJ0z2yOaYlNWQql4PxKSpccBmzgVqS7
WPB2c6WuwNZfiZttbP8UNQJZMcYPzna8pdK8tD0kkKk75f/NtqmBLIB46fhfknpHNpETeZH3wUmn
cCbwSjumPjZaHUV9QnatEJhNv0Y29WBUaUixImlpT/86EBYtOhyc3rOn9QOxzgn+XlwaHo67aOVe
J1RLn3sKxtcBG527AQtYi9fnl4Z9/lMnBtLr1MzYSjIysopanFz4ctHzXK77E53zFTu0z4eTKHyU
k5w6B0pl+q2IIzHUccVXSR91wQBWVntIAtfliqy7dHw9qNG/uQDikkK05SUSTGA+hSbdSliSn2Fr
SZGZrLUpaby3avfmQOrEpKiLdRiAzPM5dkGPS7pxkwnCxcLtmOxIX8o/WBE/EN97b8gITzzEIFM8
28gBJp6W9Wdqzm4D0hvME4xSCCHdVphlrpUkaq316oADUaJ789shqKNepwuoWr1HCXB3rsusEkLi
8dEOjSZZeCjdW3euRz+3VhLhZ5CpMS3Q7M2DUbAdTZDx+5M+1RWnfxc5v2FybhsRGic9IPElhdT2
dqFJDjM9B4ZzvADup5zQWOWu5zqMdVt/XRBlBNM+i/byx+nPGFGMdOAbGWEkJD60yQ2qfm4inktK
Usw4ZaNx1CSSRgTysc+0Bqv7luiyd6Pe44wV9fOcQL2crsqkbuYF+1j9VF/zAw1CuxCor6rqDta7
wWP7+VUU/PsWvV+3e9hQb/Rz2vrvvYFe7ldpYmilLNxz5uZpaXo1NbSfwnk7rNFZpAb9UFbsctdn
wkBJeOsidQ/pXdoB5Kb8GXPQoGy1kWFvqIV3FJJShZVBLuCzgdYTrc78LKQRjkVhu8+YNS+CrycT
KY0OHmopeK7vy/LQ3xF/EjFwttl+a67BOIO9vmqPEwUO8GGSrMW3RvWH7ApNki0uoHDzzXe4ETgL
/HcxB6NBYC7+6dL+1kqD2yqBiZ2VblgGprJQx5AqEj6Hm77FEABFFr+sk2XA5XpSy9zO4NquTpc3
QBKDJBVQLsMY9bxhb32iama0HxEMB3mO9sR44/n6bpgflHu8P3ynO+Ylss2ptcP+VlzjjBuIUwAK
y3D6pg/d/Gqy15SV9Gss4FHkpZ3ZJ4tryrvEQS/O6qQOQmabWVC6LAvMmwnp15GUrGJ9QOHItK6/
sWUuNBMF1zt8GCoTlH635sVmyTCdE2NKswqqjzbXTvscyiU3Ah49DLDQmI+avwTfEvP8Li8KttkR
IG2x+TbgV0GnsXxbOLn+1LmG5l/jb0wiE7C6pFvQodYbaHtQJPGQp5UmqrUiNmgEJq7YlqVS0SH/
/6TM2rRXtbO+CmkRAdYAq+2WMpRPrFBwzy1AjR3APX1rlWUUEMNk1NoOfq1uysNDBjn45NQLmjk0
WnjXvqs49hz3xexazMpGUHziF3Vw04YzRKASJe6stPNRUnvM8finuHjlAaFYz3nzflA+m3gqF7Jp
YnC54Q3HzWNVnjwgJM0KJvDnEo8e9tGn/2rYTwHliWtZSbZIjOSx/htHRzeuIbs56u3XbKtB4csJ
TVOBkiNadmqUQ24PpxHE3AG7X3YvLS1hn41wjzJ+W22wuLgIuaORplnjfXX23gFQjKD9635/AAF6
XOtyYUqxXvD2LNgZs8N9RjPQv9Vb29GeN53DBSN5NAH7ornrEU3Ap1rIVen5S7MQQoCD4bPbC1fl
ck082MLHCGzq4dRzYaUs1BXh0AisuLb1KSRPlkyCaC88rfj3lPwLWy6dufGkhhRsFytW8vBYfgND
2sCci9T4ObuDDaJqPTWgyXnHrwnYLjMlr4KyYwUU73qLUYCvm+LCzUd6H6GfIAGC4GdaqnCmfHbW
dBrn/D84RW+VpFiQn/dVPUdJj2QC3u//DEgfcsaWoVcSAp9FaE21GzgZ64nnJGwq8VcV/anqk6O1
/ATodTHeH+GXuGPIiJKXtLFFUS9exp5MueO79OL2z4f0XpcEiOjbxCoWCgJWPQ1ENxsE8vdYXpXA
XgbUuaTjb0K0n6kfConkVL/xFnZeYyMp/LR/dkYMLeg0UzRpor3ESmlZoJVyei7v6vw0liY19G4N
tJHiQDYxsL9INVWuUMsqSeAdaJ9BpjsSmyvQbZn197WquYQ5kOn2kCmHUTNAifsgaZsp+y+EByp9
f5gWNq42Wd2wGqoSeozXf0wLKyIHY3CiJJNVdkuhyEEz+SiVESmgscFLl2ZnVRMDutsllD+ct4ad
XfGAPN/4zwMRfjpIPZSXQW45EFn0DJevG92fgUFDZAEghnFQldU6tbE/sQdIUiTN3cRRDfpD9lK5
EDYZcAxOSvPlq//F6QwebHFCXjtT42sVxR3XPMp66mljgrD3Hx9RQW4ZY6XQq5TQRGKD6HM4Pb/V
XlxoIDRXTIYUnhD4+ycBWRM0sma+be6H4LjuwxwxOIYRbnpIBIXJ3YRGPtwSxl9ghkq6etSRo8zt
hv7eNK4lx/696NLJEvgDNmJ1h/rGp94IBnRrTlOd/q6SGWkDTIK/4dtDxYeJADeRA0rrAcF6IjkF
y5tnicUV/IOX4LbNhqaoPBy0kOfU5uBph/KalhreHf+ioIr4hubTekYJFXN4xC50SawctCBZKJOr
mpIlFK47RMxtfhaSlQo3nr/O0TZN5VcoTbJEEcxzAvi6AIdpa6WB2Cyh3J3XZiVrSox4z+wTBKMr
cY/D+N0O4qgOAInGnzz4Yi+SInXws52ClZs8KSNvBP+quepSKJFusEJJjneQiXTq0EF0El6q2+Zy
dGsrXrtbJDSFXxXofyPse44A4u/ncYwDCePx8/lOGDVWki3/Y1QSnr6LmtQiSyl31GQnvm4hGCqW
pwMH0Jelt4gb9vbTuuXIMwQQZFF1eMiwXm5iMmKln8y3IQ2U6r6xuG30n0x4zTpSuOc91/9FlFA3
t6DdSqYEDTEupmYZrKUvef7VmiBknXkH0B0JyfJWBOKcyq3QG0oH5gIXe8lR+SPq5fXQBP39Nu93
oMe85+hJiUnSj32tJRa8rJngl4Gmtnkc7p+PPzS5kzbo0od0+6VbdVnw6MXgQOn8usYjJ8IhzBP6
vqbQ80yov4fpO+ye+ip2pomhoraJyfdxnXCWnlqrYs9jybEBWNeihNw8PIXmpK1v0Hc00jJHn/tZ
AicwzTbY/8SBQ1TJtmUksGCsdAQoza8WbIJWnznb7onyaVgj0X6WSFF5v5RgOwh1ssGKdyjxuCj8
fHnJvvyMDOHZJWjrdH+gynkvjka8uDUzi9phaZ7uh5yH/EjmYqWjn/NM0AkLZtWCInow2u4IQWMo
cX0H0z8Ix0rIMWtovFhrswc1Ck3mpEbd0VvsocJyC18lDr5WetLDqOBXXy4bHGXmNkxJ4cxayXsX
CibHMI5CMp+dim3TNdoxUZ7Sd+0mVJY37+Thrf1voKuZvWfga43sOVigI0sWvTbDbc3MFXR4j1+2
ZcTTngG3LnTCZeBj9+mVcGuqr3pyxsjlfj/aTPd5cEXHuMphvbljM1QQltE/5SXbL1FEEPWbAwe3
nwrg+dmjF5g1iQ5qJxdzQVcruTreGsgBp8l7I8kPufQujOVmac5NsAbvuDBKgnuFSRgUonzIa+nN
eFeOFeFVASQzt3SmynPGlrZtSMq3gOmBD8AIPli9HqW/lqeO8oCpXlwy6IzEcDDo6pKZOy1WPs3p
C8muX8Ym0WVATtnX8osaJ+F0J597bG6d86AmA/Gq4ET6MVzCbWLMfU2bXzU5/oz36lI+Z2y2Om8j
AuLBzANAj41znp6JGqnWoJti0KHmHexcMCu10k9vgHuNmq3by8CqrMStJeNiqzrJ1OPxR1eYlxgB
XBLaz7EHtCwtreEJpPQVY74QXiFq6R4aJbm3aknazzp9ucT6tZKSz6M0ZStOFBGPDMnFyLkSLkt+
GXBjtpsTpf5fYrOJpEkWUQyS9fIbfqW/x8uvsnC1qwa93uh000dDa5w4cw1M8QLKtLR9QGlwL88/
MubjVxI7QF1k1e6voEU/Sv8DuhPENBiSC7Uk46/rTdV7hODLXJOlCcSxFDE6tq/sCY6EI/8KVVvG
LHuRWwMglimgHGvN51SGQS/Eod/65+2W+ommPTfh8l1zlPzCTyWkpS+8atvdd1G0QHGNTiS1mtY2
xj7j03nQYkcU1fFjnBai0l/rgrYoNFLkvcgXo9I5PqSdsTkUW5QP7Syu+Pt6nvE6dnDjAEpSb/ZB
G8rNt665i58tUkxqYjXkaYqBBoccJykNO7AxUerP9/1ZF42ud9x3X0HZmBlSJzHR0t9J7y6WFzsI
hsoCiuHPUzTkXYKMQj8/PqHpDWHfEdRbY8g6ZmOs3mki64AMVxud0e9dj0g8RtftcWYfTPwym5NR
MWu6rc+P4zSXedIuoNaxRbsFVwJs35N2hRRwepcgHmkJ8j6U9w/4+t0XaDFZMz+obkqIU84Y1g9w
j6Nm1CgTFyQ7aFEJiISmC32YJ383bHtcUq8ZCQbwgbf+mliyLh24Ue/Jc5Ux3FKDuDcfPxJs2OxH
Gc8p+iTtlsXD/aGK9ZPxgPT9qAIVdnu5rGPzpy+IZX++nVnFkZsGm1WibdamWv2nG1bxEHbHPXxR
st7R4mHzv3K8pbJ2bxeY/jMAmYb4wXYnC/yXSvKtCAxssIV9K1/cUyy/FuGPRoTZtetGIxha32QI
KHGdV2g+HwDSuDFyjGwqxDUnLYKBDNRUOmxLbelHwk3ncK+a2YB1VSHCBNmL3m6ZmOdrMA/tXN0G
P7AI15HoLW7MI4BzoDYnHZsOK7f6jVkG/DdH4B7a/ml8+F9wQyntlqnoYNYUfLILfhA9eMmUYz6K
X/Mn5tzj9RPWM/rtxc9FeR0MFSUe/5P2fd3zzzJuI2qiXf9UNxE/1T38KWuuO0bzixwO0CduS3nW
zTHxLeUnoM3tZ9j4VlRo95M9oJTKlNEaAmSCGbqnjqKEDeUig2NWYeGFBJGL7gqG5cYTUb4t3C3R
80XWYw75xugm8k6UCEORMLXNjk4qcgj4Si7dgQ1jxqe6aSnyBP7r1l24syrZEZ5ercTVFk5L5MRw
LWuBd0vhXpvsqCQjhTknZVvD0u3Z5us61MQqQFJQYHT7+ZY1UqCI5/qlm44yGw+voDmFI1yFl3fK
HQZNsUjRmHeaqT/x39o/Y3zaYecK1XvMQI6kDSPoefR63WKImO3rILsda1CNXSA4BC7oGnx3j9RD
LLL1s3igcE2euHkQha/6/cvs3oeM+SzapoB71jwZunM7zMppXnFjYrLOEObCpgppUFJz20gvLaxK
zLgl6hsmMqPRlwia+qfaHz/zIY1ijv/HZa8nMFFTbGsiVIVRdOwlI64eMEGkghhlicTh9/7hEO9A
N11stYOPWZxUdP6ESmqKyhvwIsw7FMgW/sx2CpybOHT4MAaGFvHVB/euvcigDA+h3qCieCaOITKn
6N3czRYRk+190xTt8cmlq+S2xZVEwRDQrKSyylEjDoktIbIJ76rRn9P21KZH5B5BGVM/c3QdJHW1
umzjHm10+Tpf7Vx3qBRBUi4mKEDmBcU3AqljzLl1zzAyWxHow6GgJjRxVnRHnbkfF+BUVT40s7LY
nusyCLDIY8LRGkpd5mBDY9fl3myx/JKt6FnSrS6aa3T19Ix3YFPILugCl3vWHBEgUrL9CXWU1FYf
rELwh+VY8pva6IkxtT9OJXrXxDMxi9Ft509RhLnkm+Sth1Z2O1P6iH/VG17dbj+FJq7Sw98kDCKV
V+LWOnXDxj/peEPjfuCUUGd1UdpJnGszoJJxOhCj3nlO6xDKgn7qnxyi47KNmYlkBCKQ2ACMq25i
PlwMDkYG+oK1J1R7JxPvYlfbvN6gnmtYSUg4zxyJdkHrmUGkvHLh9l8qTv33kBIDIGP++rep+Bu7
wd+aLV8QEdfeYI1JgtuKwOa7+/AzcBeAOOzfi0cv+YuamYbpE1dve73x5rG9OdcRiUCFu8qDG99U
x2rDqoEJBFSpPDEK4wP1YMQkWtao9b3SL7DFPQloIAXLgehf4lwkAAC4GsHEtjdXVi5ZZCN1GY6v
NAz8rLXcKys8eu11DOezch4JC+zKf3LPrkreTgo3C9kaywkyfwv0Oc8bJBiZkfqVFfDbgum3GRpE
dyQYrQPDSEsyXVDtJiUL5hVwdwkZTRGVpKRnbSlLUazi1IlyHtOCpRBijqQB9yj7I2NfleZBTMR8
/x0tAPMRgpGASIx7mdHRy/22cwD4ak7d2HLmI57zEJhGI5jSWGjyxEbP/D/7ieoKOho6B1M6di7f
v8a5ieR1G1Sioo5+2TBaf/OHsRHB4cdYsE2Uj9gUcxUdD/U95YcBCimLO6yWzwTNiyow4+2vgbPl
/xKt92V58AwliD/hpmeAoLP51fpi9wvvVU3v4xH6bJFjeZ0ORBMtxlGvluo9/8N8E4n6S9Rvq5Hq
SVxE3XysW6uEpoUodvxhNA60wJslMpTWqJ5K1x0rj7P83/6EkKAbQJVJdOn9F7Zszg0O6BkNTz0c
vuMex9lUQ2+RfLU+0ZZgGtI55Qvbm2FFIL6Rrf5wOuUQVrYpTiszMqR5xvpYpQSSPWfL1bnOUK11
lLn55f9PRKaLsOUsL4B2woDrj+AR+aDT0akEfOUaK6qLk1DCkKBt6UGDL4CvDOwzEgd05KmsvIit
G5sgngck+tssbPKNX6ZjGdOYuogldKKC0o3MkZcKWhnGM7WRvtdSU2zLwZSh8SlNiIoDztyVequx
blpo6aXck+KmQb6QFK7D37cjGuzKxGSmrvGEW4BBNtGwi/HWdsL6MqJnW9Mij+wnUOt2d2Jx3B9N
0vSwhOzFqb4yN7L0hnIccloyagj+YevJEKporKbu/kl11mC1D2cuKpdnIDClH9np9J8eZQFy0d/R
DQjYvUy5tNgdlcZXTVTJaeSXPqtnOpRpuiTqHFyFOxErNNxmr7dYkQQQNq+vtbyIUNPRf/nePasp
eCAYfp4itVsvRqJ2VpB8XKIz5TUvPNstDgL3N+2DcYY9yvPvJ3cS4hl/zNoneN1QDI8zV0qSEN2C
jK0N5qFr7mgn22rsY1kFI6iv8BbpeR86rwbJ+v9dlmU/fG+zqEbbTbtHBifyjJZ+dC96obQC5fvA
lJcGDjfrorGYwRgTpNah21JupvUVsfzHlfrhrqA1IFQbFZiV+Z8+SVcUek70ZGz+91oD01lx/+bD
UEmg5SLWfeMGr2qfDc+FZudFU3KyfT7Y5CLhmWazqKvpSCObgsjZNCSd75V7tvY8G3wwkvJ0sz6v
e1BaiiKQsm+rn10BgyXmZVZK//pNYXk6k0crX1BJTgsExNPEq4Ss4aId8KPdfzUqCOtYJo9sxD5v
w4s65f51MsCNV/Io6HxLjqUQ3ogdpuTTeFPqKHakiNMvz70gAT8N9vv15OThk+EIpe5XLrEE5wWQ
lxOpqfSKQ6i/WJxdwo6pXLPt9o2s3i1SvHyE3v7YumO06dSzhQsipXAGrAv/2Qbc6gMHsOW+BlXc
g5y46+3sbw+9cQr6EAosFeX+ZWA4i9u1e8P1jWvMkm+0vyfOWIS5n0WZJv10ZDYnW7/S1/cKJcb1
Bk099RbNObsq6dOUp3+gFfTNuUWv2LBZ2uFQauBdOsDyeHShB/EPFf1o/vUfoVFQlN1ZDmjdqohv
c5g2BY3i4lqGlNhl8Ym4XEZT+ywcYsMnELgwLacWdKz+d9ZpMkNXyxUzWdgZbfA7clFbApMoJdBR
eVWcSHnSgI0CBTeU4FMR1S6dwd9LU+yFdaXdtZ+a5aHeyU+yK0Md599gEVt5+II7tEKjy+jThVEr
PEIA5hWChDGW8r8Uu245/0f7GkpXnSgc6N/Gb/+HW5r5uufsrt3p3FP1RO5cBmj1yUv3gHmgwnYh
hsVIOgVKwW1o65lGYWqWa8A8WR98ZphgKbPhXvShKUZkj8oNe3PWJGGpEtCIA/Lojk3gxlPYFUef
efESPLbN9HDC7swAa6Ry3lrO0/a/EKzDPV1sqo+7qo1OdYVEWe/I4tkSKBIsu/GhpSqgolqDmhwh
kiY0IWtQQgY9dBUy8TdPyuhYOgAfBKPH0T5i4OVTrLttVZaBTuu5QVJ1VfLcYbpeiVmRwdZ9pN/l
VCISX4p9xBWr/Qs+IN3Me/l7FBT9LQ/OSTFU7jPdU/+3L+UCa2JwKPjJyp9vcxc6iQJC9b8LHq02
Ac+ZqIVf6qbLNA7ZRfHKSnWth2qcxq0KWOTzCd8WHYoUJthq5jG+d8wvQds5vOLYSL9Sdlg/shaJ
ZWWX3WiYknwsKDJ3c4Fx1y8vZRcgoJ89Yxz4F1lAciZhNBK5aC1xSAAHCXxy0w9ALfVD0rN0PMT4
yg1kM0e7nwRoBfSHLRwOvvjbloDXWtqjy4dnWQ0M1EsXzggrcDOHoZN8fUuhEwmOIFDnoyMP2Jgd
8QA+jn2n6W7kZcf1cG7YSYDZxmkOHLmf1aFmxciMrPMOjxi2P79xO3C2K2o/jqzYg2VNVpVmAf9U
Pl9JBdBRs6k2oEgVb/H3yAfyCt1cm8UfeEJGv/SU2Svpz2IkKpQ0p19D+WO4FgvSE1fJwVF9wbAT
gYpx0XRPlWTDri0jhPQQiZ6WrT0Lf933c9obh+iReEXaR2EML4caVb34a6fdTg2n75LvgvHvMbRa
oFqsT9GyBV6/lA0Q9qPsS/vBmPQqfWQ5O8z2WSEQyItfjpa6M9/1XXUSTw7vowD/3CE9N8ZPoySl
IFbm6hv1OCIv7uJ0iFyOe/CnM9U4oC2X2ZQNPbuwx5ihLpeUvhCyhH1izdLLMSj1NABi/fRMTxOt
eS8E7U63KNo6Lp9TGiSB9g2dPK0jx+fcpq9pnGb9xaGt7JtfNh6ux7gUQjjl9mpgqonqFJpylauS
ik1dwOqeRTdnn3WjP5T8HIEVjxMoGKJT9TqboduZcM6PSOBacD+nac6hVGfKx9WhoisWS5xIJHQK
T+R+SRc79d0Ty2k4HkuVAmNQQxNJ9D2WHI37UwiovtjbmonWwOy+BaHzhgMiY0rI/EdEEvUc5kwc
QIwhzYgpPj8qfTG9zRbCS6X8+jDIgcBugP4ZBT1FKxiFoZRA7VhUvAU0jQkaOLonOuLk9/hyUcIu
LzD1SbV8C1p1D6bSzZOgydtUAo8clmoKJwjAc/Mcj+unaWbzBON/uvLlqylXS5NNJzKIDzIVyrbK
jizhSPtyt2T/Sa4c+8xPcA/QHLHfclK5/FDZ5Cv/40863LMGfzocMrCu+idjG37GeeqGzcNlwBL3
QMvTCry3CjottGGLUskOWhOliafRjsmTVQUNxiMityZlZtvmvnGT6Km5pEQ/HNWu+S1w/5YpopOR
OujRGYSSy2JQuevDYIwYMjkDBC64w6yEfG4HY6jlEuV8moEO3xNWCdyg+Ds+sfyy8HKPaSBfbOL7
hVDSO2DajwOFv0E2uEcrMnjg8CyxD4motuAXcu8o0zJHNLujlOvjUuCO1R0Oe+i6tGoAvDL23Mm0
QtfqU91I26C25PSFFP0l4NCBsglocxJtkP9yYfK+v88tNznekGCnO62DJ521nlxLwBHXIkf6FYFI
hZ0y3gcSEb1dnOO1FwuS4enSmDCGRHiu5PJqQaKtgBev1nn72hAABe5LTnMAwM5hibZ34bAFlk8H
ugax79pt6xyYjxQAKB9TPxWOvJBX3oa3OXrjLCgshU87nnQEbUDx7hFAkWloVXWzot7CUgQ4nCrP
fgWhA+Kkpyp01r7z7HFnPVZs386FYT9guYt1Q2PsztS8NF+DHKcnArCBEcyMMd6IZCYjOesOGH1P
TUdNgqyxkTIL06yDqSlktiUJltm90A6ML2VKaIJbvQisQl+M6TltI5un1NJaQzALeBjb9/gFJg5c
4R8VodAU78F/c9OTgMxyuqdtdV4KwQ9m4xd2dm3zFn5mvuOjYyCfMO5XoRgAjyb7D0UGNcgfirFR
Dp8hcNYPBzGaVNPUl46gc0pZEO4rjTMXOYGGbaqIb4cokBCAtrPBtphH4j8h24jo+nBqPeIlaMSd
DvNkSMnLxBPK4M9wqNL9LLEX3H65EGtN0SdiA0PKyFlZ1tQvsVpR68PC/LtbWstQX8fOMSRJ5QT8
FPZHTPV4HbQHPxtSG3Zd2mPpfksltxpPMaKt1WPmsEjMS7/Hhlqa7gAkXuDZ3reLDhnaFog7hGmk
9Nsm/r6r2d3BAYIiEBGmCKeS82rVEM8de0b2OmDfsJ4+r0VZYzhtaVgF3qXbmtA8/gsGi8tFxFC3
aljecwpVyKjuIT1Gi7FCtKjduMb5ajdYYD1PBHGQ9sJvGnO+Pv2h+2ED9jmBjeh4wU4KCYflH3Sf
z0AgMw97zoUKRgDWMgiDdNHfRMcQW2aRjCSjrJX5u1bDLfUS6r30u2079wi0VL1qjcgyvi0hq/F2
QzgNYPRgu4e2BN0m597ANSC/wE5IwG28ANU7D20IKhPCfZJtGRvZ5qkjPx1WwNijBGDGoQG/JC3f
ZJ9G8qG2YdoChoFNMEdK2JKvxkWAwNnpRPjUOZCaR44iVHLVQXURj5HQRZbjcnoxXT3hrFrZDdr6
CSTPy91eiQPzgoIa58Db5OkMiwU8B94PyJTj8ZIFXdjacp0Q9zcYSqtB+XgDSzY7MA0EdVAN14Mp
6Grm6twi0QxREDrelvmuCerL0ywgsbZ28MRzeIDoCu/rP/7Ukg+A79XhmPBQBs/RwfmJGBaEjf0P
AmjMwZ7Jma3ezYCvrgCbu9j4HMECTiXAAjtNOEShZMQW2VHxLgfRpt+rZtSfyJCUDLamLwxkjGMq
ttsKlauoFT9G/s1OptCUL/A3F50badSkAE+xrZQzAGUmEC/7+k88C9o45o2YD2f23BPy36UcX20M
bJM3dqubyAHBs2FlNd5eZIi2Qyh4gaMjnnolov9fw3bYQhJ1/fSDctjrtHvXQSz6VxCP+83ZPhc8
ouFzaiHvcVoTFRf2tNCKK+22q5k/CoXbK3VYb/5JMSHPRqH8z6Ekmdqoxs1T1G2ot3VY64qusTJG
7EjRLP88VsIxRUto8ZIyoWPP2M/2R5nFNr/ebCitD2LJ1COjOWDiWLhA2tuNGVkG9R5HTbHmnS5k
L4KlhFkIIv4s3W9GC11nXVC8UOC029AFy0cEqiUzkhFM3Vyt7PttxkgI1HCe7O/Ayot8Utrn0FC9
QlmiYSmF+8RJpen3awIcBAvZUZ8LYODojRSp6QFYm4tWOIEd1LssBJvmgS6ASj58of0l8sscONJP
Jd0XECv1eGnarfvu6jbuT/7zJJT1GT5heTVFJ5snCUQcEFHR/dCLCO3eH8NNRTMguxm87k1WEPrb
lNwjcmpvZtBmpcJS/kmMemouPMk+PYhJLnaLYIZOhaDVQHRwA/kxfeJKRu2AdanPKCa+nAt0w7We
YnjfnuFHhOJ9HQxkQN9pmz9AZlY4r+Emja3W/KmTDsr53gbkgCuisAF4pDiCQBvMxjzMpsYCd81A
gnqncw9E3to3W0kQYVsan0LmKQJQOUqVKhiaaQyATErgfPbzJ8Q4g8YyfKr1RqDZ/a6uX3ijmpTz
b6+qt+Tm+ddtAT+XRd+6BPaQCipYCp+d8hdeN/YcrEwO2+xP0LfrW192u6z31WF9U70O3kfLe2O5
7F4jGpIL83xv1N54ac1Oi/Hx/sFfdsE9W9/FkZzMWMWU7/wDAkp23MO1mOhQexETg02qGn6tdaYt
HQYX2ax0SaAcEWEWU9ps+nCCbLVI8OC0vI0+wQC9uBbxbr5q/3iRoGnYwplU2rCNST95As0omi9k
VatHz0Ttp9QbrevZlp7FPuI2a8A8SgtPZnzaFoiFQEeha7MT6fRwjdGpQVV8JdUvTWn4RrIoGNMc
6VbIFIHtQrV6NrWyQVwydjdtDMK8cYRaHDDoPVXgrRZST5UxazYhXpXgasmuJRcJCtFv3kXLbA1Q
cdX2c3ea01TunzoirhcwKHi8wj9lJWL72Yjjlo+7JQIoAao33rSgw40FqYDwBHw8wIT1pRq+3n7R
dgY6KJbxQsdm/Lo5ew7XLsYLdpSRcpSu4XsEnyrqskmmcjfjon1DCuF+684hfBrwKblz5isQUd0G
mOsWhvC2Uw5hFij9a5TLImhiCoXuXhR6lThbdu21BRG7VCG+3jv6d4I3HoNOLOnUOLrAOfTCWree
wWXdsN94Fpec39wfaMdTARE5ik28kbyzZIxDmaUnxreL3Nx5hfkMQVeiZ226GYq6SMEtOCGrmXsG
JfarPl5OlHWBc+xskeUyY6EP8MyMpCjsKsYN0P8IzRGizyw4aVqne9IOopfguhytSS0VpFPuVWwH
lFzjX9TX34TjkGTwxfeuOu4MAUAEcD2jo4vi0ixmqekwC7fWfrlW2DJjs91cLVNcE9KEYNByL47g
zHJI2p9fDsk+YdygpcGJdPEYyJmA25FcO6pL8SFxUupxTbtbGSCRJ0bjz3ZozgalO1vvP8gQPEF4
1qlYmGYY/XgG6cTd6EYLyZKusW28bw+ostK7HCYBNj2SfDV7FEQooeSd17DMh+9VEkVMdGd8DzjO
3F/HpNxemJ6b8dav+RWJDcpI5lCdfygKsTIeGACPl+8y5g9dsp8Fdd2U7lbmv9XCIm/kAJlLizzE
S06OoX21qQOliczuLOM4tbCpnnc8MEq/G7QF74CL58E/0E8kFFNc8xs3VM8kA60dPW9LP+eG/0Bo
+d+94T1ZPwBJczqG55nCEUiIC0XZAUVI/ZU/oXYerBi8qASJ/hxSv277dLgKtAr/hpSi+h4rK5fI
NHLN8miJ9xsOZ+607iOVoDZeEl7mRqTpGGRQTfeI6J0fAQ/vh4+ztzw62JbbaSMeGSqDGX9SZV5e
vysjevFhoi4wYGKjhCyVN0OXPvBCmWNUGf/+/6LF93ZSclviiDa9+A/UQjakWanOabi+e9eVuvly
sKbrViX4fk3XWhu/Mw5MStIsf6Bxsq5xC63s1+Oc7ub8q3gW2wPbZZjcXB6LLTrsVByXKG/5rIJi
B6ZLT5fS3LXJ/DVPA+fK67Gi4ozuzoESawa7zjUUVsTgwMwBTc4qkbbUubKwEjYirKim9vXB6CH3
Teb9YYbgXddLKmyT7uVAxAC36e1qYRDNamAQ2DdWtG2AaVOrsaoOxoKhLMB4w72Ju73o4J6TVFKQ
WKGeDSMqHeRuDLM4/m4q5blrSggyBEjhTUawTpJyeWw34eL09+/HwM2mzmkCqgGgQK2JSumqLgNs
S86373EGG8QwOe7AdyF3nOn1sEFuXKfArHfEpKEC1a+ytELOct396seWus5MLurB3MYmhfQcOTRd
OeYJZp4OyzP6r+/TkWZm4cEi4wfHORRK4r2Drul5lYitM67rFBYY7LhpLtyiRHQRbb4F1HYUXbJz
+ZmZa6DB7SuuRi1if7UHoO5x0qGUchYHKk2zAyCjOS1Ba+c7QNFjgq5bxhxu04pKPNFs+FtjelPV
P5gZ3YCx+zCb2kST/pXWCvz+geFjR6LCMU4LvjiekH4QNOmme6tmQxDNbPUjf2n0ncNBEeGg8UFC
lcEfLAhMcBBLXyyBFEL4L+aapv8XN40n0DqRZ8NZh0I+okCwnQexPMiuhsaoRnAalayM1R8kRneo
+tyXHmd7+7feLr8pn/p6yAUhssxe2PuN9yoKTAqvLNnu2shT3yTds/yH3cjEVKEZG8gSPBhfRfkO
CMNdNjBl1h380utYPF0UXEkDPhZ5JsYZjJ1dzX9Zh0qMdjH7G0my8nLb7AG9PE4XSua1hlr46M/d
kPwfufwe2MSoU6aosHtMcpxq7Ao+IzIX1gLsj/yxTubl69lAKqeVvyFWHS38U0ynjD+a+6bPiRxC
ADhC15UdcQBbG6dqscMmfcJteXKKAn1ZI4qxWwKM5ajYcGvOAJyUfLqBTM5u6xhmjVvdehAH7G83
AR4QdZYwAY0JmpUF8TpswplhXfVh8W6UaoYIAxJTYHP0n05e8YZHstsgZKdtnp0BFihzLDOPgRlK
VQ7HU6j5teaSZdwTHv0uFZaIv0IaVaAxRQtQJXQyF0OeozRUwzaqFtl2zqRQVk2no//ssQEjl2Xb
XFk0Brzq+GUSF5Z4EgBsQ1a9gr+Q3WVfZSl9DoVus6I2TNx9nUwBxojURzw2zp5k3MUVoAbS+zBX
htL0opJ1gcRP3lnyfE9e5RaOZzUbHfRqVEMRXzqvEVhHGvP3KgtvBF679OdeqZJOabfF4tYBTk6R
I3ff5OXChNGmIjU53iR7JwGm3xcOznZ8LLopmWbvNkhdx8yGvKHBjBK+qvPKI2/jHVpI/SFpp91V
i8Oex23VFxZCKNYmDJxMf2fm4hU3wZXT1I15JXmRyo9m/LSdNEvQMIsjzwzuKMr+2ru7R3yYWQxd
1DSMsBjaT6Fn87RRmJdUcb8lN/guYoYj2WLfY4yl5z9tLnR/lFn/F4xPiYqfgTfeHHkmZRDukS4r
ggp7mgG84mmi32UWY1WDEoKbNPwJnHffPlSXR2qj1TgzJB3ODL5oKFaAbCZ9T1Dynx0uC7br5OPN
w9wQqzY1q9cGtweikWuCbV/c0/4Mf0Qcq7VAzjS426FqKeb0QXWAHXYMz8ywJY/SJ+ZBiKAYWM8j
WsZLBlonzETR3/6ZFYHwl+uGbH357dJtAY6ZQ1xLw+t8Nv/THyhEpOSpzw4ki/fmoGWxL26P4CAV
+gQRdOWZXsCQ2LM94w1WmNpQhwOfb5SRhV7HtFygSymkiNFzMzG+w7zwUsBFUmBmv2PcPl4xEkM5
mzr9TIuEvF2q/7ahqr5p5aoLyDDdZOFgGml2tpENX0/xNe+zjs7dLNHxbQa8NjBmHTnNh7/WwTRz
RyU3H8xvcydpo296MoKFmnS/WlZCuMC0YOBa3VXnK81CqvutPfalQ/gdvtjBqIyP9Ws9cECC3gjP
38QMrhLbH6hhOuLMskE0RZqCensXNI5RIp4g62zuPBZqSDGLdoIRv7LIYIElnY2/S2Ga4dor6KuU
UkhottLnHkebZX8j94SwXaM+uSQ9YKyow1XfYQdtPfSq4U3v6cI7lPrJwenN/MIEbTQIzJ0Akjop
s8+bRygdhlFIPp4rqbCJUcVL5wWx/KHQw7zNeDYvcMJXgtEWPYzzzuTi9wlTx+ai3hSKjxblwgby
K0t2yu6Lb3umko/E+plaxo0RQTvg48LsEZ1OIdqZcHBBqcZo7qsEecJwa+rcXRVHgn8j+MUu0d2C
fr76Nyg2yuStTr+nQyzAxmj3wFsy75y8HEEykrhHd2EYBBItHTyrj0wReJfvCTYgOHuQZOFfVAj2
/uxEtCqScLuXkQZTwQ4XjBNLvUMSUGZRbyzLcp3LMVybac33XjcCYjEvF9wYbtwVYkxPwbD9AdX0
yqr5918QSheneAIskKRXschFXjJY/Tnd7MnXxsJBpJukC4K2J3fdbxY9bR4RTZ1pYbkJvW6cFLoC
vGyoAASTW170BbL9mA2TB3oZOGtfiCqYH27hv1b4HJ4ACBxz3Ex5QtCknNvPY3QGuJxxV+hMDCA7
LieS3FVxOvHMs2FHZWlTHEJZF0vPFn6I09ICF25iu9P4IQiw255Tc1CuQNVjqy+FJCe55Vi+ePKW
mx50sgm3Gz7Kz+MO6hwogVAGtpSJ+DERHlY29vYmE6JC6peuUpEIBHanH5DoFC2mDRAY0rrqPo8u
aikbqcVwLo6HAqYkp8foC3OcD2ci4A837MKZ4a4sweixsDGzIdW+EnINtBB/AUCXJW01N9kCaHgL
1b6WHZ0Kxy9nYiQtK9q3o0baJTrPJ5zud62MYFkQwD6cWoGC59X5bqG5A+913hXfuVcTCkq56fml
LNWrPg1L+hSOVC9P1h6zxLKy1s0JW0UPEEvDYdK22MKDgU9/8Zsxs8KIwNNn4xkeS7Bls/q+D6Rr
CyE9VEt/RiDEPePgF0zkcTgPTicVCwnY70q+3Wk4toCUmd8T54IZHeQOTpKjgJEBdJZ8iBuR8ef2
8YaPCh6uh9ZH64Ypv3v0f6Ta1MYtRtdqFvK/cEAla9mcQMZQhe+JQwe4r0ecm7+wgPK+HHGL8x/j
LiIZH2O2HXqfCRtTg9ySCIBNLzsilyK9PQiqeHLXDMB1GFbgp5AgEaxt7i4alk0BcWgXciRM3ECd
YJy+sU3Qrm9Hz7BN5aD8c/+v00vXg1XVbqkuwuP2nJAUZeZhqb9fpQff186as4vSmQoS8zsHxdtC
J8AB4/chz7a5lG7i86/YzMjN5BpY4RyRd6VQVYEvRbBreS+ta50Hu30SAxOrnpepOlmzlbV5uaqY
IPXusxlyaKGouOmgZ3kC4JPEcY+3mOx1xjuIwg8EW9fgAYqVKcXboYgrhT96v2F8doolHhoM2LJv
O1Hd7guOXNSRv7M5cNmvxAIG0aJT6rnxDjuMpcctFmCnLlymj5/a8DY5KV2RNzckJ2C2P3JAarby
S9EBOnbKmhUbDK4SXONEUziSHPcL01sir8EQ5EHq4ctl/MMTTNvRwC1nzt9CFfvW7gE4rKwmhwat
60qo8ziRnQw4Jb0i9X5E7PTkxEeT7UjgbijlflzdqvHw4V5eW9+DwtpEhrgaj8wsOG3Z+hYmIe8n
4YPqggIk7RIoupZP8RfM8gG1RKZdbVDxeGqsyaV7junMaPbLM4ACRPFdUqw6VTwViwBMeiTAJ1M0
WI8/n482Mj9gdoO5Td/snuX6xX3RYdL4rMK19Yxo9qC2jOxTthznwYdHua6eDCLi6KpR3/Oy/pOu
mXeKh414gPkyxtJS1ve1O8T8DhzYQswLCG85e/wFF41GN16lkDEQFwoQlz3JrSk8DVRNafK0T0jz
mWvcSJfv8Xcs/9P+1JEunwFwLs8HYMq1q9w/q8xIGwK6/B7yLrsHDYdAi2goElR8itXi/5opJG7V
YDfXUZsGyX87bHQRHkPdDnNPaGxn4pjhVdN1M5ZYoOgzg9QXroyqJtnOwobEPhs8aFHtqUYZUcRc
m4AcqZQK2PBE1pzbKVRc2sujx7DVnl3PeoMzt4ptid81EPM4CdB3TCqMrrEsSCX8hT7K609VBZsg
cPNMsUSE5ocakU11dokPQlrtbFi8JMujXgCxr4T+o7+uANdJolJrlshcYxQ5VSBaNSS4UcHWfwR7
JSAFP4fdCY3iUo7DCLyuiTvl3puAVbWSK/ByaBnEI5Ua64+o72964mN11ZWFD8QVMPDARFNxSFsI
eNZjZCMqlOOBGt3B2I+sNt3VfLKlmTKCCaidFwjUlpI4iclUvGnSHMGg4bokrvTPoZouOnRjmD6I
NtI/2yUILySTGdQNhBi3HZZ/ms3bTqalL/GVE7aCNiw08wKd+EqFnJQDdssUNmGLhEiV5yYQX8ry
mtkdxXiAhHubZxo86d4sT03nHRudd/BWkcjp07M3I8dUStFyA0lmqoGPcJUicivChNXvxN2tmg8c
u0PHcG/s43GUTqkmeukh0jTlcwF4kCB6McLg7caJcJ7Ck3ZAi8L1K6F7V7qm9IjEG5shI6hWWN6p
XHQZ+Nt8DtG1Kz7Mg9xtiux9lx23PFbOwU93YG9t7wb21xgXir8rNQpEiTs4fQRnnrhhu/wunV8P
CTRBKo7DSjByM6P//BwOIB+/Gi1xleGuMiQ031vI9M/5vZNfMMxpIqFb2rwDODRsPit66CDzpEVv
NKAIbhvAnp8FABTXNHh5xkfgjoDCEMA7BILXyZK6TWvTnxzwie1pzV/1IONXgscSAQySbLCbZE/S
7A0GS9JhIN+SytOynhWTEMZAcVwlx+NdGx+SboWv7FU/V5fj1iIm+ZMoKQbLq1dBjHyhUeIUhQ3t
6js+G0X06A62HQGqXTuJeuiIPpZDX7Ha4RMsfjJKShdvRPhSZp9c03pASG6+ic6NPisxzgM9hd0C
iNCyadC+JIKTp3AsmQhhY2TRAEQDEO0hvIGmm35IWo5FYDWerktfRSKNgnw5X/QfR7C4j2BTl7AE
8SkTDaBhI0dQQKRqnx4/WyYHePUGZBqwclvQYQClxsMaizosIPRjrLw7IrwYiZIKWokakzFPphkx
K9/s4MdECy3qBuImbfJJ37MzNZyWlDhNXn3HLcBRHs8kjt6UZ2UVkQ8Xyg/oKXhOerCnfaxBR3UA
Ap+u2O/op7iL3WL5j1bLsBfC0Orl+IszJm7ynUbcC0nAImZfu0dF0bBO7wMXm9+Zn7zG4lSGh3lN
Rs5pUcwoiDzEMiK76m7jViLZzo2NHZ7JpjG31YD4jagy7VkYX3gRSkqo20mDwYm1Xm11lWpJl9e4
G+me7bVj/2/D7NeXe2BvID8E2CTEYe17lARvK3gvY6RuWGb3zISrr+j9wW2uQuEYIFDyPSgGLrZW
FOxahRSjka/tWueBvbx8F7s1vXSg5+6IxmoJUDiTYJYy3/gwarLcbfIZ+Fy+9EZkBkVn/isZNLMR
av8BScMaGm/VsIkoaSGKDO+bj+NIWYtIMWgC17LBk+W8JBHJmw/EaGzTPJ1ujS6vzcgGKUAzbAcI
K1CoQsdzV/xTegIFOVKPG9Dl9L4mYx5msIFYCbemTyeEJISWr1jn0d5kprZG3YkrENbe4AkT7A/T
gP/YjExXmIVhnEYF7tL6hLHQlRy68m3ER7+Fod0rMb+CKcN3WF09H54lWvDUVMeEPlGB2+ZMiLV9
qlQ6NpRP1/Adpg+4HaESIC8EC7/32FSZKgEhzxTsmHl5CjjDZGhUawQbdpUy2NQmp7dtr7zSAqL5
pXX/O0xBX/MxFJJN762ezVKwFzaSXg7v1Dk5vPiS3K8FhmddODYuImVoPmnCiVz66O54rI6dKncE
w8YI/RDZdhPJOUZbk0t8qFRGS3XQku1J9TljcO2A6hWlD8v4TbSXqO1CLny//kOpfoogUFkBxI5s
CUlhTSH7nIFV1Ne+sW2Y2gGWiXBMvraE/Zs/CIc5tWnBACMYtH98sjpId3emd5qwZ4uDaRjzOLuN
xldCgW98zQcwHsrfqyzF3BNwySdkFC1f9CUMZR+p2UaGuASY5o93IzIX8rMDROcnUe9zjRR7zQ/2
gH1xGYmWbodN8aw1jgjaLuAkVeFEp743gPYxLgTRCD52wr5CKapbVHNv+5mrjwCOmv8ZNfRUpOFs
2HR+oCZu+i8OYDILvnu+pwyvWd6Nkzsexu4S+ZnlEAMDUlCww0qyIhVlZWmYDYAiH1srJvHd5P93
sqlHmUB9rBtKXZpchjyhkc1XLfkUp6yyg/4U0AAYr2JN7yYN8qSHp5C58bb0eIe7NkKRuc9y71/3
9+c309HLfifCqGU5E4NjV+7GAvNQ5EjBVkezr3pLUU+wH8QPx+PmS8tkggRsd4n3Frrg6Jm45bh+
fS8N8Fv1hfqFSs0VIZAZWA2keT4RAzz1IHcxUkTKV95yVIpfDE7sviT84yPdOsbYTjArjb+0y3Bu
dwH9zA1KQ8zFbJRJD4WvklLBFhjCrLS9shwm6UqUDnkNVatT4VKxFVXH65Tllac6YhGNkpBBB6wR
Tjw3IDIBmckG+NKatjLoHIgGs1DclzElZMR7swLi9Fjt4TnS97aE+ykdjR9TTgFdRdVZaDJWY8bk
1l+B4bQ1MLc+Wtw+tMoJkc7AOF9TQL0gAjskZ3seMMdDLM59rh9gZmZW6tRNSXHUQRj8IrPMOUtw
pMxVvt3LmumjjAugqXLFwRWJCgHExrWxK2puUz4MEDLumqO0BSOE4f6D3aBEnXo1vHWjfECnVIRq
7Ji5twbdSQ8WNDOst3Plyl0tpZCAGMOO1ubO18RIaJwezLhmvVxG18fOwR+R/qSSX92zDAimTscb
+onhQCyuZaGh/uuJ8/Ft0W2OliIN3JKVE3fCd++AfM/e9P3mROlHpqGL4COaaYwz7KVdBfdLPV1t
o+BGT0Jd3plDdITIvwtOdRuswsbgibMXsrM2VCFtjVT0XX3TucoX1uZnd5sap9FLeoMYoeXxfji4
XRMJs7eNDqa8+9Q90sLpni+lbiWwxjyQKNuLbWfJPFjBLAFuP370tud+cykH6/2svufzHs0rdzTX
VOh0AYppZ4yntJHfjwGfLbZ3W2bV3mRFCSERBkFhgg88lwW1FJ9rAsDhFxfaDoUvw+zolmYehYV/
pVBAiqKbOyHS3WzzXPlTBSHkq1i7ZUYj1fhc4uX7rQjwSeuItco6MS6wG345BvgwbKYJCKh2MMCC
ag2j2WvewViiYACN3qrAyufw/TRbtpWeNv8H+0qovdARHr8m1ib19e2+iK/cgbcJh+3ZNAsiceu/
+EtYqHyW1Y5w8bDSE9fSEwEEZM4TghAMHnECVrSA3ZjZIYCBSSYPPmqABKqUV4wlN7N0AlQLYaPY
zB975EkgFSpssT/who7fKcRSQjDNELS3zUOuqvR8SHbqWqnhRbKcNGbZ7h0hAP8AXDyO/paC9ZVU
cs/EKqPWWYxXJ+HUjKbAwi3em1YMQ8saFwkKaLAYf+hEkGICw5VAZj/vTpDrKV9ihahwLSyVib2S
LiXwlgx5uVlIKW+GKV4J9ImHd/WCNej6r4PfAa5hTHVS+B34n8d4ZPv8Z4CxuHP+ql/U5DoQhDB+
BJFEe7hEX5cWsfMwPlQj1dTLG6VbqKyrH1w5+vQ/WMB/fsED7Mq8qZ8eZxgEz7rn4fbeiOyaKhKV
N5sHTBKdSp8QfDS1sxTzDU/RuRkLj+LEwyraB+q3WugdKeKyass49Ncb9SfEdSdPvY6IJU2yimT+
DegYrNtocUIdZQTq3SZ1GrM6/cEFxLz6GfHtcpySQaHBrDolObjZ73dwVY1RBFJE74Pub39Z3JzE
J19N8Xhw1lQrDAjHnvmZ0SMwWPT+ejGV/y7u+uMDco/8RnC86ifvT4A0AVGMXcP22hAl7wxp2M/9
ytSTyKHusSQ3vtrUdTvNPU8aYkYPaTwN+u+LWtPp7+G2J+bD8Yqhlmsd5ku/+tWKudJiKI9wPN6F
P/bkhHYe+JGPI2YhPo2Ih/29LR2wZa6yFi2zR5WIpKiAJ1iKb/i+hf191XsYZIQ3MFrTpQgQ3kui
1j+h97Ca2rcx6FaqWxdbsO8kWlae/BRfA5BFIp5s0d2zIYO2DX4EGcdqrtKMju6Ng46UEmzITx7j
CKx2BngaR1cRAI5q4ZJ69Flzt/rCMBtJDLRFuNrw/B6wmTjBPV0tDBVeHhB/XKuTQkCFlEYa//n1
l9/MvMZeARc0Ym6jZT0GwhAZ+BaIb61ECmZJINNSmgGOwLIUFAvzkIKNVHMVfseP5OuvbndEAuQU
AsmFp4nrls2dSF8dK4/8cWE3ghSs4fIJa8mBGEQf0uj63hHv/isANnKE4csObMP08l0gi0FbotK9
zVkWBVb4h0Ta5fzgOwItgOVTl65BLQRH3QKwSaNJwZ+1UAfQu3qhTiyz8RzzweAQOK0NUdkX6/BV
0Vu1oNU4WmrT/0rstciHDEQreDgGPRC9JtMSWHqAslwlwWIecqT0WN1GVu3q4RIATV/aTjuig0WS
0l2Xy5LFg1HhWAA+c+3jYAWmgyyJlynKekUWEKbRVMgEj943y67zGg7LLgCaJG8yPLAmdWqRvTUA
al+BIVyxQDZo8VogobD2TNHerssjIZws1XVHUkn5MCWkm7NnK+6L91FctYak14FsDNAn1b4y71fN
1WX06nLk+opN4msN/tsb0px2jzUsdGg2wxKT8t34mwo5GRCbh4dYgOb0b3JCozAkTT5HgC4264g8
Qh2mwXVy72pdHNyGt5HFsJMFFnnt/wFGZVCCydfdb2WNQGyAOlcCxCR5aH2Fo0/Mnh08jtnclmId
dRcYibKvrtosTVchX0XCLVwH4lT/VvMjeSfqnkMap5u36IDo+6KwrYt0np6/hntYba7gcCdaN23i
EBEbRoDYGFEfz6UxxYkc2L/cy6nb+4jzSYwvzxaxm37Iw0zWmOMbKaycwpR1wxHnW+l/b9+zfPbZ
IIxUKQaFl+LG+kP3YzTEYArtqOvpVDE3u7id+t20ppO9347xITMedArMneW97uy39Zqycoiru/9a
PzhOTVbDNlJJYhWVLT8FZHhqey/YwN0fX9oQDQKJgns60TNA/GTPxpSsE8n8HN5L3gkkapsOvojs
H95LRSQCj9SyuKfI4bSSWzQbR4oCEwld0c+Ga4WFr01anesuu2F3W//eJxqCY+nlvWoDOW5VLJiL
73XnnOp8YV2BxDJPLejzhOtaeAFkG6eB8sNU16+JtmmolkMbbqf+xgTq1YnQhItX+yBDwi70zYuG
oTyLe2Pgvf3WgXr3CCpeV06PPm+K3wOMXya6FielhcT3ldSlkvG6Uzpkqus3hIDDzcc2mzh9ogr3
wgrxQwtPJ4HqeS4+57ri10PGbOUM56XKMAgRsIMcH3kna6rJOWUDYM4ugFLFBhHVGE47aISVlzM7
SciRnNtkn9PArAe+4hBJY2sNGP/dDcsGypb++h4xY4s+jwbtDngb+ofAoIf7mGoC8ZR5XyuriTZi
3yYiH1flHjc5jhHFPq6LSU6tddGebFJOlXkP6V93FOxcYtEpC23agB/qjJ1z8Vi2tOt+AIWrd7Ja
s2ib7KpjetWZoVVXkKk7MTdilfDVlCKCc8/1Aweh9Y5WoTXYWXAW2w+0c8Tde1ociPWMY1owSqUt
BtLcKLmSslEnHRJ175Lx5652c+Q+PywWvFnFCkPwVog3+u9t32tR1eAASSUUEBuusjMIzDKofCov
2W89G8luYAhpDyALeIJCTGQLi5EqqmqnYXOBDz0R33Tokv6BF1BVtmaT7Pi9YesddfJPPxlowpji
qgcvGzbsu3m1xRd5hDkCkKK3y+5fqghZonYbYQxu+D5Hh3+0W5rHQZranSbZ1jbjr0MSU0GO2BcX
AHSQ+Gf5VtekJsp4vyuUUbqYwI3UZ2VzadCBfPrgE06UP6XARNH3vi96oZI9Ts9wYf+kxB9dU/b8
00Cq3FoxAUvI2V5OERwGPWKK7bRLk4V9FMrhHCFCRL/KkFpSSI6tGgBgVsjRXKpG3dKl4DYSVlxo
ERthJVissBNYt3blcCGra4yl5E7RJtool8V+rOYkT2Wyi4OmZfgkUIIypa6f0XWWNNqql81sebKO
J1zsanO2ksFxA73GCDjllnsPn1lXy9UjDQaJtOzDxe0Grm+s1DggATPDOBZGrIRoyX8Kt/Eh57vW
xS3Q2tMbA8FhMqTu3dUz85E8AT7IG7kcb4eXtdP6cMlKGyvpNwyCpJJJsMCADXTw5OrnQlSwtyhG
Skazr7HZJfPBcfsmX7zXCffZA5GO8lR7p/Esy4uh56dJXE+LD/KCTBJIctc5oITJK1FbBKVlNHKx
FBkmkv4e1DEjd9tpsHVupxV0HH52ZJjPERIXK8SLlNhrmnW0TT2BahWEUEyoWeOCB+L4knndanm7
T0o0dmiAfbnIYmx6tZ0O5Ag16Fe9MZF3PJrNvBWegiBtapNFesYUcvg51tNFqEzE3pWNbzT1DSAG
rd6ei+OSLy25jzdnlOImZ5qRN0BwZVd/mRcuwkPEM6tyCPk4NXb2N2a+vt3/2RUlpeGM576LfvB4
Mgxq5Vg6kswPRqxjmo8gE/6bea8RA0+zUmgD9sShtu9hpXPHkxCg0gaS7QWkwPzpVCVDlhPgmMfc
4R13JekqaPjelznRimpiESdsiP4/hY6NMxKrSkJx54La/gXsL7K1o5zZOVjM/L0VeOmp6RlmKGmV
tVpU1JBGXyZz0ed3ETvERS3Gf8CQL9XLkb/4XCcwBlOi6dSbaXWP3S2qU4a+t7ePmzWwexqxqz9V
atdaqdxJWfFuyr1l9iMYuQBqOjmNGYvsLYeVWOsmLcnAXG8bIVSwhPd6EGZaX3v/Bg8eYFy7EDI4
41f956CAzbsqey2OFiSXJ1fYlmbmP39UJS1RRFXlfqNdihiM9qqBEyVpFxKHRyXup7FBkJdxaLnw
/27vNmsdJuc7My+ZqHphsc3T69YYUX+a8cNYUregXBDbbcgYmFIcotu0LUg5Ocb8RAqLmYo2h6fC
ueJOVvudn9emHuMsuv7fQnFixBkK3Tx/SN5WZoBB2ma7SmY36JX3xC4DSfH2qDgP37v4WVxgE5cQ
njL4+/In5c6h7GokNsfCVftbWlIKNMRrDA4TVzyBvBBVHEJ2BJ8pHh9hUgON+MEDSslNMoesX3pt
tUBZG40/SF1ggnlpKMlGumkhnGJ1KBErmIZYhZp6PpSRGzHtaIkjM3PqYrFJcFbdg2zyeJ9Xe1fy
ARdykgYcK9Xno+o2zpHsG+1BSeJvTdzWqFPZUpyYUjUImnKvY4xTj2G8j0lCLiXI2YLHmwDDRRWC
Ni3w+tmK89/JiexLiBc92Y1wW7IbPPj2EV0ajHpworCWwIMyTkA+DzpvtaF06xBCGMhRH2m3ibX+
k345Ku5RqrfyDO3aE+H/DA5eoGwmRou//p2DF2eJ8K5hvPBzgbdMTyy2JwXE/R1pjCMwpKwgdxUM
VXhHTGG5wh/YCqZ6grionaHJpxNcwin46hxR4PQ93i33O9jC6vMQB7QFBvf2gxka2AAMkqDHrgWx
qJ82cmvKN5qLd2V0UPVX+izd2VGeYwoPyBEsa8KDUgkTzmdxiHazVLpb0MeGDaZ+hS+U6L82dcop
1MHjx2jg+DjSfwJ2jMGy/YuVl31KFSavmHgZcTmfcGrLu+gmajLoGUjz51cSeGMlKhKE2VkLSu45
y932rECvNTPhBBMBaOdHxeFI3kyBMg8BOScKqqRzocGWUin80Wed3vsDtD9aWTzHkBBQH4qsNw29
4PuW2Oxz9MatxGqloiRooVbBVW4+E/bo4RdGjqPrr2hQxmbz9B0IPA30piH4UruOU2gA2JS9g3sN
+zZPVdHOPjpqh1cWVHHa4QZiAB4OnnfjHwcrXXDz73L3ZdrSo73XEf2FZys5bEm/wUhDF3rs07ky
o1pGTFIS1xG4bqjuMZxk786+Lefk7gW7/oFMjeQ+LKWnh8zxqAX8D8sLLKPtXDvR8PVSNDcbH2+i
1Ei7nsaCurP14W0xO3LkJbOL/zq2FrFiIjuYkaQM/NecMRJWerQSwELDEeVGRhs7aockZ791q8LS
DAOKAiQwND/PwqdjVHi4DdOtdEhix94XDlp2bzAuJGM8tz6plmPDWzR4Vp1ATXWlLtEbk77/rrBi
zGRQeptw1XG9ogEKfnYx6wHPyyoCWUnAf4pr8ti5kWzU7aSXRhWH9dLK7UxBpxpa5Zg9LdJHTzqO
wK24C5sAXR/SBPLmNpI6+wTA2JPTjXwfu7U7MwGZfCtmNeBh8gsAQnW4FuCu6jUvvDRMiytnwhBN
pBqLCuY9etsnR0JEt5djmFyA2o5W9SJE1t2hdxWoxpN2SHBrFwk1W4Lih8DfnMmDzFgt8zUxVPmE
KXSqx09X5hqSwgBMDun52eki2DgGjFx2RwkeeRhSe9d+jq2iUG6cupVNiMHT/jcqxywdWdAkzsZV
p1JfR1eIohCykENanasY3qwq7hiaSauerFRO79duib4bgH/zZOKJHN8KOGfGgUI/ldiD5nXvpXJa
1E/NPVkt2XlyAXuaRMJb+mtH5WlqikIu+WFxwnrw5Uygsm/IjKKqpIGB7m/nuu0h6so1J5Ctai78
rzgMeV1Kket0UW8GXZ9lkN2FQkA8E4lm+CBIusT+a/VkXAuNaNRFiG9eK1tMIMNUJzomHejGAG/e
6ZHFAjX2AuiZ1WAuck0yTshduxas0lE0gAmmtSyqFayjXUZLJo83bKtirbKhcbbEDO2lKDZhqR55
pvOEUNiRBagpn2brJ1UbxYN7wB8CauQSNJ5/W7aJYQwoP9lZCg1anagsyqFCtGPr7EifyjBH/Qgq
LuG/S5O7wYYDpoq443xdp3k1iNS54J2oYvWT3V3Goid0B4Lt6vnCneiPi/H43X9bmv1XlAzispMw
kiPo5z9o/iZoMraNgoIF1LoAhOA3SqzfASJnTy6lEWuxLujPdYOYP0H2lu0IaNoSDIiPyJw4zDWA
A41v5h7zXdvh6ZWLSnrk4+75DjO/MnhU/uoNnzu3o9ZIyHxXrpAMfWYJ2Mq5FllJtcGaNbYQhxqJ
c1VKtLO7UWEvH9GBP892mF3E/0iX/zn+NuwQpW1GR0A4rVo8kT70ZbWNQ6YGdxwZPrp7OOG40+7e
qM9d/qXN+R+tV/hWRjd/kwl3OOn75r6EokG+GDuTchOwLm7Pb9bKY8UvUVf6sSbZ8pyGozjpDOD+
sq/sDyvjrOoLz1OUtW6znsBehXHA+6Ttau9GK2xUG0XqYuLFwZPhJ+GjEZKWzvox2dAKSUtHRkE1
M3TzCxANL3C3axHXiv7a4yQot+RVKjfXTs0RlKgUK1mawlH6i7F72ZZ82VrrAb9GOMNmnDLErJ8G
yR/P+nMBmzvDC5ZiJPe3gay8tejUf01PfXPj86JX3ZAVG26IHdy668IJJLAPVauFO8NkaRdHseIU
2gz7mcTxy+2mNSyxDijo0+4IGDZ+U3Svo0rIgNj7g/bqcBBNDQvqySlIbzu+e5+nyr5ADE+2QETG
LZRixY/rFK4S8741N0FCHaXh9vVjVju7dcRoG+N7Ir2XxpQkEI4+lj5rVBW1kp0hzGPWOcAoB8wu
elIPq2bJn3Y/Lhsf7Vk1vSCrD++CiZiqfOrR7NqN5M2/aqmK0jp4Mf1X40IQKxGRI8mqr6afKgQA
V9zpwi55OW6UFmABZjyg6KUnZkVlXCkL/jldSB1JqsfLVDZD8x7nnOcLAesn/vzkaiNuDiEKei8j
h3bYfD1qS9xpfjtus07uz/05dFSedHIs3jXeywQiwr518nVrh187hYQ2c0xrD4nTfJisWV6PLlgl
ihi6iK4qpCq/JwE9kDksOCUzvGUI2fwmRU+5G8WdxdJYey0+cHeL6oK60U3P8UXuGTzcV1F6ITbI
jmPlW/1d8IiDJo09OOqi06FLRt2PYzgetVTseTBnU00eLgiQlGaxnfOe+NBFTBnyxjfURO7K2Gqh
2O7+4G7JVjuSjdkiJ9Bs3er7GTCh5tNrYym4+cW+ZnMwxgDnpGAEN7PsskrUOBZtjG0WiQuv0BIx
sDh6TeVWIn5wwA9Ho3wgqaqwMNAwQwaB+Np9MfLxYB7Jtwjrc5rY2bCZKEOhofP61Sx1yYAqLxNw
a/mMb0xKMTnHMfkH8z71TfubHO+ucjWut6Qp45ZwFXrZwu5oHWUGuQVPzrnBBJK6CE8EoBycvgB3
XbWURsk1PSxgk5HlBxJH7ZHEbMm0X75lblkH+7iS8L+fH023KXv+xfdeqUA1AYmg9yQY1Wg+KV5E
xfMiusKbNxI2OC+Ik5Mm4AL2Z35IhbKoZIvZefUaO4DTnSeBRBS3lSENPr2qgsJVfYdu2qL0rtYa
FOk7eEfgm9MuPrxcVXDOb35Ll0nGVGExmvXupBTBzQ1cPoZe6ITHsIM+AKeu6LX+i2sNhPAphAko
StOzOjKK0MP7miD/pIvg8Vpy3LMTr+zpLozJf5+ZZhZPPOOtWzUcjRCj1aRnPKyKHaFnwvTZyfUw
ab9WZkaYhmCdxjT9CMzyfvDnkewijMv+JtHaiDVbSBgdnFV9qPkji53R/0SpLTyFI0j/lxRV6YLq
P4DSM3IHOo4+jOAmuBKwDZceKH2ewfliGrC6nNqIttsQTZ9L7As6OKCyD8GYZ3PRJ/pv96TpYXVL
n0zAGfGWHmeST3GvQP3gshGbj0hNqqSGYCzCrEEAKMUgMHa+36iFFmaHjVhJkQBh8fuXbn20OzwZ
D1rIMXXiakuoBe8T/dJ8No55NQBhRnEAPDbO6/kGpWpfcUnNyNnSU0QnE7uxniFOEdTsvKrkermE
nmkcZo/gFEO3/ZvJs+vcFFkZbR6nGynrquevI+b7Vxhvu7ZKxospZqgZG6RCsqIFlpVo2AfX9b67
kcZ21+kEUqnVXqJ/HaBCiToaIaz4vOA1nLjLuT+OG1qyeoeAhRhTRi5MtQ2WtgytbzHZiSjq7kFC
0CvDDhpC2v4KtSO79iGwkZF3z0OSm/8CFblWe/hHswBkEOhKqOq80wSFE5XnufcqKMAx9a7NGW5t
z2VxFbpRF3hfhIcY8n7f44uGEjqaVdTDWD/FNn+gRBcU2WOEfYYPrUzFC+DDLrY1Wv9TGpVQcJse
V94vdTdoHi+21jE0WGVbWJL98VT3beUiSyIG3zC6V5vOBXqnFI3jnMRRgy9gNsi6+XOa5c8mjZ9r
ytpFKRJgFIRce9+OZgIDyCXXIDJYfKRRrakF7AaCFKcFYV/dd9KL2k+VGhJjtfqVbxciD0AXTDrz
vr48j2lxrn3wO1uavuPnsc4wygJLcT8E/+0pTj4i52r9R/5+gJ8mxkSNE7JcBzNNEdwtoZZJ6C3n
tFk6PrFMOraV8OYwa3rU+RxsCX20owNlD8qJ3CyBaVmdJNWWAGAA8MQk18iP5XYWSV90FKsJhTz/
uUeE/Fu5thCRy5SLtQKYYbt4gY4B0emaOi2ndi4C13pzst90ofTggsYjoqQVTJmqkz1Ni/6gg+YM
e4ud9T1MRIUk6+P9+TaO/49EVJS4/3bIwP3o2LfFc/v9dpMPr9qiUvnRCUpL/FDvuEsLNsP6ae3V
cFLe/m87QqLp1wK6/KT53hr3HQq8jv4FMeGNDUp02NVDMewgbxJ6xGOxpMk7KiJym8yE141ZmrS/
u6U0fLXCE2PDaw8C7sC/93bzKm2B4gmR+hKAbDF0PU24v06SMhIEy2vST6ncBtcggSI87nV1L4WC
B5/PTwc9sfj3e5FQgPfwx+D5j7JmfGFHe2h1xNp8OVlnXG/8T0HZCwkgXsMhs99RLUuuVzvVipyz
GeDNkjJOPgOM1nqihFRWZu0MF6K0tPYOiJU4gvOuqxOOCxYQ8Nn4k83pnfcpQyYiGFWl1oDDXMKn
s1W0atbRtbAooF9kK6PJlqK5KWkBFVg4Z3gYr+yTbeo9J8QKHtc3593bGrFjg1AQDL9CR3M4I2Kw
86euSOmLW3vVKgoMJqtjPlIvJ/O+jcB/kKlmbEikcX8W7SLY8/OHgy4Wq4uuyKN68vCeU51+LZ7q
rxM9sgVmKtO1taZadua0IgCRXxi82Fg75N6MtfzpzscHjV0vEJOehszyx/Wv98s4colLPburAKXn
eTb1FxTPc69xjC9Z9tqFcixUmiiAg0T4ZJvOJJ3Cu3NyTHcZD7pnYOnb64lY0+MBjxWI2a4nSRWV
/y16BPR40vDJvHlCkmQcSaFJIEBYOcnSv8kxqXvyzdWBKLmXobepqCTEKmUotgC6fLVuRdOrxPP8
66aTzW3C58PWSZco4LO7A278OOlkFEDrSUM6/L23MKOP8PXsHlwiK9UG1xx2tHabdhznqV8DDMat
YxKVkLkF5ec94MabHF+y1Wl+6i4PiwYiSpkrX5/3ZUptR7hREhOQLLfX/V2JVc4jMBX1WTbd5CnW
oZW4cOwV2Rz9MKieMCF29/ZfxEk+kmEy/kBTpLRSt/LerDz6b/vXpRqMnvzg2Z91JLz/0DgDZ5Mc
eA6mOqHLqLNTioJw4HjqwJQH7+6qjBeqe2hM5G9mHIPafkBggX1PmsEck+kmexo+ZEcSlYmrjbj6
rS3eqD1e4UmHZ4bbzrTp9qiLGSdwgESL0qxM7Rpt6rUXf6vtJVs4vCoTQcBeGSN3tylnzUTzxYk7
zEM4d2xw9CoETbcS01GrnlJLt7XAhIi1l2bq21CVqGUQA5k/oddhZaJeAaN7ZXt2Or321P/+dWiq
2uL9G6P65Reqntwn9F8Azgw/uH2EDIPOlZw0i55I4EQ1CJVwghfi5+r/B+iHbrGzV21hz7BPreel
iKlfYsMh32e0Fmsre3kkMelSpDOyaJXkNWLIRnL+pqBSc0kA87TMe2QzA6Sh65Zeavdwv3YcrXEt
oi74oIZHaXMpXTVwHSFVlopyba861H1vsLx2WqE6gqPX66K8clVGDjQ8MQy7g0/n30Sp3jT3msJx
Tt41rwFHl3bY29jAUUwr/3lTqzHEr4oXykoo39rUUmGMiILke+fn4+sxx5r50hqQ1QKVnq3F8QeY
Qa9tFkDdiJEYSUMjeu5sa4gpZ7psZKhHcillPj+z/ZYEqH9g9hNiQfk8C+pf71mjeB10fX2VSRGH
8PcvkwYxV45nL6YG9vhYhaiTEibVgaH/TURoSJ6Nhr/+KRNqNqOXljMcSFmLmtvPUaClbPYUKoAE
Jr9C8YcpHjmNYkxo30v7Wgx876sU2xd9XWHhaIcB8xE0MYRe9XVEtbfojJRaFrOt7jUkmSJupOom
bM2lyp6n3P07uK7RE/ORzQP63viwdmoxk/Mq53MSNY8Yxs1weGGIIOz/c9XXjvIZ9RhsrjsdzMft
6DxnoYx/E1YEf+6P8v6SsPC7gAIEcjk/+rpjvtJGyNv4gfUM8ncF025Ok+nPQADv4DUV86jHwz3w
HZuACxNQfOmZ7ape8KPaGvH6w5vR4dEu79YI/luL6VcpYhYKNFf0YKU2kIbbtCZm198vpu03cL0S
etwfFZb4r0xV2vqX5Ge4SudzL18Wg04yqWVMD3dOBVcuqClIGSwQxHPwfjqPBsE5OQIKL08xPCBe
NzPjY9rdK3te5ZcZ4/mqUAtirPR8XkL+C4og3oyl8n38oxUdPHSa5/CO9HiW5j5ZkOyhQST+gw/p
Nq/uUorxw+Ll6YLbkB1K6gwYBZCCY/64kg/oX1lPfgRERDNHgmR69WqKEkGnyAeRVyk+1XL3qYmp
rhkHDgXsoaBNfX5WjzsmW6EjZA8pZLk4SeF4dBlzxU+Nb6h8R+eOpU6jhbkvnXI766K9ppSWM0Od
wA3hyMgmyaX4gSgTVhJZiRtH3ICCqymlPWzKeqDzIkSvFeW8YycLZe8AAuok/TcadOcZlZs2WYyp
XXzkOTrQdmsveaSFkMIAVSJe8GadcJgL+OgX+o281WfaoYXOMLBIWh0mH+8ZmrvJExkkjN3mw3kl
AxzoQEGWwgjrIaH5EBYTDTiKxt/GeUhgQrPD8IRHuvAW/CfvYYzBn34FN1Rodi9W7FsAh87JuXHX
ScpuAmeLGTwjBaYQuRKaDDGB0VUfmaA9bgc1F7O2FbTw2k2t8ZLf216hoWBMpM2cmGG1e0BmkdMp
yUIiAI9IEfBZQCjMUBxRYS8HMvWzlc2+vnrkYY/4f1Y4mMzWjkomHLaCByAd166tCeIk9Woe1c1Y
cIyhqwLqgj0WQg2yF5n0f3nZcv+4Qwk4I+Htd7X1Qhn6QlpgmSY3IVZG9rV1Rg4pvBH3ArXr6m9n
ODgP+3jMMuJQao2yc+91CrOd4VaFqs6pE9gK45gVO6LSjqM+C6yFTs5YRY45MOJJBjPLUNVQ7bju
KaejXEaWK3xxDEEUcVMxgaDQZKCab6v7GMdAWF8/7v2Ov59WMViVkkCzwnRmgadRLHYqfFLWShLi
VAeyLSqvTUqOKOBmDk7Ocu8fVMyhnTL+sa/KJIR1g8ktlNhFGRL456LHNiRpOqE/x9TD4uSlhRyw
GDcyyyk4hbNk+wBw1vz0nFEvr4Rg6sVo3dLzyL8rklxOFLLkLJl/ahqRT851hpUChF+JGhi6KhCp
QCxyOKOSx6JGr3Z5PxN+ENSijYFPs6i6Ydr4S+doNeoN8WO/t66Rx3SpB3Z8ZDP3FAh19kzR6bbs
QScM/gJb8oaeQo8eYadjn2PAWw7FCCSherK/LH+FDyX7Gx0LhR7HxnHvvEvy9ceuNa97AAtXcMUD
oeRnB0tmLl9ILZuAynrsajooVnWH0B+XfZphGb61cntJPkM2nOyRAom2aeL2QQKULEvLFRZfXxmH
Gg5XyZKpVKPz9EKgXsFXAEVs87D0n3WUM/EPXY3HTxg9P8IV8BarKUYzPOq/HUsHypySyT6q7kFa
zggSiPowb3M5OocJq+EZpgUAGmtwCqjCmPSkuFzhyMdkK8LA76tAVJO7OxhOdG4owWmkwXHIIdlD
KDq9+1TqHEHvwiCRxFuKBFP/Ap1Felj5vBlTwkPQ0s5mvvLVM7wJjieCxVt+/YUtyPLo6RrT39g/
ismmZbE40YaT4KTXWWq++h2+SYes5ez8Rg9y1tnKgJhMmuobY1ckyqvm3pwEnawXNrOhaYpDR/KO
zHpNwVeLJxZ1+sRXg+MKREoa26uSgRcGbTlEKJbgU/V/2dShjpuU2Hf1UML7VjaavmGurhtyymHe
BVH4M/ndlOR6yYY3hzQUYIW9L914dkzx8iuMAptGli0eGGoFM7DZKJgoJL/CQrL/yMsV3piiPCoP
9uQkoRVX+8PTQ2prfhfbX6+drd+0+yn/C5ZgKP56Eaq71s5p3cwA3k/lnekH05YX2Q2ME+su5EkA
IplFXhuQ6RYmjEbQDcTkklY96ZPG21F3rTRu37naDDYX69fwW3GnmN8APlacVEQlvjgHvb9LDiIS
oqbyWyx6+gcxnb6Smvxti4heMhKIDMxY2x/JhR9aMnMyBPhwmzcWieApPEovgTYSQXypHvdaICa2
pZZSlqwC5o+m6nVPdJ9rsXkU+RSoNOBS4G5brzwm8JzTzGWfQVIEyXv7JuUUoIT4Qm1iOJnkQeP7
XHryFyOYi8I2Guef3uAmT+ooY4M0TbPjguWYC7xEOqcVnDj0/FY3sdnKH64e4JnPzKlee/t7Cgbb
HdS1o1DC2qIm+R2u3i559ZrSe+I0b1MzAts1nhVS9o0PMypcRaSpy2/3sO8SJcrRfaYTpT+i58pM
S7feGXQN4lU86f6K/P3L+Io2VqFMR4AVnOA5XXc4vwP2iLHNKxlyu7+IF/9AV2KtGgQPVIo9LBea
ymhT6XrrpFJMKi+4c2CQG42H3S4JfDdMoPrnhMl3o57Lu8xS8ubZ8OOXrUn09EzbsUL/mQr29+LU
y9PPTnOPaEm2ijNH8g4BEww3YNrGT8wtn1xhA0/myUIQpz7uImXPUr387Tc9t85PzswaOYYuvTUw
SgTv4DxJbpDq0JEzYF0kKfGK4lzXWpKwfVp2oZAFTgDgN+qy9YIia7niy1Q44ltdFJo6OkojBwim
tKWttwb5DgERWhydp8zuCRUMlJiMRcC5UEEU3Oyjc8H2U4pGny8sRvJOUNMm908K5ziXmtbSDXke
BtTjROcf+YS3rlA6gRksll5piUMYDSn0TuOw9aF27EPTqnFJvg+qc79R4dAJijoAXi8OQkOQdAmR
ruLUHcz7s11UDg5SyTQIZNKnDLRgffSbHa2/peblLyaFyMxRegYwcBxfuVegh1IKIeLgWUDiXeFI
HI+RnAebCWqYe4opXJCRNiUm4h1ORrNPGmAzc3XqCnIMpPqYp6MJVueucDTW4aAGIm1u/+CFN7Zq
tpjmgTsvJPTYkWffTGdM+lwHmfvnAjCRjMAfRtW9Vs1Ech7mHlF+c+FZZRR7lUUWIMrkEvLGDGYp
cy7Ghcg3h1lBPSJr4KVLavfxSBvUkhxf7+XQdxMq0B1Jj9T8vkHGcQiUQ41yI0oE3tla/omkB6O3
7j5u5bSxKSW/XOKoo7vFRldMxNTZVzdtYzSfr2Lth8YosmYkxO7FfXFNU6o8lIP3vuMbv9/Jmkqx
YcwahOhh0M7m9HsjzgUuIWbfdbTw70URxGh8yNVa41m5TjBHRo6IackKSRYj+u7QlO+kMlRAci8i
7flM6MHU8HSN9rjksSezk35Ilggg71dM1aDY5gU2hddUBhA/9ClhrU6sjMWxS9vcOJy6xfj4W06C
pGeZZ4YpMr/vkk1HYClmlwzbrwuxruLc8Tcqtp0uAWsXzcLhdGl3s/K+22EvYfvHAr70glOoQeEH
ZCVTlDWQ284l2ME7MlfyBjKOn/uTbUfOsZ4OVBMig2mhfTf40sQVnRnIta6sQL5nwLAo/h0N7WtC
WckrZD7U/9QZETfg2KQyRdMzg2S0xa6+uILqlkFlh7rsX/E6oUzKz/aQ0MZG4wDfEaCgdlQvWDu3
svnbo+vHa8TUb5dd6l0LmwRpyXfhmoNBcM/fT/kTUOyPoTGxyaAX8b7EsEk97QlNjl64MlTXTaSw
zlhauLaXGd8X7o7jrykIoSvET2Y6Jywp3QIOzJILxiADMGraAHBveE7vJ0hAb0RjL0N4IvorA/Tw
OO52eSb244J/ZFMK0IUcd58wrlKcACEWJjXVVphwmJLTQk4V53HJ7P/5c+6AtcaKz73dTe5yw+YL
mvz26qOkGDZiP2+dbkMeXyCTpVCjIPhfQolKOYx606523P+OEC82+PivGjdYY0dCeAgDWvm45A/q
JRvxWZsJoKZnE4DJ2g/X01aeA5zOg6LMONUT24kQ4SehZ+2N/z9b66p3F2F1mW2AI19hngdHvGuu
9mSnSJX2sJ3DxGTkG6SQl/CELXEzvRuou4PsM6EcYMowt3p6NWKEY/JliiadJ0QybsIOjI63m+jx
1KFzAW7vCvRNlV5ep5x1yIfhKiE1LaEzkOKezYkuJYn+0ZYumj3P8VHzm9fmRAPox6GD9RP+vN2o
9z0auL8K4BdU1/vePi/iVvx5ve5tl7l6xmOtDEbzwifA18YmywmIbIhGkv+5bboNE+iwr7GXTUil
mwDHgjMMQ7y17zEmT1lcpz86kSA1vYtP2TtYNeBQ5vFqqvJngeThq4ABfVoyIAoGPd8727qucyfd
ei2wwstTAJED9+hblQ2/BAzVkhl4Y1uNeVP007e5QaRpSrLTdo5g7LU9HDB2DfZSqMMk8JeofCia
mh7737SBixSd45GjOnBgisZcOTTghr9ksiVlQSW7AR61PeF/5mkiMTOlKgaZ07t/1m+iLdh8+4CX
w/eTibbq432TKYIi44M/USN+MevLAcs+yvrWDG5YSLmk8U6CzbFlEOtGeqzv4nKHSEmcT1XUJfx4
jApk5WbwmWNO+FRcbBIP0NQ8VOIz40af0oB8Ez7zJndCzOFweOgTr3eli8IZ+fTBPTxWzsWlyLZA
l5pVPjiKTIjeYfPYqHckJRY+kq+iYESsHHXmrRB+zXL9CLz7sCFLNvixKLiN2fMaIZV3L6iwKQLe
Fu7t4XJEGtrCLAo6hw0m2DG5kJjPUuO4goTj6guOD/oQMufDz3FMzp8yDOEjlaVUKrGfeaxzeNcr
cNTs8p0jNirDPUYpGWSbkhw6NadoncnF3j11Uw3/J4e4+ndqEM8lzHkdnm/LckGJvqMnuQ1u6H3k
UYWHUm18nsAeHsVg11iivgtbZYsh/09NexbaUdvMhBOUcfC7s58PjcZPbjI1kJzDtik1Xnc9Rqmo
555cIVcTql8GbZ5pq9T8kNKsYQBbmkQrLr33tiHF3MJz0weckijCSgwZ6PK6ILD4jWu0y01+EHxb
8BebsFeDWlksW9ZQ1qgqdTixxJksdxmnG5oYwbajPGfV10DGzckZdx6/KbsizzCLla2c4kCMNGC7
1Bp4q1isSaijTEW4qvi6ftzDPPiJ12hccOTralfNBcS+7LPwsPLgHRRSt+WiEIzzGlx8+RKu9t7n
jdIpAlyJEHLt6+QEUcLSrR2oKPsL28ME/BT4XzDIZh4SwrY5plp0U2dNi1nV1X9fL/s+OJac3lgr
hw/880AFjU+IQnuAGJE4pSCHvt/MBmD/C+TF6PWHnMTJaJ7fjjPcF972sxxRCijtX756ncFup6Kp
Z4MDirru8tQyf0PKEpkxQx8CfD6OcxClCbUGTZ+jkGZVcOEL1k4ZCxzwDjZ/8L1nOXQJK7VgKTxM
9khV3NAcPnjx5Yd4UH+ouwMHOtSvIiPBO9SL3T6es8jpqatr28+p5AOoQaJ9tKfHp/33+i5yTXxw
zDEsjLt5oUSuFgrKHfDbeuA7lzgwkUbG+EivvMzg440xOhEmSnZ8CmIVguw3fSu/bz/ZG41TSn13
M8D9/sVgfghv9LgiT1ms1Brcx2Rab3Dx2O2VO68m1hUqv4o7VY8JNAhg7c71FPRWCy2hCZjQfNtk
/yvmDr8SVuINGY9ODwAbmSHDvrKl7Dgz8wzpqu/eJJDucb9DE1NfFvbMMrVSr/+4SN6vfRe/WCPl
uJriY9+PU3LV3WDEi0kinaqmYkbLOLF/h3n8uxS9I1T9Ev9LySB6gQwDIiX5bSWOC4ZMTNDpVyk0
MOjikdon9w0STzHbfiDiNLscYju7dGZsxB4FmpjqGx53exuJHPzYQl4li9N6zUs858CNwggzVPj0
wxdsXpQdIEB3t/iHYgQCoFQjD2GI63Et477Nd7C9Df/I3vwb2b3W+OoQStDEteqKuy8PJiZ8Z966
HRfFpS4F71C5NsjqsbA+QZx1TYH1Fwov4YnVl2kxwHJuLNXr/ODm0cX17D/tAvl58aTq8Cpnk34L
SQ7rq0XmhmqXcT/lDMhuLCbJ9QYbfGWCWgGvw8WE6GHkZEdZOqtuQzMYne1DtdVyzM99LlDBgvI7
odFMyqs6CTl8jrSR4KNwA7IdXLSRHDiWI9agWyXmeTcqyYWQIwVq1RPfB+mTPKi7JirqZhFYstNP
BljHRTGQg+hmKyVs6TBZYgFEHsl5utT34mHU4PiRHTjVs0xqNcwREu+N3DFPcbvJ7XHzi0tKZg6M
n2b4dDhwF6G2eTJ3nmhYZm0BiW9JvaFbAk0cK3JDRy/VxVedzb0PbFwOhpsyOCIwS57FiG8Bqwue
QI1Zzi/cxbbhv/dg8by31MaVwaEBYiEApEQrfqYOMon2OQtyxboQWraT4QVZMMIugQkyG1HTzdtN
BvL2kLZdMDqD6nqcoGCGqPbQNt1PeIgcok6e15B2yoVPAsumIlT8z3USg9J4yhsPwFZurvVDv322
OsUcGlwyLmts0LaVF5FWZXLIHAxNS9p4YQWuoHLNRKhIpJyW2Ew8G9T+8eVZFkSEw5CdRTD39NM2
yYUwNmnI0ct9Z2dTB1/zxU7Bwg9/ih0egWKzRgVr7SdWt9tgGd+QUtSq1KLPPqOe61SVLDk+lhuz
UqvIbNm2ICzpCymV+BSEtqisyhNwX+QPyX/flxV2W2YB9GAzMkD6E9ueuMRlUgltbgCmhkRdEFef
CP0hWP6QWs5FZEn03QjxCaw1RlCN0QMS7rfrUEQIyIve2vr5e3JUqsqlVbjihGrFDJPqqol6posb
QupRHZNARyiUFSc7DkvrgaxCN4JhyZf2RYZCqEEAmmQI0n1a5+OvXsNXZi29sRgcmqkx+8nrCOi3
SNbfkNKfQVcYn0j0xA80PZz9ENIi8m8a1pO+3iJMWVWx8OnAiIAJq100HpF/9W3aVBhjbF3Irl/b
qjitiRgiFf4D0UnWEmyf+ui4IYWPi8rEH8h9YejhT9rDmqNSPJHFw3Qbt/ouHjJLYM/nXY+6+uFR
bzswjvGjoRREPWAPQkktb9aATvf9/8jMAPzB526v4lsHfsya1JGWvnWsKmE2Qu1zpY0lFG2f/D6B
6dIFKxvYaToOU8X5yyjnGISL22JCAwFeuiaY2aBsjgZ0xcQ3xRXdhIhmrZmmyolFx3L3+fwCHFhG
qQhgNISA19i5GqIjo+PSBbn7OjB3N4e0XbQ2WExp6z4lvFP51mA6uIS+EmJCSWszGkeNgsZkyjm4
yMGRl2BgO/taxOq0EPE3QJd2ERf8maK5dv4EWNEiv832gkF/nQx0srGkNKSylK8akcgEg38o0NKE
G3rkgAlrL84C43EY8YwfTAwHU6otXJLawrmm3nYC2BfJsco1d1Ik+tyyjCQtTUlRoDwVRtN/sNQQ
FKGJjGi08TVYtVpuqFZahbDaeeQwAl/pyRvalUKB3iJS9FhhT60b0JBgSvTXPyhKj7Fah5FIwHYl
1PYgM+JcclQo3jKFK2Uynyjbpv/m7YStkU09hmz68jZZhBYC6vKnQrX7jiD9JsoRURk1O0Llb3sv
bc1O0+AfQijtpbcGAVlo5LtypTPqACUJo7pQpYz7q201R+DmR2vHNwsBwS8JgIIUihBidzqPdcWo
Y6KSuSiMR9k6uRJ7bLDosPC285OXC7CtjJnVQ3nJHqcluOiS+YAtIMcH4kAx8s3VW/CHj44/n+i0
GH17pxBb7ZbSDHyfLIeDZGXOB1Fr7yjkIlgV/vdaJ06ILjBSR//eKMFpcs3VIvzMiOeZhImtHt6N
oq9ce2MBzanHw1hZvL/yZqBOEWsiWMrcH7Lsu9O3fUq6RYEMjLc3rpWFgfF8c8/uA9LxfTdagaKS
TMz67MQVdfH/hADkwKXl8i7ljoPk/wet6YqbOu2tQvle6zoY2qYbm2rckBwnIPlyd/u7KStOqx3W
/Nq5BL3z14y4l5J5Up9nh12ACGDbYShKNNgbIdg3DypjosNAKwvXNpY/BbE7dV5prGIMvL3VQDP1
A1suV1DIY+Nf4Kq3+VhW/5G+ktYKaGFv2xFtZmaLQpwXpXISA6WemfRBVnfhGzPi9ToU+TDV9onH
VcQbdueyasMa6R5O217CCk3orEQD4q1PFO8H5slPOvtXU6xoRTI6xNaGU+8WusWGlFaJDRmpzGDF
U55p9X70TJg8d9ttPOLroIsT4t/Kw93taUMJNtdEksZ4whECu2+QK9aoT9/d916lnzJIRyiJ7Tr9
3rWuSGQ1nTLZHlNxPk2eGXQkFDo07JHoGlDfO5GNssanAIrBZLMIf9jPCr24WYcVNKDlznGtN9Js
6/u2BJeZgqusBf6j9oWJve2UH0w7fYXBQ459Q+vQZpHdvPeijJvpuB17uAf8tf9zzvzicp2Mrt45
vtv4onInHYANXU73Q0pOkEYnurHPgL9dfOfkmJX9Ex+USKELSblpw+ZW/c+PwmUnHUSsbYln9NZP
t5Uvlnab0TUkh7q7UAPB+0MSYkkV7PTVRtKBIvDSuwTdRS6vweDgqlzrn+WtG4QbN9ZgPh8dWjv0
rWKAFUXulrjlrDXhZccJwklPxgXB5/FYce2T5q0efi6rhyH0DAObyZydDDG2Vpu4tJpFoh7F+7PG
EnFMs2t2oERqhJx10lQEou2XQ1FVg+Wx3EaUOaf7UzT2b6mDIE27ENLuPqaQpViIYTNRVTw4SmZf
LFHTJpPL82P+MDtj6idI6CcEycZH2xCU/sdA8eyNVONfrzVL4DB3VEV8Es1GujaKg3leTP2Dvs/6
zY/SUCc4QE0qry3LgAqCL8XsMBDyS1AYqHFd5VXMAY4YZG6gQeE7QH3yT8UAa31Vo8Pf5YA25PPJ
kLcaGuP2L+tXOKg+QFGu1GOnMNl5VmZoOkOIjL6eeiEHUAFZ0iqqhuSXoJ3c96OH9j3uomXLG8O7
qLmbJvetOFJ95GOaH1NhpvPMvpOj/lK3rtzAi6sdtaYKJGMOEuKtuDDW8IEjZc79pEQ6TA+2oinx
IySiJ3CL1hOLa6+8kGa1O9ZGV+3GfrOXZWsmVb1FRMe0gW473v4Lh2U4Q+cHjEc2PslRjIWUI6xi
bmlq32ji7+yptMAGBS5AEGH5SpnP+I8xdVvem67vBbRER2sANt7ZFuwRYdO2CwJ5JJ4WggcYpUH9
CRjp8fZz7HV5501DAksj2oeVSTb4ZThCjwZ4aJdtbySyjFwxmhF26NcV7NvCmfw4w8N2gbkFqTY2
paqZovcBQWGh4oXlWF1oH6+I3fxBTKr4StRFd/QZIogEIrMEWARpXqF7FHZpMLge3fbL0y+nbHG6
HxmPyX6WEYSgGsGIwTHCg7BUnfVJHOiVXRl268JPgmPNVCetE4yMyt92z5811imUyZC0rFSXACAs
ypkC/ZFjdk61bzcWf23d/621x+tbbDTkrvanghYjRHdGQZAmZPWbA49pXUidR1yDvmkLexBlDjjj
xhD1ufmqiva0jzoKRX2iF6A8CA4VyErSc94Hq9xfsgjWzQGjDeMdArWK37CD/q4YUmwP0Q8d00RB
LgAVKVnQAqmln2gjQFImp6RAq03WZNVIsDm6HsTAYMDJ18z7NRwtDh0WF4nHKMVimXrvKPXXizEM
fmZXKKq2e1rSK6yeKyaZm4KSbzqaOl5BhkLWA5ZHxCcBbkugy43y/ms3sbJ4rUR03E8C168fSzNU
qoJdTRZvH4KuB+0es5yewWs6u5ZVe2dqKH2jfpeFLxRzQMauDbyvgxdDX/3JzU3hKnv/cYVyMYBN
2fD3iNB4LcD7PIq7XkI1p6miX8/16X8ySWmbg1zmR4VG5lJKdvpucndu7rbdK+RRUUFvXZbErypL
LaVxMw99PdN6mVqwCusqeaLcXZh1xklJM34mWlcGkr16c09bQKn2+cbvNdfRrNcZbLgCgUV4ADaA
tnqlodhLcObnaLintWAGo2X6AvHyNUPfWWWkvF+LjyEHCIBDK/mA8pGKNLAumpSyDY1keSpPMK03
KtqUQAzI4ZT58QXdQ9szwocWJ9iOqM9akS/W6LoakYMTduv3GYotqai6GZTv+4TwDUrZO261YyUp
tJSqDwpCrYBWBhq1qpypkk5KUeiyyDZ9rWImjxjUbgrMN97KPUb4+aeR1l3jcscfCFAsb0Emg8Kn
Ty+ME/1vguxIv2xWRjDyEzEpoTgbuwNU73CveDyxw9P2q6zF9m2b9j14seyHKoyq3RFp9vJc7fEE
jpnsCCWEANPBxMQq9Be33W8cww8NTy4ihhC6SDsbDNOuaWP1aj62MWnIHcysXulU+V9t207JKD47
gcqQdaCis4UxCffOfbH6z41eUBz5l72Qvd+NYrJNW1Fv8KJXll3Eh/KEhKj+qESjsWtEh8zBi1ta
2LaKwbDq2Ar9v6mnWTRC9dbvI4BiuuBK/ObY/3VYZFD9FN2yiAX99kdWvLaSFDSSuTNcBK0/2P3P
Xyzsk93VIEIl/f5llXmgso2kyNKfvvswV9PtkxmV0wAmOU+Ggq2xI21/5jw2oZtp26aFVmt2azu9
vpI3+u0aZY3WR42T1dVx7ZEnv8j+DOo2VTZdG6v16b5Zo+v7H4DLyfjOXyHMUfPPe6TGDZqcXSlb
ytpsRE5XM2atUsOG5ZjkY2FvVIwneBAKfpuukQZVfClklfmXB2f9daEjwVruMMGiJLZB8IThf77X
oZzLbMozh4JZgCS2ong3YoZHIJM3S7sJ2lkh64CEJFMRT+iXTYeUNJVlhlXV/pSb0OgqidLyx/k3
LtJCQl3aYP8r141B+lrOVGSTdk/QiYVmCRyCt5y08kCbMLCtGktb5ZP6HTxHnknkQCuyGejNr065
sDSmghO440tlYcrWCJsA8rtzlodIMskak4T7QDR+AXgllh6vszYXn8nQdJXxdZokm+A3aWZ/JMMY
ALGlJriDn6F32+J4dBZFdnAS6uxagpa9FLQMrP/N+55QnMAZBoPcGMd6qbZevK67EFgkDxxoJsKp
4j2+VO+Rt6hF1JlCLWVZSpdhPR2/dNPHQSYMYkFjfR0NX02v/5Y/U+cGNJLb24fP3IO2xya5Nrmd
5nEfn9g+9qdvcTsWId5f8Se2p0cJV5MZFDp3A6T/WJaIAbpt9M96o6DrSfz25tXzCdu+GIxRKjy7
DitnhpFM/fbdfguNL1z+fHsNOyeJ2NSUGdYJIokZ8TvSB3SS0+xKwpfsFUzF7XBniI0wvUU8zNdG
aP1us22kfR4eYFqhF0VL1EME6iBsXQqxEpYBLO/GYn+aeRs6RcQianIl3xTI8Wd8QgeG13lruafE
rCt6wckVJFkp2yT5PjPRGhk26u8rdXfX6uUFVHsS6j+JyiW8Li2cs8FXq24gg8I5AMfBNgyJ8Lzv
fNNoyJZdaRWC4uabkCw8uQ9Ku/J3o3K5cgYdLIyBkpfv5pfwCAfe01EhnGivQ8Ie4j9m0WpH3y2r
9AKFbSU7eke5QHapdJSXuluGE9ununwSyFWG1f/CI3AbzzqFp33qfRheM/0fAOMdCq4BOkKEsqh9
bk7tqJF+cHtP9ecx6LeO+/oUSOc6c2KCzFIQ8nVAuELEQyqfGVps8IbrQf9GR47tsW9hV/6Z3N5K
K93lXCmdhFXwl24o/Lvn9wBNxeEUlvpYm7JqagXQ8NunvDxUFI8yAi9Xw9ZEDXSsAnnVT3vuMXa8
nTZ75dtTlVl+2Ee9T2JsCloDm4R2XHUpTds5l9Y4ZNg+jyRUmSQ3F0SFf2pdlEeeelxYOsyy6ml4
KuNwgEKoiQ66BCY/1qA1AWioo5kZd86s68rgGwhNSBpZws49QCUe84/otRVRrZkHxFMsnoMNZ/di
1pqr5JylJR2kOP4bI1MOsOFdAAYKbTA+jQ2KvBuSTmD2BjFViEIQukBv3iyz0diEAmNI3PQTb862
obymr0H0sURzWxAETQNJVZX5MOs2HFthrbFAkCcvtBxDOnNS+Y7lo2EGXCmxU4dAfelsvMnnLXp/
Dvce5BgsoZXzCTWSkz80PKlnhXAAruOiPE5HF7hiGDp9uJRUqVCCxiRsgTJF576/3n5m5yHgp/SN
zCjwuy9Ho318q+5T/+lu+9OupvSdSAkmzI+l26TEwQrz57r2f3+nIye9cU3vC0Y9MdnPeSHeEfNj
JP8A6NRvW6PHukmZf2hXKkWQ0V1mJXmTK6dlSKAw17YO9R3RmXyGo7M/kyCTgFYP8JtwVwvPFoQW
tbh0Tc2OMY+MNSZ4p0H89zfx05KvfzjKwom5M7Tmwalhs386ZLSJw31pGgzJgzRIWKeXxSZu22Ie
CzMuMkQn8174g2yQxuzVkzkFa+Z4zI7MUSS3u855RJh+7ju4CVs9DPvgGf4Ls8Znw75lJGlYrVzq
JCtyaPIDB0ndWlTxz542YtABtviwVb/nV4yWkmjWdwH6tLd+wl5kbq8mXBHOTBU8CuJRK/Sv3skZ
gaLox9ywZChN8ezcbJwNRDfLrJLppcwYxbZ2N22dkMdI8WzCriBN2K9auBWfyBlP0+8EW8/1sjTt
/6QZp7b56J8YP5p3XMiK6SmthzAdpu9emscqjd1DNQXASXa11KcCImLsDne7/hnubuBy3XJ0tZYi
46kjGDg+kAnbHoq5MhuMrYmiY5ep+305JIBy5/LORshishGwmqwErpV3JtEYL9tHqafqdA/aoEl7
qHxWqIEV8cXxIv08Cx5CBLRlGUD4iNiHnIrsWzofLxh56kkfLajz8NaUVPqYH5RQBW8NgnRjyyi+
1d30L5H/GAP0V7O6OrsYJLBVR4rz5OCcy6K4bmegd90ybYQCFgZGNRJ72Appr1VOC7fbs0n7iC50
kZgTCLJR8Ij2qZUlibUIbj2AZUlOsURg4qd3k95WT40wOI5fD/QOW6yb96Ns/dJZy3BVJRGDb/4y
p+PKy5d6tc8ya/Cri8YXuzjPuYHF+BaiYJp7FkFxs5ZgnNdVeMSyExcnmT4FJf8vOhObd6JG+UuE
sqb34XvyAJ2QvTB7r/ZvqyYzXfcFMIV2CZv+m56ZcKfrbfIE2ZuZKR9pzUhh5aK/euyI1rGDYmnQ
bTOp+zaH9askrJllXUrBSTso8+1WuJ3/yZcKU1J7ar8yyw/FilgD0hczvhoh+DRcH/c+3cIzU9Wi
dypPMiq0g9rLF4MwhNMooMtiBiu+dD1dw2NxDDLrcZoscT5zTmycIsF2p7cBZw/LzoEKyBY3y4BF
9/Pf1YsGYJ6ojvdpDsjcDM91i0piYODyNYGw2HOqBcvoaig4dJTvWvH7W3qASAXiRNeADaWvMhU9
SjdA+KMOdbDVQmczuHUgtV/O6MQ5y0KFLo46OXso8ooQlHzY5FtqMf+cHT9se6zk75vHEai4S1zy
H91BfC2PzKFOGMU/bp7sESdzjXCtVJmq3wlXDIzvEcGj/dRSNdTWjOwMa2eW5ZS3WfjCN4tDqGMm
Svh6WzFMiq9en/dLu6qL7I3K1gVPfssAfk/lNex/XOM/9FVi/ziOvE9kT3f36owkUFuzjM/5f1O3
7A/WmkNakIoe5m0jYbXh8hv+f6072mTVIgk0ngwo6I1bFUpbuTl9WT/cy9gCxF4mXkecHdEbMk9U
vldADNr6Rmr5+jLWZdWACY28/M1FrVu3JxdF65XazXQ7SLwphGUVw/XqhpsZk8OZ58TSi3F7pYTS
EeEJXf8fBhUGJOzpwTu8bvnWberg++7KZl93QUkv/TO5nOadzIfqHWPPSDYekkDzM3wWicpyDx+E
4pT05QKl6osRPQqSMB98brpLj8YOUNh2GSxyQ5JX3W6vuxIVUQVlU+3P7TevHP4NZVNNp4zXDLzD
rMwNPTjskP9XQzbvpqmW2et7tOvpi7YotxA/O5Kt0BZny3rMwHOLPvBuHi+kmr3lQZ5zKdOAp0vZ
NmVGR0EyGudWQ9R+hmkZ4rWphUzI4BoGvAIQ8WSC+QeWTGvScU1oMwMaYiaH5qpZbtKW3aNJ0U33
hBm7TKKuDlJzJhcOQBDLQkhAwvRMey8r/u82tX4hf1sg3QZFVlKKzVdXwivzBS6JcmY5SvrjYexo
nj7G9lrWjd0FMS7Zo5iHq3q7FQoYHAAKCDX6ohOUWg+y6dEDmj6RADWOIoRjb4cNFWRHvoXc9idX
StlSv64kawfDBlQUh0GtS6p+rNWtTtGVLTGJjg1J4FRAsbHthxVrSx3Hp1yWv0AqcU/3n2zE9Pq2
XgOzpteizaSGfrMf5QEGINu4h/VhDeZpr9NB9+MgIj9VQTOgh3M+J63gyjoojTpgkjyr9ShA8dyZ
Zlm6YVGivwPYQlQznY6bMdZ5s/h8ydJtwCmp3GrJ4ljtP5/e6VdcHtacs9f7M5IyB87R1l4EgnwE
m1hMum5i6pZvDSFP9xb79XNs7ACqyf4CIhxWhkl19LeJlj7WysvHup8Q5PCaukT5NmuFjVW3K791
Kk3fEXKLOBf0CrEUneKGzxX2hVhPiZbFCnJDtVbXSFBfzQ7gEXjLxlZVdDM0cSrg5GJlnsUXMbZi
XoAi6ddH04o6KzjuEo3q94plYX8IrQSnXMoOxBKtiED8AQ78d3OLAOirxn05C80OnYIHPb0x2dNx
Z0Php+0TAe6Ck2nXFJidpcL3IKa89Ov7n+tZSUHLOpG54WXX73CmmEgPJ0YupaK+5h1PSc82P4xn
8gsGCPynHdy9fruvG9b7QlaTOQh83YYRgz/cr7W62o0P5hCkbjLIlGO36YPQHA7c36OfTW/v/CN3
CzZKK6/Ll9gQzC82BbOzJ+hlNe96gWglz6e9nmEHngLKO7VGbdHVOAAvQSVllcKTNSIDnKtbZTWC
ftpRPNNrCSxC1HgweHZcT5uj3kUI/Y4PuFo8bpk6MC7OAdJacEZHxnXfpbLy7sK1SQNSaBqc1WdU
xsa2rMcqaHbXadVzACd3DZqQxn9glkuFo6NwTXlTr9XTDE1sbEi+BF57INpAVRL4Wb4aFjj2pqFG
ezDcbAnSMKeyjheKnbYT7rWFtboHOX8Bq7hyyO0oBWy5Ox1RYyTfzVttodcZ1jq9gEw4Xsf9LSBw
wfNNTtRIlNFQJc/FVhgbduetJ1aAP8u/HpworQANSFSq9HZzybxSALxdi8gM1rOLDmWVveDkDtvF
JflLzEubH5/WQH+BowwE6fxGwqWOY2ufmHFIDLeXGYF9Xh7uYmYvaMYtzi6HEwu5c/RDx8wEdgQY
M3f7WRrdRtG3sbX0QHXbQmy6p8mBUadsMB3iyzq0mLoVp9H4i/IlXrnSpV7uKmvzX7NjHO/Jc1Aw
V6SXxB8dnrT2OzSjmkbtvBkhEljhLmP/y62SrkFDCuM4gAi6m2WdR0Q/uBJGxyBc2yL4/j82NHld
0KQj/2k99cSAFQEcyeMyJXQy+2qAdl4FQRf7iSKVthPnu6lhnShiCuDLV289MDn01aoYV35KcmZ5
03IACKlvO4dUkW4yntdHVPOYNCuzKk6Av0jxOtzrCHN8C+i50d9d3v0m1V3IVf1oPdcF6i+AdfUN
Ir9VtGgfDWXkh7rEdVt5bZLCcUh0FU2Vy91ETb677dcMR4sd+3QE7GIcYt5+rh5c7RySVtVpmmRC
sFIiZAfWLw2Rj3xpLwS0aB8Q0JoVpL1w4f64nGoG426ssChKh3ZrKAumB3NP0iSAY0apADdTxeQ6
z2FgO3jX/FQYHQxreusmorga6GViDZQN8KrEAJHTQUYCfXUcEWSvpnZJqDVDwzbYUFGCnHkLeRef
sL81tpKwaWL2Pc6V9/xUvd685kGOl0GHjMpOx9RW7hRWSphDdK1rWK7/LwrpXNzRBi9F0RAMe3PZ
93En5MsWQmjlF7vwsv4FNuqZTv/msnChE51k2NSLUq0L4EWEcdC8AI0fEq0Utt4LDJZ0vhJRhp+X
ysWu5b9wXaXRci+ZJHIRY2XJ0QJVhRDCQJ5sfsz9tr9p2A4czvEqQgEqxoCjZfVQVI2F5yaPD0cM
Ae4JX2u7d45pcPL55pSBCpUDIScST2D21ZOvjffoAdIc6V3cCpWXJD4HpshxVDolfsaXUTBSzBUT
xTDREljRxYX5VcIXFM/ZBCiI4twVhI/xs+xcmKvhukDDkzNeQevblZHKgQ7k59dCei/TtbbSBT7L
yhxuuztF7eFt2jIR4OTRtNasb3zoFxKSuqQkf3VJYOklpkrLHTdg8W7NV5+rxNde4SvAK+0HEE5A
Eq+PN3RnR5S+frGf6Q1z2s0CRNnvo8cH2twUPc5/9nyMfDmljBkvg0EYqTH60a3a7pKnigRbkdTw
z+Y/UOlYWIx8DbB5/f3my//tBysLDsTA9eHHBREadal3x5v5GlFLcQ0DVKx7kBnTqesOPwQM8sZF
N4Vdlw+OUDdpkndCCsyNXhxTAwHx938At/Ugub7ai98NPE2jEWqGwG0XUII7/sU4T2q6/2DhNE9x
di3X39TDKDM7FBDrH336CT/I+nftFq7sICfcDrjE/QWQzDD6+1ahVMTwbUDbeBJeiKLwNjDRUMq8
mhdZtD2XsaJ4qJnl4HosWK+5TGlv1NAd1tB2hnTJc7UiHGs3ZSRlsONOCR3o7xnwbZi1pRZWd2hI
w97nB5V7XK05XxnrRH5/89MpQTN2nrNDMPZO5YZO65FRqa51aUEFefJ1bimR/wUHyg1drEN28Zkq
KkEFEpL11O+0Ai4oHbjvzE5hY7MWJW0nUNdsi8nLCqCHNO9x8HFrb+lUNVZxFJtLy8rxrV7WqzPH
BjCIp5WdZXQyDx5xiUI0LARt31kg7Xkx8HvoValojum695I3bwXhGcj2kvyqdOVK8BL0v8SZBWB1
rF+H8fwtldrigywISygaRT1CJAufC3647xU1xHrNlonVmSUQx0mvS6hleUUlsTQrT8t3Zr7l7Kkc
PscOKF4da4CzRA7KbtSMLbGyM1NWAysksUL8mioE3Cd1C3qJdvhhLaX+ytiUV7CKQrQ9T3hcOv7k
Kksa2Che0Qt/ZrJITJnjJ0k+vULPZ4lMDYaSJ5gfg9w68mW48wdpY+IVKiA4PF+c1KAPGs59cMpT
cdd7jDOTduUoCGosk4lsmIWQ3GB1TtjgjDGobr7FZf8lzJJfbTNxT/hRmDcqrr3vvTLjUiG4DXrV
t8npa9rto9jFwEtKjaPP5IP8t7kTQyDlDGwCqG/kNmKfHrR3zexBvQTcE1jnDSAjgJtJm/EZgZVm
9aapm+sDmlr5JJghqZ9w9MCr+vNYlydZ1H7ye/iLQkgQ3qIZb4iZW0+gPDK0khp1ApC3FE845HU1
tVW/LLsLnH2OGiAUP60keZ/YPsa9l9Qqs+/iqe0EjJE0IzRKZO/ONmYUQVYtkOjcoP7Vhb9UDn1L
m/Ws4xtwwKQdNJbdpVqcH5INch73GxBh3GBkshXeBIaZcKvfnKYoAH7Bi/vTBrJBXBuPZ+ciCyjU
/wM0MEkqx8uIIFPl0SKtIKjC+lmr39iHw7w+QtF7ZfwsbkfGlh1hC4EGL+wk8eHIfUOPNH3MLpsj
6HcbeJ0j3Izr2tP8HTRdETjzJPBtYuPED9kGfXij79LuRL7zU7tx38YOaADJ++4x+6sCPeCvQQnp
N1uAXyxa3p0gkCFI/yqri7ZLylUg86zq+9liZmokER2tTk4DFwTexJ1oV4sZfmDFkzbgW+pqlUOI
FilYNNY7xy6je9D3B6EJEJrCOl5mmvaylV+SN4wubAVQS77Lb7kyKEeOcS3inqWFsNRXlkHXLhzy
WrOoMyIq5RfCKK4zPQECjqrfDZpidwzpq1RSGYLKMkGO+tiV6ClEQmW4cUV+THPcRV+dC4fnpISn
nmkarYBLKr3DhfRWku+cWx7JPtrJ2+yCZt2jSRQbP2Utv4BAZ6PonmSQlX5HnpQTe+oAF8PNVrPG
dBI9wtoCkU/BX3CfnNfGwXTnw1uObzV3XIl8OmPCR2rSjonxfLkwhYToOY0Oi9SacYz/9wt63v0r
kt0eA9cJ0TTw+iU4WAnrH7IQDEk4L7H93r3uZ3c4tteXfQ7oCkD063EaVGlz2/u3p/dwmj/c1J/l
EPXPR4R97ZddHjWa+G/FYCFwi5InU4pIYJyzz/QQE5zpcQC+FG0mkEnOEoXlVYBE2uvWP2xaUouA
1hTRazu+NDuGRIN9Ctcp8QXzdbvanzkQ9OobngUT9QXEsWddSYegiPnuWlrOoSMEgH1ctCYZ9S0F
VYibVaiX10vjAF1JHMQQI6aERJcejbum6WvH4lM8NqShvuf8/OPGCaTo8E9RP21UDxCn67NBJN2m
/jJ5t/gH8JpbSYOVV88DkFKCSCLVrIvoXXNeSZ8sSYtkFyDcVFFCjAn0sRcA/iaFGtXd4dpq/8W9
cPcBy9jAoXO+kzKKkb8SMNRolvdbz7iBiG9AvTHv0ZESFNV6TKGbJKHwCjyPU0oE4Bkw92D5xQz0
v7/OiXKst5+5teZhL7quhH97+99l2ocARN6GbrJJPJIc1g6sJ064LmuAttvI47sOdq27eO6gdhEx
wBVA6N8lcphSAcDfoj2zWHs2w4Fiw1oLtXCaj7qt6MEOX5lrVMqUNIE4buzQSU+jzbm+wniIM6fR
yi0xkj2KvLsOF4f6Ot4PgCi5EdI134Y/BT4I2HyqlGp5B5o5Zn37uk4WUjAQoAD5m0rHjQZT3ljj
7DKkgCD7vRUJbxrRncOHxiI5LyKXrgWRKsdNBaz8R5VWQ3HsPW/XLihTUCuGgnFXoP9/+PgM6ZZa
HE5GLpq8YYtJIJ1Hp1qvGYcK3tovkycNTU0xyryJrSJGTsMNQmWo9OQM6S5ySciu64T/sHMMcqyc
W4vmepRTQsdjjqXrVm5MwsHDe5HyzCIbYNOdTT11UbsDA9FO20EW9FXqegehrJiSETyDivvb0dYC
BfsR6jh67MuYBZk5tK5lAnV59qrqHIjeu+gt/8LXC+VJUoFvBPMZ6BV42IlFegKxkBi4nME8ntf6
girQWblC20Yp3ZRl2kAx6n6jBavJn2wN7Cm8r7+REGDs/fisYwk7UM2n4VpnxH9wLrF/Wf1Euatp
HaDsFYpYdc8RSBom/YcpbyqbckaIBHeDxKbozEsXZpY2M6PaaKwc6HPDsALUnOLv3zNlj82dyCL7
JCtj6aLs+QTlc6CmE65alpchXC5WzfwhmevNZEdvtWD4GmQi05k6xyfV1Uic1+agf0euz+hJ+8EJ
vD12EulpmatZL6rmtw/iJ6Y9vHaR4GCxtlHVwnUnLuea1K7ANmhYprqYSz/2tMTOL/EUPpWZL6QF
dU3ZYFBFOHkTJnpuNG2Hx19z3/bY8ARzjC+l27IoCASUf9JTvOjtnaUiv86Fy5GcgbM5JezM0uTn
ej1YotXON8rqeBFGAaUmNlNCPMblTV47Zm2oy8+08eTZDE24xGyG3r6J4VJPFxR461GNXLTHlWJb
Ebls6bjstlEaWif4YLMvPMz4cmugvBoYt0BC/vDDCPxuWK0bEwiU294MhC7/7t1cYE8v/+ivvxjW
8BUajx0wX2FnGm8wJA5hngT/RijZB/qimHhBZRUbtrpEPvw9B4j5WBGen+mydFH7kcvWigQUQnE+
fjvfJndOjZdU1ekEHGD+N4b4uh41RZ9j/l7hvbZ2XhzJaigP/lPfcFC3KsMRO09oHkK7OkdOy5pu
MbXG7Wgk1DTJev94IeuyDbkkwe011CmWhEdazwqyQp1CHIKtIHwDuwdZln+H6pbwHgrbvfqEppQU
I4namIC+xjO6nzN7NEErn6sSFdS8FnUlC5qNG76Ay5dl1E1IryEI1zoF/uqeDrdZfHZ4c+QLYT/y
xJR0lEu0bMmkKjw/JKfc4w9kCIfNtBN9j7ampJHyYOsTYw+Zmh2oX783EKaYe6mcdWvsJcRj4+dj
EP7NtO5N/+8pqPRtoxdzYg2502arFq3wdcmGBVLm92YSjlFS4+pCGQWUeLWbleDG2a/90dloK5En
8LdXwk9ZQVfq89ELCXkTK4sPpjn/e2UUJAejteQPI48sRP/RtoOQfMixewaZ9Yr9mcCramk0ZVqP
vu8kZ98wLsO2t6YReBghPt3lrjkI4bb03D3TvtppgSxwBPRNxuAKySq8s0njtTPSbEYlTyyqAb4k
ajNLyAWtfiyg4BODH87lKBNU7MU7BHAOQSNQxmg8qXWeInAycE1XVgnDTv26KHlthUJrYKYhPLfd
zz+0vWBlHb9f+TbUAs1iyIk/FokCgX2A5SE89uvS73PtCfr8oBmRl2iSA+XSQC20K1Q0whtZiS3B
EWnCiVu5pKPD2NpJvvtBykHd+5E53hzHDdvNIPk0G5JJEWBH4Tz9o20QKxzdgCg7hWbpr0Q2bz2u
KUNbnNfrnC9RwIhRFJY5xm5/hw4ljx78Ga8NuCY3vFq9I151P8vOmxlNrIl1dtXY9RSOZ7207HdW
a7Sb5dD1Z43hc6mnTZVaoUzjUeeqwepNqv3g7N5kW3R2DS7MMT0m4YepiCp4YsHIBjBlWEmNdb0C
I4wtsx5hj08dENw8VZJVq98uJSedsdNtQTyyKNbqnfgsNHLIEn/rwFusi1qkAAw9BIo1nwOmMpSm
NCCod8rV4Bayi1ItCvg+dnFw0IFWLHpEB/9/jgKYFXpHLiN0qXCPbsiOHQDdIQI+vQMnbLzjIh6k
LAwTtAmuPR7rwSWCg4tQLzmRrRiNgo1tBxRMSGZbbw/W8cssJh/No1BRByydAScTOTX3KDR66wwk
WKp2Z/QBuigBWsBkJtRAQTKQkUIvdPDtrdPGNgrW2U5+vIIzGH4QYn2G+klJZPQrMmpRWHB6aCHR
4oW+iec8miofrU0BplOZ0b5sT6x4aBXpN+tchNuun8HXgLY4UTLdPKWCBV7AaWcyoR/MpyRt4UDa
v8+3hT+rFCd+uYOK5jjikyAA4OXNEZ0YX1vYRO/ArH85cMTx5cRObLZWUZb0SmgqlT1pJDziLRWc
LRq84dwSXqTaSQUNSxNl1yhEScyPVY7IkyyIFv5qQkdrcK7pOdIGg5MJEALU4LE/ZTS2a2tfbdSV
aS6wiLESgPiSHAjhJyJ+AGfUD/7h5iCNedZlFsuMJvAWtu14TFeogT78u5YesyAq5Q+ss7+XWPSh
oNFwVf0a+7vO6ggpwh84kitD0bvkZNZe1zlxY+xBB39u3c1gxqXlqzDlY3x7hcXGaa/SCdHhs10w
e/NZgeK5Pe+lKUBOM8/xKUBo+xDFL9Mf0dvJNaU61hhF4EppI6AVtrOXjumM++4LZM4yAt3PhVXH
Ub7YUa5+EEqnkPUZxreLZFuUdhGn62roSaI0lrtypuIeSOcCuBUE5lsm4qC4U5Fz9617fIDvRYCa
Q5ixa6xDmMljlesEA6dPUg6TlEh+SFB3Nim7g0peyfk2yGSAJeAFB4XbR56LbvGOuLs5ss3c7xyq
zXorDE9WrS4w6AhaJt6Wxn4FaQxBgKb4qFT++kgZTEKrV28UPyiqTWJdU7b3o4ervfmDTzuaeZLP
7Yzgzj+MvGc2MD41QtBVTaNOQUQYZQkoQMOJf3e06bHGlMbsgPPWhSffkdp5iRKFIOf3SkRoUirS
K2xdInBJ1rpQP27EQbqYa+5a7FQ2QpNRkPwwxZhcvpJCAcwyM/IsHx5jZcyZHACI8QYbLH5c/ZP1
HC8j4J67EMGRFjuK1O16RrBxfyeYIE2BPesHn5QEojeXWG2A76n04HfVZUuPT5iZ4GDxltE7RHxR
rdhQiJtE/7MzAsjl1Lc+071s/ijVVc60ccD4XGyPiN4chhOrHJx+lS3TtapwCBDjXWddKGz8eDIx
R1SPhPrV61nUV+zUC50w/06MdoRoq5Aj4cXdC9EK6ssD2Sm8piTjLJxHYaSqJaaKLyIBAN9XVfNY
iHbh5KJmkRU8llgwIcGtBaQ2HlXU84Hztev+KGo/pHf2iMHUfMMORAVQqsU8NyfB6OhWeL2H7Apn
6XL2cM/aCMNsutxiShcLPNDhmqpYqMiXRykjlgK9y+yKxBTzFzk/klfooGdxS8TubGtJAxuIwE5R
wKAUhalshaFLcNDfFGpfPtVOynVuUzMSueTqr77tLSJvNLNHL2MAS9wuYcD9L0b0XqFNU5u06Ult
34JevDt/5d8w+PZSGuiIdoRCxH5yMnFIT0JHkixXZvJ1jcAU5f1WsUZS/ECUZQxM/lyc6a4Q2QtO
MmUljsoa5goTH3alRqGn8WyOEE1TxAH/TyBu55ZHWqQ1CeEs+y+LrNKopCKKC1ESF0zgiCjrXdxK
LbZD3WRkHH4HkpAekOK31QTaf2PoJ81kfPQ7JLIWb9P3xacTqS3A02xhML5lC8bku9fC/UQZW/Ld
CRR7BdGO8k619O9olK6ah4n/WWgsicGW1VHgqbeIaRCvTZhKLtEReOW49ty3E92yf1csYnR5Yi9b
x8ZLTyVdBY6LPKK+xVP/QlAmVw6SpaPYglvz0VlUqjfXPVlRNFSg5np8vjxNbo7m5Ip3nJ9FFd3y
WSXTWkZ5SVbl9O12DYjDH3D2DDEyufwPsNMssp9/CqBIvdgPItZcsCopqc+qtCBBrM/tkNTlNKCb
8zK1jRjnYX0GuZqx4GlppkYFSSMxpPGc43ETrNHCjq3DzQzd4UH//Hq5uYZmYQOKetxKA/Vs7oFQ
Rq0eSTQ4DhcoWPqFwZAQwgescQT9iOoIqbtBpqUpnU7/AwCv4wtKzL3GSBnPfIPYY0hKPWHSiiW3
2DAlh9ngurZthoSnfWCYwH721liVZMc9cFTwjKg776AxYAINs07LuvsCrglxXuyBjeiHTT1ExzJB
FJftFN4B89iID8g6+SBTDCjjrKU4zjmGwGi0LHHr3NFw8C+zLfmDI2K1SIKNDaS9Xa7jdEItu+E3
WYkoLKkRR7T3G9Pm6ml0s1FKVfJLaXaIe2EwwtHxhOwjf5G3gysPaCEW/WD1yX3kx/RaVROkWx4D
8mYzlQWglTJifPS8rQquieIgZwb1PeWjjXMIlyxoNcJRRZt665yTbu0aswSYdX+p7N49d2RpP3Pw
a8C2nanGpHTGYZxyjfBBwGdUR43yKWjaakE4OUACM9aNk/kEal79GjDhZtWAq/Vyu5ss9PJWblZD
OosUOs2UTAXAVXv3y7rDyJQkusNEmI8Z5IzMaR0oG7Gd1c4gpKkLSthe4gYL2WXlSeZKaWAePt3i
pSPdy8mTtmI06dJEtDYNOX+SPOK/ZErL3zhRVMjeaq9vwx5RcFm8sjWfP6PqbDrowCLHFWGr1mqk
J4AAV0lDwLyl1nEH/lkIZ0klmk3KTs1ExUGivIheX/CINW1YQHvdUj+k+WsSmlT0V5P78U6d/LKU
UljsDrDiHUD0W/F8VxpA9+bi+QEOQNUhGavOYcv7+EYr6jECCoLpstmgpz2L/Nw8q6dpIe67HnOG
/0iXM3gpDUI//ra7iv5nIV10EqQGkPvm2I2VC6NGaBelQAz8kN5WSh8ikSL1o2KibNgkdnbP6mh3
nGmbmeXEBiTQ1l/Ke678QPOfGotFgoOtIqYKFF6VaEUumuPyTE1bW6yQn4RXcm6mF/8+dbaif419
qe+/KqBN6qzWx9Jwy0hirqhOM53EPDElSsDk5cr/vXztNDdViuGH2tkbMho/TPaKVvBXwCZIBxa7
JLWaF8L6CpC6mN7r6Lw4hIBtDWYNEouUPJJ+gtxLFBfqWso4FsxzGwVJwFFrrNBlfdnkat889zNC
9nR5nFRxYPJCE/FkRaAXKZqh6J8gYeSqU30cfsqo0EM5gBpGT4oBsL1V1kK0uAFjfD3xFjWGMKhz
2m530rOEUgmBmnfFqxmaGHoH3Q2z2ECdAVUW2jUXBvuzSI+FWY8ReHKPvhi8OfA3SA8xG4DWeH4Z
0txUV/5awedQPnRNKaByNXhSMHwRUjzQeHCaNNX4s+81izmQlmaA0DGerEy0GrAEF4Nuf4gk7hOP
NCuWm1v51CHlYeD66ecw+8wE5Fyar4qfuMlzJDixz6B2FltJ/osFtPCeM+ubUGHYcnYOL04YAF3R
rqKa0D5/ZwviJMvWPkQ94e0SDS5gEwCIS6kIpP2n4COyJWrC0gu2x1nM+c3wgAia67E3HtksF8/N
JPvOpF3Yr8S8muJvkLI+NRXZoFjtPHhNDalfYNuvZodjgPubMivlbsw0cBc9p6e1EShKYJpfyzYW
0rbtiYDYFffgjsoTjDzmyeJboroNmbHPcNVGhYhJ4KV22Aslet1py5NVTN1dT2c0wdeLI67iBcTA
P/J3lLCrnI96m5VSdI84qhbcssUzW4IbjbMinTJVgMzarOHPTn6o95SDgdsVbQFtb8SNWgcc4ewj
4fRy931krvUeFWEnvMv5TFQioscRsAqmCnjjAF6pKmUGYh37PK83fU5CpVobrhl8kThzaqqKij3C
op/eaKvb0n03fh6oWmPz/HiyxHXzwShRSSPbFw4N88Q8b6ovlxlUtI6yT66occ6OdG5GoYsGzCFe
q6bQ/CRQeRkS/iePKJdxfahCBszUfWGtgD9EZ+8+39u2bV2KWMcFOrczxAxMdiaGkHuOkNUXlfR1
1S5Zv9/oeyfFSuYlREyjU8mCbjWRhLpmy/Sccl1CdUkfGXfUVMf3Bb73kjrH9N65LhF1iiTdZodp
D0IH+68oTDNLJ6jv/2k1Umuq86eZGeo89oKnjwCW2zcjOOb7d/cLoJwTsqqXzJ2TobQIlpo2ffba
+f3JlXzXMNPAgt3XpR592dDgjsyFSXBGDz2gU8HW3WSg7E6hXtCzbB58IEzCAnlLfx8IYw18c9kr
pnz7+ytIpijvlXNcJCuVvnjLvGeY/Y96lJxDcYu3TvwgBDpAIBQ69CuavPfPB3Vq29zQAnteWFHc
p2cuDiivTEKITQCu0vpCyFYuzRyQECaKOfEAkAXYBo3llcHCD/0dfpC9p6SHPu1AVxUQq0uHy29E
21MBFSemsMOw7IdUShJyGpmm2mBb13qoErIQiTmKDLZ5QVFYb5Q0M0PZ+dZ2UBpwdi9HA/NlmnWb
/wa4QesUl9cpgnIBJ7UIQNySbZnJnhEERiiXwz6OkcQ+c2HgZ/9fRcajyu3vlZr7+9lphOYYlC93
qhjTkCikxOgvmRai8OIP4ENBVniXiw4icu26lbolNQZ27HtOtn/S+s3qK9YPAkHQDRr/jtLPvkAW
ym4rZBlROQl4c2FUGhfAPOa6gcZoW5eNHsOPpsPdGjY1sxChybw8K8b35xynt6w3uZrqHZ7SVuqF
btbHEEV556n3tqmHqGH6KKvo3ocMUIjeVYATuQKPovLdolSfZ4pZKpgXWkNWtUtZ8Ja4tSG/y9Tj
UB/Y9GOq+VLnsg6wgvfBnoh+6gZm8ay/mhBkpoJL6TgttWzzagXrvMRBYglT5u/wpVSR0NRHdYUV
NiAgdVf5sD+enAHOosBhEIAS3zBRqN+W7zu7LyJuMfbMk8okbXhCGxcsLGHWW2s/CE/CM6gWNvwD
X6YUTkYcl/WLJwLV0adQ7au3/btqkAKPQO0dbYrCr8QyGs/wVJVEnkPXZ6+wOi1lM7YTAPvtFgZ4
dtHb3Tz2fs/3XAtrkF/6P97afJ/nkmxYvDSCEPvYtExrzL+48xLSnN01KsDoJ+LLlbHL1g1IuEZy
rZ4qD7nz5GsBGknHMmfeovgzTa2hLJRJHj4Ujop6XIZ1l4Y+onWgeB/wPjySImgb+5O5ed8+9Xz0
RUWyM+0jKy90LxPPczkocNGilg92YRVg/oGzj1pwhFF81jaKXUYuK5yz6jX3SrCG+ogHGzD0QIEI
gq/zyrA6AqnrjWKCaKyIRTsOs1wll4wrTf2gTZ8So2LpU7wl2lfdBgtSg8p13eDSkqSp4A/7jbs/
UIphvX9aNpNNxbnLjw0c3j1wheRz0+fq3FV8rl+aQw+wuNz67aIwJZI1ouvBuZa2bv3W5svntVJe
MwSN2agmctS7wSXq0gJd0sPi/8D+Ai9jFShAAui7CcscX2XN3IHrHlVvtOUlKtEdsHH+Nnjd/Xsr
dLEesoFH5jHzrVUwaR0Wo8SiL3fGDaXLCVlX0pgzarrreSxWFZKxDCnx0Jzq36C1aX5ISXvgvI1T
9pDJqwh2+vlZv4LpApXE78sCswRFGX7Px8kd3BJLe1BH0fxN6ZFyb+VWq+/TYsuiygPOnhOJKjOf
Np2wbyEcE1xqKJ1jAshUMBqIPfAqMON620lC68CSeZHmbikCuqQlgQlIgSKm72GiLaristQ4Vtia
XS84np5roYDQyE2VJ3KFRKC6t3sjy66xxc0uJ3N3Mxi73s26ABBxaYs/i7BPYIYc9EodMb5Rxxpm
F32k2SXwjp/GncKi7UwO6ncse3TlYOpySXDNkr/oCcEuRfEcF/jFdGHfOsEScI1I5oYPE9s5Omq0
P8gq/JR1fsaOnQ3uxQsvqzPGFG+HDnwof8QOgbVJpqpDKtVzGzIYRpnQWyVqG2kFfCXB8vD2Ogum
e0tOW4soHKizTfQMoL5cZYSw7SFdwOvctAIO1XGGOo9p+idwZJ1IIHGXl58AHzpu39WkOV8eSUM7
ot+UPqNWDHiOOePM2+zqI1pk5p/a0d5jPMsgIXOwStNFP8CcefWtENbRrzKVuM0envenu0yJCQAm
l5z8PIfAJ72ZN2MmJ0rXCC1k1iDZPnleAY8F+BMUrgysdjGUD3FA6gAeUWMORLnmBI3evKYwkRIv
fa2PeMn2Hlo3BVlaT8qxoscucui2nEHU3E9kcryQrKT2K9DWlSKPRGaCJ1HJ+SEhRNUVeNQke5mX
iWrqFhs7wKaIAjGeWYBcJzfwUbc2kTg8D+gIwZza8rg+arMI/CjfK01WroyDTLfiF+Ix5rFfJMnW
Qx5TZzUioXqq8gmfGbCC8VSmVHI8XZOHjNSMmrHOvFp3Kn+th4kEO9EVZARpkfZGMGXxHlOqTp8M
e+G8DCrSNa+E/Mh3Of6mYoIrVxZr1dEQxLSG85J/Y1JIFCB9o10NYS5dXVBramai9/83rKuFwv7i
XWoP/RPUciecQ4lFwwxVAP4kLFp55zvhZT5HvCj5nySq+GCK6Q1vQHRXrycv5m46K3WfjvX3D7w1
sXmIoKabSuOoh/TCbP8zcaGt77Kv8+Shiil90P8RfHtyn/Ikll2ZZkDG4veFXqaCVLwmZPkymc6l
9xRQUrl0jRGYRNTJ1AbOzEGcPbKOdnzGfxBhW1PUrSbz7Ax6EepWzlSKZIa/YndE8xUW171W6s7v
ecucmGWhot49XyADKLLv4Lehaq2l1v5lVpBUGI9vu53/2jQxnd1JHgZ10ElUQmUMjJziw1U/03BW
o1Q03l3Vg8j+YYEFA1NEyIoz7xJ7yPAVlWWKe1maQq4xQfsLBzPa6OYNVjrne49cjGyRlAyUd2aN
Hk433iKDPbzOKxBMZtEfzy5/+KBGEOCrzTNL6IR+QafG2jlO7SgZh2TIMn+EUz1YgGNSqnz1vwEp
L+gCbNYrRzEfDMbZpynOYeHuHJVdUipVIBTvEkY+fpb4OUEjCOEtg1pLn4jvrq4unVrA0Jnhr4Or
qWjj18RhokxWpDz9SjPKQIJcdtJ9AreUxj5PnK+/pdnCs5YEsXatDzUrdyhGcfdohDoIRDDV9hP5
7nS3PYxofe1OiLbJjV2SIHJ+Cbux2vP5fSYdMX9Jsab+ve8FMNtBbPphk2cl9ZQB2/JS5DGUGg4W
uNGMxltcXgL2PkhjEP5ujmYAVBUIPFoQTT5iP/vm6L7zEJgqE0xzfa/b1I+ITFpYLC/K+sbIs0Ow
54L9y+GqjdSkXNUlRjXjmmEyWJWSe+famsz2Q/D7mRPa/FEqXYWOd0SxcNkoDgJ6OsqGi7/Wozb1
dOuyNLec91rq80MvbFsMzmidyECGt7j5REX41Lug6PC5LWfkVHHlp8qw876TBuy3PyQcJtxGbzoZ
g7bm6M3Ws4Cnh6EO2t8aVPKS+cbCoxXTsG5rSoDqRyS8XoAHVt1rAN+Tqb8cS/VFsmJDArljc5rg
4HyvaUvK2FveVh+9DuLWtKWmFjkvoKvwX9BOcN/eBgGL/EbXKXQoSxETfbNVtltsKckQDZUFKzpZ
E0tWLwEa8AISCPwzfysOiBnkXZ1XoltYW1OTvlXcrz3J5+zToqNSbkLI/KR+hxCelSi7xiO8ZZGo
TVCrUCihFVolxDwvSm1FD8e3EkCUhlQILq6Ix6cY6S9au3AZn+mNVMp8OqfI4OQPTHFVZpcC4cTj
pjLufcr2ObHT7y1s/+ahG0bkjJ2wqqQvh57u8RQVlLd4O2Nw+5RSdGUOcqpOfUO14kEb2DXxDSCh
R/Ax1gnbrwHc8UZFQkmjxfsKHk5mrQ78oaA+1CFTFDWV0C9fLQcNN0sSCDYLuwifka9w+8ZWH+ad
Wsjek59Fr8bm7l1ZqyyguUeOxslw02N4zfNTXqA+WLXbkczeO/IwVsjMh1O73o2ir+tI2jVRTjzi
eQ7T3IQBN5DYiahbwXCLdqlOALlhIDQ/WC2whWlGZRrX06LsS/1sh9DJcxbpIdVGdLc2JFdeaR0e
RW3bs9+Wz3w3ApUJ8Ll2cMhSLSns4wipBcPegrLLDsVwjFc1YDZwsf4zx4sSIFcl58l9wBx6DEeK
7L+QfvQFZ2JCg8IQ1ZShp6kJTV+DypJKr3vuZw7dHVzlz+mY0oIWnZGySfOVIXSE+p4JQrO6EGsG
4N4HarExxkSA3vOe7wVyvgKf85bP202aqzAE2BY3TAjNhu5N6QSsxoqDMf+oVfX/Bu6sUos8+9K2
yxFlR6VDNI/5XikmoqLFTsxgbWAJbvcyEg7rlVIgpmPt4pu/k1vHy27bQb9kN7T/zpmA71RRTs7P
JtrpDpJ74W+L2PiXZ5+n2IFqvVeE2naJqMZDbLbHiYk/OO5ovLXQAAmtf4Ibsrbtl9DjCfizXKZ7
yBzyZgZkGvH4yAcljZKQ/G72wNDGZYuE64F61FAxbGWW6AGCrUrbxzlDSgOorEAxiuth4kBFHILE
dYZY2ttt2ivLLJIgMAMO4V3wq0Toi4wd7fGbq4SHIBMVf7RJTBbxZLARz6uzPT3d1FX+HWe8s2bE
l4FA1KvnW4esT5TzCRjWAXwukamjDxrZtwe4NoDoRi6eERJvmQUARFILgu9D5QthzGgzt6cHIw6j
iBX/TbOhW0ME1K+2tUlWqo6jTxTdMNZBx40q4kH/zwe9uGKFEEVzBWHK9sYctR9hntt/SPvfPcUJ
jkb0Ni+6rqsIZe1lpLR1bjaivXJ5vEPuBHnzIZ4phi2QBxYemkKfjNp8SrTIwO3CQMhAc0J0raAh
xw7DrxZ/MrP7QSNI3GLrv91wQY7EV6OnjzKKut7GqFmw1duB/eHHvYf4XiarjFN3jaVGuoO5fl9f
GTYEYmvi1YaMGeBsD55MWjL/o2EpaaJl2Pba4++IXUSPpoh54PSoUQtI55myQHijPbcHl4m2E0iA
p9gRWUav2Iru3nAiOhdfdZo0T3v51r9kNu2Ow8WID3reYYbli2oL/H317Z1IssQMEINV+ScFvqnF
hYcCuGbwDj7Yd+2vzGT9JEuOhfZw97gsfRd2C/KX46GJtzkiQonMWapAWagY6dv/WB0XM4SsAPqA
vdjZm0qwPbLf0XPmYjgh6d3jNXjevlwJ717+ufO8pvGLcQWqgVEJtGhYAH3KfJkbnFjBl4v0ALpu
eL/37ux17RtXkK/EDJYDZVwXD8GVwOoIkzQSL9Ev9URB3qhbUy1MTpwYqMxc4d8XmPscEAXgHN/A
kpDnh69BXe0f4Iv+0vC1N1l8KTPe0oaAo5JqYgj4/R9fMCVdndJq96KO24QcH+rAQbLrzmKWzQdU
0gMhA4skYOQph7ryQpD6ZlslCGNX8Wp3ax1yJvdmfUX7iqUf80fPhIV4nsMmuEcWcozjGhVkjDoo
9Oww/RYmUxALs7FQtkbycYZYRlgWqvLotpS/mdyngycFUsT7WQQVdGDgGqHQayu7uWas7p9SUbP3
MA70DCMBD0g0zzYadxj7jmW2qokkmBHTvXxVJwoaNuTfxlXfgScfcNzR/QBiLf7ilW4Rxec8xgO9
tpoy9TgOSRV01ZCD/0nlqcLBoX3b1D3OyrC8xcr80tP666tg+qnu8gDZBnT9hJiDssas9Ef57Er1
2bnIMHCiMwPl6Cvsb5KU6oQxFxi/c1b70xgwKonxqeZwOuWmtmLArJJh6CihXRpZTtYBsqWPpQtU
25sTVaE4BgPlvPaZR4zQoDPF5hHgKBgPXMW0s/r1KtbNWU1l/NLXO0qqEsedE5PT3XrPMdm0u3zv
ADoDPI/q2cCVLbhp8+jgE20KaKEeGhOGrli26boAeGYlWMsRKstG/RIKKwWcC3gzOm4HOjC9RDKN
yvFrSfGg8NdghbvYfzBJjMMlIlCS2a8gKRUO1RltFB0jyHzg5DCg+gWdGIDN4OJTvnG57M/aXEIr
9fRMVywQgxINhmHa66zwsZ/VplDytNG6gsGzhORZK6V18IPtudIwS49VeI/TyvicUE2ykbCct/nk
QgxJarKsLXzm+W0bB9l4znyq1WWIcynFs90L+bbHJKPFUuP41fcKVjsXzNuaeqzpaBa0hwVMFGvN
YukZESjJoULync6tzbvXXd9kN9yj3o5x+zsLPz6GMpRNcA5rK5dmeM72yAOHPDRJVMn1vbiVrLUz
Tezm43v+g36lKwxKMdlgNg1z6t7P2bAirooKJpo/w/jwQ2P2yFHFQreDk6eJYa1AdtiNOaLdGwLm
S/1joYItubkWcF4IYSk1VrcC5H/nvY2ICQjcPIYzyOcXeklh65EfwdQIP9BHmdIKCUfsnvHHlipP
U2j4u2k73Tdcjsy6C2n7sMysrex8btsgIgFhkdZLLPwhccJCCKY6rb8KJINpWCJIN/CNBixjZTvq
lY0TmJ6PDkx49mE3iJWIowJlogdn3ZrYSvUrK5OS0eKy6BJFgAEIWI3zK/Z2nSgyv4oJqG/T9ZKM
jMZBHPRdJc9a5dYek5J4OZ0dLl4+Q2/z8Ebyd4xqryZ0ojNVh3x8SbHrV6AVqLYmCqoqhF8dokEZ
VID06DiFowl2pQOe5A1ZsX63qZJElOg7KAFFnqi2r6gOEK/yeYeWmSCXVKhbsIQjMwQvVnpOiwTa
8K87z1WDnnuhZdNQMqfI9shMVg8UWwKCKfFHY7VLQ0rYV0o0U/MjaS40GwlKWWd+XcKTcSHKFAuc
qgl09vbFuJ0vwyijCJK95bShzmIfNODw/+y4WR+2MqSjgfvwXeq3IpmSoLBtQHg+k80YkWzMdpe9
GRdEEdwOq2enB8LLrGrssONlnApAei4iu2x0XRZzsQN9WXbKbE+5pM7TuSP8KrNmQF1Axq6b1DIl
cYdvX5WARs4r8dOSJEByMlSljaWQWwbFWjQ5dlq6m0faxSi5mkMs7ocUkNd5Vf1eIAjGb5PHFxFS
8TRh3mgGtl6t6I813cFq3uiSBX9nJ0r3ldojv8QPQHy+k0VRtmGXLfckvQxBsNS8RDRjGA+qNJ/I
DLw3tVOMXToly5/caDPIg/wyiQjALwW+X6pY/8MJQ19xWt1F8TUXyvkcNnEsGPGompRObx3nk9v8
zqtEifObWXtYqcXLLC7Uw/LZISnT9bvxXKi1Uske8PLZB99/q7FX6ln6dSILebn51XL3eHvzBUa+
PGQFtkCBMk9MJWqcrsySHUcEmr1U4uN7cM/fC8gqIVvB4tgd25lzVf9aABHRJ0ISsTK2h4y7bP2/
BApuam6oMDWCXO5Ba6jSbF4k9ROfNGg0lr+btS3N8DldYp8rMdFMc3kjfsQKV7/rqeDiudetVgty
4Rl7u4x3ImyIt6y0C83bPGddUe5ZlsHc5XgDKnQl40Da+sFYBvHzCwe2IuDGMSvO4VeQziXFvFVa
tdgR/2GknQ1SZhn9b9Wav07dbr42I4fcWzg1Cw9xmoEXyjNFMhHw+SMukrTmTh2p/7FUhLXmtcLq
CxdFHAV0mb3fD87EvrAu+skxnN/HZEtGkvelVuCiOaj9sIvL0s2HsGPbolLQJ+gFYp4mvjxBadze
0oJkSdLq726XoWfwbtUV9pYHXgqH+hyOZp7fRTjuAcSDRZFX+fjG9Fr2+m0HINEAE8Jpm5YHK4PL
iPYI1wRERYIYv/0pQdsB7T8SBF1Aq3blCJTmbR7eVaKeVfcqcRlO7SZ5cqIW42PwIiGOTjluFcSJ
Qbl1RnYnqMc1SbPwaHMZLjWJ+iFecj8gR0Km4/iAezXTQcMMswiEmpX6G1RQagfp/gNxRfExXcAj
FNAXvXZ9g//AaPDq4RTkftLcQfL2zooAVpoawKcMa2XlMdRHMkWHzPAaOiwnIedEBmt94lVEk7i9
sZH1EsqHSl9iJUgDiE30fnwVNMz3iQgX1Ep382sF/GPm6srWBr5fUhaPgG+DiViTIe6OP+XjR4qg
80SgcAsslO063CSDuzCwtpuiRkyd2OgLPFLEJ/2opLaWzdftXq3OL+PpW+fJ6bXBEBClp/Zp9/zv
wWE8VrErvTxLQip5Qb9nES2+KF17vEu8GH5S5hylT5Zoz2h5u/wSAVzQnqLHiQwjqzH3a7QcVmBm
/ef0qcKJHzNG82yRgg3fCzJm/r2K28m1X+YEy+1fd2PwfwDBMAVqc8tvB9DhXZLs+U0i5yxPENPe
+tBKosTHNsilDCL+cRTwJoyhgE1gsjJmW7D1JWDkFng+6wFHae7Tq5rm1LXvnnFqMW+cuIrLVhwk
agX5KuBfyuhTUv9f+ufcjJE2gttzGykB6nUGUDAaF2AYZ/TOHzFTTuVvWGFTRrNiMc2LEhvCpukl
dPVjJeKFdGTXf+7NLThkNmzT9e8P2FDzI0WBRl4fPWtBYqwtsGfqGpoIqidapLBao943nOWfP0j3
QqGeiFHn3I5+J/rj/Fqyg6UA3EucORMg0Vue4MPWxESyOx28kAjmkP2lYMJJJ+XlhaYXEfuAE5wo
lvW4jLwjU/YAeKpprbiLS0jZlGBkmRHje4wijSYIsiatuz7EoijUxwNreWQrR/AR8i5HBsc0LmZ1
EiLMArH4Y5vZMUCVXTFKUh0DgixorurIiH6a4mjG0rXj4dRgK91UDA/8OCyUFr5iN07Q5/uT3hLK
90Y+6F0/WwItb5EDAkewDttmVMI5dY14oMF2H7lc7CwIcwP1OM57yl1QZtkr1S4XTgiTxj3XsZ91
LHZ0yDjfB6iK2MzdmjlBoZL8Zesc+tYYg9OBsZFmcRJwsIbwwr20DEwJl58m5jIAe4uBe5lVS9Ge
SR86+JYlstCwr3kFvVINFpkqE+sRRalg7BDgjn5U7onaL3EMH8yQq3GhHoVVZJhbgUtLp0fQDlgq
2RmWqRwX407wP5Dc9v+OIO2HFrssauska2IxSqpqrA+vw1rWAhgqnr+jx2FC4GeHL+u5uB7QViGo
uXFYXx70h/pvUUj/7RO5yR9nLh9y7y8m5U/jc6vumo7LUufyRHhONi/s+NVzuB2K4GVxoVl5p8uQ
zGgtX2Q4A1T53VRpfwk4dAcp+8FeEXqXtsPSacMONC3LeVsl1bkdIW2ujkQ0Or/QhzFF6UpY27uE
Y/xErhlJGBkToeVYSAFsTQAH15gdTdZcxRlpigny5g+iY2KIL9yhS3qT0Jl+T0IMIwBRamSkSScM
ac7ErEhAUckp0quekLTGQtEWNQ3hq3XuZRyVpt7FKKBLEuTTDAC7Uw9oYf1tiFZs87n7L3ZpU+3e
fRc7VTqibi3qmTFfCgXmO4MDgesI8qICiDo3paeFBXs70Kphrz3C76eYchNMRojqC3Mtwxxugzem
xxX3BgImYxajSgfVEuXGGrmc0uHcbZcSMGXeD7dY1cxhLIMk3q7iPqXXUGBUph9UpDnz1L9AmRMq
G605BueqiKVHfobktNBw82rN0YxRm4kJl2gMK46xnOZul6E6mmxOyYGaRSH/m8/qRx1XZajH9xgB
frceMwiSGoqhwkM7sg/tJZhAeeLrmowFtJUOg79rf8Mij95j50p3lzOvihNR+D/YUT25sQWnfX6v
o6ZKWGaIxSchIsElkHFGeA5znm0xN9uodU+SfvenU91n3f5EOkthjjH0ht8ZqeBMdgvZ+TI50KG9
11uShHBdTYNMhCI/oLtmoyS9eub0DN6jp4B1dMBavuFgvsfbo92Ffn0/R15OiXkexikW5JoxuCSd
WKqvNt2u5SsRvoJSRhOlpbyziRNESZpaLwO3KMwwRKOLc9VBGvYHrUQz+UaNfIxyKLRYzPLMwXmB
RSHSct/l5ku48CJNLl5GIevu6sD2GfO2HYWnwXACNxkb40tl92AIDNU2TIZ8HhN1NDqPdhxsaByj
KIrBZOZbscY+hLa6nCDqBs6vkQJsSL6USSUwH88pXVnH2N2ES2XqeN8dE4Tccb9qatYKujky8fSG
FFLRHZpLjI+6Z2g8p6oQXgxprpo9DHnw+Tl3FvXvd4zZmoTCOc3l8iSoWL8nvsB3kY2S13vGUwC2
2YbPijvK5oC3BqXoOAs87zNMIHnv7ilz6Qao6V+vxqFEoe5gcDaYXuLtMNavRnTHaLjw3SS+eNa6
wngS6GMFZL7DAJ4JYao4ve1UnKw7GEbbQtlER22bohk2+b09DNq3x+XesOZzYjHVAGGG1zT40kuP
EYsWYFb2kttI0+yFlcsMHUtzHLlYwDxOSzIJtxDXhOMHr9Pp603VxG7r2Eu9w7Wr6vuuZebkcjjh
pbQWGluLC9GkWjSVkAFCY+Hr65UUi5XkK7LAyuQ6/J4PSpvUKD+mOowraU1oKv6CrxNQg6WKb5s+
Omramn/fiWh3WdRVH75UG7ecFkzOETFko7hxGUkVi1/jRbrMx6ZHnBUeWL2gldNfZwcSD87kjiSd
2lAkNZn8YM86WlYIYu2GN9fVwEo7XY6unSjfo/zNXshenv9aGSefypcSlvHAhu5A3uk14YaIhQxU
jPdh159v2OwNLmC9Ohq1FEWUrs/mNj5JsRcFtEPGnxGIK/+ZM9fEhex+GHse/WYukYZ3YbfKis9o
Ele5B7vv0+mIRAvWGK0CC82j91IrHJYMdpmfpqwdOmq58DGGAzdYNP7SlE5WYW+rZvmg1xxMSFOf
MsX7Zbvoz6vm5FoigkX+xLkmpB7IJyadsH06p5pmvqUF7RXAEEAzVmJqc1cB6PtmKGq10tXXDhfr
6lS7IqZMmLFZ6r0Vlji3Tw+CLtD8IgEXkz+GD49x9UxIVhl18yxuKNfohFZEm+NBVgvmotHh1DA+
I+E7BTSJDwoYbGj1ALr0rUMjNUXUCpoy+qIlEQdb8aS0uVYza3TxoenOLSZ85CqF9xB7xvD3URE5
8BsN87sWMajXDVEdFW6qIEVhH8YXVTnPnuXWqsiIU4AwOgi6B0LWDmWF+3RQRSp0ZWCBurC/Z8sd
VsCTI0CLRepbpu9n5Yf4YHrzodad3zLMHhPIwUKH2e1BFGrGYQHla+AvGLY5V6WfNYg01q1BuurF
ucRtq0eIEfdKhGnjtJZkZkAlNayJzeVvrtp4IceHV1wy7tjz3SlL5/ksHklCctn4SqAVZR/pT59E
cQwx9WpOWqvonzKMSZxyc4mx8V1ZuLyVONvApnud193nJZ/TRhrabCclII2INPkEXTsTp+V8OQM3
kBiawVw59SqBECNoiAE4cWWjKl2iFjyPOm9zPLjcptpWmxP4HWhyd2GkqV0i7i1EdQ/rNQ4Ju7JK
ilPtAhqgEY2TnFvav6GzCeUG1ki4/3JHx9gfCtqJtRhAggkteicVVO3KopZYqxbFktbGl0kFWxts
M+YLcg6O/IHrmnWc6GeYUbzEYdJ3B/GZz9kYYArakAw8rqF/PpCUb1XANzpJtPWoblI9FSwanExx
5urjwV6RLh23gcvoj/ihctZUncucb82Ik7/FRyocYSu9E2kRgrIwn/CV4by3HzA91XYNKmrLQFAE
qfGlBTNq7mGjhEP8dV9LJqPtwtXcSiXkfq/Z3VT642Pi3RV/piGPS9jXnz75aFP3RvkxV7AAdGiv
bVMZwhydL9WVlJde8kZkfrP/yTx0NodRHMo+PHLQt/2z2phKcJWEMlqFPVku+IzQhg7IsaLj5+U3
Zu+Jf4VidIwNQXs+zs4n6XK/dwTqxHJ6N2ML2PBRMtQ2YHgHOPb1mjJ/N70znKGbwnnEQTh1NyPm
R7f5sC3BKgoa/Wpcbg8PlYh6gyBDA6clydGG6U6G4eQUJ9d1zMYU7S2Zm/U4x3ta5Fpe5ntFAJ8K
6tLXdty1Jt3mKw1eodWC8uSmz2ThHMlgvbcmr1igsWUgkfCOd6UBdRGbS7feXvoYRNLYwBLz1lJB
LKTRq2uypELCW2/wJx++QNzBq4GdD8mLqtSZw9dkiSKVjnWrUXjQdmYd+ObWSiIKQ0vZEr3D56GW
E6d1aPxvtUOqDQMvkf5mBFPMN7JXqj0stHi1NIkPPF7UVouitj7Njsx4P4fgf+vHmToeGdLneNlN
047ChHTBECKqqRfKVeLgn4gVnt5Q0x8oG/JscSJoCpTaQ6eKaWIpOv1Z5dKHYQa8siv8Y94QbzXU
Obvsv5fU850U80WcVNsbb3FLJQ5aqteuc6kQRYADVgn4gsyDSMi88mdXDqO/6GTvtTrfMtE1TQGR
WYLC9QZFZHRBzdd7ePJ3GaJAdWaEw3hLHEluA7dNODegG+kcnN2XXkNl4QYR7arGCv5+WtMKYD8e
0Kxl+nHOMDiQkq44C1ui7pcm1micqjYTvR58657xzV1axMZiu1Bzh8kW8unkUHXMKZuig14OYL8J
+rfq7vYJuUOkETsqIk1cv4itK2dmk8P91eyrG6tqPzGqoLWe6UwlEhmfap1nuYxylWHoV9izwM5f
kX6bBILpdZ5bxitmT0hooBowjn33nLyeFOIvKLf0MMk3I24nLNGiPZrYiTdC8u4mty28pduG9oTw
XN1dbKrww6oq6z8JfpJNw3w8GvWL9bUg2bbbZhF4Vam8hY3jv1856dOvHs3vNYw8/9g0YkrsHanj
YMsM/CmpKyswhNYXpZ+KuE6ZuVtX5iNBkBr9AXZR7tkiwR3iaZRBrS/ZRNXRFh1DY9oJubPAgPwC
tq5POF4sqRovasLKGf4hLswpq8vqScwhTnTsJ0ueCNf63RkPSme6g4kTLbRkulBlm5KeW/znEbO+
9mFYf20LlAPWUWQ9sEZJsLMIMm9hqarVaWeLCazF/sePn1u9DnFYWdMvluYE6vqD6kIFASTC4A/J
jAdglI4FQGkcJvg4qSwjPLof1nwYyrcPQttoDHrfgJpnEjSYirfkkz6j60DmFZjKXSm89YmYPaOA
xsUEw1FK6WGnWYGHc64DcA/4PJtizMBYJUh5Do4y8ijXiv+u/jbKnpsJQxaHbXtlN/cg4YpHg08h
DHXGxQPuWWkwQmBvQ1PxlUQIy/jBk9gdvNoObMG+mOwlvoCMDe65Zcm3d1i2AafTtNN6x4H20xNe
98yCVjjaSRqqA2uvD1+tgMXwemX8055SLyaaTN5EsBupBmL2jvfB8S9vmTY6LZP0b/OZbbqfp2Tl
NOGLXNx2UuwGXCSaGNtpk3oAMolhlgdAFLB7RsLi24E1y4mCswwykzXfhhdzt3h74QsXpXPNYdZ0
AlKEHCKnkrLg/q762NCikGRpgjkJt8HVVEi046Oz1oXnofabP+u9mKyWjuYRNqOcA7qf4l0EqQke
GrrSEGbxHxdlDHWO15WDXV8Isey/33PnOt5GwDSHAlhpMwwkgCDB2YBP1aqC/HLYxsq3p9nyIlS/
LzNWeYVpy44LaSYQESCANsjHDrvBIu8RGUVUS9rgm9X7ezFYuYuTuszUKHTbsjYm803BFKq//qfr
mstYYMt6nNnbrXD+vc4LZAFdQnoyLOvs4WUHgjB556ZYinMVCLokCyR01UVZRNRAn3hcx/7Bd/bL
5FM8T3jZPDi0wLQiYS089frGYMsqZlGJkJEQ3mSg0alI3HRaQeffaJ/mv3IYvYxyszjf3Kk3o8RE
fcuy4e5PjRLTRcfB+0N7hWBO35lVDn4/qOu57M44U+nZHxSCdm2f+Iyd4dybs1I9PsqcEa4crXCa
I9BoyMSmNjAiWs46YLLhHhEc/sfqvsVBq/ZDU0fpMFO1uJwtVDxIlaE6wSaxCu2Ruul+RwmQbjEN
TUb6xpezJPpCwR7nFuIHa2s9sltBDqwq210u/NBTNKOGXZblO3aEjp0hMUdWvc52tRnGUTFPzZGq
ZnbKRggltVvS+jAzhHKmCbFiCVP7+1gf64nKqiLbMtgMRC6xx1ER8+zYOlHwu9W2q//Ib36EbIaL
OYTwNuk/1MEo8AcGdU2Ece4n1p1QdyzwLNumB/UpYkqbxLpz3W+5kkJNrvEBLI9fshXdEkKWaCqy
VZZ3j/BlqqjWWtwqFzyhv3P+KnH9qjLcr7i3RJSDz2nikTo8bERF+07Is3UXhxrylH3n8PQqqdjf
R+8Pwt7b8pAsBRpQ/6cXdb/EG5rcQuL0Y0qCV+FCEKnb1qZnFmxJiLE1SZkjSf5R+jV9GxaY1Z3e
eRQfUhc5lZ69j4tW9ocDjiEiU0VlouS87NOhTBvl5ya5RD5DonKZARfLAjzVQwj/sMb6S/DNjlLZ
Afn9YGgLTQiXne+RdfO8RtBFE8kk3KR6EMm4m0e/tMGPLouM1imRzh7EyzMykrIjFXT+kXClzaFN
WtpgqYfrlKcxo7xrZsFVeayq2OMHuRPkkhl92A0JvV7R4SfdpealmLAgn8m16H15duhjMp2svmrB
fsvm13Ll7KsAYxhJEAHwyNcm2GzX0Z4o4xWIJ+zhWOJN4c6VLCa8jaVGD7FJ1zKXTpjmwMTjNCj3
TpecU8uBj23iQMv8h29ZcsqQSgW8rhZlqYbjwG5dckaFD8UMAn9ATkZfwPp/YaOlbvZVxg0rP88X
L86ow+dFuyiUGhMW7cHcrWuyNytDiGGHr5h8CfZTZqKa9q4LQWZXF/XKi9I6qdNbudYfOcJosDS2
0abLSsHpEuGgSK3VUw61nwK2JVzXEeiCEMtMJrp74fdIUPFSThZm2e+kAoacdooob36Sp/dKTxs6
4bDGbYrtMSNAgLm7WEGLmKZHvQhbaKhmvgt1+rDmgEbQzRT1zkqikIWLM0wr5o69pI2rOFMNP8n0
FhSWvZwEjFvUHK5rBWvq0PVpyJL7KfMNEQxH+tai6qYqtjTMTzvQLA0pZhVFFTt7HzX640VoWaT2
Jo633DUQfJxgg7i6HhjypTmgPYXcsDykGjanO8jB8kcQWSYvGgZT3okSNiPwtPmfZGKedXKHT/sm
5CF5SdBY04Xak6WxaHVsZKqhvpMvsCvWFf3VlqbFgH+iuMaWbjtqftPzb6dPiqNHMN5ob2fi/08k
Kb15ft9BXkz4s0tPa7Y1HLVDnJ+COBqWvWx77yRjywROdUaEv0b8o4qDWeSFyAoOLo5iW22LuBTl
wmaVIB8bVG++/vv/u69iK/Sa1hfWmW0MKE9AFETPa8NP+o5baoBWE4LURTvq5o7Y36D0jSBBHX+d
W1IJB079UpvKva9lCTIVyxF9tl3/PTWvzEzKPWpFTmy7oaVvIQa0zmlgURnV9KLaNWBGVwN5khEV
nn4GE1mxfgMJz5++2NLzUjnA1hauskVwaVfeTZAIGBzJV11QshJAxql4KnBUhkdsMaV5qIeUEz3a
O6yLYEkJi0MOmgkNzg27UE259ZVvK40tvvmOhUWp2rUzVr2+V81IjQHVa7L0jxaNTPwMxw0iB8tR
ogZ1GRzjYZhDSmXGfliikM5yIGxp69fQwHZm2MoU62Ispgh8I6IirfbHb9oIkswSu/YjOe7qw5wT
FfbdUgILaCoJDxvQSDApJFGTlWu5gmY0faWCmEin1/ZGWfx3CWsAz2jCiG8iP6C7CxO2jU10Qnq2
kqpSAXD2a7xUlWYIWp+NesHAxZUSuYMSyLIXMtL45WB8Zpm/9tzP8vmfW1ULf9s2HZiCQIMs9QUX
VCquNIZ+gk5KRs+Vn/PTgeoKWNluYcW4yqt0TE8IDWKSqCLrrhtepfOhIwDZeWBJVRQR+51X0HDI
Chqm2zMU7hcvaII70YjG54Wv/FS0wnevcra1m+gFmqFwI69vyjnoi9XVLAoV8U/etgBvO6Z4Iqui
dp4aAVAEOs/en2CIrGPNl9kdeHkVyeDILtjeYemWbrqIT+GOFeqEANaeEgWdWyymzTC7/IRbPg6z
1GiLFswgyd/nWlPOqt3g/se5OOuE1/Y/cxznuT+SPgMJMRyggTSpu3Jh9bn8hn3+awREtJ+W0ulz
iCftsLnybypjnU+pNJ4HolmNkcrlCuwIra0wBLPYF0bHvuyofv2Kp8tuDUEQg33mz3HZF0qQ6jVX
fMiiZn59rJRc8bTMAKUysAcHfrd0Cgl/I6pji7iXmhH7rD0QaqOxw0Ro4EIsx/1me7UUvkbpa9eg
NVYg41uLNY+qZP3z0C7O8DYyAZKd4uBMSWy/AOW8PAHjnWuPSMJ8aK/7hE/TNAdlFZVSnIMmbREN
WY/pMcNwNHjBPjWujj9rJuhCo8CUg/FyCeAaY8kOTtn3fJ8xR1bRhidEbtUvijhWnGNeZ5NHbdzk
flR2LZt5nkphzuEuICCkyta8lcHHWHsxTRwYggXInWVFZTadpIWAZa8WCEoUZWOd3h2sDaOBmuu/
bW4W26GmLovTPsD3OYfFm63mOU23ti+gxENS7DXXeYSpJpelGyLvUPnPl/bHDnU2vvP4ncB2GzXh
DeRFPcJVn+p9L3ByfA57tO2it3W/9GP6L5TtXq5V2RmfXY/hyU1w6hHIy2cyj+ojAHSmKgXmK/Ao
gXxMj1KaQ8VALtD9HCnPmdXkaTZyOvWC5frgucYHV9LOB7OxgHoqITqaQOP0mFQsvZwssHvLuL5V
Z0b+dYXNydIo++MGshsX58IEzLmg8UndwAYL6qijFcMJ0o0CKWlVcCLyL2SBrPYCj6cb6E3SHGuG
7VI2trBwZ/sFKNmwMzpWS9H6yVUkF51BaxyuZhRKd6anZNItRqdsK6haXbSeQDWCRkTln7Z5BLJL
mUrroD4BIhpAoBQ8erd/S/43JvmUCJxySry2YDdUj7eg/QcTKkLaxksz012XEdawF7dGeQNk1PxS
M/J3eHNt5MoQXqtAa2+R3HadLTtAoEE2vtwAhANc7XaUlAP9AOghFL8/W3MQhiOsNAevZHnguzsE
6G5GdpuUIAX11GYRLXM/kCJiTvOa3ADIMjNmmP5KBolVsZrKzO94wrTOvq+Qu9HjUI75NMMOU9DV
kumiGQ1g8LqZI/M+E6puPpANluVSetMIFzDZYs8nNtci2bBLSDT5nhg6aLhcsi98qFkxJbjVykRK
CFgh/W+doswF8HkkSYp8PZJZeoKbaJeLs5+6iQ0X5qlUreAmNjzSymwlqjDsnucHQLjPjWrtfvPa
T+9zyVHvU0EvmtTNxhbmLr9USyD44GtmgufF/L7j1mR6t2kzR7vTx7CNz1OlmwSYpfE56qeCB2IN
ybBnTvJM8OjcQInXzv+5WE8hy6yCA3QtR6treb/tPKGUAemqX/Fnovuq2WsX38FNH1rB+3tk2qWF
vDITSda3xaRaX1FL8nSLR3gbZgQC277g3g7z44vUAVXYwM+wMKS0sX3GrK2mmS12MhjvUu9giNQ+
JWWyxHdsNf7qE79xXvw3Zy34MhXlvKvgpyNljB9wNITK2RdyxBcZgXfD//rCAdfPQ42mesHImdZi
EonI9qAg2S34WR0TcNtT55QbAMyvihXd2wlHJK7KFVVPVDHwN07kEVbz/y35HY1GBylDBNTlCdEE
zhL3iXQvB2pT5FvI0EnVJyK3+DX1ZtTYmDpQ9yEtKgbv6WjMbdm+eUc/E9bSjwXkOWp0pdVMVEmG
P0cSjuBcRuk2xa1iq3vawuc0kHvp2X5vWPKA8c8BZ9WZcRy1GzAlUQcK3R5b1gA//GnFlO6i5qba
AyLV0+niJ+1Gz+ZBgWOSYS3z0T6xGgBthpC3+RShPfO0xe3tr2VBkihxZhkdyn9YoU/+GwrX6uLe
r/wVmfiJOmx7pz3ecHGZhF7svWSehLCMpIrypibeVGyh+f/Jyvqq9bMxBiA7pGsJFD/zvf31nVCF
99OitVt+U0HRHXQ+09tr+3ML+l7/jcTRbautS+9CcDTIgavtkVmGcr4EUTWkFlRPBYA1p7NM5o8T
bomDRjqpczvw3bCqBzplI5sAGQ6cL6dfoFVWV4bxfDKtDJWFJhdAckFNEtpQ756EpSGf6Ugji0Hm
2AgQGf9rI1LDgqxe3I5cg+1wRHWwoG1iRNJWfMTsUcjSrjTWWt9utLrdlbohbjyAJjZkdBx2PDWo
liTopXlPTV+guzHailkLCYfMzlIjczk+Vc8LZ3MO6Qlt1Nk3NNgPWIGS//Qzi9TwAPfjEfCw6sgt
YdZrqvsP+st3+1K+bTm2dw4ZVPulXDQ5fjQMnNrIeB2871v+aqbyU5fi879qLA6HG4+v54H8iq8Z
QW4D/iIqu4ITR8tACuQnBS+i9iPwpsP0wDDjyBsp4lfI9c1JODZQYl7+bqT1TbELReVPE2QKX4y6
uOwYRpnSfUhoKtZqiJnzuBg5jPafvKVAiYDe3mUyA0z6k8PP1dln3UX1EvRYeuOPBBAZgVjHCMyB
8QFx6dV7ZKYvObdlEaJiN7+ABmaoyuxz5At0xMxtnU+PHc/GxzeFet+ygqFlpdXiSg5BiY9sQFCP
JHy3a2G7xTl8VJEqencKPvLcjk4QjTdG+CMCODyLOfcEDdmdfVzekuB9gaHkHEgGM1BuIX0JC3N3
Uimok43IAcgNxghZmRvwSdYkOMxDXktx0hX60aOKB4vqKNnSAyCHErNjmyJRrQjXMNDUVbjhkQcg
FaX6pNUpGHsb/faEocmAf2xUmKmfQ2ZQajUqTRA0ewZSKOF9n2GJYxY5GMqyrz1hx0bZ8XEOVfs8
JLGvPbd0S3BBklRcSi06apRutRD8gvUpDR8TsP32CkggfziLKlDd15n01SYu1Kyp98f9LbThAHg1
btuwXRjl6j41ruvaePZPzp83qUH7Qlrkdy/3v92YoXG+bvF607SILI7vYKijRnjgM29NAJKAOgJ4
BqTyKccf6LGPWEC3V+LKWqK1pm4bpYLgP8ZhnOcemydwFBC9iJ/j6/S8FgMBmmdCzdegtFeby1S1
fqPfb0Bf5GOtpfJTzO8So/1b/SonTCTi/iWzO6fXDvrkEMWg3Ne1J91gP7RkaPS/7VW5LtuFl+MP
H2UyTNRGtc6A1ypZyHwAH4gHlA9gkiUi+Saekmj/1NQfzQQcVTTNLxOeBgyKH/wdFGSrl41EYfTk
bGeNZ9fxyeacfxmgiJK2MAnNGtPICg3fA2Q5PRj8njTu9ARLlXZetZkByN3Wa1naPuOq2gL32f3G
rFM4wjrbS7yXlMBhIf8b8zG5dWfZh79gJl8aFcC8X5CLahqkPQM5UxBB93YtGByBZkGMerQepZiA
J0Tw5QexgLmdN6a9Eo/wrBQ+efBB1/F7E3S+56X4aCunD8L0F03Rg3Q1kxHGLqSKgHxmbsXQqmfC
le/ekfYvXGFexOCSoIcGzbwNcP1F4BdNthqtvb/gVjj18TUUHyc0e4C8EZq/bSiro+6/IyP7MUL7
5C/Nyk0fR99HhpLx4eCww9Lmc113v1ll2+95ZVrS7LxiVdDLG+eKbWBbKMnWdDA8KmMX54DcdZrk
z4iPYZ1W8kuMEEF9ve1lDHyyoYBQ8QUdnjPHxBoAddvEHZZFiJN9b+zmhYYCnTRiiE5aZAOKYv93
qNx/j+N6SUuokExzPAfKvh0Jqw8tTobukJ/Wvnz/uiK8MFxNTO2Hd6p0s4ELyF73NPrQGKy4pISw
XFIGr0TJxj7L8n4jKsgSwTS1ZeEgJtcN8ji3ZJ5ejIMh+tiM2WYvqdeXO4FHwl6a4byCHYk7tg+f
piMjEzBAW64bVKdX0xSHuCm9skrQLmudazY0NssjFHvXkUbPGrrlfJIB5uGFuPFo1Rp8n28FioD1
HakoJ2EDoe67cKj14lWAKgOAwAZ+OL/qJRty8eZU+Jh1SVhrkNXKZfWFnmNM8am+mzMY9T5BP9S8
TfjIRBRHDxecvyHaKrC/w/lXzs8x51ItLVsfyCAF5/mxCG+BmtS8Yy0TQD80d+QmoucyXWbp+ZY1
LRMEnecD8R2VuVzE/vi+qX8M76TUGXpp/RLpzChMhCWpgvddvCW+ZNz9x9BuabWVzLioBOMSnul3
4rfY6jElHTa1eruqrUYjt5t+vwA8KyTaRKfxzLhnPN3x097ttHorNrqrPotrPbrPzTVDlV04Wqg4
wZrNJJR5y97UzUNGXmPCvL6UJ2WolwbT18E7h0gAUEurgUWfetpLXlnKBoEjPGWUcPyOPTkObJdU
HTfcWsgXl91gFAiF6DRocCW0Wa4ct0LZir3N+Q4Waa0IOsqSZHonS8poeMe2NMI6aX5OouWAUvTo
AztSqPAl4xj6HdaQSmO+A7M23aC+BAt1bcf3YgkHipd+JYV8IrXgYyiEX7CI1y3xYmJF4wjzwFqz
2JSJsMGQQtAVEUPybwRIkiybN912uGM5RjcS7Ux8bIrtxWc4bul5qbcWakAhnAx0pDUlMnH2+ALu
3qHICv50c382N8RD3GQFcTL8KcoqV0fhA0Rrty8KRM3yCmsZXaZIFISYaw068lJLBx4n6wCwqnr/
hZCNGw8T33maiwa8CgVyWhB8rfPGKgAaCM2R+RHyFruXGEmYfq2oOuDOdVLhDzkltbLmJyj1b+PB
s3msm8PIrMwCGMo0P1VqSQKoR75FhHtIzw1rivicmSls906rGvZEGrN8VofeqanAimPipzPGPG/S
uXwh+8wqj1aitYab691nCcPwxQ466vJSProo0cauRmkIPJ7qWAruSCrvE4xabiNOMx0ycijctE68
XYlByEl/tytMJfklj9lTcyvXOaJxgCeOLo/aHjysEDJjDZcgKcyGgYw+QZsa0qLBqEaGXNCNBVtr
8nfDqD1mNRxuNBUHtl0Syl10TK4kFt8gMhyAcbT0smKUgukiToJx9ekFboXjpq/vgd06LI5dPiQO
yaTKz6UC96bgO8lSfEuM5Zv6mH0Y90tbn0oD9BQNFtIt0x5jN4pxksIWK36l3jBU6czLJXwZc8SG
2JEesVmdM1yQ+OrHi+lnQ3+st06pFveGOfq/Zi+Z2eMyCPgrvE4lgmsskPymJqKeFe+EupdMcaU3
EqbXYlZ57/SD2KqzROGZNnuO0Qm/amD+B0sbQFQm6SjYp4bZAXbGlrkzdnRC79z3mAKxeUluVprA
RGPGNzJVBdI+jEF7ICg5ruBinNaEHiQOUeOlO18ezWv9gRdL/ToI/yGEZlCMcBVnqR1KEl4vNo0h
y6pvGEiM+pcR91f1rIMUFMb5A7jd1NivwugY73KMsaDp9rbOzwdYmd1l11SfQwNPxVcmZW33FOyK
OYe3GPE/Z/h3q8YkRqPr2lTGB2O5uRa9xIztKWyHVy8+YbOfubZS6hKugqnaSJH+O2UlQUo59NXg
ReLN47lrhYsVLEIDfYZExLMDronNFN1Z7WS8lOvsPKbC72JlkQ24yipO5ltvXnNVEEucfAiYY59f
ttwYLxi6yAnESWEbp+Vs2vNE0joeo8vdw8lgMc6JKj0YfXtPHmTEafL0UPsSPPOtbNLEpKroVbk5
uFEkyeHwAYY1RJDv1l2qME7xkRnbHk6psz2izvPL24MICZ6Sx7lTszTRA1OuauG4Yf893M7ht9sL
Ki6a1gJnm/JjAlb0rJ4HdilRgFcsOG/JgVbdFduvioVF82dDTHoQhukZlKOTf/cMf56wkIOdEa4L
O2QeaK7eg3wcHImTAfuVAsuLF50LW105gV3E8BFnDYY9qJ4XXj8/sTSyMzOEFk6OpdVQYJmZPiqD
t8MRCuv/3zk3VoLtPRXLLgGsvUJSJ+6Y7smkvfXZR5UgHNZRPmUsqZ0i6ysb8MVgJeHzyAOzPQo3
w8wQFrZXd8QjqVQMsUAyTTDd9Bj+XNLeqPg9KW4AjSwC/3Z/XI9jMJxlyhqJL3c7CoOBsFdPtzgF
BzRv344gT67esN3wMMFYYP7Jb+HO5mRghPAFe7LR8XTPWK2kfV1nHARHO8rM3Dth4u+2b4bUCLFK
+L27IOapAA5p0z9dRa0dG5DkMzd9LBcUFOBoEb89KERAa0SAQY3xJt5ORjEz73jseAk3SfRKUxnK
aw0ILjzjC4Eu4TQAMlyCQ8jCXyyk1CVUzyEUh8+CAIgZNJ0SROtvkxQMpg0zWAch0UkNYOoXfixm
RZ5l/49eg4L5I8yTx2ubApEohQJJ0hW5FEEMdly0TWkgb2DJjXwtoPz2Cmh4/wkPFmIdXD2Kld/h
Jx58CM+CIIMrckE8AGLJ0uk9k8SbtLkehuL+Ma5HN/jOB6GqFbBgRoDnaRyzZa9Vfm+ZIbQCNrFB
rO6bhBctuBLriwqz2w/weS6Jr45jQ1fRZ7hfyoP6rhVeCQ9BCZYFglNRF3Qi88odJbJTfe5TqIbp
OWeA3ClLy4aBigq8cgoprVYBFiDnnm7C31QF4rYOEKZKmzHgN24Wm6BsfxS88MHAgw7sc6H97jGo
XixMIZjDNK5Q5kUN0S53shELwvDnv8+OZtMAjb5gWTZV9tfofU5FG6uQvwjUi3CpifoCOWj48Zr9
yq9FvCGbtO3lRL/HNWDlj7eKYsOoyavNoriUuOKqWKemwVgnkY7reB3yVHUaPmYYcXi7p0aVzYgk
vdmcuA8SEUy6c8+SdI42/fE7I6v/fwm/NGkqe3PEObVoj87or83bz6ZAIWx/ZUfz2aPCjMAtgApA
dZitYMhQakPx7YJcOfxRh3Xd5DAKxXFkrMNjG53F+JtDsOL5HiMG1KDW5QzhVBtrchkxeJcIfL+J
P9u0+rtSWBsUar6NclCV0tTFEhBMJ0qoZ57zjuqURR2WhXsf9YkJV+2kQLblSGYwQnnpwrDdG37z
cQTmx1IbEd6v4yr96EY4zxG1rvENQkTlui6wYlXJ1Q7NDU8XYxKul4r1r96ruacpJCbjvXvUl/7c
F4vz+jGKHepJuozYPXtt7rZAyDBYZb8Al9bQlLPZJX2+6Z1wBV+MiXFvfOUIjCl80VJWtZXDYndo
wGp5EslM1EZg/MA6DLej4C2W7yy1qQ8W91m+dmaxZ42hXchAf+wdRUYzFJ2usrG9J2ksj0E9uj9A
nbKguY/SBYkguuFaj50gJGHQ+1mCRcYBBOyg12eIXVG1rRp3wrs4lOVAh9G3mVAiTYMDSzkAbHvU
L2rgH8SrkauMcypUrxk3+I0XQuLXatz/TUsZ51eEordIZq4SX3XUvufnEm4nbUFbIPIAPZNkmPyA
GE8BJXV1h7+3ctiWKB2ny+CXSEC/+b23AdnXeNOpmjtX2iiQU6CgDT9/rK5PJ64EvuEVmR3xAqJZ
zaLAVlIkdIE7K3MnRkNX9ND52DXicocpEEerj255XWKERk5Xrr8+SBb8/EIAZIV/VlFTBrj19+hQ
5gb/R4N6Nw18zK9pbluq/uimmNyN7ZMIXnlqwgerL/kWvleeznMC6/BSkjcZuPqi859ZUlf+HYsX
F69bIJdv+JKStZbI/Ih097MOPkGoenaVFMB3TX9xaQ/8V/ZdBmO4y46KMa7LM5pUjiwHDmBlGFKw
fIFR5Ch3xmXsHmN3x+5SQTe6GuTrpCKckDqUPz0qmo++upTt+NiIq6wYdQkJNxUaA2PtsprC8YP1
22n+6SOaxsl7sqxUX++wZS6LwLDyd2dYFhbWZLFN5kDkl1DmgHOmUev6roUOwMmdTszZN1MKFH+3
0pkeKL4s1lJsdvl8Rzytv5lI40Bs1LlyOpqg7CJTcllBZfTnHEFexxa1NUDgXvZTML0fGb+/NruL
oqE5atqvpqWe33rz4K/sA00VqhvhjSEPlwCyWnPrB1zz234ZuG/tC5hw3P89lG6ZSfE0OR5rQQq/
3LAHrvFAlJVRYhWEoypuHT8jvKKX4Y9pQNObpcPbZwyyD6ekHEWDWW6MGJAi0wAJCbVIeIt7sxRO
PZgtaBMbyqsNbLm4yYCB5bFjSn8PHlurTtqa+4SHOOZWvhah6OVkGZqDbTTIvYzfsuEiDtnTQRiF
zlUHCnvEyYlbpA6tSqV3I0CK1L1pTOZhdNUm48TakU7Yfn+bdQUoKQN5N6med+Fa6NhBVtyuBwF/
veNyIWCzrByYAB5mxV81FtlnRRk1d3D4Dzy7KOS+uUxfQg5MWL/doLaU/3muypu4cxswN0hsz2tb
ZBFmuY/MMUW9FSLXRFzw+o/blF8jv0kCaaJASwsm2X25rDDTov1a6T2yR55PmjkMIsuEegdT4Mh8
NhQIOe3R1oEaig6GHyAHaZjPZxgfVLfKkVfF+VQk6mbe6xyoG1YpWDH2L8aOeZataSACl7BNlX20
XfU4Spa3gymnV5a3h2EjAWlfNmr0Fwns7ajkyIbQSz0IoNQlicUkoTfXVDxBKThAN9TE3PMu6oH3
1xzgUisNNM8v1cMVMXlPkEbsvDXmMnMhli8QFQrZlLEz26UEFYnsR9RbLd/KlqDOxRXyCZdlAqhn
Z9s8o6GMQbozY6sXLDlVA7SSHL1TVi+CRbfvszlFYIVRHGFTCU2M2nBWSL2ZJTCIMaajBhk7dcXO
4OPZDfnIRjfxo3IEXwbgEAMB3jrJIDhT933wUHNxkVop8mue/un2tZIPzzzxztulHV0LRUjqR64e
scNzo+utyunDJW3JpLH8sJ0WM/RviBrwNy9TYi5llK/hIsSN07TtM5cA8c5nkTWNCin1Yen/tlCs
7Q0tA+lPNym93WhIsss2fAAXscpxkyQmA6psWf8BAoQ6Wo8ts5KgtoFkmghJCPBkjjjIvHtVo7Pb
pJF5mnSQGCsh3DOym1BrJpI+EgAsTMK/UmWtVrOqG7LYYH1IECLtmKDZVNxbsG7abYeKgd+tehd/
2DJ5vTqwtAUZ1Mr9eiVNeV9pm+TA4kc3KWEZdKjsMGw8cdZibnLSWy6oBOR6Xa5+qLRKHgF5sHl7
++X/wVH0eXoMcs09QqAX7qqP+RdGx428Qrz9teF/0kpf3kD6XYMx9eoKifxWOg6feyz8a1oShaiL
jsYOBunJW1vRNIxrpcAojdn8WSWeRx8ERnA0G3khHBbq5hRnvqU9jINBeXRRF0NlG/UHFzdcB5Nu
/9YTHnNAk/LxFRps+3tctx/x0NC7HYVtLG3NLcYHdbbv4P8lZ/WzGikiEKNIS18dWHMlmdQo+EWV
Ipdj2fOIUbDy7Wx3G/Z5N4S0TE4v5UcJLBI/j4KeFLCrX1E5TocRRea3UhAIkVmzEgJk7oXL4pip
QbWnVA7yyJcRLU1p8rYXLEjCrxZJBDCwpZ3DEcWGcuqzy0csz9m1PK7jrvGvrkJSYDdhIurR6SN1
2Te78grhnLsZvSL0X1WzWHT/CkaNn6JQpIZDOBiq3hWF4RLbSDZoZ6B4VGQs4gLeHDXo6hoxC39Q
wLGLTqoz0KSjClfqbZb5koYloyN0VVwzgP37sFxlNjijVCYu+3LpmoZXWcxTGksTHRevhaGp6g7j
SAiMPDd4GTrbKW/T4zhoFuq35Y8yMLIMXrhZ6r98I3ZKWcpw5+1mh62bLKmjRGCGuGUg9jJzIZNX
DiPWExSbVhnPD4Q636mUSSKNEOjl20p+G9KWEKfeWY3xqb2VN8p8xBBUcXUd/4R5oCR/LZkoi0kb
1BPnPpp7f6AcAIEgkFm6Ceja9/ExCEAmFCJuBVvIVUqWZPwPg2Ovlg/JPx7SCw5QcD0I0us1Ik5J
LUFYDRtIxVwQYXxAdyDeR6Zp0Gaap2Jn/2C270B0yr9ukfRlfuvIZVKJ2f/RzMl5VppKDT67bhP2
anhjRjk/nbZC22l0V+i3+1/QgmySBSVgbmbPtidGwWZVl9vxkhkresipOiyrE1yeKuKqKwhQicfx
6TIWiy1rKLiR7EFgw3ojcQV1BbC+Ganhj/vfDdOVnqoq9RXAp0967yTVR6jNX9RAMSs8YvaPFps2
yVv8j+/GEBLa025GQUQZxq0a9uq2kjuwn/OO6AsFE1ULBrDY9rjxVxzYDStz6/I7vfUxsthgPr8N
Hu3o/rFmBTKTBb8FpO08XduNsGhwLv7ik5B8XiQOQfB9Jb2zbA3crMdLxvl9Jg1ncBPnX9//iwLU
cgSGsBpAa6LhW9JqVfCKHXuxjabdlFKN3XK9RC92AEdZmLyLLQIKiJWk3MD4Otpc8cMQLAkZxRo+
9LM1vKoGDA/xYScR3Dp33xYq5knjZwJJzCsH7p7xpQjVugHizuFck3DP+rPh+4xWDUDnTLVPaQDy
Y7R69vNtjrpHNG3+gZIcjyK6c1KL4xtDj/F3WYI4m89iwucI/pR30ToUhWGSloXiZlcYY1IQT7v7
PMd8MNbkx7r+GEc5cHgWAPpPn3oej3H3SplULD48w4qYMWW7eoKrTRyEHvuxqinDdt7hlCFi8znD
8W2jpoEsAFiutD18Lkk+zMuES9XNvkYa5bgg5ghoASVdXnuEP6FNwV8ddzHLX0ug7yXSoCAZ3PID
mZUqUP2pFyoYZMonvpGupIZxsx+2m777V5GAYja9GGM4HPaqCEM16HDH6qBWORzx2WB6LaY6y5Ey
5x3sQhX5BPuFNDkmkz8gsRmVEv2WTQ4v2D1A/bvr0XSfyAKYXE+bHhV8xf+yLJrAo6pT9jLaUMi/
1qxxBji4o/34amRAN7bC4qQdHaENfosTmHxoENiWXfd44NHzR5nx7scPZxmRx1XTV8vkoPBQwtb4
D2EyXRjNUcxcgDj6mAEb80lTVREZkxJXMf/QQVVHJF6+QjFD6L5nZ0KA7GGV9XHOrEAcWYoN/qg8
+zEaUm2MAmi70hQ4M2wGcGtvOE1J2Zstsvo3YSbfySc7XyJKjbWG00aCrIzysl5w+ZvKq9aAYdp9
vHq3kdCiJqZOzHsegLC/+3YtcrKw2Qc/W9CWMatuwI/dgb8t2grFxVeosS7oJknwZwyqv4bkf+7z
fg4pNCMTBmz14JpBhUaGVznXFOGeXT21tgOoI3lEhPL46Ikg18L7rqYwWebnuTGBOJqzCHGzBsAl
tyd3QYa2xIz2p/7HAVsyhaQmp3+nyobyFWOi8+lanyq98jOvcrSyjsAkoNZyzVwH6WBQYKkG5ZTG
jWuAjpmZkgwr/FVE8RvQQORJrR9wwASeqlAWsUSZkE+p60eGqhGKHUcYfZTSiBU2k3KPoYhkOokT
HaYy5HtAtfJApT514m+RZ3MTvbIB14L3BDWtkSGjFQEHsfXFtxjWr0GBSS0iprXU7XyUzXGwuX/4
Z91F6vGcHi3EIVY51T7varL+HBBV6wzKCVNQVkL/F7EPbHc/F93eDJOLfK2fI75M7KVy44eDmUY4
SanCyM230bq7Cbi9HKdiS/O0VtRtxQbJQ9YPD9MUUjfKKzKjifQcsOMU4KMLfqWGcpO4UgCzSHpg
3wY/uX9zNYRYI0dEzYS91W5fFIr5zz+Oym41AlIyzJIPHU8Xvuo7jz0o+qy8mDQ+RfDg+lTf3ezl
bgUAIcc9r3JLb1wjPpaWb7HIWR2g8Kcbz2lIEuD+KT+jR9aWL40izSDYOjtSZxXGC3PVAvonfurh
oA3kJgOH/l3Jv0a7paGnRsX7PStMljvKxl0GmQxGMZVxrrRskoebgHVIWPpsZspctYWLyXUsMYQ9
9wLBY3XfB1N59Ud+pxrAMeA3PQssvaYhPZTj4I/vtserHOx4hXes4MZy4N+EZQ1F5dTiWArCwaVw
0xqR9/eJEBTccipexq9wGW9BU5ZsliMVzVE5Zu3tARtoBkqU2o/5/eOB5dVJ0swrZJ3rxnnL6bm0
aJb3oHpKHXfMpCRTRM453MOtmLzkjPhIOQAY2UYClbZjo8rndRnpeUpE+ptGY480VmV4Fatc3Xb5
nRmcMTM8lLePmsAk0/D+DUlUjeAPE/MDPEyZ0RyETe9JCAk1+rbbbD5Kh1BzakVLS2HqKLtHMrSZ
HlJpUoIxxm4MyKNlW6k6D3OyN6DUljz4TkxntuvxPjSzYJwlupNV67WIkXBjmdbXk6868QIco4O4
RcTB/4W2AdI+LPvOijd336nqm0PyeTQal8GAFW8+fztDIBewL5S81svjgyP/x8ZAKrM0Ui92ti+A
1jUJ9fiUFCYTxZMfMQo7wPlwAZ7+TLQdKslX/TmuVY+WxP9TVT0P3lj3gn7DTtSyJX/vTfO/0pnK
mjbzetsuvpMWg4G4XyqcCQvVfJQIuX/Sc/wV/nI4tfoYqZL+EMZT8vbN/BuDvbbCftst6pSfIzkT
6N+vkQ1HqtpuFTM8zYeSp0wY+Bu0nilZawsIFIeOYeeRWy7GY+KaMa0zT0X+t5UkE/nziUiUzE7Y
T0lBAgypyHqetLTLPP5zyGJCVdcLVKaz62RqiuLynS/kJoqZYobac5lXwPqlpDmlPj0lrAqRp9zJ
0FUbs7tuy3HsnjtViBzABjlOebtaqczY7UHcIq78N8Qo7LQXP2Cwb2KIEtB7RMYT+IoxbkUkoPUu
3kZo83lZPzc8cgtwYWREYvNsliDsINr/xw3EiIfDyixykQHYaXbYt+ybSzFqmKaoTy2yg+tw+DIV
54OKVRrjKlzSKqVo0onuaD0US54yCTXPP2aJb9thszdSJEB/zZYVKW/3Rupa4RLcg1pJG+IkHRfo
ES3z7kHcpxUdRaZrOYuRXwPxbE18izbNpA3FT0SIveGPpMIbC9WHqyBl6K9syXC+8wN9FFT3dR6Q
f2bC18OpBDt7JUvFElMFa39dlRB14m+KdKH6kkQBXx24qM/EH52tdcriFCxGRUc4uPztBOkh64YR
qPHK17eYKkzfSeK1quL/+1jFThut5rOConrYnLYrPd+1O1PMTIJKmHN40eB7mgGPhbcH2c210I5h
6hSY5rFCWSML1cdH201a+SZcP34zTzAQeslw0RvAM4N6emp/iz6hSskmqBLY/dw0wRIOeIOkWXkb
i5UOS3qwlTT5dXSqbBvZcOMthBSZo5IfdvTi/IKIHdygioK3dkr7uEEo4aCecR3Odqayj5bnuUvl
a2QnkBpw29gXgWT3yxilEjw2fE2gzWP+UnZqNAwmLJet43ENx3JeobFCtmD2vGQTHPCg4OTs2Lb/
cHvyYNhMEW8oN1fu4vHaQhb0JWTtRyVTvksOMqERsLoWLXy9HvkL0QKSB4Opk57NhPXydKRGsABf
N6Y4qqu7mOp/2ecM5++rGkMvzHUL003pu0f8fWiRo/ZdLDDy5KD35LPvAQ8sbOH76Vzm6yyBBu1P
K0vdO7w3qAydAhd8dDRkvpvuSDk1avZvzPSJlRukAo0PyFWQtpFW4pZ16oWtApvlNCn4a3+LiuNG
U/U2vvxf+u9wTG9tKW9P7HaIv9olIs2nrsUlUruxCmKD6wYggU5I9ijjxKSarS22TnMpVDAOb90s
3PQDL2DsmJic0ysHZxGbLJ6vVtOXOCHtFTw7PVXwhPQ/g0XT49fmPo/ZNQjbdzSfWKRyBeq8ti1N
nOa2k/4NPHfDDeSccyRu+0r2DLGIs+2kLjWUpr+27mUCoeI9PjHodHiQZUeRJM3SRHzGuXER3mGR
8l/LvV40OPKcO4bFl6eAibWq6hAly45rdZ1a/loFdFKtBZctxhMiVaaSBTEukELyJ07vQXUZOv6z
Y68BFDvnWVZW8BHwjrMBxg5LvtxKJauRnTWRsn/GTwcVsugCA2v3nZXxl3verBC/nbp70Cfwjo5k
qaYcFFdBMcOLV5QLI0LgYESWHm9vCgbiLXGYCl+OjeBWMpbHqiFPw4DLP7v0enPhWf5z3rBPMDFh
GO8KWVtzVwge8dd6wo2dAWsvoCLXiXUCASTaYJxUYDfiQvrm9HC2tBNFilqyg+ewyALpEgk4W+xJ
U/R5R+ZZZfebN3dhqTIga/cbdK9v16FmJeScs9LawKPx/eAFBb46KGQTbzA1vQrrhOE4LGbK4CsG
TDND05A+a0pScWfIl7meFeg7GIt1SpmKqrymkaXIEB2ftMiOj+lrNeBvknpYtc5M5s/4LEXFZfx0
P91vjRLJSs7/wghjZ/Ab9bpJzkxkUuibP/R5wq3EAHXbMXnURxbXC9umimn4CGwSK2zviJEzSaNb
nV06Gfq5L6YvvOex4Yo5Ej67wECFYyBRT9G3QRMd/QX4CMyC/9XFgESNtOd2dX1T/6lwWJUAglfx
byBMx/BpPouX59dwoM7H1G4m3xpPm4QjEYEC357hgS04dFkSkN2zHAx47k9nKkJ3AMRWyGX+EaLp
JW0NtykvOtat5cN2ue9SvLQBqCH/WNGwFPBrb4dSJ5oV7vp91zGBFne70Ykw4uOT7yHOr1hV4m2D
QYO8FX2MZ35IyDqa0+e7E/Brmv0BYwE7BvBAzRqGT1WJ4YmB7uvPbiBKlJloLyGf3QP/AyX2JeI8
SQonAzktsRILOPMFUWoxGmHDGinjBLSdnosJcad0jGrECrlH5PjStNnCFEk4z2X0ZykgqqZqPetu
lavnjoo9vR+Pcyn7IVQ3r/vGoM05P9YiAhvT05Fq/OLsy2A8/SVYLzIaHd+KOY6h4Y5P/jy4k5Kb
Ln7GE2iuhugKsSgbpTk35SBPCwB/TIXSuKe374WNLO1M1PFs+KGAWYcSYJAKn+7uLGy6RXyPPPk1
gZ+ArjZepntfxZrp0xn5Prx4R3C5Sffej0uRiHev4AifCpmxgl4OOPERXpk26UmGzMRROEFey4/j
xY4kWmACqCc4RlfMf+KoHucFgvyn7Ju6uIX5/xw2bGtQgyL4VIkkkTE4iSuIgQrf/qgH4pHqxHzi
y1VTNTnMR84+mEEBo+GuSRIWPwRMDP8agXLJUmMUKoZiyAZebWAI+XfVlZyrWRSOon63ATsNafd4
LEXyt/4GTXoBgLHNI45WBVMWEEVtUz5sx1nOkC2Bme31xuvG+v8QHi/FBPPfdh3b6YQ73P0aXGYp
oU73XuQL+bTXJGpo+NefTjG+wCH0MysllJcInnsCrmMXeOqzIjMTr3cvqIH6YTwX5UT/dkAbcoLC
BJRSkATwoEhIm/7LOGVY6hOQ+MhQcgK4WArTMkaqraeNB0OZ0ZpwzNk5gT/Nz4mCXSbLzwqfPQ9/
Xa5Wc2G6l2w6+ilRQapnnK0KRTjNAOgYheknghZb9UZGMrBiqWP9MJ9Z1l6zoKM/9bWXi3nspmPk
21Dv3icd8PgpO/Wj9cQbXmd8eBW3YpqyVBxV8Y3qW3bPtkYcmi/ZfBFlzEe9HdtkNoPz3BguOa5H
pPrnbCi/VqvVBCuzK35drclLaC73n+PIJYUT/YVIEfJFZKSdoJ9nH6NYL4qT09b9JE/XqsZ6ngea
kTTzNG3o4+1Bx0Na6J3f1mmXzESf6YR80pJxgQZ/V5ItHFzpnYl1eLDtHW+v1roxDqIiPJrUmFmc
Qw4d/kMMbhFShIBVgZ51zkK0jY9Pnz/5dj4orhl7ha+LTmt5V0SydmZSjw7nulqJ54Fn+6+GRchE
t3BQ3HhenrlDeJjpQshuKJ1LpwkQJ4hsHromiIChNxE6DgBUlwf8hT798cO13qaPQGbNQLO3+E3J
VSlf5STm5ufAro42RRQVbJqUERX1uPD89yC1F8pJocfy/VpBxTT2zdwd40fP8bwm2V70GpMUKYGl
/s9+ObLTSWv7gkqgo3Z9Aflw1FIbfLY05LMTxIKmB+qb3hqRH+8PcFUETnmRHyIi850EgHSuMKWT
R10+ZGjzVneUTcHNplR2wGcAOG0GOTYq3xe6ePv2SN6JUpscnnOBPKMZ943HsLqWKsILqiIyMi1v
Nkyo0hS8zkhm8QdNags+2pyBBdIp3uojjMgajCVAvxRpkU5l2Rhqd9588g4EMCUH9QzNa8bXz0Qz
anudmlJXlge/TZVRCp1mchjCk7D8dJe5dYr0g6hhsE8eMzZk0kQ85SJNiYSXpKRW7ZqydmLxLAH9
u+VrK6EHx/hLDMcweWIJnILRV94IPjP1xh5Ie8aLJ+gXgeQHjuwUrC/tq6VQjWtpArwvrfd+ufFm
qVkyNsd7cQn++GeWBiXZ5E+br2aW983Oo/fGJ8gpE6qDXd7A33ONfH0VF3AcsxM+Sn6ViwOKs8Je
/uV0b6lyjaCih+f9DxDjx85D6jRpxZM1ouQ/Ri0JpP2L4jRcySqMmDUXy0EPhNZwEO7UBrJc9Dno
0iyH/uicxLllbNs+RBFQNhpa9tKd2vqCRaC1kvb4Yysk/oPhBAq2DIkifAF9bA7e0E8aSuNdCR/c
VAlX5rnvn1reo3A+nP6E2hmuRHTmGtnfrAVVGkuLlgh8b0L4jCOZWoByVoiGCoPij/GZUyAZoWm3
qqI4t6JsdHb3+vyQzvsaXN00DwBNMF9Vs7z9BuXBHHXj+sn0AwSceqhLDoeXzz4wAJQk76dKoJor
vgVHvcF6RfoYH9EA5F4jPZSFX2AawuhdJQJp9YrTonSMBIYxzcn064G4LvslblNWNmpRa99P97Z3
0d65tYOtOtQ5YU7Ms6CooeGzoJ+WAjfQeW7NN/fyfZHpuANCNEu+EQTwkuMNhNL9298/xNxavuN2
M515uvD6q8ELWeIa6GZNwVdqI6Y4t/myoQLnVfEQdxcEKf2kPHJrY4fhC5TtyxKMt1+AfUwt5FQI
UaYWyfr/2+a+8cxRZkj5rrhDN9CXoa19vae2V0cJyotdI+Zs3JXEQfuTsuAQ1GukMhSTUyHnRji0
wAOG+3jTKMfDaXqVGwzknKMax6XM22H6uO0KKdzb7dlS5fq0bdyIrBX1oFuCEtXNY9Y9plFLgjo1
jyRBtIoNziVap136Pritjd4KabP6oH/j30ec77OfLiJdAcIQraAk3SqOWMh9iOpYDDyiiRtZA3TL
aSbjcrS5eUzQhU3TmNLzO+TTVif/0i/3IEXg7OTmpkpsc8Xzzz85uyfUdR3JtJz3Pn6ezlzodrGX
g6doTs7VjrlHLB1KQcX9DeA9O1iqFVIftnv4J7+T4JfIsGi+rxJ8RTf+hW5YHBAaD2j3nu8XVD18
wKbrEgYz0U5bc6rJ11+kZSvWqZ7liy3k6OX35b2e2tHCkeT5BHk/2Qn6Y5Ylr1eDfdMYkDyvOqtx
nZpSXVcthWmnAkhVN7YbuSPb/REnW6vHY4w7Y6kpVyq4Cuun1QLD2DhQBiK48ILo/iL5OJWHfKKv
WjkJjO9Fohu21KlNe/wPIDtYuXsNwabvSEWQXxDeTLqM+tcVPKDctcYjz+C98jY18iRn3DU5UvqG
7s9Nn6+kbJw7AH/L9EHca+wb1gWlro9u0K1v4w16XqEZ4a3/KUYOsvDaAXufVdMgWuYiTAe5Zso0
hYFGZKbacC7DsjwdsPkxIv0DM66qFyPBeEOJxHqyAfjIY4L76jVv47pQ0yfi3lNNYnnifBl6U/1V
xH7mfkd4TlTxz1HcxWusIeZ0w5LtdK1ZTqXYx4D4UhVyzFBReh3OcJNPxDw+gSpyh9GknQSLm5Mt
mvT+8x24CcpszlwImGHU5YnndyyqwdmkcdF756x60UZj41i62+/Qdg3C9LzB/+3UWcwnRqq2ZJCb
ZYJtYfLXsq15uw/yzEpe+psf6fkhUnTQgbOdY1vM2iumAiefBL6zrnAB1VMBiiAGoCa4Jlx8a/lD
W2tWW7Jy06nQTvRakz3gvM0m8E3B3tBPa86IgkrvlVPEpuH+tRc6Ol2eb2MpPunlWKBkwKkGbEHI
5UhLCW2Q5V/bxkyWJ0P5yVGa6u2wJb1w4MgFakiSkw0kk+3hHyPkjINhifZLpe5stzvDJSD+fAES
YyrgNpUjjRz5CpRXiInc2AQZ3Oogn3Hvkr7GWd4V3Iwq0rMjQx1G0CyUubc3tc37POH3SA7cdKko
7YYT1jpxeKKBi6ROX71SV97D03kFVGs4dX4RnuTBZfOieeAoEuMNIhdehheQzduWMcFoWzndftO0
drVyUaKsCRflBWSnjPn/FR+PylLIDtodpr0W7VUCqGLI6P+J4QlQrC3OWwdc9ePF8B1DyxPS6EZj
S7Lcnu/m1ztEQPb/vbUp1tOb/Npvy0BXUVkV6JoHryP1z5iF4JHCB57WO3Qy9LiH2GVOmtuIRoDL
yLQVAAKZg5Sf/nbSs5dToTKdk+AfzzaiNIxzYFCB7JgaLKBlTKf59V5vv+sYqCTybUiy2oodlvy+
o0Vq9cjjm6ZnIFAS6El8HnvlRN8+irWqDR45hJnJsfJy7L2OoBRucmlXtl30vo0jmS19xzdJtP18
m2ipu7GfG78uhre2Fr/lPYXwvuJOJHhBreAWzLhAY2/nn9fIn54dbk+KePF79RWYx12NBZws+byb
kXJXObADnGgwGSZAqsIuHieNDKOQREbAorE9h32W+W4ZjPTp0ukyEdiMrNicgQR0j4Of+WleAvjQ
B05K9bS28fYzIj+0usKeFn0a23Jx6bD32yUj91Yfb1Bj+QAY769HMe5vcky/7ne7R6C/VTVImwEr
JT6X9eD1yDc9mqlusNWVH/9usnPV2TNCDHGbkkcd9m52NL2w1zhpvOY449EPUXNkSNWaoiewZQka
ha65+haYQVMLYM8bphzKSoN+LV3h4jfEPGHOEmsxoVBqqtIOMI9Hhay2ahs9PANcQXCRVs2SuUk7
xOtXy3VyAiFf2i74dc8TztT7aAZVKdMRkEIddlQhtC1gCnL4WNfzu9qdgeTTDz/FBVf/WG6ppXb9
WeGzpR3dB43f25pkK7A/sWQ3+ATb1USc9VdHfDAjNewA1i7UoyryK0TY4vLnBPWFFXreoIWGmhrR
VnFIeP1V1U9FTGCSD9mnN5TDJzkvfs7Zge+Xqk8YeHGsa3U6q1/j3216eeQHGehdT1QgWFo4SUYi
IuwCwmxz23A+pD9E2RBM0CJExKiGcp1o8jW3iFJxsqIm/BBQ4QFGky6kChK08umLWr3xGV8DHxLf
N+3bmx0QwGx8h8T18oWH7/oAgggN7FWZTOBDHn8lzTOXHtBEiiaQZMFegzA0orf7QMNqwleo0W9j
1pJRSIC4L4LdTPmgv4ojfIxNmcpSYpGN4UmTI1xl0/dFOhz7yUoUadbjg/hIu4Lsv0Gfdt+c2rVM
Nei1KwUZANmfPjfkDHWar80yFBTWbvZg93wlO7N0c9kOAtB3/G8UVrl2+ilK5/jjjPl8OEoWeqW3
s5sQCtKe4U4FwJPmOijmwM0XhPqavJ9MoVKpAbDa/A1o7stLqNvQuWzV+S3gMrLMH1RV4fNIn0Sz
cd1sVIMoQZMraJBywKhR45LLfQSzQ2be2Mn6BiPilEbrAOVakFlzE0fhcxvNDV4fE0VuuOfCU2Ve
LrpJwThlbak4dhLHCSKgX4B8XB6MauRqh+yrCrg+1r/m92QrSrVxS/WbIF3z7586f1xmv1IKmjIZ
VxtsExTgHrEVApQ1oxX/FzlXpUwaCIKa9ifV2bkf6bC/G+wvBZykgM2ZBoZ0jbwhvwYgJlNmZQ6a
NFA6xvIVxMkGAOajew2zwW54cnGrNGyqWMtemhW5ez0N+8Br+3PPW8A7AHgeeH4ZqQYKVnDVxcOu
lWiMuDo/0BEB0hFM/WSvUN6YOK+VNQZTe6aum0gYs+gE67CRb05ugNr+OoLjTQalJlLy4Xlb7aeB
5VCetU/Iekc0lJs4TI106NCngthifppRRPGyvvbzMsSzWeIXFQUUhMyhyJG1xTNJkK4S1cHUw77i
bisF9xTxw9BepMqumEEFdX4V30jU57W+3vfgAwvOcXN9/6QTkDxVV/vBFXHtGxsa9KxB6SHFbOnc
4JjyoGXdvstRGhIPg5JAmjUjBQS1MgH5bQ+2c1pYS+NrL9Bb2qIsakE0XtrXez3803u32pGq/0y3
G7oLPfmCx47uAUpEbvHD4EyFDZyqYqKPteJUC1uAjPeT/YtjNa0Bz6vusbxlp3enLal/G7Qk32dY
jEfgm+5QXEVGywXDPVkyOD2xeSIv2Uggtx8qDmaT7yrQqKqc4sSUeb45aW9+plk9Zo+yKrsBBV1z
Ba2wW+hFtQXFF/ht2k7dIn/1k0N1yIG80mAyE69mdt54lKLfb7zoA+4BZgyjoteZFlzDC2Xz5hM2
Hh+V69hQ3ipXmIf2oL6lXTi+YxmUxBAyXIzxv2X+zi8upoZas43l0nOQ4o97cWtu+/tofQfwLL8W
SD2n4rMdcM0M1p8FrsX7QwzjG6lvQiRYYKcImy74A8P/AbiA2sikrMq7IhjMNrkecQVmqp5lyAXT
gQLYirOFucP/5noNmxerEClvnoRB8LfZ/DsizBwRpN6dMZAWJsvFMC+RDP70OZRTtqmgQPSWnmS/
ijR0cfcawFIBLCAzWfRzFJ3EVnz3kMW9DfzS01K3arIvBKQafNV5NYPFd5s0AWQivgHSAF3lvi7T
5sDlBqTThHnWVxLZzsIQUV0rJypSlXV/mxYSv5ww1Ez2+FTVLAI6K2h5azIIR5bbIosJhOCWsi6w
AXGLdadpiZGAfd1eAzBsuzKWBAqGrU6f3ZxZb2beQwnErnhwyHJTco2iCyhYSqhnpoUpxFMC2zvq
lUsMSWUfjERRk3mii6jioX3v03cuP90Jp2+sxATzpTGp6lV4oMDlKDs/n6H5uID86FP0tZMC7wwg
Gbr2p2n0Wfapo3hihwwmi/gh1Vraa8/yfnCbi1mm2BSdSK788vecZ9DuRTk3OArOAgs/AsQ+jpVG
i1AmeYDCjFUUcUNBocGG0uiJ4dfgB5Z5qvtc2U0wtWCn5HoCPp1cCjqS3B7Drr6mK/PNABCeJViD
twQKRvKY2CcGtDNhSzT/4qxZXzbq7ITXI9choEH9OayoFXEPiQnSX1tDQYHY5FvfhPdnhJ2JtP0Q
vh4XpBEAQux5hLd/GHaQ28+71Gg5FiJJGtZoFyKsMiIpq7iL4A+N1WhQLkDKzZHlvZcvuQgvZlMY
wrTHWeR4tERXcdLiYTVqjDcZOa5z9oWv18U+s+9SJ0pN9fQ6NKpsk/49uadvy3c8rsvura4UmMiZ
JwCCSXmiOX4wRHxocWj7QZhJRp6TUqBfu8is1pLmFbOSRPD34wSOMrQFMWbTl/52CBzebENS+ziW
4lOIDLfEbtSjCBAX+SdHWXnRu+HjNMQxmM3dFoT/Lxij/PFmm1z3r3j7HMMlhyHQ2QbwXs4vSBF2
phmbFqOC8oiriHwxVl91/dgtbCKDCvljwdifaoBqMZiVz84i9+mbFErh/JVyktFp/ux6D+091nw9
8MWZhEp7wTWiBYa2buNMW7m/0NRerPJVoC95J6arlM+13UWskY+24vp/0mqe607ilJLaHdRkbm4L
aoj0gLGeZMoQwo84nhBvCtsgNbc4fh68DRSNxUd6P2eCE4pVqnX8PeyJA9QSJmC6VBc3s5awFhVI
vPiUA2vUCGAXs8JXtdprIA0+K+OvuJLTq4quLFQ73K71rA0VpkmV4DgjUnJoW1pJLvgbwWtJHvaQ
mvtmz9wJwW/G+YvLCVqJrYnN96rutJM9iHM06oMtJjiYIglW/3VWJ+NlkKu15GDNGv8ceYgI6Om6
thYwPURS05mbcCT236JbmbhmF9pbUes1I1ccsZnr+4JRQYzfLNmOl/AXil08YclgiIRkEvTXOLVm
2m0VPivONHlrNqUkJcQzRT35b84hXLd8IYQevSRw+7+Xr3vfeQlO2TxGJF9hzdQ8D91dJEvNx1zI
QgKwFdJlrj+OaE0LeYMLzN77lwACVDKkGCweUYcORr/TLLkEww2wde43S/J2R928hkQK1hOtqUvt
WaO41SmYSyYjJfHL+xt56aYMfsG06pJJqhvCw11aSAUs6lxBNmZNTJ1IG3MA7o9gDH1UB0No7eDJ
VxJ+UbkRxt3sXGq3skJkmAF4PH335KjsJPC//ppcPlLTVUo73rcyJQw6nJzKCuj/HJNWORraqn/c
FhhI7f8RWiACBgvsqPqIckBwIsNxXLZb+vAnsSD+rj4hD1loVtrvuRczROu0fSQ9QxNz6oVU1eN0
X9qkKFjMsfAsu2N4syt414wvJrrzJ/OjeHHKciiZXQM8sVrGRtloo0bIpHtnoI+XirHFITfvrvrp
pNsR0eKLLYLa0FW998vwappz3CQrB87OKyzmE1iFp87bXOAxpgidWODKh1DY/gpohv/3cRQ6coj0
ZO8trHJlMob7XEwq7TcVg+MpfBWIv6vv2n6RxzgwFzDFX7lenB1L+uli1pgPe/vVs/mAfAx0IWPE
UGbTXJzI5ATuTpG6G1NriVLM3a2owE9EE5Qh6cBF7Bp5+NV2qTmKH6oP2sgRZwnSLbvG+rYat8fo
2LpZv8J8RPZrhAyxN4L8/x7XY12NRl/gnxJrprogBAuewQ/61nczewrHpc5w0AfMG7NE1dyrUk5e
LaZuhlLBZPjzV1v+uunFAJB04t61kiucb9oA+Z7EsO+5EEgIXR41itjqtcg0ya/iWuIZ+DzWNXN9
Rk0w1/D01u/k9ozwQGWXvspkpgGC3ArafXBFyVda2ZANPonIzpHb1De7FtMTjk6cx73fm02KniXQ
1udW+zp7ql97kZQY8Hrb2SHZwG3ZzlCxQ5b0O7o4ElS4KHz7uXefuGVlZFIjhj5tAhoAh6+aH8I+
SJ0tboqK0FMuMYu3cVxf4rt63u8+hVA6IpPIBgy2f0jHKNuZG8xhDW6oqag61E9z9oA1lG5XK3ZF
rdoYpw1HVty5nTAEb9l5ZMj4MSuakxqBFCZS6kQcrpc1FGx0N8vW1g9fDE1vqiA6pAb7S6buZtOg
AnupY8B0TmEGDdwdgJgDn7eaenje/0qDBNlO3JeeDwvCMg/tIlHcQB/uQs+9nYXaFTMGpEfWcrbH
dI/pQyd+Ky6zlgPycLCut9dTzLTDcIBkouE4LlUJfkqprFM9jgarduo2q8OY2mffivsR8VtWeH1l
LykG3SlDOoauVlRzNhZ+GsqS62hIZn+r5b5SUlP+kGDJ7yLQR1xCYfxdNHkXECS3inCwVQZTRGdh
ei/iOEXGz2Ro7qnsLu31S698UyTow7W3cAK6cikwWagnVzyT8P1eML32a78Z/srVu19c2Q4s5o2H
L1fyYLdxbYjatMMtKQ0Km1UbqDVweo14tmkc6NB0TCke5/DYD93Xl7Kty1XrsvKTLeMpeBIijqsk
ed6CypmPOehAn+bqGKWhb+JKFYVeySlNLxvfuhnqtGxfOvxEJfyDxsoWC4YnUCBjdgmavTgdDof9
RbvJsrGktCKNb+2cWaIIGnNce3QJSkFPD2Y0vDFSKmng7k0M+T9nqlhzBfZotu8l+eZrluJvIGdQ
QwJUcmrExjxTdQDIUMO8oFIGtIVpigS/YEs3M27FGQAzVWrQ6663QGoulU4pd0yxf317ORb+FWro
XWzl9m9gjiPUIaVrm5QVjUnjD3zpmsILKuXqtFBYbblFP49MkKCqhZbxI9Uj2l0YaIOBPiN9V1QE
MCb5Bp1gobG4jUUG56rwntzL1eXfmKEg+gtHaf8V3G59ajY+6QAcSPjwGvuyac3bW2Q7RHCf+DzV
lQFdQpSCPk/J4bXqttJhUF2Zgw8eubVYuIDj82JEiOWMyBn3CRHi06EkF6n11K2UJopVUGxNZLPW
fauV5P9aNskGdWqzIXT/Dmk6VERnZR+/htZ0hjaEkHV5Q8/W/WFs+wr8lFeLnazdMK9Gp2srKW7j
nLB1yLxOYPhKBmI7cHzpH1sueQJbzUcTz05KUD2Eu8tOkT/sVjQ5lDvwEtn+9qUj3FQOCpu4cRMl
Xa9xNBaHqByyrXKr8brkJ9xUMAyfRDOrPzVf4Q8+LfoRQ+v/iZqB/UIq1RXapRHJ7pPN3rOUFR6x
URJcm4YvGxrITlgP3Wq3nq0QAOtALxaWxmzPmpREgQ6HDTe0lVXTVw5aDeGhNZ2lou3buKBV5GnT
ilUJM2hDHqPZTFWO5BPDKa/+NHJWwwHZFZYt+oH5xmjJF5vDUZn3aliY7P4AQtVNemot58bHw0+c
qp404L/0//wfZZO82ujIfdydRyzQ4niVMhA8ctFgxb1W9ZmJdnrtT+5Cwu/5+fgUbociVJoqsfnB
haDaS+SMiHDqIBnK4xg4327OIuCUm83bLQwGT9DwHjU55fofVPcTfQa8oUTn7sR0TDjQS0e9g+/m
uBHvzswl1PiqXFQJfO1whqLa4KoRTsSe0pTxqGXi2g07xwBDH5flq2mUenz6ePCUJZxlK50YWmAG
C00zPxnY4OlkntkYKNwPWaWyYr1Bx3oBfzzWD/gdm45Ie8eAFmBhJ/2m4vkSn36xEo+ARnU+uTGi
GdOGa9me3DvKcdfqOgm82QzRDr/gVCMcexMsSu7xyu0eGmdGhmGOtXRuOD7SczVV0usg7xfCER9j
Rl1HRGa10coqXV9hzwPJHiO1qy63j8kvU0Rsecg+tTexCT571fRhDmKUnE4xyqgbEJ9LSK0GJss4
qGSZX5LfKtWNyxFtHAMLb1Kgfv5cJfOPHZudBI+ns32yKv3yPLmEHm1xG5IjxvAxgVd2mXlzYpHY
WF2sMgl0NN5VWCSXny3r/wqo8XwcE9ZPnbEmDpzfT8fdQ7bPKu7QMcUy1HSOYeIWBnp9m2xmGM0h
fcqgqMb9RhbFvu5oZZ73Yn/7AWPS9M1NW9n3j3cPHmm5rapEuGWWq+E/jhZHFazOePlNNKv++tIb
6DcrvWqbKAocIGjaN8rsBCoAFUBrmotYbc6N3Sa04/DxJep8tSiipTh5ItvMqLJ8ZYT0whysJK83
LxtOYILMEbTlodLOclObg44asCeYkArW5ffih1dOF1qf+om/0/6fb/ihNbLL2qPAtFd6n/F4YmTc
ifrYMZ2GVqUmWk9rNPsuITFI4HKDFoy7m2M16PxENrRzffydGtchFK6qUoCbjlxSbNXab+bTggrD
GynnFbwJJhXAnNd0iYokzzVP/dWXxvSUY1AoXjG7XKANMZ//LZQOG8oEshOhJb7mgcl3mALeNH1Q
qxhf5iSxtDWRGK37Ys4X1L8uxx/8M9++7YTMQjr7RgKzXyBFjtwpjMLMPuJ4PtD4DS7Tqw5jU3u+
LqQeD+nTh0LvSCaMVZc5byyiJZtfdhy/hH5kLZWsdopthPAv9ONkClo84zvyGP4+bKOVAHNdZM3D
E7sLDfdUar/24KU2unDt/Q7dnpkLGpgEechhAiBaYC3JV/6GZ4qIBthS46TU4W4SlOXZ+SAV6he9
eFAn8JHzoB6UyaI/wYe/r1+XN/L+jAWIpnzfBwHctSPEQqQEvY82/RhywTjixfL1Ig6XCdxZQeQK
Cbg6RXG299WyZpzz2m18XwTJPhwusxJ8geSSjOLYtMdiIRKhBjdlGp0RCekcxiLP9Tf3mclN1EZ/
6rX5TurNRKbdZHWZBMzUTM98lvSsdDYYDJ8aCD1XEuxSFfUXjuTYjkQpmQequC6bXVOKFeSRvf37
sXI4U6imznOK9A9bDl5OSE9kEpUTh/3+M7gXPD1wXaxtkwHMQwCb8uVGPWa6bqXacvZwkk40Vrb2
tjsrQHU//so4aGgNAvXB8LtBvNJzAjU7tAyhEDp9KXFDb7kxvIbgp2mhDVROSLXkvSt2pcmIRWO6
L7o5NBZRCRt6+Z2x1C3bNR0OPh4Buy7hAvGf3+v3o5mrIezzIACmhzs+axpBHy5Pv9mAtTxg4dEh
b91X0HGMm1fDuPoP0sY4GLk09gw0JJ2TAlml7K/N2XXG/4ybn4A1i4TBmg6dB57b+jpXqgnmG2V0
0EwFiBe3SOTNqKtNGIWGlh+jLg26ks4bi4+3I7q+WuTE7Qzmnw1G8BTDWfDuOtSjUVxPNdAfxkLC
jHOWq0wpJxyCVv+yYalH7Lp3yau4B1C6qT01rqoS75NiO9bXqkqi4XqrHQDjXThdpBdVYLcnShKs
Xm+TRam14zSK90rs5nHS3zcmU0svFDZQVkC8TuYihqmcEUHYY0qSByc9kmNjj4RFUJOzB6Wz9ftb
VA3pVvCmQbNvRy0toNgSJdXEP9VjAETKgLTHAQs6+IFm1Gyz03M/X7qdz+QgVELIevyoiHh+geV4
3lRtYenkZWS0VoghdX0pdwoGIFewBNE3Q2ph0Cp5zSCjci7XI/sWafj52Nt/7BcxtfCsN1qYb2RJ
+7VYboMK4kY3XZOPMVKWffuYtAQZjyWnLeRS2oHge1QOFOosU7YM5Wwwcux+lMhxGeVwmb088K7S
7i8WuWdtpQDodIrNaTAPeEpEHL4+v2iYqql2EoJ4eHVCGOvg3jfbQWKz1Iy4ziryzEYBn80QUqQn
HmsZ+1NkmoJL4MVxCXYv0jtU9I5gJ//E0rDMAygxWpye7U6h9LbFKxKmRE23Ky10ZvoRRqlgQA5s
zrjergLnHyePPlTV5vLpREl96kX4fcEsKq2CC37ElD1JzqK0L5UYXOlLtZ9KxMCRrO3r7+9VjD8d
TAh5Gx3vl0VVEoaC6reS/pU5AjmPB98y58eNAVHVBOfWvzmNDUVYHnRaKPWb11htKxc8nYoRgdKo
IjWpX7+lqL87WFKVbrV+Xqtd05333+CCal/C1rsoX5mctSr3hfVD+B+Ef69qtzlNLBWP9eqv19ee
tBdTQZ58oRzJwLwyYMV/lTdUuJd7nR3RCTTiQ9aHsTmjjuElMqoCUsUZntZwA7hnw0D+kNK3wsd1
H9t5DYYEh0LZgDJP7lJl7rPonqmwjzCFHi8ZXrmYgVLHj3w5OvsNopaFHW8pVVVAFgtvqpcumwJv
WQw9ITTy34QjFuYosk+43rvCcugnAIn9zQUjw4liq1/hgh2ZTifwd/gkF5Tm7mYo9jcwauMaCwAv
NoCBSKErwHHbai1wFg//WjT8K9fZz6vdjH85PhIRCC7A0OZKpscEJaKg/IlyTQOuN3Ol7eLv5YQ+
IDFwpmnaXgsErnatv6fFFS5MNHzMPBlNcjMFUu8hJjClNPfWJAhxNL477/76zkB2AGCBpestjFdp
0MQpY3LhXWSqejxQGENNGbuNkxc6Jqn2mXV6XPvnnvgQ/geXPfWfXF70nMpo2dt1g0U4rv4lpFvp
ZWnqpeOw894Xe8GmYz3OopaOjRPmOm14gnSwsFEVgDbYSGPcIyLGeXTKUFvarO4Sx4ypYOtkkyQR
dlQARgp4oPhm4RkgSpUbuPnegbso9UW5oP6nB0x9OP/1xWpgHIZr8K0Ihcr0JFF+JqZycaHvSimf
scpYkYxDMNCfMeZA3McD0Ij4xa1YX8lG3G/YBbrnlInY483Pv9aKNtjz0X+R/mgicEVyV+Kk9FVl
cjsCfBAzfik6Ha9kCN26XYgFXFbT22hPwUPqNfzdPfjoBhjnc88B/7Wegb7jlZAHNcz5YEeM+Ob8
1hx3g7LNpVZ2SC2GXNtEjkAvKsrlgEhHeryEOYbVl+S5INwt41ac4FMJbDdxuKkUISOCKdvXh1lu
8m97WmftBz8+qd7NZKlpp5cQejmIqlXfuKycgioIdOxSmlszHRdyVEDu5FRmISunGGrijCHjgPZB
fk64Pi8i0eH3NGQ88bRfL1N7artSMW0Wo5cFJBy/urpzy0FybM/ymgDGv4zMtxBcbYxDW/u80ZPY
63hJRBw7EZCe1vM5Uk6sucJB78EKJe+zVJWlFC3Evk+0WqGJxdI7Q6jS0yjP3EOalYjJ4Fh/4GSw
DVTvVJ1DTvP+pDO3+Jrx0JEcma0AruKJUHlYY4FHbFPTvcaxTwW5osgVJZdI5yNuF2ully3O9iCC
VvkUAoaNbNpeZ4mooQDhmIs1oa9abrdto2CS9+FAuvlSxRXFrjHfvqV5dpTXK7clTOMq9BEHgJWn
zQbWtQEKRGdOYRb0ohZEZP5wDAblF1IG6nsDYqpLsz1+JxXeuJFRPfQbisIZBk2v+4P0kB7x/0M3
wnWTKvNUSBeWZbQxlrdf5+4r728tC7c7nTv74YF1hQjKWL6yeBcA3MhW61ywwyLx+1f7dY+VyTDp
/6hlu3QP2yK2BxvkBV4IszeXHCky95CUV2qb1be+YngW43+HteouGhgNBmbd9BljOeQ0mDld4hkR
lXK/IqbvMeRbIKXnj55kEE0r0dbfG98x/i1C8ZoliyYVH8SI7WILcBnbQxbc7H0Okr70uNYVeT6S
BttGBsyHcG7UdtUV1Fygr9skNoybeNorH4Y0iCxojCizL4kV2LCvAEzJ8O3r7adGzmtj3P0iE90f
8b+zu+Yr0tkpRWoL7PG9yMSUnZQprmhQePX+87ixRXHdJKygis7fiMfGd33M5iosVwRw6enC4mbc
sl/HTxYqxSZmy1a5lnDtP5fBE8+/HtIA+kJ3DWf56firYTznMSurX3XedDLRloYn9c/NKX259Wa8
IMvcQO4q1f9sgO4/k9GCRhQ53v8Yxz7ruKU56pT3Xy5i4e+v0bGQ/JsVmITCSJ2+GxIVyKhYVReF
OzJPsul76rkOzk3wHx2YEXH3SfgPoBpPWEAw8hOoJOyeHy41Cpu+IMUiupBHDSr6ncanJoMM7ypd
Y/MwiwWCHIuUCumKq/f3jlvdMTf272nNaujyAmyl6Kr9tRrse0ioGHOntOqH7WJUhSJ+tAKynkqQ
3DwFHKSSdeQMAeliVCyPCZEhmUcGrhBrg+CZ1l/w7SG1yOqLAedUVb2ADtAqUgf5BCAB+9D+Kb2t
WiGdV/0K0nP+tUQfOfARiGkwC/LR68dhqA7pLCD/+6TPLSjlfpfoxOjSS+zOPTsoSdbz8AxLp92o
VzYcQTcI7NNrmffKbu2kCCs1tfF6S4RXhfjLActpFGYq1xgC3XBIJ1kxyK+M6cHWQw9xDl7t/1aK
M7Wsb48QnIhSM3bp+p0GWE5E/Qjlwy52FJ3WPwvCOQdE0GvbkPovnAWtOK+eUvbrfieCHcda82Ga
qSxk+7Y4guR4iWmaoEp/5V41rbkVIhQMHvXFmAKj1RouIgMNhmcqJFF7NTNXhhawACgJDbiQvOTF
oHBmzjJrdcKFq6TqApCRlzDWUe5mLdl1rio/jPUgwK7bRxbV0yy2oQYcVdoWiJuIDph9gG45J9BD
WnX9cGXOW5abchIPbiT6bV7aWuQoW1aXq6yF90uR6kY7riEwfDRJ3v8PXkxlikJuMXPabvUNirVB
BZvpO9vlZrtDhZyMRE073ygmcioTzbVbQHMRFjHznPHajlhgmQ2E5FfVKNpEZnpKMIfHtusYj6gR
+Z/C/9R3vLFv0kW2abjBiGuSWaSyxCHM1fL3FgrLXNrC6Ym6S5f81tK5P2XH/gnYCiYWINT0SOkb
44B82Lzcc2LX6FfRasB8VPQrQuqqNHWU3I47vjm7x5VyaGZ5GlPJrnN6T0mCrNdNKAM81olRRCCk
1JM9SJv0sXPEDrRJ2OFYo/XbN9WuoTQLn6PN908rtrkL9VGRb3mUjEaTK9FPXEgO9oBXArPjWl9P
xarJ+CwEb3ZYZoJs1LThghols+yJN1lbvtqBb4TwpJGco8P8Vj2K2Bmym27/UHZLG9kT3cmby+6g
HJ8wwjiuCDUH3sGhjlp4XWzomkzbIiIlKghfhZH8psgfwieY2Mp46+cj9RP3BHeib0MuRlXA8m1X
LDqyRPg8f7q9dUO+qmeIQSCC+Y6OLlabB/NJeb7lS36s5ZssPd4J8EFuiaq9y6Vd6i/4cNcbsWGn
fUYiy3CAaPSIM5uar8ylMKeSrqIPFFUDO7OTclSsoIDrd7f0qxCQAVVo+AZ8SXOSP+iegfX6QLAF
vUVtaX82tWlc/zZ64Vnx4uR2buLmkIorBhuRy/FWdkyKAJ0+nwxogO2myI3uMhhQ/Zm5TClADpUn
Ss8Chwz0QkZul08IqtoNHyNx4es8Er9Pl3k2pG+X+uG9pkv1bQZ0jbBPFqBpMXYVuP5+cZQofnQ0
kDQrbKHDsVLbd/bejCo5ORSZAKfjYSrjJCcWMR4mDEJeyB0KjyINKv/HOgdq4t63UQtwe9nnurGk
iGA3As29XtaiobWL3CVuzPhFQM/vWdAVwdkWyFgBsBtlUcApGm4Y4Y2tpDtX/bdc1Mp6b2lztE07
HfR0V9nBEDmU3qpuHtoF4Z7DD1HusI5Xt36c4Uh0w4PbYsv9ANJeh1OiCBKelA/rSBaoOWBnQ0aK
EgiJ61EPDyX6wOsxDj5k00pIesJcWa03h807/Nfy28SidvaQB7eJmvagijvBeS6ALeHoWxgPbQny
LoEN9gx4jxpR6cB5EwGK3nJPzbvVP+Y5TFofl1RSRRV8j3GLAbUFeFegnp1q1stMO4uNDDyZNOXI
oSS8NQwhkWJidStMcofHjx5vyl9RuO6lnW3RJdrAoYyRRDwEkwfvp2dp0/DYTjDuLPbly5c7Ky2a
Syq8T0QN7HxK5KuDpUCFxBm9uN+C5xUxf9f1R9l9m1KkRkx57sPbvtYq/PacSzebj/p9mSYIUTI1
d5MI8S6VdkEUOVVIhtzwAKjMm6ue+7u1UurorOkgKfo18gcl+pR8AonOIfxbpTAQ/qQC8JCjLk1b
2+OFCD7hEW4gbGdcLQd83f1lVNvolXosG++9AqE7Ru+ni12Y3rrPAxTmgfdM7m66rR3yFUtmrjBx
3d4SMFcuWwZaVg9enZza65/9UnmkwXcyVKPkHYCNruCeNGTuS8V1SmjJHThXHSieNcsfEkI3MxaP
K1N5FhNbup98qXXsmhVaqqyc0J+XlhMt5qLhbzYeFxWCvgoq+H501BCy0MTSkMqN/gHcSxcijgD3
Uf6+AJZ5mZfPCzjbPLzY/DMPZPgble4YrysmppJzj5HHAqSj+WlgUwZQ1N+7xp6RkUFs8AtvR09R
MPWLeeqIVMDbaQfntzFeyXjbTRHOJwGDmqrd9O3jR2xSMqVUcXX6dt8+xD5eZTURM/6iFPTpa+yP
49snjFJJ/yeyt4cmJ/pg/0KJUDok0DXzP8M10wjjS/cg9zV73d/5O04Rv26H3B3hVuBZypia2X0R
8sdgtzaPUM4RpRD3FJUZYpkU7HCzgqR7dIIskZswTucvIPWFrU5+fGcdL4dkjD/FbvXKk8Le9eGa
lfUVr5771G+CNYLh5xYiAocii+/T0wG6B/SufFftjPFWqMIZx7fBE1TZDxHyKy5tb7wenAWZOnQy
cwYA3HXBMR/k1Pew52kZIgwOpF8MoY3KjrRwexf49bSWWbk0F/eKBsN2L5AmfGuCwFDq+K8oqnPn
l1wM3Zl6cclxJ1a51X3Ncfrjl77IaTHyUrW9TAg3bFgyjHTGP/tsdWm+86JLXOrNF5LcdIKdDAL8
fXGAmCHh7iULRWsmZegs80rg2moNpOjckS681Ql4hv5KAVrjmPMyEH8MdD00IvVxdWowy/BGo874
FH0ju1nxLVUmqdRxztdvuU4uh/Wge+8jW/m61WpiylDwczbtYdBbV9WSx0S0w+pUGAfmAko/r62A
PqtCMBL5h0XO+fUoPsbNKnil28VqhXrtlzz1H6QeNXocznx6vXNi/XD+HZKJfUfddYY+kjE0A+Nu
cQBjyIsbdnZPJZiG4hAeynaqU7zg7Bpm5LeVU50KSAkO0mu5pY5q+ReDHEA/tLSfkOmQgz6QZZhM
zyQbxlZzeNVDmw3QN3NUBTahnd+ikg/MelEamucuY8opWeC1X+pffyVPfs+5ZfTJw9z5eVzWSpK3
FRwmJ6GpDAhMZVEW2MiBfQRdnrwHFtg/Y22wQ6Oo6wjGWwL4H0KP8yFFLdajD8Tlt9uhSlxRkhxR
iow928eNx8pBUmvpBQq/5v0J3RAYSBQugZJxB8eskn0iDapQGTln5NuYgByTgcf8zOEtw344joXB
e07VEnlfeZ7XT8RwjkL9h7cVR6PJgGy2BS0nQwUpMBBfA6oHIgEY2re8RVStqcfhPiefDJv0wcF0
04GW+8dQcaGsrt/xw26y5fI4rVzERr3qXx4f2UcngldN5XH0jrOuB6iFSWmMrUzs07Rk7h6ZBxUz
3t/RYv2aHZOgQ9/joEWsOLS6i8Dyj+YGmM5AcMjBmnfFFbtnbOZ9ywXFhCQlj+UhAkcGGF1BX97b
YLAP49cbWcPSKhgt/wUeKuPLV3PEiA+yyWPLbgwiW90D9iTwBBJ0A4z50EQm1kHUg/XEvFoBQjol
Q+TwCVvhTmNncsNG3eLu07oVrK/git2/TasAEk+qLeF+DkzXq/6oj1OegBMzoditPHVQeVwzVKZJ
gRG8OcytHVUS1yc8U/VnbTOi1A0u9ZMh3PICmqn/95NMEVkMT+v1z8yZAzEm9QrviZqPQk9yD29k
bBDQMYnh52TFZU9+uKLaglxv1zC1AbradXPrR10RtLH6RKb6ZykiDKtl/xB5syxG4VQ91lzFF4Ki
k0CCG4A/DGPOQr6zFhvmIzRkb13ulDcR8PlHhunKj5NCXdEDt5HC5uwprdrwSMSPXuMjbF2ld3uz
RGcqrGlOeRbWhR1QaXd+uuc6VXg1y/Y1ZpxWjYiSQ3xR4aC5/EA6Q93+pwa7tDz8C1h6/RZzdDQq
wKgwJRWlxy6B7S+5eOAVBDv8jQ+JVK17gLsfAUkULuWZJgpi/k26+42twrJk5F0RBPR0qgEPPT3n
Kz/Z2YkywgSSJDs/zWpckCDgWjPs8hwBqzT+6It2T1ft7vJzpkOjAkK65+Fzt2YcKmMYUZ9NW58T
9H1X1zwyb5GZMnwbPvO1qJg+Z01h3vkR/ogcd+NJqDamygcSb9S/nW6sMwXvD7rO6dhLL1/YyDO+
/NfQaBeRVofT8KHg3menIeDxeI4Hoxy2UtjKGSlCOu6si+7EZVyIrfuKNilLx1RpBDHIxiiOSorB
Baaw5vM7Cbv0/XvCa/u7LAEguewAryC2yt141pYcWFdyvzMwc0VIoDGtR3z5K79OdgNTj0uwBOUJ
Ev40qGDyCAM9WbKsJQ+mvjfT41kJ9u1xE4Q2Pxgb9lcx5W/MQ/KnrqahPAsflYnk5ziucU71OuHQ
scHHc0xrBpHnmeh95YfYDpLxJwJ+JpdKGsicrL6zYe6bcfQQwn0y8v6QKssokDoIaZTQqs0qYFwe
1TCk77+Izb1rkonnLh/QiddHY7LOCnfNjy44GYkHjgm7kRA9R0cONlqBpUckUiilzHozTxZRCKqs
+4HZSkK82RsuybvC3Wt9cltmtZmgykZPrJ/VSFbAPMV+S7B6rAy9nUJwz5/RYP4XYzKrvqO3JWou
Qck9bLwaLRA9ThnTDDvQmBQ3iH1CYvpjl17UR2ppjgy0KJVXHVLQd0/+AIh21ARH0i03+HtsfZYh
Co9TgCZwE9JkEfj2XGKgZPz5FbFpaZfOL3Ge0B1xNjZiSNeGBjc1mspuBF5WAwWxRjxPUX1rab/I
r7IUxz3FmfECIUcb2e3lqUwHv50TDrmKU8aZZdXWCdkOlVimVhaRJyEDem5dEmHEj4SBltw1xc5K
4PeEsB3LJFPUAV0H0YcGYZt6fji/VHTfrWF1fQXRDIXLIvuJrLuamN51Gx0GYV2smYS6WSSn5/5d
wmaHUDiJgQ0C53qqxEEac68mBUffgYNu38mEcjQN4jk++JMga6rxxWlIFX4UGonj9Vnl2m1XSzzZ
/TmaQUgxNV6ntyUNNaCOC7BzwBnppE6lZ4yA3EO+oDG5fo2odFnEzA1tYKotUd0nOR2/2KZBbiU6
1bjUel5fcrsJqu9SXCMejq+LIoKq6mGCRKkajsld5Is6L8hY1FgUgv4dW6x/cu4gBzx07oW9TRJ5
KJ9RyVBEyCGsPyIygOQ1g113vkU67nwZcKgGUSb7eprPTYkXrR7Cizogwg3kEMxS3mo/dSiZUe+6
p0N2oLvDaEVWOeU56ZEfjfQrwxAmac95J+CjCIQHPRmV3WSMlNaqkDViRYDnusOv1o7vr2NHQKpp
zsdPYBTHG/HloaQg2qiPzq1iVfQu5SAQCWtEtAN4tkJPhJr1hafGm1YzkYhybdurNiiU/jIb8++j
3NZKcGWubeRMSd1QMb2MjLV3d1pGB7Rs6EC4513AvLop7UE6p63YRDIgAsI/Ql7bw/+mVSjCae5z
F629K4nV8ziNutLUYlAW1Rd+w7pLfPg5FzI17uxqLggppUVOGNkqTBzSNeNNL1aaATEgOT7TkKtg
w15GLENEmPLjwJouE8P2B0u01CkcMT7UANjfwlSaFDIlQy/ZEi3Urx+zC7cSl35hUYI+NRyOZG9Y
bFlPKyoEKqyTshUljFByz5ed/zhr858TpKxm+pxgsO+mt724bZYWKnILAloVQh8l+AVaEOYoCACC
m5JHZYFq+AYkRokdznzh/ljLKUdWmlobe5vylrmMyKkC8bpFY/LtaeuTFM1KdIneFdj+RBmbjvUT
3Sznb/lYUU5gtRW4qcd2T5yQF8AESHtvP9mya9E/At5dYmmV7U4Lw2GAk1l7vNK3+tV55YHeAQEW
vCrA53QuZqtpLqPatk2i764ccRRcXka5/+aILMbXQeES7mdoKVtEUGGKbAIpdZcYZzAMadXcsyDT
tFdxMF1/kmQvV4QiRwhKFd5ZhzdvTuTvM9Q99sYfHj3S9tKVAXLFULbVtZyXoYBfrR6wgRrwn8sw
YIgOC81UbY2uzFykfwNIbeEsYArS7F1xF2BRhbdui4m/PBHede0ljd+Eemy7eDhMdqm2owKMKhD2
cGv6LPTvQb3ogT7LPGTYSvb+LuntPftnXAKeXCV4kXVZwhi+vFnYEWHs54iwZ9DWAcOcezS9MlKn
qHnCHhSchTt/6VKSjoU+RrlF4v2uxCx0iDnGPQUwN9OCcLaU6sUjJeP/ytPZu8/T67Y2zNiiliae
LC9vFnuo6DC5qjLvpXhcqTrwTVjEmcJZ6odj1hXF/wCM8jovY5HttysbeuAijRnNTdl/A1fiO5/o
ApWTOZqTEx/gJ3+h+edbx+52Hirqrp1QHRL218nb4Bu2Oo56Pg6LyPzaHfrNMaMnjIwwF9liNVQf
+NXrgvuQh4ivzxsik7+ewHziUjCD2cGFIPFXmZqwHZgj6QiQ2vdj9rYUy8L2hWmH0rbc3a2JmmR3
YXrDRolyvohAOlifEwZUee1tmSFUG2t7ccb8ZtnZIIAp7JCa5/QrCkDOHIPsB594E0CjzAJ0TKFG
ZmX/qUMa+2d+enuJ8qIT4pNao3oHhcBco7Fphe17yPSD8JQRwGnVAWgu5VX8Cag9juDud2OfrU7U
nDJmHTzyRza4yEQIniHm2UgJSp5wp/5Hcm8mTFQc7VKPjGBMY1zpzPffFu8MlNLp2+xpSLq/J6LO
frZrf7Ddy/2RlAxX2qxn4Ayuw1uqIuRUe+TNR1v4T+nu908A05Yj/VYm1HDnlb6yGUzSVUgNxuCV
ZVv7y3DjvCe/Sl1/bDPiCVc4SvTXr/zzWAUMyKcNyw3PXkCpLOiv++rOF3BMzVFSXD6QQcjhfJEp
kRma3eHNusw3eW6A2rnHNmJvXBYAqcfykIwO72JSx5Igt364cy3UbENoeYxNeb53lr3t9c2/OfdM
079yiluSSOTEGRknOsedngBbWYFghmK3mzJO4Oqgx3CyJ5ITmugwh4m3fDYdivgfmRKySU7W1y0s
KOlKx3uAoYgJJ3GrZkne1zIErv0MfJMx09aueJRB7cU2og7Zd9dWtP0MIjKnGm7TnQ26xTDlw0E8
+KaQfqLD6m0Yjk7SbzuHBKg+RahGNg/8ZZxtctg0+pcjosAF3hn3RFry7d5paftQkK4gR9YU9M54
U3HB+X6rW+XEpCCUKoARaLBuFFr5t3QDFr3HfWbgl+BSSiibaLUIWYYkvvsN5jHLyumOvnNRdVUP
08oaTXqr3WQVIDp6NKoq5Jq4U1N7L+n7RG+VAqA/zMIz38/Udjr/2G9WfNA6DwwJIsDdc2M6KKRP
ZldNV/sPkYrAypOkDqoQ9lT2k8l9qVdejevvksGUtAIp64NGJfpBAmSzXumaElRDsof5zzdDZPur
9egOhnXvIkq+kNchnWkKnzmN6VLqbKm2NSKMUdBefbfidPSX86647um0OYs/xyAli+mO0bQP8i6l
7gXCV0T6wYekRMAzoyiMhh696zGnlhhVSsh1PyQje+JmCk42Hjn9aNor7HqLhUqOlwGfvcSwaifJ
WibYmSske43Cd984+l4L5E+YCQR2af2Wbt2t+eefA85K3LeIX6228FMQAheSHzfac+HH4kn5utK3
UVFXfFUIXkZZGHZevGkiRKdw2nwJVnqL+zpHlcNxETWQ41gGgGEfKAhjDU2onuJHmFzZ7tACRmbk
ctyqriG/3YWMIgnFftg1OKzXxt/6z6xgtZEWWC7xKZbEK5rsNuLAdrBslIyPmO1Ze9kX0875nRJ7
Fpji9vYiW6hfQ2C+TaAFVCLqZEWhG/uKePs61KeWnHODi3DS+CzGvUOmy9t0Qx15bPkSyd5RxBcu
4yMQaooRz7wPZ6GYurAe6usaIdqABv4uTpy4dnkwrYDf6fyyF6hWqsD/lo5VLjHOnV5iBszr6LnT
slPG0i0b2rTU+P5Rnt1xlrYf3uBQ+vQJYWrGn9q/vIywLv3oR8Yom52u4rVXcQ/XgVMyA8v2DvLJ
AFjQszZQiXeR1Lf+M7551jDyqonxCObIc6QuSXkYu8ZyCawet9X5qet56+LjLSA8uL0rQxupcGvn
WAAwwudv9TYszhw9D6oKmI4TaTsTp8mlKE24QFB4Nut+ENPpwtyrDUoXJIx3jRfaMGn88QryhlfU
aXstfQNCua6G/wqCn9xh/4BaqcJhk0pn4jyDrMntTRfLQmitDSSBcRiftADQMpNvz1omNlO2UcSR
zaaCKbzzcm+WIyMBUb63EN/aMnpDn6z+lPddkCOU9/luDZuwUlW3QlDV1mL9zhhC9xZ5LwoIBHgw
JmVgHKPPIfo5Q8lzo6/rKICE6p7xSDZXcvwszu3LNknKUBC+sr+hYAKFpdtXI77buDKI56ZsVb63
Qq0xdZzKZh2LUS5cxnrFZUpVr8se1pXkhh9hTC9wz0Y2z2w574hv8jbfzyEjtq1+ag9hj1IH2VaA
g43Th7ybm9FLFcD/g51+utB0kU2c7OH63aCKA1QpQjoYo0bacijK1KVbVkcG86VaH4QXE0t8gtAy
Pxu3F0wT7tGpJemUwG1WiwUcMWPs+upjimXjwtr2tjUSI3lzk/xmz/hdi4e2hYHCHlODoKtL0KWX
3gDJK7Y1M4v0Fxlx3XaAlJdLsiuw5J72JLqm+sAiZH+7PChgwMNurwpr+HZWrl9/cmU8l1ELzi4T
K5Yz9/0iePedB+dq4LXa4cepPqMlYeABqYwaxR7CkcsFeAGcdBns0VoWovN5beyiKUUO5wQ+eriX
QL10tGbmIAQi6wXNIkCoGIIuIJQ+zPBLs3E58flSoo9ngktOQ30u51Q8NYIwbptWI6ey+4uPi6+J
ItDG2cpDTY4/8x9yr0gcNT16uaLKnwbvOQ8lKhHSI0iuYA3N5qet52TQan+DcjwFLFraYSuXf40o
mljRvYxjycAtC8lhcYGZsaQ54whNKnrsRq8RNyecC4FE0gIzCZdX1Ecmos8mlETh3fxxBE4JsE/y
vVpMI5zlMgBHhyyVWuy538lbouYBQcvqRBvYkN02lsapgbrVO4lIebcwr/GqU27+gfWepvZPDRx2
xJxyDjcejMd/c4rTsCe9Z+W7kgvQXHSln8xgKwdtBBAS1wT+3WIbYgC5QU5TPD4j3NpIO/QH75bt
ep+YVHa+sGSyEMb9/7+eJQq3EwYsd60nl40UtjdhoSplIq0YF/0oLYYcGKVc68i2wdkwdFIvYZQ4
kzh5sHOaC2RKv46DjhIZFivbGsWwxpLYzqquC4jOpFemYi55VvPltCpk8jaBm0mL0Q6gtuT1l09p
1+eJoB7wWArTdLPZG31VjCyvScsiRaRWpubqAe1gparoB16wLseDgcJdwTASpQqlP/foYI6J5pst
h8/7GXkRfybTwr0LQcrkMUmQJ2SBK8KA83bYLw5CU2AgEeLFZ0AcgCVdK5rywUk3tzZG7HPKaMFG
T9i/YkPVnmMmoZXhAn29QP4uHy8TrkUcJ+62xUZlRjm4mk5qsl5wiHrDprtlI+XYDUEYDJPuL4wL
rBhPOqHyBVT5ithz1d/kAjQabB+PwRb36tEu+LDpJ2DPFrW2g5o0PoAubfNt3GXusUXISyjROt6E
noSomm4yVA0FTucyfqpJc4tIY/1cT5tCHmVTUsXqu/ux0OdiGfRBCBOu0iWkNdCZDvh4FK8j5u4I
BbL+/br1tfg3E9oR8RhHBipvPWEUaOD2G71NMJ3s+Zbe0XG9FcZ3QCs22+twRGIeQW+3pAqFNwuP
YYjOCYolWEd8I6mOttKD/AluO++aQqwR3bRL3+9zRl7d3Y4o1mytmlfkd230VpRdhhe7gzLf8nEP
Avy3Eqa5WF0DxxNpRQUNzYbRL9ycctLhpsUkblauHpXtAYnwxzwvfqvlOhLHVAOEGZeUUZ8U+rEo
72tAic6pohK1bOeuojl3Hh1QELjOn+gjvwYKPAeAgT1ymBaSIquy2NdSI4ESVfVXioeJwa/hxxl8
GCdLdhlrQ0gDA8cNeLY6wftAHj4qH5eDuxNNMqsOrLxzq6FEnYT4cAaCk7ohnv4YWY0zuYpGSDR7
HnjAZ5UyumeoTavEy7T8VHQCrwzm4eJcXrpye0ZaAj63k2TRbAbWBc1MMv4+FNi0rdnGbArBMgpa
DMfcLO3e3kTDXRdYBS9KzPmLqcYkWUk3O0uc4mu3C1WOHwPfH8GXwhOR5tw7OnmAoqjo+eX/Ud8m
+YNHnv5ANiWPFMwoyvYN1BessZv1J4MwCt8Kx+a/W6g/6iQnt54jZzxrgq0gvczHaVyxrCFIZDn1
r3W7RsBozKGZua1diUvLnHhsaDghg4uzbak+6lGU+Pt6776ZiOnrGPCTTRYNNWLfZZRq1BzwBX1L
E+WhkcaOBUUtxYkNGEwemvgxuNnb4zlagekhNc4k+kQUywcFAS/tiiQ/p4un8Ziuwn6mLX2iK5Je
BnPQk4naw9nT1GULMxj4PZsr5TkbDrRmte/s1gczc0A2QdXuXdwPONU9xA6r7u6osTyAVVsL1xqv
bDzfuj0oYco4X2AUIvCMLfA81CWibo1oFS1ugPizMYiIaPt8RdFYO5XGosxaI885FrznDaYi6Ajn
ITAoYRr9JjEYBBPqu0CnQS2kl9DA84f4r21fLfDmDGhlkFzUXuiGf2dMIC2r4/7X9nTeAWRnA1ye
xO+5AADkK52kZ/aAEFsgANdj5/5QpARovRRmFB789jJs1F6kI6bG45SXgUQyrufNLhD0xiEEc9rx
5UptatK/ULUybtuNaeve+Y8LIfS1QaAViHj0xO2Mh+at7LMREsd2HRWRl5Pqo4bKc5ohWHZCItyL
66sEhNRchzR447Ak/zNoiTNZY7LmGLZG6yKolYYsOFkHBsHrv+W/JdyewuaQFDZ5FEDAxPHWouvn
3Lg03tHlmlza4VGfUMexdcoYtKPLaxavRQlxvMI6SdWHU8M13bhjG2JwstC9D4THLjABputSCNGC
mVIGZeFrKNet3uff28WAMJjPxE9k28ZaN+k1eYSVHyTAaG4KrxqXrdwHYxu3HFam2qQnLvewfNnL
7JlER2CjUoEoOEwDJLGac1qFXG+HHJxOR3945f1VVd3OGwS/vZol5c7ZXwpbV5IUDaWrmMvG8qW1
FCDPIVc7kLGw9DSTgReIQZ1okBIuUH4pPPfsUiR5DkCyGOA/SbDgpU7k9DZe3K++0/JjdeJU6HsK
huAw2nXwky20IZzIfsl9PhfKIjW49RClKYuL4yKlonREY89vkrYTq116ET0aC723B0o2z33MCcS5
WGhaKSOKD911crmMM6ZTOw2qgqYtp0M3cJi2uptmudnCnfqLLsVTIQYvijSJ4BX6OwksQkOX6AkH
arU613AW9YiQ8/iVzEgb402SYpi3lpqfwVqHxZHV0gtAY5oWxMFSEEn3ySVvnxNUYNFYKNAyEkBM
rBqNw19VRl/5KjUCW0J+sl4apTvSx5EK8l0jxKzqVWmMiJCAq3JGALmaInuiaqllA7+QBm9W+mDz
f0a0tEO1Nghlkr7qY54JNycJqw0Z8Hua+w6pxrYFb1PDe+n3veYP6435X7H5IHW8RUU6g9cEtVW2
mQiYiVJ60SCzs04qq4sNh2KXvVY4ypzhBYykpjKLB65Gi2Y0E1G3HTSf98ZN510dmqosA1iCJ2XK
Vj5jTvrAFQfetf9z1QWVukNAPdtWeMJFy26y7LmqvZC3Zf1NL2MoUWZuCjIY9Lulpc+tYC4gLQ27
PX1g8W30fV2ivxvwdbgl2kcisRcdeNSDeCqsb4Ud+jrZNF/1/dZ/B6hfq96jd7BQzuHtR/gmJhL7
hA1ZkfD92UqWCkCEAKFMvKb0tOF6AH1ZB8ASnqIiL7MWLJye+ZwcK9hrcKHUsMCCk/fTRCPPHrQA
xIx+U3I+Ss2GHBAy+SqBRnkNp55RYhvoz5OTXy+jMjHGIlWtnjoIw/onE5Um0rGn1ReT1FMyRXnX
sZ5vFZxajUlXI+vSBzT6Ta5MXcJWuTy1sWUb16fvoi/GpmcFY7SZVpjms4Wkb4vqt8iMkJpyt+2X
ZGBqgbZNLE3kBpb3jHB/19V6OChyE2P0Ftx06azzfQ2IZLbALRKO9V2VFfV9rFP3L0XT0QDoF0ZR
EcJR6Nviq4mOdPu8akMPlwXadQc+leBQ4DS6bPZZry7KsoZMkqWMUIdZl3PZcXxyNLH4FH2wlGMR
2YUodwZks+gSf7UG6jw8AEGG1OonlvVZ2IPowCYV0iF7MAZF8umskFL+2KeT7T0EFRe9XmDsaFch
pJRNxCrhPH+FkNZhAtABOedLGmj8xzvwgKv2E08UVn0ixX8HtQ5YV9ArfXbP9PkmcpKwbj22fM7H
G2YQAfJRQyV0C4VOe2JUuZEs4rGqual0FVETVpADBaUoJ8rDtg+XGgmq+e35Qxmm3pckliLR+b3J
opRg3oYk+Z9HJUBOzckgou4a4eVsD5Q6OBnzvKMfssq72RL+S3LZxxHSF2tar0XJbAVmkkOsSiMg
a8+WrQScMaQfsdYuqb5/2cluaGDLqys321RPCqvRr5Y8QzmbcFu8hcObH2MJdfguvbWa0cgfQ4lH
CLIectB5pjQOfaMREO2XC+bILKxx+z8eepYJwTNn9ahnHC3btF0taRBzI++m3KlT9btA0xutBQGG
4Iky9YN0z6i52FWu/DmYgSKtJpQLSc9Wi/02z3JoT0ZCUIzUm6bWTLrkiYmWg7YPFgmLHk5DdaOs
fhk81Yf/25Wkhd43uvLtp5tJnbNoz9TcxCKIY8lDYMKBCQZgJppI6FyS0FV41dVuS1OnbUdNP+s3
X9dg61GLYRyp3yUqFKWjesgF3gkibH7Irvlxz76V0tKapjd1QhNRD3SjajiKSCGbgskHxwsp/sj2
HFyO5SLnAEwSpGGj+hhJlzTS7jXv5o8wCMAfMHnGmeH7/CCjRRNxMO0z1tC3nNvO/U4GOHRrvDrv
FKaSnPB/GH6LcEiZEHYclFiziakR8bsd0DZeNUpL3b2xwvLFnldgzFeXd1GZXQLwrZ775qH1pjb/
WgEsqZHI05gCFEBlw/7rAnJ3pHlLv0EyAyNHPGCqdvytw5i8++8bL0E7MR2iEbw2PczJIibju7dC
MYIZyVeCC45VIXs8/Eth2U7Y8HeRiiSMjWW2RgYLwMOquPZSrz3/4rpOAVZH8UiRe0o4Oa/em+Go
7RdrWBU/BWu74VnQeCmYSvAlH8PhhbDnOLtkjcjUo3v9bXhfpHlO9a6eV38zDygsFQXz0hVG6fnL
lKPaBzTeoNXJvN7hiSxnqU8KMMLiYMKysxmEuVi0Q+0vK80+t2tgVQDCLnutKVoG3BOlsbdvEBig
NkVTqZovjyoh07x1boln3DXQSihtNGBmSV/FrIOaLc7vqXmxt03S89pFwa2xrrEBkryZBhURcw21
Fa5ehf0xsmGerQ72GpncuQgjdvMZPX9Qp/0f9up2Z7LRyNfQpcsBvk3FHaJhnZgO0NPQw9rfQggf
dTLoTIBGUsAYoN5ZJgdlDrylLM6p5mltf0AeSjOLypk5bN2r3C/g0YcR/VkDkMP65H8Nr6adHIxi
i6bsPsQz6MXEEl7Y22liKyX2WOdbkOr3e78apWsoRlXJY8jvexs1ax5AHzPcSGv8GP6TM9OyPqnv
dNlNwH7zHyURKusapsL+BrPI7VKzd4Fud3p7WZtWkTdOgEgBv51WX+fa46XSX6MOlW1tuoZAmIRv
fQFqQGH0fSPBrzyrXrcfL1R82OWwOXHfnNW4swU/VhEAxKwWeSIEL2M5IpCpRMOOdkHbcTqWMFBn
1fTo0RoR09yIy4xcJb12tr5bhTbLO7o3bkhL6TTmuszQyiHSZVCl1EfmbZNtzF7cS17V8jeLNaX+
3/Y+eIZZSTHFGFU/kWb/6qmnliOG/B818Y+95xPt1bRf9OnG/QJYxf8MIQ8Bx9E+Gj5zsZfJwx4c
FAopE8AGjZoQWSfS7mAgf0ClBzldIfUUjfzpAvszInFqxcknPNQ7C84ZozLObT2QTuUCVtCqvjo/
OXm4lAMKuL/CvqWrqwwbWbkMB9M4z3CqaF5pyfn2WZxy2qA15qZtL9ABuLDNrbzxRP5ZVjGajBSb
IFWCFbRds+oRCChSp6TMWatqzyap52IfDZPFDXTnQ5VjOd9AIw+JSvfGpIp+cLaAYePg8/pMFoJH
2MVwEjy0Wq4y3unUqQN8tYPqWIjZoY4ip49CpVrokJObfItmzFcIeF09SSazhIV7J5myJr94WbZJ
2+Yny/Lb3rMvQULXglWjl+AJ6qiZAeQR2nfYJnsghn58TjgklX8MZ0V0CN26/5hw/BX7n3KCH9Gq
buEC0kw3R2FESNbIm4/Ru+PEEa4E7W3NUXdD9H3PGnypjuUlK56fLo0ieThdpue0TvYAQp/g4kjO
VJ2Kb+t/FEBEEOS+j/yLdA6D20cjQbXLRLLBr6FhSLHHWF/IiIYAkGdsRV2SCn+BjTsqmpGA5Tt4
qX0M2gTtyAhL3LGV+pjHNTnOrrcP7nvcNPn4/HBvVxP7QPpRQe7ehDzK9eVINdNzfAau7B1trxFd
8wLl3n/L73AIyoExKFHd8gqzN8Km1zpQZWShRzMzkSEI5jDAmhFhBtk8p8Ge+iLYIWq1xOvh74wy
rtWKQBLDydTFRSoZ/5S8D3pLq1kQNpAJCiv6gL3dYydpn/eDvPw9o14tiTPQ2qI2PgxZ0B8mK4Mo
PK0hSLyKcMeCU0pT9lb9xn6Ad+dWmM5C6B+m/u3y/8/L0vaT91bwNx4OHYZ3cxaoEvNfXhGAb5gB
VGYgUwgRCRJCNZUjfThNwmL3G8ksrHRLzy4kZSYZAQLxR9O0LwPsZDNdFzY/iIQtxnRpzEa6iNaO
s9fuiKdez6K4RJJWSIyKZn3kItZlKMMGhsW9DtVBBFHP/kWjYAKLhyFXPUORZIaoY9RgGoZ5feOb
BG7acQAONYYMIVgxQoDosr425OnMx+i08geNH200RFtIOFLS1rjw5jIMfvAsXlMaO8u94vpHrSF7
eNqZbCfXmD1alelHwVqoaNbcbxkg4wV4DQOEQD8emWxcEWyfBbRlN8wX6l1EcxNkYfy9GVNVmEo3
w9qgK/vpeR2TuYVq0xc4WBcv/XykNno5ClJnGIMUn0xEvVXkUwQv6dGo7NhYpKIP4Badwf7/+y8T
2lAVmps5t7M/dIaX1Go5VRzPt5ttcVBQYT+eZIIAdcQEQfwU6aFM/pDFkhgW+UomKlFnAXhSMKv+
2Am14u9m2BpVXRT0TwIGBCVjQus2BZp3y1pP8uuBd+604wWIQGm+u7dMHqfUt8ij5D2/fp5ZWHqZ
7KcTZEKJUja8Mgvy/tK0AF1EdF7jv+WEFBCEBy8nm6dpUARfjvKWmvNkHb/ZR4d0idypGVtYHQK5
aNKVJe+WyauY/5YzW7jWAFwlPb8zz9PbMlRJ5ihAoGjCMQjIwncwiBDeMg2pIeqwJnPrLaERUaXV
W+Ptif4Bs89YPnhsc/dQwV/bHklSiVqbPxVpo1RQ8DxUheVAG6s9eDz6Nwyy0d+aNMIe6OUCe7ug
VpWwmHPBoBSod7x/j+qDK8Ar5CcGhuPVYO3JDz3YT4kXXlfpPfnml950Mz+0HCsZG+eRQViqe7Fx
6tILEJHRFq90DDwHLpbPptuMo1OLd38sxdFunxXryMS8y6MqdPQCmO3sk//euNz//cBsa11TnBpB
8eIUrPgyvnq2hOEpdKritZmW1tdidFMUeh9Jw4PI++5Xf/aXMx9eLK53Rrz4Wcugbojx6AfE94d4
MFnjPB7ZakszcUtSUhU39/g81QM7Y0PsL5GsJhO6f+TKN+e+15emutXLwJJGypbkhoxNUo37aiWb
WO0rCv3C5tUSLiAaGYq8wg+rXxxuiheLeW/XZ63Aay2HYBcN5xRlbrXRAuKCgBwz3kyR9/HWCIlO
XaHxkoM3pYIDlGM7SVB7yYBq3Y5RoCFwJcZpxuRJ7uTnTPIX0FfDc/AZZ6986oRatYBauRoWBQ3T
JgpeDno2r39VDwEs70EPN1PDmG9XzXbdx4mAlOup6YXCupInxhHvGvAAl5oLCsfkbfnpGyWpnssG
lboLgbSDBjtNNG9gsgxwhBBMEe5KjpBaXJj8FViHbcNVCu18CGf5CNZXO1m2pwmfbCZREE3HVX/U
7h4dHUp1mBkAxAvoRbfLnl+AYlcLDf3nW9UbX8fWNH7LCflrO5PaUqjocsyE/hO1SvgLQm70WIfE
LqNaGG7TY4vmqW9Y3Yvx/sdHIxgNtQ+0uX56HvV+4rkx4MAk44g5dOqrmvkYQO5Ab9l18xj0V/VL
AtS3XEA3xfnd9RAdF0ffk9EAAbiIEk3riUFtiik6EAqxpD9lWGgSkLkKyXebgPkOrxOTMDIo3OLZ
YMb1x0PorHnsxQqysUBKY8nrelYFSiodPVp91BDxOiSKtb5dTFoTwZzbmS3mKYQnIpTpPG6CAsE0
1imZBlq8Nu106PBuyJ3vb4f6anFJ4WX1+qWRV3d6L/0cZJHgEm4CfOcqm9EeIgcsMtsFiAW1zHdU
OO2JDLlZcz8fqhEUPgFzRdqDQrVueaX6gLHFUR0SBL+K/Jgu7EhYXzrsdXVUEz7ZwQopLRjOeIwU
GQr9y8tCr0sqEgc+CTCqIng++zgvhnxQiJuORD5itcsI+nKLyIULcyF8BLY1XWUXZHTwW1RiyIsy
VKw1p3tiiM5ydC4+NL/HhxGaQG/3IZ45rrqCXZobjXTdbx3sUkT3vLwcLGCsM6Z0KrVL+9Jjst3U
CzdDz8MwfOvtQYAoNvyZRzxKXneRzkhhohtStbqbHeE/K5cliwsmB49tCddnZ7FM8fVTNiUYn4RH
I1X4J+zAo1xSvwEaR1A/xzqccj8ktD0Hie+TYGLbn/tDJLz1JiY08jsJ5d+p7mx7qSTd9V2RCOo2
cUojo1AKewaeWs7G5oxKogpmnobd+MCr/wrFJ/paVPn2L71R15mEuYDY9mHmaEaokstlNl6h6tgG
TqgrQ/Eu1cnfcEj4EOpCEBp0UR2ctUxSrBoV2tL7H9SRtWmvNqTmNC1luIPc9HIO8+4Zu2VF+mSy
zjhcn45UiDDkjTiB2iKY9QOo5ZUrL6ciTusdVKg/ldeP73CzxrBX9QItXU0fbpYy/pfZTS3F50k5
J8aZjTZLG+O2xW6JL2FIlITMJYTB/Iw4er9R2BJS5MSfFY9RbsjzURM64xL3yP4cAVCU9mDmZOzr
JmYGKm08c2MEsIlKh6hb7MRZ40vOf/FFiKiUDQ/XovVbJkrTu4zIcmN0aJxlA0P66Y6YQyBfUMmF
VKqEgn7yX1UqUsMxGt3U2yLUSUJI6mAjc97sKAWGMA5Myozy99NpbLW6Py9rzgrk9o0m637aKuhp
oGBNcYXCPHclFn3K27up4/HwJiya/1jSYzT0gj5ImquxyeIo7OhudJgsi6JIu5AfvcJQYZV+a8hj
Mp5Dp95Ne6Y+nLYj8lK8ysAzL+hwYQy0e2m/UFySQqOHr3/unl6XxpdxU4wxz4EE3CHRy8jCsTu+
06BbjC2NOdGeU0ryF2pMnOiF/GOjdRaAS8styL3ox90jPwIvKa0KOl4G485JKZgtBuQLZi10lTuk
Xsxm9viKJix5G4zAkloTyF3pLhC6NlXguZKVgFw8W44WZRchPXK0+H6ToLmmD5icibRyiBwle2hg
V3sL+UpMYbe9NKe7Kv0VBebrypn5ymCSsVnWULlMDmm/++K/nJylcaNqm8n7xkl0dU5DzXhb5oen
XpD47zeqQsomfjuIIY97mXr5nQ5dvr0i/Zju3HqvIY24au0k+z65+xz6Pckx4w+gdTNC7RjXyh3P
OBw+WCvgtDn3v8b+S1AM0glaZPaKZECp/h1bcYg7ckSbG2MVm8Kvmngn/UmTwmI5UU8sV4qpzE5b
QkXpy/4mf8XbaVXYgJyrec5e7q9oJhWon3fyhrvZJnJU9qFqxXLpeWJ0SpsbkKl+Efppo3CJ9W/O
ePfpyi8j4tp6Kk74kT7xEeiM5MpdiTKFl2X1NnTMpdE01QepPSR4TiPFWve5NOWRNwLPi3MJzvzy
T9TqlBA0F1S0qPvDxbfo2xypKTkKvgtYuI2YctY6GeuraJpqGkPnA9e5J9d+B4eqEi5Iy94zYm5P
yUHMys6oCvPag+vyluy9vwgQJ2Btlax73z1XUPyMwfQDNS/vW5b6STYJRfAZeSbdd76fevlQKjts
qQf7t+1Wp5zY3n0UPVQtxBKfwQhI/YBq+mgSeQIB41EXsHEGOic++NTg19ZIWA6jWrFWgsqgcP/8
OEH2i3wcSSI5TflodYVm5okEZonFMSulAimSzZC+Wh9/LfQ5K3nBqtnbEOKZuClR6ZC7WNpSkDuq
llwts3npqMV56KyjfTMPs4Fktz2/r5CVzlJAKAEhFLUxSmXpx7BsGLidq//bWk0Ak8iu/rKMO3si
O2q1bcQoF9bT/CPGidaaDlDxLo+JDvKRPUL3qwxzZf5s1C3UUcilX3KQdfM481k7qadUvjb7WiWG
BPvLWCYslpdKeaJwCZm2wOJoW64FwaKto5YJz9StLY0cfC1mFwwRceCuqstX7cIZ9DqkNbKacfzs
s/4m/W00leokUdlsatzwdTHGEk0H3IcYEzK9nHdptOODErs4gzsak3U/yuz1xsviUAvFhOL2T8sK
Xs/Oy0rCQJNJOwdCSDAw8KPv7120aYCpnLlFE98DZjtPoefrXWq1ffDS9Q9quT95D9Tco03nFxh2
HLYT9OsecdA2ZsQpSjZP2xQglcs4MlDTe3LHQBMaiJXdUGe8XW+h2NesItPVita9iWn4OMHqYsCY
Nj5ldh5va/EzmP8jjWzpRV/1son66K4Q32RMNiT1vL1mr62BuxJSa/0eUGdhXPQxEZiT6VXb55zh
bD4YdmprKUFu6WKPyzN1lBKNpkF86QZBB7/L9XGUMJaYm9bMwD6uNvtJvZRQP545XVUuR6vOLkcN
S09dICMoxM4qPjOHWOBW8mhVB/kLWhYrxl2KAK6Uzzpa9rmaopYgfZSwyJ9QPtPwEu9drJ6rg2u9
teUC0E9tNl6pvC3WZ9xaFE0Z4hPBs6a5An/F6bGxNfRPUAUzf2PPA+PAnQqUidgsA74yZ2XwI8DC
PF2aMRCOSsiScBgvULx0j+mlgD1jFwUMdLGXkFs537gOZxcT2CJiPxEQtvs5oBdt1UndtlAP/dN0
B2W//6f59YEStt4Iv7nWmD5lFf/+6SN7nNrfmUgI9xsVMIIvlcJZcDzzmsTQGL9675V00zSvCXAL
bHtFsF3h6RI3XFShpqVsTBmcpnKggHhn77IPB2ZRBxAhfOBy1zznBDfE+EU062ynRfif1zFjb5Y+
QEPz1aA83lZw5VVaQ7p47qPw5d0QXNoeGHcunxf1z9YNt5me+9nqcG8Cc+8uJWG6pTjVU6DiHWMK
+zV3glHQw+kxEvDtzeZMe/rzvj2vf/Os7REUS61fcrE2+/xeaFQmwZce3nSiL0nSs0q//Ez7rjOM
AFPnJm6vY+xYoG03Dkz+HUMolWJDsEd4tHeQ4/mf/8cZKft0evqel01023iq72ucHarWlG5J6Lf0
t2vbeHk/ICBxiKVHkS1m4WZWh4//pL3ehbQ0TQmBIwgkG1zHBdGzKEyoQIqu8nzSDY8auc8eXz+3
8Ehg0S4Y+2gpxUGhnSuPbN7ZH04JNTSigQhKP7wGm+cwrBqjMu+XKT0qhuF5z2QwR964cJz72eBq
XqeHYYIpkDkEE99zZGC0ILny7QM7bl9yLTA+rxNmxoFvkhoxJPvuqTxAjrQLBB0FmYkIQuXxJipB
v58KauKIct+2kE86IJQEY/MuCBReCoVmIGaJqdj/k1h339mkmXhFhVma7sX80apSJnFN1qsbHl9X
GvFGpDkSesfmX+qgfxIzxoQiH0HXG38utb66dImlxco1VRraij46tOKqW9eQKLyicuCQ/21em0Y/
yUS98ZANQYtiKF2+qaE9GT4rchx10O1ALzkWMYSuQr5pb1Kvdo9338jdnKMbofOZjZpImuUx4yKP
j0hqBmnFlNTOxTVsmxHvQMJYhO/oKvf1UafcMoWbQpC7sMZntLrPvvuqbo8kz4Jt81yTxlg1IGti
PD/hCm25iK6hOe6Nuk7z+1d/UyOzVeQg5KTlTf/XnsJJ6htK1hrC4GY8gL+WbQgoqO79Y1j8WxNV
8JBvGifFCGlG4CYKx+Pbt0ML6/WXjCCqkdReRyHz2zRUl+GjEtCUPbF+HuIPyGrzhGK2Wfr5Oxaz
gxwV/aA3+TfUUYL5jjo0d1i/8Umx9sX6keuv5C9HO+GSWvAQn7eoIwGmbCeg+mGoTNQHaDfaw7Qg
UsLJ3TRO4HrBrSwP+4LkuMT0bzqnA9E7jprkww5foMajqrxFgbdz+pxUtpzPDcR8WpiQ1R5WojzJ
yS7809+yKcR2G7Tj6bkznnYYLaxFNxOyjD+Ah1hyCFfnF2eoIoc6wh64ywR8cBF5hsoes0FbDqLH
+QzflJg6hNBeYZl4yz4KpXxnukicDhEC41Y0wHBLx8FIx8JIKXOxkyLAS46EzeJ4nxTBiOfgwESR
zjh/48McIdn4AOfvGY1uLHNYaGSMkFGREYI2b88es6zCaVb0B7Xc8WYNqH+Vhp9gK9fKmssd2Vn/
C2pD4WhgKb8kXy7OD7xBKfi9s+L9Fj5Q/692bF7mOt/M6mOlkxFUHpkCdfLsl1oMZY9eJAO9eqyu
rcdSrJlCCJuo22zp5XdOXRTDFWDLTA53rDCXo1doNGN0igwCzZ32Cd5AH9HchoMX7/YVNAvyID6X
owvOTP6xPh5ego2N9nEy2F5aZ4Y7n5glF/StRvBX8B24lspZGjqUWunAPucdXijCekTZgk7l2BsR
nC2ho1e6fNpUP7t6zgwcsXY7i/Zwjv8frM27+42N5EkGkNiV8osrQICUcXy62L/y0SRo0eeYQYVO
ijoqJsLy/jJy4A0YQTp+I3bJGAtMPfIGuMGnJT+HgFHbSe2mLfcWu7VugsNvHTxQFln/2+sPzxvE
+3Ea6gkbGQBHuj8v9PNznHQDP+pAe2DovbeeZ+7QqL+82EO2KQutfaR+SbQj7+1syXlOt2F2NIcl
QfJ7WTB5uYbG4wyrots2LqzcnreLD/yZTBi74NdyOEJb0SOR0Nk9IqgYuMV2qbtSQnBSShzz8RD4
H337BU9RHRFZLV7d5iYHpdc0N5cKpeLoH9GuwdmBrnZPhbk1mdrAIqUByF7hXsTBzaHDMJFVZYgY
T/mp/9Cm8hZzhI+Q6yKfDelTGOLO907arnq80Be1qNAVdcf23e043yOI5jTgxzB868Kgm1xb8V/Q
pZqUZrK/kSYqTIFqra9ByS1MX4lt6VDHnb8A80MlrwHWSiD2IQeK4d4a0MWffH1XV1n3zaoZdcdi
Q/R+TJcSG91VCKfhNwOzjAT3kaVR/wzjoIxoJ3cWodl3/pyk6pPp7uAZfg+hGhv0aVk7dJQOE2hY
EeQq78mSR80GG3yYifFzlwZvANSNxjk9a+eZi4/ELjikQhC4OJE9cbWhfj4nLsmXr2Y2jwgmyrHi
TX+JUbb4Ssq4fCsFwASOjpFtz6Gk95sOcXQyYHBWabeBAzHJK0E5AYyNqG/Bn0cp+U2AcpOb0XHj
kpamLXC6Bc6tze0K5WrWVIBal2KwlgfNzmE3rKwhRCTZNAOxr4xdaj2M2MvFVJk72WzHdaZyazx6
2NtagXy+R3ExdlpQAl95xbbXQ4joQG/vMZst+UtPKnUmazQvKB3b6pALA8eDamTEupawzvKy1mZ9
fd9RJ6IBv9KofI7/vmiaJD+zrsPfkKwj2qzoGWmWVjYsdyF+5ed1ibdqU+80uUqQAk8wMIqiVRBm
CXWMUjd5rqa3pVf8iQKIlzPacMj5zqvhO1a4GRhd5Stip2C2jRNE5QamjpJ33rRb+/i/yLrzx9bF
br30+TdNVjeBtUY2hSY95zHMYxfa71rxJYsg46AmFOoAbkFY60805a+I4/ro15HuXwO9O05EQjL3
dlHGzlQuPplfzrW//8Vhp6/lCCP2By7e20reS6IsSDXiYAWxY+CAUnlf/97vXnSNmMd8j7rBdjwz
jWNIVVFPO/ZkLNHPLXws8gcray5JSmoz6bbQTbpr8QVgXspMaw++h21HQcln/Elcy0BD/GLu3CeQ
B335fOd3trkMjNpdFNffNEviLj/tusd4LfCu8z8opIZt2cBGw8UOkEs6ntUXvjpqOwx3cOsvlbUG
l+v+rEtldIqH0pCrxoR52OgCTxJFcW8zRuO0c3w3NyxaZiclgJ8FFy2IZh2NfbCf3QLqM1+gxi8m
AdJQF+d6CR7T5HkqQXG/VlTV2KQZwfX/f4eHbLHDbNoOTTKMkzgBrP3acqcF2+qWgiOxrap6llI6
2bwwi/to7TrQrvW0DcPGwNODkGTqOa901xC/NABGfGe72akZ63CINzYjI6JJaiHfn8r1o9tsAo7Z
p8SADDIq0ResgFdorwaJGQAwcCHYvuSJd30EHU1/UnAuSg0FVChEVLjr+cTkBPaxjjL3Him6rjCa
I349FggVWZMgbiad97ebZVBtWJtagv6SAOr2kEM7oSjpKeZky8GomzLY3mJmttnhSdfjJQACJZ6t
Hiykyk7w3ZGlz/vF09FRcl1fspMm/zXbqJT8MNfC3d46EzauokaFqgedbIlmq5hyvXV994N3/Bz5
Q4hPUYS72oJbzUUFkX33DrRJ0OC95gyGAK7neNqTZKgDl+SmbIehwidOWuTore9nd6yxBYJ7+Zdi
VifKmRGwE1++XW3cVxoYk7aVGfc7y/0ifuhQJ3rRMADaAobb4vAxVAT7hX4pmiHI9nYjPMxqAzXK
z5df/UEfeqvp+M+QW6IenGZcB5cW7S+ZeBlUayx9x8eVLWkygjQW5OP1DE+qMJkOvyOXUtV6xnxS
3/2cBY49Y8PiVGnTgz0nXARt/BMbJPjdyU3fDMgIUMmmtz/54oHRvb55pj3teEfPtRO8VycZhBvd
I3VIA2QJdhuzDoOMHzav2Lf+yqpgrZyAJ+7XoVQ4wyXbwqitrO48hmELiZGMfuw3IqFIS8CSavYO
tH8MVDoT9abKpOzoC3UeGBqpPqQR0Vj4KHL78Y5AqxJrOxpOxWHNBNzoI17KjL5r5DsBowQ2lFKl
hKVfnRte4Ig3BAlVu/NP2FX2RKT6eJTG/fharanaLrWyudp8Ori+TBtVhVNWjSDICoiPok42gLcg
/K6VoQsg5ERuEDigxDhxk7CvhIT7vPfSEzc4EvYrhAaSu0SHvZBlVb9T2nBJtINwhteaLSmxE4Gi
YgPrjroEXZgAh1epIH28RJyWwMFCyaIrGawJ8FNa5wqi4zhOa9f+CK5pqcy9JIr1XJfTJM9gEWo7
ofZYguAUfNZnFOn5jhJqMDtVy5Y0/GslqHdGNY0daEe9r0I7+SLWMlOIDR8WJDd3XYhG1InsgKNR
VHeAa7pPhVNg37eioup76/q1RwGNeRtWJctWYv5wV85eFJJR+QBWSDliqn02VlFmsB5pNzZhRSAW
GG60yxbxucXgxZwWqTFw48Pm1VwPfFhFb5EKm+Rx8b8rHFdo9a7Zvzn9L39Dx3Mcme3gjGKZ3CHM
M80Effv9hSM7LvGrKJ29M+6U0JQXlZU5Rf+1f9cn7nLMH8kcgg+8T6OBHhl1qXdnPnvIc04ms9wS
PCEZSLm5R9O/BHNhr3PX93p1sNAQ9kduY9unZ2zwD+OscebrlpcFFLwl0HvQgW0hWKh6ey2r0r1C
y1t9N21RmyJKCbCs9eckjiqLIkPV0aCrYxUlnscAx5L6J6W633cqg2kbLmBsbWk9Tcy+qEnCyf91
fRQ2jGcLUeCBdINuclkbA0XCWA6MpkJKTwVQQ0kvyYTZVoLU9PEvHy6KO11fPCtRjgSUQt1iSNyx
1vZ+xEWlK8tVU1ffR5LjzgI3B0Eo3K3jusgYvPKw3mJU0mQg2dmJt8zWvo0gWz1AkgzJepp6b1U8
cyzYFuTFcWlDBU/ddvuV7BpdSswhJJq1BQlVCNoksNcdm3Jqd2TGPFN9E+Nu+sctTpOSg1h+1VrF
Kc2smSotOrLbvrcsiIVKsmhp97/jbtISjHg2Z+Esl0jNndP0IPhmLpUDmix/O5zJ5mLDI9T4Sf3t
fz5ygv53cpQvpeuTKFJ48cZwC1zLrYheOpDjQmFDGtrsYgVsFy9FFTqIgdy7ft/tjmLpYcyCKRG4
3fIge28EH4Ke/TOphL+oOCYBHDwh0OD93Uzq8xfTJ7p8bEWPyrdoZCJJxtVI001J6qsSSfsnktj0
4N09hSYRp6ZIYRPUi6RZ5OjOVgrsl2LcJwcwAIEwq+u8YDheEp7nqLEzkUh788IzxHV3J1SFRmVQ
BlXdOgJu3q75nNO0JMxQNtfsMFXGkS7uMeVHZfKe6v/q4QeDbCU3s6F71TJSiJxVGup8kB2vCcGQ
o2MJtctQnDN3jD+W46K0+Afq8/9/2t47lg/MCBvssDjxwBgafxflD/n3rU3wEXZJ0l7e0E8J+R//
FAlSDha4Ek3RurG2iFxcqThBr7Ley0zOzwV8FpKwJ40W9gr51iNTpOMHA5O9ssvugSSFj8qfGQqe
hpkZsSLr8wDn2nMoPxrwnWqrEhD+2tPyp0FhzhjZBlMCyTu30edF+Tdn6LpnjzC5n1h89lhJTw77
hdCC44Sfe9K54oIxRbQSumtJqEMuW7H4D68cxoSCFxzgCx0y94mHIpKy99Z1zDuTVIem+jzngM/L
9h3Mpe6GkB2elSZ7qGAWJr5BI4mJnjsu1XQ499WF3uhmV22ksb/dYY01zP5kqXolweFSTExZU0kW
kPLDpEfs+inzwanW7xLpiS35tB9gXFjyj9UXoMfRjNnJn+nSR1qA32VfkWSgAOMehogYV4p/nW9v
iOQmXeZo5w9ebHrSy7JFklbbSzIgdt5Os2ftp5LY55B0bMTr5kBx8InrM01nLA0lli70v2RiWQWz
jVYwblotlXKjEDuckBli/I4CID2JSZ0AUshJfY/AzX9hoK1V3AGmJd6inlyHcczeMVMI6WyAuPrz
kRvDjA6cefLqF/6Pm4pyS0rAq5SlJ+EGyXUZVA03fwV6v6zs3GbaoxgSmfc+6tejN/iFCy3y6hvm
xsyvw8VMnzQv2namHPOjPTOaWVKyY2NPFb8VhfPs3QUGGZYeNGV9yxPjdBBz9UPhkXkcZRVNaws/
C+t00a7S+GRN9dm3fpUXjLBP6j2EhBmLsBn0Av3w71yz4+Q8mwwdDqFrpklWEmlhssQzImD1b8Dl
WMRXnHJpgAlR48OZlq2Q7vseW7JK64ahgfRoWgaqud9DSpd1FLLtUdkl2NtwTKofD96b1JLQcLEZ
xQBl2cuVAUQLhA+8TrZM0XECm6ShlqJUhEE7RjyfxwIBVseJREXYIAiJOKgIhyUjWzoikGPc+Sqo
6LP58x9BqZzJ7a85096nSXOxpdePQ/KqjGDjItaIVvG66KZXuoOq7D1bSmx5SyO29KU7klrwEG9T
EgCuMMOcmg89pecqi8rvwXzPN7ZcjquxxD5loKRnyiOJnKfDL7ZKV9L/87Wp+xx+gIxkvRSV+gUE
CiNa5TTUrovAMEtWE8DxgoGYUTLcNEsKfpLDAR+EftQpAqXDWBvic9xJgWjHqgs2GJWOpJUAgLap
Ch+a1TpVr3bKTSYg4Cs6QJZvfqzDBYiJWLL7aOmdTWHEu75Ra+Rv1avOafsmr27VlYFi+SFN0pKt
kuf+V+any0UrvFW1BZU+QgM67fQI5wMJuvnEUjr1bE77ME1h5rg1joTyb2ABKD3z/JGrgQpIUdra
NOWpHapa41NJzJLDn56Ja+gjPibNnwU4qKMzwKylhKTj2AnLl557wfvDyihPErFbSkH7YX9wHGga
uw4qzo3tsFo8satYkwtmf4bA+Ipt+gjLoBcp5d3PpDTBIJvRDyYXesB+H4IwWVFgbDKSAVJEJc43
VnklhIz5SJ1VBrjtUTKUI669sG8M7p1sXFzo0eRBaJPrDziOCEqhI2klQKeVYm+PiM7mwxdK85A7
ic8Cj+ahB9NwAqOo5b20sv5b876B0CFSkKQYypV/mBovfeclMrTOpLbW0x90pGPDqHrMU8xVB+p9
sU0HlZVEJN1mpKN1l/XmG3en26/dVF2dbiuDEKJ4F9rUuzkFa2k9X/xDxKBn9nis1YaeIf9J8eqF
Mn0oPDVuzcPrS8RYzKofzkJrhYAzJIfy0ye+5XIx6PbflhoPSebW/6FdT5amiQmn0Egk26kT2uv+
82t+1PgqeyxIebL8NSVphT1lbfCm0vXuY7ssfx8ivIpEZTMHUUZcEEgFWulbvuXB6/QGbpJ6y+tq
LnNNb9IX/oQ1gfb7nNz/JtENFmIL3D83fAVC4zBA16tAPVCSw/SoHwrhQfN1ecK+cbldHsvNayKi
4eOnyvLs0PjzFkBLILK3N3bdTUj+UBvj/MTMvbkIXcolp1WfaS5y9EjB6bbNumRDYsNsN7MbNTW/
Yqubba4Gi7X0Udaw2T7Xx52aBPOSsMBf7zZr3uqPRtgjc0/2S+NT7NR24CJTpoerFgVPgjFWbMFl
fXEoN0jry1+THAJmI8W7clegNWl7Qo+hwNEhidyx9V6Z+YtuYw9TljV7OtbhC2SJi9oApIfZxJ+B
R1h1jZgaJinz6tonot/zdXOA1kN7sjdLPoHlI07x+mCIhBdHALJZSrRJ/eDVBi3wJFNOkHJ2vv9m
17zlHbdl5jaXu9UfdyNGzyj3oXCcwf5tEX+euAKE2oSV8QLzsBCqh6NTupvb6oud7pc/Y0WlCAW+
/N+6Ukv6XMUms/5vK/6S2ZgFhWHyF5CQ2ZKPsZ/bv9q/BsPmkihUCtwpjCwTS4FC5SZigss3lHo1
zwpR10Iz21HUFkdGBUa+3U0u3fgI+02S4k9f6bXSbq+eSgVWrscbn3VXrlDjU71qAWICWg2qpkPy
gdJovNCnhymmJ5nG8xWlR0t//7cypwiZbU5pTNZ2NJb26OxCkeEbtOIbwpK/CqaHKxrdeVX7OK/H
ScxH55c+C3u1MYxN+UcmMgRPnweKEzf5NY295Pivu364m8yhu2OhkgEr1uHShpDCWf2mVDzMVQbn
t/ufZlafO1+9sLM+/WrTG9409tk5d3qNS3NWk2n53GOFG8sqZ8gs/ojMHpcjxWCpGtJJ0KVQ+I4+
VokdX9nMp5iQboezQDfYKmnfvwtb/M0jlYxvVaWcO5JTKHFW04ciBBjQjjNZWcuDlm+2+g4xkPzW
8bJil8px04bwsHiQIPBcHxlhB36VD1QREefvkHroXSpct7qaqENrMdlNg19KVNrnecIk3pxSGDnC
ALyMcaiXeWGTJaEa+Vu7jVluI/FM+9rbnZB7zIjmoBxeFCXWQVEPxzYszJHrCBj346BuonFTKTdT
GO/JwNQLgZRHfkY44uCbXBknyiYevGwqLesgYnWV3hLgJjV57lHfuf9ZaqYPnV2a0xTB54T2FZ3v
lnkJdXroS1UZhPU9IlcR9bXRuMj8iI8n+mTH7ftUg5Hg75SiA1J3uYxPfEiZir8+EABvjSYFFRR0
+RF1MQgKPKnFco2zhpLFHlBU+Bd9fsZLe2fQ/yIGVZiKtPPns8wp0N/1AfTLTANAKtjIzV/E5P0s
KVufsqSmh8uTd4mTSaxsMhJnKmspy9qoOwIPHE+Zr2rae/PVZnHx/XBlwqFUqHCh4SSuAhuSdQ3D
IL5VjWQ3LlImwS/Ok31+SeK7SzvpFWaXUYpC7Z847pil9JN9cXXyXqbaDqydqyLjuCR/cqltzziI
Rc1wqaAO4dQvDKf3xg7ElEtIy/zMyZ2iPNpUDFM26lf57dgIzhJI2Aps7L+54fMyp2lxXjIZ1E/e
e5t6IlBVRGze3fu9waBF6mAqTFlQ+g9DrOKjRz6Qsa0mHuutCjJNM3raDjL9AKga4y6kkNpDc8Q/
n1FUPj+usUdEJCxouK9PQyyflO9vOaRVcwVnPKSAm9y1bFVqMmG81jCM0ST0imoEnlxMUgWrz4iw
Krwgt9uycJv0X+K8H0S4mfJJopXUir7cWMuhIHLiX+3qM4nl/ttGQcetI9NyZyeAQYyjBNgUwyEn
3cBx9ADCLu3LNQLzkrNYP4WzIq+q0wJHO+56SxBE1CHe8tTTKSdHIYuY+ykQWhnBWFShDotyIHQg
sCcVYr/6RC2+BwoOBHvtNQfdQDNvgRSQIoy4pzAGBD214hmJdnOsOu0dFC644TP3VHXEsynYa0l5
bDfmTLMvA90oaz3lMlzFhqxi4evJXxpL06zcucyUyVsPB38QE/XXf52UwIIGtc1qAsPGu/+9ZVRk
i57HQ2QJPZ+aGrxgy9f8Q4gAUZlXgGNpwVCrp2s7E74RS3TSl/qk84yJ0InxmEOln9RaaGGdfSkY
4WdODOaj00nXVRQj0qAQ0w3HXxVLpFz5QdrewCAvryxVNEQdNJ9PdL08pRSYe/jPkvKrwR7PoSMU
Aa+jp+qXr9CLQBdL48HBEyww4o9LYRk5a0pDeFmhqzHGXHyIRThxTfjoLZ8IE7g+Y4XdPilNNe6i
eMsjQIc/EDQ7d1WN2l4PlMMRKsGjyE5u1ZlygF4VG5Rz2Zl1JHrmdHRIO653Ikkz7W9dE8O55xbA
rrpM1oIbNXh6j1HI6sUfqK2QE1jgTOGbR9ansieH3B3KA2WO1UT8KIAJZgHNPPoeGCrckPush6rB
v88cFE1/O8v07KmbIw2cFsW8KsfiS6oJdWDL3y/R5VmlxrxB8cRKrf6xga2ovKAf8BPx56gN4ICj
VDwSzZNTZHtdcu9mxiByPH+K47oLGo0tjbpLjF9kSEVPrqCmmbDxz4C6MfLWmtFjb31BD4/Qy9oN
ADRnL3sJgZOiwHlM538wtXUiKhuqQ5oHkJ6HecFimh/45vfoAr7GdqNYAWQkFqa7sPaT8OgMSS2+
4ooyFzoNS7azU7k/kf+6hnouTcMdETSGGUFOV4s6k+9hlzUIDmS0fRy5wZOEX7Moc6ZE51id5XN7
hM18tiYfKcB3kmZ5SmVnUN+HMkEiIksHBVtZBaBut5097t4hWgnJgf84mlj4tExZHeC1C5Qqs+4b
BJ7aeJ229Cm7KfA9/8W2u9qGv4+MHsE4CrHMQXrMs+rMHgAZDBETn46FyZ/AzQ5vCHlxgu2AftoI
QKc7n34T3yR/1AYiL0GZiRM5T8/E59T8Q1jpetfak2Vv2iWeXA9C78I6+8oGUVrRoNm21kpGlnVh
kGreaaafMJ3CBpikqFCEUWKVRE5IXXMMZXlwGlX7Yz9I9MQ6R0emiXUPAy4OsGMnIwojityQOf99
nV6i6zKNmcrK9fCnNMyGzVnZa/LgiEAorV68c9yEfQfXihcOlxyNXCdTR+E5ePx+MZUfxIMt6N4a
OaOXgjc6aaKe4nVF732svkWqy4i5ObMR1K91todJYgoo/gO7FXnkJF9bG4ukXQgdkhm/DJ1/CPEy
I1A+OwuH7i5xI2734c6WEY4fy4rj2jhw/CyQsbHtD1L7/h59Lf7YwFU3Fa3JR/x1UAMmfDiKlnJb
3EoFt05LFySzGbxrinuxHn3zB0tdRoGnzgo9/UKC6qdZOiJZg4TjfWhY2zrcJirkOYORPJ81EwIS
HZeUXSEt/BuiijJqvJGA7pfLcZkJkBsb7z38OzM5v+gI6zAOWLzFif+REGRhh14pVsqF5okSCMc+
seqIAo9EwA+ojgw6P4Dzh3wqrtuMuwQcclLJey3qA2TkYWcK4GtJ6Di8l8e7cR2sQGEHyL9iGQIp
bDQN64qVA9T/oi7ueWLfuUz5p4SKypyyUZscyMs+1ZfxidMXhb66NexMn7FYeZpNdKCcctLfJM4v
yDRA0oXxNTHAO9upaLrA4IUmZSts19DXvjJn0Iv+gN2+++YLuzbtV36qRp2BGEK7MfKFSFW2jI5c
v6zQ6SKpRO9HwkFkZuSZXT2qsMUATE6RMFN0N7f1hZWJFRf+peVYhL5r7jDsHzB/D464Bm5qHw76
uYTcUmGCdiOFPOMa9UbCdGPJRFTDaFhpla/wxv0SuO/UsiO0v1EztNXdJYjIAcC54N1Ic2gnvjNi
XQob1AsU4kWybRw3Zs3TBtaPhHNlhlOwyne3cm4xA0KHB8nV2rgjCu1AaxM5J6jfMAZifoaU7rhy
y8lP+C+VsOJWSA+D67Scxs/4bm36POGHyCKr7tcXcf2QsODHBbN+IyCauWWOHhFjImPrBbG5cEVF
3CVKw2QwVrTsddK2zLlHArjhQInKzdKTECEsGtnmQkZu4FWP9CEerlkoPW6GgdN3AOapH26r9qGC
SN4GR8S/fII19hxo6KbVxpeFG//10zBG2K+11BF6Ig61mP9kJsYrAvDmdkjrDTsYZ2eSXmx6HWpR
n36VSiP2wU1IJq6LkWBxunMACiSzqbQnS6pLBoLtoWF3QtxR+ZoDEzNpvezLVZh9bokhfkm/VJxU
2pu/WPHfDxLLTOAODoaZZHpJUHi5XkOOCIU+yF6TvvKUMDk2C/bGhVYaBLWPspp8Id99AMhFdLMH
3rR1W99jNrXI2aPmp6jwFEdONIH7mPhYtm1yKuULEeG9biVJz72VF+iz4u7Pf3XnzHH+VQ3byPOT
su8kwd4evF1pVKMT+aAlLNhf31lypkphGW5zKmKX+d9JhF8YFVIL/qi2IegPU3Fr9AmWVO9+8vhw
fHvN0Rio1x76daJamvZzkCYuUNVjgThFlcEbYDi8JnhS/Lkj/coOS5F5wwbhB2XRs0u44mbVRAFa
U3Oc41U8QzwY9P2fnHGYABvZT5Gg9BZAu/nVvVjZcC18jladxbnuPm5ktQessXxlzeYw49geQgV8
lhFFeuCU142qIRa824qTONYHTA3/SxyK33OlrFZ9n4zMKmp5lSdwaar35EPRstTEm8ShLQnsA4MG
WBAGZbcqnx8Q0I+uJ2sIpeUIQTRQu4IrJdPZsW9C5wdqU85UqXsVTyZ7qgme6GhZ/x7TDL5T7Fne
sgoTeYWpW9XRrWCw7rcUiQo7hKWz1haY+KZla7BUgqyS0nobigxFe4VLCHONteV+96qY7XN5IgH2
0BUImRjM2M6OxG9qlEOSxTzAz6nWlBk2uE6b3hIS0Ugb7Lrlxk/vJvYacLhppUNeiPaWUu7o9/w7
IGbsTSw4XscuJmEHTNbCAM4jxtnU5mB9gat8LXc195gDgy2MpDTlX+xh20sYN6zlgIXOF8qYPqxj
TUkiwwcVLTrIfJHxk3Ns3CHfS+pulU84sy7Tsvh/2oNyx/syLqxPs5HsYgUiaxRfL/hYJ/DuoXIH
/eXFSBIqf32kluPhVIJYLvkNxBS3h4FOANbyieBVkQkFRY5LYOi7T6hsYIl2tBqhtLr8l5EtbaCV
8XZ0H91uOogxctX2QNiERVXVo+e1YZDUGyibCNgzEjQ0vfkpbTJ/FtX/Ph1+zff1lbGQ+Ix4UGzl
G/YdpeSi0FzBL1gdiyPJL5pQqX528p1vMRY1EIPIW5TDWgi/TOfEQ/GcLwOJFLB6wU30n9xmeH1a
SFhU6T5NmbJ1lhMnAfEQBU3zjIDCByQ0Z7eM+LYcXKRFHFUZZqq0dDVfbepoZ99xshb3nS829aL6
BDEEeKQ3+XzEaA7qtgEJKkh3cKmp1sJAGNFPbDLgA7OTejQb+Io3+EzzMjCcBR1yrrRj6YgFp6Jy
yIxbwSM2foVb9RSz+cXTbOxZZ4DQkQOvfrFNi4fCmO1PRa530tv3Kg4pykdL+crHbj4f1Z2z7A3R
w+2urMj52vxumoGF86ZyD0QgnnR7Y04yQrMSgaOp8+P5PjrFGhkFkfwlZFrUM4oF2ZIVpTKAJvYv
F6HsQFPsNfIpGxxBpw2cD50/7LGMAzpkfqBsqcjDVT8GqEuKmXPufn7CZl+WbDJpz/QxKYMBiYI5
WX4sTNND6VoWV8R4++EOvzWhKzJbqMK/a0y7He0NZrvx0eznIfzJze6t4U66xRZuMbcbYa9shlX1
0y0lU/QDfbd4cHIYB8DN2fSyDb4lmbBW96VTNk8liqiC/VRKHwX2hNIGGhfgQNw0hjlbstu8VKXH
jyliLQNZsmB0Ahnz/CNk4kEpODi8pgsq254E6lIRSjSuDRwIb3ZcuHS4W+fQieuwBhkcCRQghiyi
638S3tJFzbWonRHneNqqythuxmEUA89Jtf+Vx7KiOoV7XIpxgAbouX53s2kIL1OEEJTFLrNnECGF
j6PqnjlC6WyZNvSG6HvF4z4LDRsvvZlcSKEr5wEkn7jB2vZgLnhqceupyXQGdrmDUOhpxtFpMoZg
aQW7FI8J33mpaj7L3SIKVslRSy/RzyY2oyALIe07m+MhMADe5iPq8mz3f0Z+VoR8SlL1kWLqtI+A
tGZmJIuZy9QHk8frNu6Bh7i2yf9crb7Wqk7uyRkfs7pZN0bGUFQz7fcEV+oMW3AZdRnfx/Fqdgsw
3BYjDVkzxGmmXYBURxIHJDe6ZvLTVduEy7zY9Ee//qHc802mKHvs44jtAi9kwjj62IlTT1mgbypH
8te7nzOGrEFNh7eSQSr925eHVyEKYJmXjStMqSJqz5tBj7JSS0HWbE3lHYr3xspTneFBnHB7Pcid
sR/48WdYxbhRgZfBKnxjjkSFcm3oWGVRf5VcCJCVvV7t1SoitR7wEvZTPGWvO7PpvIQMp4FuWAQ9
ULIpJO/0B61aHJ1sMA2gu8uS8xVpDjAtxXGXm5Zs5tbkIFGVEwnhjj+5B4EKIbajYiYv1IXMEODE
/NWDdGWmwP+bKAmVHPHT8shT1qZTvW2kcg8uxy7pl+SC/e/ryyo98ro8tBjvGM7qnVRIr3soCI4L
Q/lSwK0oOLWC2ODi3JmTnJnryvy442rvKxDgVd3K4UTKbm/i8qkeRrO7JYT+Yl9V5Ya4+MNfqKOa
p9CY/dOSc/yAW6yHJNEk1vdLIBBdqxxojdrlI5AYYlFYiTkBLFztVeQm27+ZXaNKvJyFhWxM+Ge1
dzqK110KVI0jhqced1MP8bVS91ASH1p55P4dvhZ4p5ok6LtpI+nP5vLipm1vtoePBS67xqxykAy6
VtKmpooZYuxNEq1/cxzNgQ++y/zEy979RLIWgdfid5CG3TtjrFOJ196vAoKy5DKGBuj20HL1GhQs
A/pqJz2YlZ3L0Z1IaPpjMjViDp+pHAjW0lamyQVm8hKfj9KjspjuLj++5EB4PP9NXq5UVBg+HGWN
1lO1sC9HFVvcNw1FW/oYU0gqDgKUDvg6uyVeFztDdErEMBU3ihPck/O8tPiveu0Hl7fZdmwCxzEN
Qy1eG/dGTISPCTI9yACnFBKopyKhdWDH/i+1uXGOP/KjCqhozcKumrgRXHMdMPuelhfG98ZurlnF
VHcmiLqK7ky/7DAxiUDuixT5D0cwbk5uqIrg1byeOVPQ2KnDB3c/joAKj+bbqwM5TIUcOhIBrKx4
092i8QHSDye/eU/H+xnHN3/A6ys39mx1BuhlEUNaOfcHAPuAWwHvElWxgDkrnGk6H5DVyGmAGi+1
Rq83kox2kJkWW2RleXywCh+q1uI1wUFlLr33wV/WBVMSHuSiVO+EXBdwGxHzsIySV+/EKmildqTM
kaAjY32ZfzMAhY1XBtSju1onnYqEUchsdNbjlobDSQRmc5Elt0y6qHaeFxEtHyr05GafJE1bGV9Z
Jts77eE9FpWOdtQ3qIAeXcS7zxdbeDQyLwKFav4fze4ZmVv4HmDEw2aBNergT+e0JuYRMUYn1S3U
1B7D8kBReswgjQM7fyDXxIOtQZpsrrBwNW8OTgDIztfvGDWYZkwwadDfWwe1Fzod8j5DqFDXFuft
/Ezq04OPF1YXYJ+uVkLmJSiOmptaTlt02rYKB8n1fws2x4n5qHRR/WkB0MQnzYT2Hq7vk2aEHVWB
swELelUDaLWUVyilXXg9EDKfCz4LnIBZ4qdkNalPBx6a32SjgAOaKDGLRGbJ239CwA4rdVDYWCym
1XKen41rYdF+G+Rm9YkrcwwPy0ynVE/gg0UJpLKaDyI1pusnwAOROTnn6LsKk0/+NE+FrwgSptFb
xSz85S4/KY4QwMy40rrtDmiu7E4KHy+pdL1vjeltgWEhOlWvKsFJ7WGi0JZ6Wgmq+E3oETGUGtnL
DLC/nJVYWsk49+3KWdnmH83BxAe9Uqd82EB4poNyArMgBRN93P2Z8L7F3cI6+b9pCXxWiKC0WVwI
a4/OdMXugtvqtCsgqCjqG4PANShFg+ngPQ1kOzWOc1xSUci4I61qEIZyE+fTWwPM/PAzmXp8BuBl
hTHqR+nxmMBcmQJkTeMqfauzzuSXHUgNU7UQV7hdbNKNJ0D/mCcDhXCFRidUREiOfDRswoQuG3zJ
zJhEMQZEW3K5FS+Be1Qrx2qwQl3BGg1/76PaNkOXupDsm17shVpzH7O7lg2DPCVYoDAlX8ceBpl9
DfwEG+HiNaFW5+LWdc9Pp9InFIvxNvnG3O85Zlei1osEpSfaU01T/CAxAYpeIFKRHeJnTN6fHbCq
rzcxeHMnGmjtLLb5XIjPUprjFiyu0LpOyPXtrQ/OhZw98UFc0D1vNM9/dLBpD1ZsnvLN9KK927Qm
b/kgdzQCpqATwjL/xReBXKWsy6BE9chFf3svqE9yPgaZfap7UXI5eCXNfpfawArqAczlHmq+/MSt
Q2uMoBAwLBSQPWtjRPFu7aZPe1O/X+pccLMlEihyHw1FBj35h6vYZKFiG9vwHABB2yfUvPDFlHD2
UwsxGpREb4vYfj4RlL/9EG334NO50v4VV2YWKuKfDxdc/RrojQK908r6Ftb+80ISCqhXCw2vIWz7
t9JK5cUqs15M+2ixzQLcJ1JTCpLnKfhzSnRU7BQT5pmNsR8XFEjp6Sra1o7xTaZWPTjTEQbm2wmG
KbQJZYECRyHPS42b/V7Ij5B5xX0tsNUp1JiGM3xo6gWliu2qHZnWtd9uIMRPy8iRpUQPKOGz9Zek
BJd2NtajgOKpWIB74oHzlhDR8K0h8JbH0vNPZetDIQZJrbwKlSLzpWj0F6VFT6jx85gDlkYKZIEC
yKYGh7P2ukTCcuAWHlL4FuxFw7KfvBjvhDFUqqwjLNyCtdBwXnGYBl/RRFDkGWYZo+ne70rRDKfE
o6ETr6bmCYF7cBL0HR+ikPlhFCQt7BS/xO5VgvfrWAaQP7ahcFGF/mmK0eIvlnqxnRxts4q2NJIS
xjbWFlqAXhF8J1mn+ik/LyyoiUS5b6ahcT5zmykOZgLJkWtSwtZuzvGBTkrPLZidMGIgqNMS5oB6
jiDbs5/O1MWdAmW31otzpKX1ol0oFO5Px3+mCt3rP6zEIS/iqh9TXQNF0SUXnYc9HbDEV237HAPk
Kq75CMRkGGYvtdfvCCKcAWBiJYRr+LeRfgPujhlV2bJlZegTISyxZDjUk9LC4KTWdNJYstr+WRMU
Dzia9DUiKNtYpaSpTIi/Vl/DG/zlKw//5fAKTv6GPa0erzVvJ/BL9VflYMASUkfAwR+3TatCQDl+
b3nDOedK0vNneJUB1M5GoDywkwEazj7Vzbc8086uVYL+62P0XqCNotsO5EkTtiRm2xw4zutKVuqj
y+njq0Zf2ZgwNR9sFaHFhv0yYmyR2+neBjBb4BrwN2DlqTiWhWVvRJUTjdp6scNVIlKMDSxzwW98
mTiL1eGlZOzxINx9y2gsb2qGBpD2HuFwtQbryHjMIteUof/ePDXEfl80NdKdmyNR0vBiS2gob3by
vSyrMTxuLx+7jCWJWyEruIT3tNru7Rs2fxEZLl94/OZlv8SAOk3yY5XKPDX/72fY5Rc5PeSe8zn8
/AlBbz79/nVANKOx1tVMbpaLpSwjGypTXIe6Bq7BzI/tMepPkNlbrwdGjafNjNdgUlLf4Hozajk2
gDK36P0y6zyWnClYzQzn3UeDft2/nCxK7IVY8xbqCGinmIdIJ43ZPteZyVJXrJ5plf+RW1JFCyOv
vGQfhj2NIdhbpy0EKEy1MP57W5fNUx4D+ADGltX+3JIp+ilRICy32MyiLT3xTflQZ73WCVI8kv7o
dF5ZhxTDvWMPjJHMmhQIbIOJOTmcUrMZT0s2+LI1K0iqt2t0fKGT9vQxZwWA6sUGtynNtJ6rVy+K
y+yBXh1ykXYHTFr96OJ4MtHpr9EYHg3Z0sXEwZWG9gmF0PzNAAO4Ggd4Lij9MBuJQcZFEOgQ18Nx
dLbFEZtgeDTWhrNx1Q9GHJZ9TZN1vLjVZ8E0/GMpOt5vL12XM5hvzVh7RQP2nDvN36pk5ZtA+n08
l1hq94OiCtCnbZpwp6GwkpApFnjpax9t0m8KFbEi1KG/NyM21XXH3KephqszxuljsSLk5DDUWJND
+A599rR8mZd0aVC+VysDs32shGCWUta8f/DR2fcLM/Pnr3QLPN1p8zG5tCJFHoufwDsiLOdvEhZV
IT87vSmJK7vZvAw5vg9TJgpLabzxQjFyZnt6YJ2HsBp/rGGX7ligwWJFSa49Hu6D6qamNZ1C3hM8
7/xCTDCGT+u26r7vKTa70xUBqEqNgteAdt4/btb13Q0r8IY2xNwK7rlhuBAzYW8EcKYzqZdXs/xA
7zLNVSQZVmV/mZRVBdyExsLWlklB46QFDRjPf4kwd14XfxYwARj7+HNW6sSnbYvwcYlaqslAVOYF
SfSv+r6QrNb1TkVVc4401AAZn+KNV88/6l+VnvdRH6FZ4gFqiFl3Rprk8v3Pya9qvFzQkekWnhmL
PwuSiakt8yHsT0D9asZ65J3o0S74BrzTT8ncETaPSJ1ODMHVIdnXzs2tWu0uR06uZESfjWqoQcF6
v45LHko0iLG+jy0n93Zxf3eFAYnlV51Qz2bfALAmFv5YLXxJkmItJu1v/cK+ivU8KP7s8SzVHdSf
5RGbXGeGqJ/TfKofV02449pzi/n9k9rBOrKvGPIS2oXW7SfGoXW3sLQCSk0uMEP1lXUCf52pFXNX
Gcx3T+Tc2zgTY5uFSs32QU/DBM5+2Y4BeOE62b2Lc/U1902SM6N0A78KszsrRQ+Y1VgD5T6mP4b/
+MTsRPi4ZnN41onwslLLb5NDeGkQTwXlm44vSDKc0PT0pZ36FLgN7ri0UcabHqmtVlpgjqhEpGd1
5kZO5Ry9SUbIoWRMfS/lRMt+y6AV1KwgTQx+2r+FtDqHqARdXa6dXNYBUUfq2wbWke5DcdNGz1ve
CqL7ET90Jvb7NS6U57iesaCtCHwPmtstUeJDTM8/ko7+MW6+Jl0n9CDCKqH+dOV3NPWbxRsXK4fI
KxGI5BMGLx5nCIhnlKw9yBZXsUj9t5WP6Sg5z+zWdLfYuQaAqLmvfJRFSPHR2/a2PumQimFeKWqb
op/W/BtWQXaO4sK5LsWIFtAg08UfSmoUJZRZdKskEz1OpiZ/hz7FGQtONjcU6AsukzJyr6Amxnxz
n3wz6kGKn1OrkRx4eQEHS5hWWBe0W+HdQ2Inv6XfSkmz9P4TNMKvdXg4O/I+ZCPTysgdeTqgQjob
SqrgSpQOS5L86thGM9UfcjMRFdnfo90H4qd2sD5/NH/KP1+5/KkTxK9ihern7UYQuf3wV8bQ+8aE
O9aO9ahJwhH7+xdIFwcmRxNWBwXJsb2740//TdsK4p6jw18nChU2uZ6u0Dg8+RM/bzrOaJD1ap0n
3mDSrhT0aSADDlJzwOpkLFb22EBGDE5f4ou5HJDtru38iSg7T8Hmyv/v1qivCOcgbpVKwcBzhGKl
Otjd6nDrL5eioTSnwzFQRxMXbGJLLg2bTNHMgdT9Vh+YWTbaxIQmmWZjD+tZLU13doKerkB6hR42
kIqYGugO7wlFYQ83WFbD12tUUEU860Gy6biyh/fbYi67q6KeR1RnGtKsjHDrLtQXT3NYgcVF/AR6
kaxK9vwEOg3zOTzPGLgjQ1S+9NN7lPEAgNz9dwzME2A/87Q/M7nU63vUAEN8Goey+ueSil2S37ra
qJl7SN2o+9eDZ71g93QWTTvXLr+ePxHwwv0a3X+YoJ78b87pNpuk+q871tfB9sERj8/SB3VHtFIB
nnDxjtVretZKHc6myZDpc/2NTNs1/Dvj2BAyQUKPsb1+GlIoAC9n7GZUOpRjsRD0AhlYDznRMhIh
UohuB1pnkU3G49Dy39t/Km1c974j1yJmopDHlemJnMKwAax/fn4WEWk6dUK9ZVFr4tgyhwGhBmmE
BWyBJA8Z/GDonM77dIO89IpIU8nl18FhUgl8ERWw/7eEEKMqvmBxddaON+ywH5IK6feFC810t4jj
/dY88rNbhXnTdc0ek0QchPF+UZKK8IAFPJIllv2djtCZk3QwwGCy5uP6aEDz2vQCH3YcUYDNWW+y
t6NYIy3Qn2wFg/CdPGOR2308mxaKNgLz2f7IDUhu8/If262FlOsMLpmZhqPYLeZ5bSTxIW2wVwYX
JhzW4ZIvJx3nymmsKGzSvJNzd3fIWmMM8XJmHHZPltrfPBYplzprIwgWViIA5nm5GaczT7NnSP7o
b6wgDzG8R1OC/Dz9pefEhD4tdnaBQlA/7d9dDHQvxgRHW5PjfQmjMSm8MWyYugQ7skqORN6eqaD6
MvfKcLtde5qp7myUeAQtrvKNJbjOKruEUI83WEnnqUSbHVuXrBWVfxT+urA5jcjX1F+sx0RKPVW8
wZmf4LcUsvvZpgm7YP3N8iM/aOO9ROdoNPeFsGG81kiDFeGpcU7TDH1zHFvlK/H+jy3/WJ6baYgm
j8ONu7HuguEOZRU7NN/HH8C7R2nBYpO4NUzC1fjKIrVQHMIYBvPZCCZykRTWISAO65EC8mxPfES3
WdwIdG7BZKC8VGA7UZjpd4yp6drD/anXMZf+Zo66f40iUcw4lW9waZBcncmU3AHuDHbh84phhsyF
9T85/Ol1myTafMVwgeOJbQI+iugbr9tPL+F+jZi/E0IWf/m1474FN/OJpB2h7Gml9AkxRdCt29Qf
x+JIPgCIgNa+GvIN307RqSVHcoym7P8/9YLxIbe5lFoQuf/EkmJdsK+UYtpvAHwCoR0Y6vmFqai9
hma+CcvaflFh2yZSv3eDRKzmY0mVAZmsflgIQEY7ucr8F6BNLAirMf1prP7xv4bEO389nf+ghj8q
knqACWrYVuAa2V4w1eu6wGn3MhRFDApIaurJiFzfkHWTko2gpYqP9hUWSvfYz6HpkOkuMlYmPXfa
2l3n6De/onxa/SflsOzradwTk+aVWN7v3M/ggGhO3cWgLZWGbMGnmFYVEOag2y2V+3JuGn9jo4XV
kNTDulvWsBM5EQzbCDMA87x+oOFgXMDgcwWv/x9JjunSXo80TkA7kpKPhOSUbCFV4gFjIrYjykm7
XyAIJVpOJ2kMUZUBIcUm02SIL3s4NwomXllegfN7K5f8r9zvaPgOGYLKYquNU/5Ptu0FuxIyS8Ny
9LuzOhGiQeCiBui2fW+eYzMbd3aE4cgPyGJkoa1u1SmO14B0WnEsOwnIDT4Hpr9OnArsNivCT6uD
j5cjH4/+Mvd5Gwu8PjUnAPnarXRYnp6HtpyX0q/NidQSe8V2XY/OXnArAZMIqPBBgBSAX1I/Gbhe
EprHRkb9P1hZkx0ka2TJmRTuC63eVVeI1mrFEycS1apDA55GTVW4sjCcEVLUPksGtfP6hi6lRBvu
edzzO1XgO4EpJWpR47ClsTkwjIV+8GBml8D9qWttV3oxps4YrAq3R3JfqXOGvQ+AWISZ29WYNJ6k
gwo3sFns0a91ftkLJUU+xlrNOk/U2kjBafTWdCZLwKVVcR9Y8XCP+jj2Do8f3QCpRPd9VcH5PcjP
oZ86ScspMRkR73/gRt/rJiG+t2Zlx+RxcdrNGTynfK22Zo3Oow6rhOc9xQU3k1g3AbpDh20e1icF
YWO1/0nsSLVMArtc1Ba3ug0m3hzRFSMBiDh/bGmjyDYjkdMaM6hmM8rHsVixWzZ/0s7UiQ/tTrDC
vqqucDeZOWqu5Zi34YhejV+cdh4Gql1/C06MLLaU88ZLiUYH9YSyWWAQa2e8GhldDNhENaqVUmPF
JpV9cLbAB5TNEmmZxpCZrQFpCT27DvUEaH1PCofSry1vOohn4L1XLnbnzz257v13CUc6992iWJDA
Kg/5cfqhQiiusXt7Lag8/TWeLy+o+OAE4Nlsp1hZNOI5lanhf/dH9NmeqZFfASF3U9tLGGc3kU7K
qqGFsHLwU4d8KyeJtQEKZV17B5qvL0YKS9TAX7epsboFsPSj7IyA0mgZ+Re1W23K0//Oljq4mxKo
qifZU7WUEWGVcZlIa+5OqFSPxxrfnTcqhF5XYnz8GbOxY58RHhyW2xxKNn1OdF+LE8fa4fVkCchr
vIfoHN2Mv3t2JRfmRcIo8n1uplbT+egB5qL8qAg1rdlG+VikmKFT5pWyyHwCe7+zDQD675Iaw43J
m6LH7Y5XVajrfglvKM0jaNhwUAW7n5nkgcdqNUfKyCAasoywXSkJZjkrbLncwty1j28mPqIRzRsQ
t4NAKAwJiSd5VDlDHI1G6Ra++YITVzPhxWTQlI9uVTnuVk1wF7FHz1wN01brN3qJvmxN56IyHGE+
Jcqx1JK9SJGJqHsfKpsW+G23zp0hxKASHcH2A9YO+fojW2uklhoJi0JnnM4VqB/8PjoTV+6RkZp+
a6FIvxX6XGBDVFK0Z5fmVKyQXkKXvUTzjupzMNIniFkS1Axk14kVhYP9eOFZ8IMijD/Z4z6ffkFj
0WMFto6Xdjj0hFnn0sv/6/yRzphx2i42mkNdHg9t3UhlLkGdaLnp1GRyrnpeTihN982JZw5QhyUV
vQwqFakUeHroiHQqjMUJpBDyANcplG28yZzw5sBkuXeb6HuX/tsG7l3Onu0ZPFtbuM8SixPWWK81
yZpupGeVGWS/Do4IOI3ER5rH6J0LvOdpMCoB4ApylGkpn2UqRDSOybexmCPyr3AQIxQCauR4R+24
zjXPTL8ZXLQtiUuOLCU15vBYYW2xQfsJSy5Wok8ch7FtOB6V5aYmzmnD7mWP9fjFA2+cW/zvxwMo
fivvYBnISlvPURwZ8TgJ40RZYu6bbevoDCvDhNWaHe4bwmFk6qO+L4yTt9lIzKtHdpmJh30cywTQ
GvVKTCbNR5L9eZA5X1rQmbtDGs96Pw4LtMj3cmpRYkJrUpCGKxGl/O0PD1GwW3E8w9BU+cP9QG9D
o269gOur83W4aKjwUsWb6pD9dKXe4WXPIVeWqb+r2tW+XOwQGqV0wwiEn3y7HdPYsIV2dLva/3qh
6/x00ThwEMx+7Kdkk1qSBsBiIGUxTwod7j/EeBh9CyJHeQYbJ2eh6lUxfh/vTWH8twgsWwaBqujG
plNJd2J+a0jgqW8agg/GKs/ULqma70coZNaGthxN4598zq19mJbvyoGPpoIyaPoYmlJOk3QLfIzj
tLrjWCzKE1AkW3y/vO71paComqrGXEyCiHTvHrPMV/SFgks1H7vJ80CZBjH8H3HCtukp+qV5oDYV
BHC/SyhOfUCbVararxFwalQno5in3e+j/mvbDbP5xJFaRTvVym/jF1LQ/1nN6o4C/sMBhdDNvjGZ
diI1UuN/STOnWNyOEIa7bkYOqJ7223c8j/mqfQs1/xHLVJOxHNWrMTHdOWH6Ipw2/yN/4dwcMUY2
tLpF31MK7QOoOhNR3UhIZ76n01qOB2zAKkGsAzQgZR1zTwN2+vOsGthJNXuL8n13Ye4khATKEHwX
Ucv5hjxrkRyyTOCSwhZIeXwvO6FAJ3vhosAoVEprxRoaPQmUTVKrVc8YT9A3v+PNjKAkVyod4xuR
+uV363r1qCZ0LjD8/qM5jZBTpyE5UJ5uoFaqMgQ47RyAFmJnhD28ma+EEypcM485PzfscQpaUqcd
QDuUm1o5bXF7EagJ1+S0V8CTSs1nCpo1TcBZ7KPkrmJh9bYQx7EHnm5PftgHMzHzYT7PPsD6GDU6
h2fCBW0QgWoXZKq1MO4R6uSmK1fHCSSGOkHt3hDMEqMFOFQ6DFea7UoRg5oeeUEcuASedDL5I1Kx
CzEl+DveNE9n0gomT+KDMYbbm89f+TufuncoV6l/KKvNMyVOvDSpc4O/hBz7WLJtZIXpzu5Hrh/h
Q85T+VFN76GfZ+HYhStlHulXwK7GLok5GJixEiAgvPaeEIhibBEwYQtAjpN8TuOcfnvFPWzWjYP/
Kj9opE+xicoFpWPkaKK5tzsK0Qemoe83pz5kF5/cH5l6oWJMJCqXTLwl8JYCTj3iBIWzywi5QIwb
AxdvrYJt26EVsWsXS+AHPgjdTcXYIcT+wjg1zjT7ybl9zVaXMzMyoBCGkqKcyMU1TPi16a6w6uxJ
BlfHeyxKDY+32ivsdh+LlVEw48uUZG5Ro/iCDHgdE84wnHcqFL8USiFQ/jEuTpfbx27MS+wi9J+z
6H5O840UHpjyf11mlzzQTLGVKWuDFw/ffXs6Gzs+ZYuK297trZmpIx/PqA9j9/atLNhSVBzqpq/g
yzVz/NMfpCm+tBjX7S4VSaY2JJJJyLbQ/YwHPHnOwaJhiJS73dzgC2OZxtR1DllzjDaB5EDYAp52
Zcb+mFrPInoovSr9Orq/MjJmI+939aDd5tMsuqzL9Ynhe+z2O/GCAQ29P2Gfb4DEjkY/Lpmlw2u7
tog41I9PtXHuX4+WSBAVAVM8HSAUUZQvFLAfmc9LDy5K+NaATEcKAqEXzVsRsR2I+OYg+3LOHLXI
xBTb0710fvC0eBXz+n3ly035lUPv2CAviUW7hhKsT6jGeTz7ApRNJLqdsArqomttl1+Kjy5vgBBl
1LYRO7dePSCkULPdG2nXJo00IyxLT5OyPkwsrmX5hK85+x3neeBKAfNAz0tJ7K+9+Mj+DmRTlaM3
tLrN6D84Q6eEEUvIBw+FgotPYWuhJ9eRcyAnUxhxHY/UhV6d+9zx0P/btcnonqMSWy8KxQ7QQSCg
2XCXEvMgoZrnmXJQTd0Ja4ULWCzlQfJivOgQANdfOyC08olDkOHEQbK92fDoIRz7LV/njEapkSnh
Y8TmcS6qoFpMGmIpmJgQSXhtI2yknpGduiQ6CSserjxaLJFSlRkL4lMZPcbdyTXfs+keNEgM7/UU
2gnv8yskrcaFTsc0XQLxoW4fiTF7kwVkeuyUcvWwMyYSAeX0flBMxnjgvUGncM+HVOPItalKEwJ8
NE7QL8qVdMg8y4Fd5bQKXGYFO7Bi6pq+yuc0K5XTwtehuaootarHFl/5tVYQzVWm9Dw6yva0Ki/B
QIZZ0xgUC9PGEA/ZOys7sIJOHRrQkefe5Nf9JVn2aamU5Lj+RRpwHiMlhn/ei9T5TG9O5T0BFRWU
nVqmRc4Ow1nSuzNLcdUVYYNBiWEvWtiGgpMLj6XFhqpA2v1Ak7HpR4VT1FqO+xORCldOVhMMVXAf
epPddZNLJmEMfIU5s/yWPtqYbGTYFZW+x7VXbD4OhB+Fl7QXo8OZFcD1b2iN40naaBng3ZQ4J6ER
noA+NwfYT/jFPFBWPunYyZ9AvdosoLeSPH0xatkDUwaftMOdYP5Tq3rbChPu68CtPbvZBZ3HFvl5
DHaNBrG0bw1jCnP1iEQDRAsmZYT5Tz+Rs2/i8tfIDTEYwyF2ezunDl9mdgqh07U/oVxLjCPcxQvr
OiRWKkwZD7zIluUVWReTh88zvGyznHVwKNSs7JIIS3iSNGPX6wHahmBJuID5bS1nq8CPNbNHkCnS
IUPfrCxTtcybGxV7H3dRCmS3R0SyfakCblLXIWK6ewjaha2qJGcXvw6qA0k0Hb3hAyT5DSr1rmjX
p+4vLfAEPDwfG3bXV1viQWv9mP7FkCC/GrnalL9rj1na00eouTJBwR9R5Z33L7Axl/MBfWvYMFxp
c8UoT+GEeh/MLjm2aFeVSrpdHJjkJoMaNEGFdv7FNRw4PWp8JaqSprWnUuWR5opmUijagZwPXGNG
GQtbIxP4dVvpmHu8giuobPTFniPdrhfZD6DgTIRpLcedTZb5se++H+1lplrXWIT+npqnb6tUuuk/
R0dEmmPW39XreGAmZ+fVR4Lkr2JWXTqVkiM5l3zTfPp345Q1Xyco9qNHWsB9D8d5juEG6BjyemVL
t1Cx4oOynh75P0AsNGHu40Y9GJtWihYLxmxfh2Z5WJlNEL+YzsqZR4jCASaWXSP4+qX3gGNCrPqS
G4SajxbxvPu0yZBOWVL105x1ZWleHHYoX+spexUW0UXL9/7olYcjkjYf1ZhVXFTV1n62RKi8SBsF
3QwBEkvW6rlFhyqm9qP9tAjN/Amjp8SSXbRWe47YJnZ5tftTSmnqGQrhodSQCslwujvxykmJQ9CE
ihsYrIRZcfDBJ6NaPy8UqhAVqcoj5sHpxF3NXeNgsNwxP6pxkuD3RhN7SWyWw/We1bYZUmbFKaVJ
OUL6lVbET9CicBpVuejIoRip+70155+gE03io7O30DyLsCLuOMsFP8QKwRQ6J07W94iTGqNYGKBf
S5VmnIWMEvfMTrkKnvgRh+Nu5gFYMAkXYjH6G+WWapSbLUMejtCkrxnQdoeEynBg1reiQ7CMTrHU
RtLQbEvtpl5BWWJ7ggWz/8xQ3CUWeNG9+2jQPoEG81eFnGxbWL3yHLhH5HSAcLPCVxk0ZRJBcGo8
2URvfjcsrqO0hOqpsEhQKNCSxmm9funP1qK4kJFCTckfoqk22rRwXdD1NisOKwgcKM+9sTCspGei
2ME2zcmJJSktLsqvy7jGYRD7sVVZJopvfRJJc9ufAw2hsFdzOjjSJyBz9k5rfT8JAru0Mnh86+ML
uhMEXQI2Qp1DCbqqWmRSaSWf98njM6MF0CVxexyOWBYOrbthM46U4LzKPKiTSqRVH4q68Hf8BAgi
wYH2tOzm/+I/jAl4joMFs0+aZWD9gYcEUDeD6hVqVBD0g4DjGpvFVoZcSsgksDTjjnMKj4Ab+VM2
csUwpJ29PQDavlBcVge3tp2WiNnBaGYzia129umBitOXRBK51PfJdrVca/e7zwmi664wYbmiEq1f
oBp39aIZ4ZF2nrku92X65z0iDz+J8ppDfFW6a2dt7KeWYIFsurHyR8vQzIGrMtUVrQn35/qFu+zg
gNleey/w3kXUxi/rpD6H6F/9rcVgVJaVj7BDzuWenu2/hzQ51/mZoHevBqk0tg8HRH52ofXc2Abq
RQtYf19/I6JQOEjII/UnZn1H4PIKpD6xoH7L8xyvQgYjFe2P9I+93Qh8tZgd0GfNX4pR0CUzbz7f
qYMNeQod9ieRnEyoS5pFY2Ambb5W4cpFdRX38lWS4Dt85D5eQ1M6FnlxeRI845LATn2VDEnvSm46
zMyJSs3U6kV+lH+bYaxPk/N9kdRpZazUQUr7tH73NI8tVFBd6F7ngS+EvUqmrR84m/uw779AQW3S
bTg5R+mJvvgctwNpbJ64BpEQtoQzYoKaYj+Bel0f6AKJOR12tGqTcYB/ltv/lpzy+wWo5dDYRnzL
dQbhcy0P1ZVHQKdQ734VJeeOmwu+N0PI8FuDKDGUIUoZPSmKoO/gzls6ce5avEs/7cox1mPmFjQ+
Tb3vO62yZOSYYPExu1zIClyGJb3LTY7fX4VuXrW59VYzIJCqEOEVWOsPBIubw7t+gu+m2T97uQvX
tIY1Knb1Yk9g8XUoHeWEXa8sqBmL5IROzUjBHVIjQiAdzSWjb+1tm2+WJJj25WKS3Tn/1WFzIwu7
W6GXlyoa4T9mrq6xKj9VHa3n+XuD7MJCNPPUMhgyiiXvvjgiKCCSKQw259WiINoqxbmUje28iacM
3MxA5nsB1EPor0qx+9ishOiayNl2Kr5yytUZPY0fRNGuMaQxIv51/zXzPyPKq0TAcZinJoTkqso4
tvyC2eCfIO0t/DYVBE1eLUORmIxd+esy56PsJJwijG0JgVBB48hxOvOEs8fbcRwmjkAPIty4xTrH
nNZAKzPlKFhXTyphJCJ8BgrAmFSVBSRDH49hloC36WRRPpi1cKg2JMAKlh/n41cdmxkq9tH8xPzb
65oxVCa93rgHd35VxYbcJJ5xwmDE3TrtdUpo56CnbyEj6GtI5d1N8rTNQvW7iGPTqxYMT1NnyJIl
ulqpsVKqcPL+zmjN9T41KpZm9yXzpXhGX+Y6K6FtErAtQosChBlXMXxapvaLU7gRrm4+a/Xu9wV1
Z0uZLuAqR9RvumIQwZNIj9evHEDLnU68zSwutxsVqyiizQjWSz1Lx3He67BGhbmafsNoBe/CiMDY
C6OUncm4LbYfr8O8dS/89YJRp3ocw2oJWvrPBgxkf0B6CiQXWaBgVyhrq8gySEp0cBW1r0TtBabK
D+dWEtr6bQZ9zc1bHppWmHW4yYKvKaTKMtZCsafr7ORaZAHOh6EKSFg+sqXdBIW553NTIePvs1jV
rMSVoxh5lJRH8TbyjQy3offSREH6mg5eotB+aukiNxs/1BILTAWqxjkjvx0yiOXRp6BpdPy6XQbr
ELDMQsCnqkGGWJpJBZgNeXDG9zznQPkhCxb3oe+cToL2E1aNs2Z1R3GVtdYC6Xq21DYXrqpeZCU1
ZjIYm+ixUCAKRiAQ0pC1cvhntl/5KmUSlmLMbCjcX2B+YnaOeMtmzwc8IcP1srq0k78jZB+qvst9
2Cb+lsR1Q519x70qeFuY19Xav9cWXgHPvh6pzJwG4021u48pouWMoBhKaXVjgn3D/Wu/isJobrXP
rOYZUszJy7u6aTMuLZXtQLJ3NM9rORyv0wdMX2nOV+2kHX7HVO18p735nIwrUTMJP0SEYAbd+YVv
LgqC2rvhmX7QGe8TAGouwywg4SGNzRjl2PUQBwW4VMO+onbpWmk8POSu5nKhDZ+NkIOygQ4EJd6G
S8uZ27IUE2tMxFqFeeGOxmLvMFsFNqGo6ccvIpFgCLg1fWY9feAXv/Y1YR/8ribbHx412/BLVP2W
aJF4wsuwp6ehrIt9Rpe6PlvV0TQ22knXP7YUVsT1SMri3RSGvcgaahFCWgXmO+AHtxHSBhhYDr1i
s3adAcp41+/co2jp52xWEzj3PGyF8uaphd4Bz+qpxOcmuEVS816cHW04dtieEay1hufAv3Jy3lxT
1ngUR+w+Vy3Nc9q+VbIX47h0NqMmYKYIEHQaaWaDPzN+2rP9qzdKt90JNHw27McTVjMpSb3363Ph
z1sb2qeO/6m7Ed3PHa13FzURJeqLcf0G+RUkNUOd0wkU5Y+giKS8QEb4f6+5BRFQq807Qb9JTmFP
jd78EP8fb+i5KM8t7nRLFEt5HKB5o37QyXklzD0YQYq0VIuHWpGZavbfC63b+WdBpm3nOieFkm/d
ztivXpKdQk86vtHW1T3uLVzJiwopcd5vfV/gsRBDOPao8Bc4utQZIHHbg0Ab05Cyc03uhMVLoBrf
Cyagpvi76hGEpP8TGDY0+FmYb2C+2ArArg2pjtO3H9yJcZoU5uW15bbBnfEeNLkbAstKixxVxB4m
iCiqv+K/EsASqWm0eECkSuIN5FH5RrTl/ZDT5vcv9E7yB5GUfQfSR9R1ag8saZ1WF6N3J5Hk7Pri
SHfyWqnqQeK46vTKT1lagA1/mTZNIiZzOVpPj6YB7NZE+lcMbxUQ7vp799AGgMTiuGugYWUp62E/
aBkK/JmCchmnq/dcXUb7H47cPQFH/pqxk1AA2uL5AGPPGib8MbHWn93nBhsF+0pKLNvK2JMn9pLL
jmNx/0hbixgxhIcu0Tj43E70l3a8+csOe+gpcROSoE5UgSOWa1THtiQ1hPUTOkPNPWt+TSAj6gr9
EVInzxRbGLr8DEJkmfHP27AjC8jcINWzZyddaxxDjvKcnC8U59QyIajXYYCFivMtR8lreBd1NYmb
l9gP23pAOKZfBvm12ufPLOFDeUPqDgWPRWsID6+SGDVtvd4/LQopVynThZz4Q1A71QZXjhhAk2zE
hBLud3dxd++0Vbd9UwI1iktVv61fkEaT5BMLlv8i1XbHgWvIhZipk1qvDbyUBmj3Y3UoU4uGLv+y
DSbOIjSinhBDPE+ihzmyK9HnWvsc9KDwmAJBHU/3gUKV8b1EFhl0IHhtUQtKxp6h19vQ6BB2iFBj
aCYxMTVqQ/zbontgFmJdKZn+Zz6bQPanaN8FHueHDhgFjrlDr9Fvdnv7+G4YlcduGgX5eWRZ9A8k
69t/Lz/85njj/Em4uArT+f6rLfQPVsUeRis73u+NaByU6t6mkXdP6MawWAtTXXJVGHoy1H7J8OMR
dC+rD5lwnsSY+HyrM+PZ3srK2kBKuWpowoe5GnnFYQxBz9itF2TLwt9DRNLaWNt8RbMUVka/WVK5
6zMXW+SOMi+UNnThKm73++q5o4sJNdBwCtVN5RMvPYxPe1UKlRkQDRkfjiT3EFSr3ZibWvZh5Bvl
QrJTPFA9LY/CBIUkh6EpNfSpl0REkOWAJiGxdhHuO6MFc+CF4hmD6NBDJgHPUvrnxiBnyHrFmtGz
rxmjSSOXP/Nv/6r4PvE1JW8q1QzpnXihGZ0rNfFt1EKtTUIzY8qlJkISulzppiv1g6rN+LTKUYzq
ySLJDKvUersGTwlXwFXUiTHbw5yoZVJo5LeEUvy4xuVa9Wbv0pzWRszwmhk4p2gzkavQSOrvUw16
2i2W7kTqzoWP3OStGdC3SsdtUbEksK3rqe502+MosVb+SdDfR69HXeSRcWOnS4MqB1ublC21IsoO
XvsVtR96yf+JZNBMK7PYFcKecwMdvensQs4H5x7luPV3J/R2KQsQIQBX+2BGaZLey1fN+pj73/D4
Ncqgw8jjy9yWmRLy5BWRMrCjzJSsW/9yQPlPqKSilgcJJB6DFz2iWQIpsSV0/RMIjTEMPriEmm4R
gjnli/6/2Vlkbbg09yQLOqQoPMNtzz7DB2dVbXXDgxEU8MyBhvV0NCKDoeLf3qquKzarWBuJiD4y
wYfe1KTtfV1da0/b2ztC+30Z6CeU1bl4etiFU/EKvGk7Et/SuqobjyVzF1qyM0EKCtcw3M4GFkf7
mtkCpFl5eHwxOO57g9RGbp0oUB9ibeTv0JxbGxNSojOkYZW0EkcrbDPEBbEPZfRw5GWeOpQRTlJO
2hUYFQ5M8OvFBP29/HE4slzIfPKWxbuAK+NgOOno72M9GHi8QGxRXhfBCcrJZQJUqWn0i5w1Y0ry
z9aQBU15NVURP1JBB98kfDHXmlSLHk8WFIuaawyUOfNxthL0PoSThyCAE4X8kP2Z3Z6aSrrIjU96
ZYfqGHdQre1MfrFmfmTl6T2MF9wh/PO2OQcPnfV0NL6uphxUGG7UA1dWFpzBdRf2upJIDv3PlhFC
QlcXi7Z9jurxsvOSPUTT+sTNlkpI3nkeRAfo1cSb15xlUGFfAUI4Vr+uLq02SVGN362OkP2V54LE
/E8+7/jp09DlLMwz7tEqzPGJAn9Y3ng7Yuhaiz7DZzS2N/bRO23KY52Z1OWNkEjQz+/i1MVtg1Nd
5po3cKVt2e3FfG/BH4eEwl5/6ItMfBtvN9LQspSrnxOc72IMfhjH35I3XdkXLP5Ap9kuI875DH7j
xtABeSfn4EKQwPJseq0tlHLNyz1U+PbbK88X2OPEnEvnT9iSWy76FO1Fjf78mFB1HQHVtfpEWk8G
hrhvu53ZqdyPt5MF/h3IocRGZS/09JzquRg6k3Xw6K+bLCWyQySSVqfrdmuQ/Az9f4zSv4EXt25b
7xEDX05CfHwWzhUiYi22MiLcSubtV1SpFjU7ej3ZHFt8GnF2Y5r95QTpC1EVJQXSgdZOzC+hc0fc
EARkjrCUkvZqgU2t9fR+mJaCz1XT6FHRJz8xZXLNgNmrtchX85AbjDc/RhRAvF2lL7ZZM3jo7SWs
Krcm0WAT9xCn+SGeaBp5+W0C874bdvres86eYVezuwRoRkrdyJZ0XugYFkSaZPgNOmK4xOk15Nrw
LPFwIrYo4N8ScXFTOeyav6QoiftkLAivwCjYoxEm8Q1dSgzw+WTAdo6eDeCKYK+LWoYsPCZBEFBx
3uN427ikWEWhFHIIsCBNLwAbvsRPOgvx4wXbieKIzwXElwbiBqlaa9i7v2yWCY3UqDZMgv46UE9P
zWkvGeeVT1UY4ABGJ8OYwsQkyjaRDA9hkNc2qf8kHwvnIfUUCcLRvFMxrWmhBKGkQa1UwoaXyoRx
NamSD7lt5WEL87PPDzUJ0mGm+aRWshZIXZrQIoMKlfj+EqpW0l0dvn6zcpkUHqeG3lv1Kk+OZHt9
zKlZojOHYUAdheNrgNEsC8zHCF0ijUb3Yr3vMxXcrvuHRHZpTydDd9GjmQglTn2nLdR9xuEKYJIt
E/Suu5UNbib4LnqUGF5cGa0R84zTiQaP6xs4vciTvV0FPLeXR9WGDiZFGoPlrVs3BBHHUQh+6kjM
+aic0rMGsooEum2tH+w/kPGen4H3dGs3OXwP24UUFw1CUKilPYFxMW74eB8FU8PL8ThR2y+JPRje
li3jlAHZz73LkgiEjvojV37Ce/T6IkZa5UtBAH+Thvh211w/ZOeVE0JlX5/BAXD6PAF7G0q32N56
K343xZg1hL2FqtLlZZ4ZX06494me2XtGeWsFvrla+gyp8vi1wiSA62TCwISfe7pTvNVntinwkU0r
GcikFs6Atd9e+Z/Vfb6bk9qKEbUAv7pScH6TRzTumYgoPmnLmchxCP9FcxWR5fQCJi0HCDjx6uKj
m6XYfLDFQqUI/RaCG+HU2dP5385Th82XbN2huhoW3ofUb3TCDtUezYSYxo4rGGjwyruUc0aVJ3BC
ai6jdV4sQeS+Xu84+6pQ5CyFSXW8BPrWNCDLmST2IcGtWx4Fmg1mNP5xszS3DZRBfH99mYMbKucj
Tib+tw1YZ2f9KaQHdfq3ClN3Wdp1GLaPrUxAD+Fn1BNngCCSR5n0AwpK2IeBV9eEEZLoa7U0Uo3q
zn+r8uoi0o0ozQceT/vAZjnrIZP/LPk69biC9QpkLg3Q3KfOfPPvLpwMEKB9yzc/PH5hcQGA/eaF
lwK3nmNsL28jPslvrn5wqLAExGzGRBr56otvHeZl4irKpngsVXfUni4bngCIh+ax0IHJryMdPiGs
dttz8Hc3de3fZcMO8YxhMOCqr0yBmaeDR0xxQGcRV14Blu4UTh3paeQWePdQj/U3S/qOFrRXxeqE
qHOSL9zXBobqqrDQ3ppsCGmCNSsXrAnEPZv1oTtfUeMPzqknQ29BDkcUoHyzFbjqKe/EQdUDoVcA
yhKVSgoj0qniSSZyP5AGkj2fIwmReV7BsR6wGv8OvOQQpy+MoXdUag/mOku/RTlc8qm6/PCXhz+p
pPT2igj5PUuUYuzwPxsGpJtgcw3ocqN/dtBkCO+hPywhWMQNW51AARWxlj/guv22cl0e8weIK1RG
mqCLW+DV9c8dONtZ1dhxIxQP96yDhpdJMvkQTZfXMRt8LngSB/+v5+lYLwh2hwSimGgZJVAv4DMg
ajEGG3fEtBJzpNAUYTD4y8LdS8jGTQk30AV6zaInSQAnG/58fscJOLVGNj0P8ShChHr3jZvhsL5J
C1LosQVyJUfuzpIB9iwulfpDj4y/rYXmsV8ooe9y7Fqhewsvjnbzp05gARQ6X/RP78a6n7sLrR8+
70K1wWTlYzL00Ypw3yYXAmdR93324bxDGYIZr+OYZ6P5p2yGXdzuSZwcOzCAjS3141BQcl5m4K51
7pbCa7mgg7f9bPq1cFGgKOBKLeFBZx/KnOwQ/JS/ynytJ6pOw5OkHQ5s2DbHjUxUn06rYOclxFmP
89yz0Hi7iC6834PBTX+96kpRp93TpSo+CV2AAHYpbYc3fHrllBl/uiRXFSOAVZIUiBf3rlfR/kD3
0HY3sZIKHO7rFTWMf3T1F1NNC1CIzu71VbJEH4R5zlDYSRBHgqpW9v148hR0YKnIYWkfQHWXcS+N
Xg7BPk2nG7Fee3T6djqYHwdrceUGpnFC/p6nBxzuxC1shk8ds9U0qNDKR/Ig4AEshGDqM9frqaTQ
hM35gVcpDcy/BCNvAaeAnhswTCxKxxSq6zJCVfuaaU/JgJwv2rj8SnaWErkvNCeH2QZBVJDvvv6c
8zWnKwi8kZT+CefeZ3zbe7jlO48CMRnaIAHqASG0dBR24f8gN5+vv0DgpComqXVp94+tNCNdxgcr
GDIejwUMfjHJYMrCHakDUobH4oUIEIYsry8S666BtrpV1iWU930xi+qxcCGHSo3IPmgyBCsFFkKl
Es2Saqnkq/ypeGx7V+5IDrS79jO86nwlaIDZGsZ0CiUzy5hNDHkcBjRzIx1W5/gwxhm0dxYU50Pg
PwX+KhpX6n4UvtJB/H9yLLOpafhNoe6j1ysRgQjYDNi9J7f6z8UUgaEH+Ql5iu71hVNwO7Nsauks
BgjIWCn9aHMQg4wylJufYNoN21Z6CN2+F3/Bh0WH5EeF1/v9kWq1ii5TZARJSgta7q66scuEZP8o
PlJom+C9etl7b1AbSmAyKQJfGObc5R7PWtx20TsjE9e24NY10WilWPZzmjI9YsyQ6eBn0U3t1Anh
AHPxTMajYy8mRQDHo1F4/MiaQ8Pp5sB3ZQ/7c+qf9YO2AG/YJhY80DNch7wEYDqjQNwLzAidhtTH
InisYKUFSZDvLTAmJRDsJG8X2aABu+9XQTsF8GwW8Womsl1XKPfRdzjQwZcNSS0nC+EyILFNyuNF
0B5TTz8XyhOOVDN27Y+XdPmcwNXvtf9tmxymHBKOtA/FjnmZ8aDGgGgYzKtzhC4mPvZ/GG+96fD9
qSxezV9fsT9VtVQxpxFMxyDW5MW5Xp6eP5WwfD7T2ftm0JWncJIbkfcyuKALQT9d7DbvrRektM+n
H+5KVcKkbtzkZiZ1e2F0VYxrYpMmncKahWvXZXl7zlvHrrbsgjmfdOx0gS7/VrVbs85vTMLvSx3p
x0wPxAp5GDxbp2jCiyBkAA6t4nKtSiky8VDZWxBqPtrgGWI7SMqhzqBTLwWIKjxP4fENl7ammmjQ
ghqSVxsfyuNamVFi/5ITgCQObK+o7DGcLAACECMurUn2xcHz4aUHb9nC5FfqAgyMZa5iOUQuLxmN
tvOPrq76ADq+WogWvgk36G1IC4f7AcRZ3UjxqQAyfR9CPVpwq7vkQlrzfoMRabp3CkAi6enD8XQY
4da2lK0wxUOgwwMTh2I5BpLhl58TcwHdSF9fOLxgzVJckkMKTDHVcabDmjFgOmIgTM7KDXne9pJS
XM2uF1T+Yw/s3OguBrr49+J/w9koKXrgmDBiV8p78g3DUDpItmzUjqII7Im4R1BQKNGzef4kxqEp
rXpRbYmKp+Uz32H603jB0IZdwrpxC14YNC5lrPjzg61jeG7hsNHfXJ4ifb70ztlPrHUU7Eqi8PZ7
C/SsLblN8+LONzQEoUqr81Y8PgsVco3qYwoNiexSi9tFbrB7Nuk8JiZLqhyLgfPxYoAV+XM3T/zX
gY5DktePy/SjcdIzmvFJ4vA72Y7epmGj73nX4ZPO5QIUMAidV5r/9ixSmywszGRGJUnewYcjsrkp
cOPj5P12GzRftaCG/eATkioFmG93Us3ULybURWCIsN8nzRJvDyOCZuY7gMlqfTwul7ezcruVGlQb
X1e+Ox7x52HZbsh6ApmTzeRBuV2tpOy4/J/t1hICsHrNWTig6iJi/BQL8IgCe49dVOxhvlsA0tdS
SgSBCSpgysH2yTIbJXEWkxNdnf6mPh9pEqMFGhmna2vaEdO6w35krM5KXa7eP1FBtfHvv2F2z7lZ
FwmvA+5x+iZLaVwYA4axfBQ3jenJFtfWPoa4SCvXFp3K2AqsAstRhrTwyIcxls1AIXqazOoTSoh/
76qIWNSqIwaR7LyFZdJ4X8QW20qAKwNDh6zPZ5PuVmRkeA4zizroETU24s5qtnyQCWueEob641Dh
vQG9jgHYBCGGWJJWiJhNVaDypMh39HpcIWIMSVCpjTWPjbyfI1VJVIFvLWxOPyeTnihKydOb17r5
3hPNhhDv/1iMa+KrUM72H1cF98DecoQUt+kV7Tx27UYWmWrZpaSgJgqH+vR12OHNmBWsVXl+SYyo
be/HxiHBfWJMSR3nIBYZLyJSj3ZpPNmYZ/Z1/mv/FOs8H0Q4Kl3GTVgquaP9nmfvH5iNeJAjV5sr
FbNbAYadWrZ2ndrRAeHTR3uzncEsnbNt76DbTtMWWYdkckDT2bpChIWeV0CES8nFBfObVFZjZv6t
UWJaro9VQpPKni1r3mTV+QwiV3v4EqMq0CovBLTaFrS16gEwUvLbTeIHM9dnoqe9TWFnnaFpk/zt
C8ge/0SHBeo/YT/KxQtQ05NcdljZ6H1PIA6mIlhFuoAaxesaVbHo3QnGi6LC4RtV6dfO+TkIysfZ
AbK3PysfKH6GFMC1otFYmp8AUTAlzFlW3ESnD56mKE9GRKj6s6+pIZGzXdZFJPZN1l+vAp9ygx16
yP08OKTh59CYsOOrYT1lc7dM9OGLEAjUyzXADyMCw0K4MQJWuYJR3YjDwfYz36e9hWjGKj6OprGB
M14aMZNxYjqfbj1aeEuZYYz+MxXrKAv2cAW82ANOyhCtOAfPP5I3Svi5qLY4WzOpM1BHe2Ke/Di7
UHBi6ZtaWkgHE9VZ3mkbdomoPAYiTyk+AF7Z6Oh3r+K9FfjJoo69i1K3aMKqii43zbmy+bXEU/qc
mXLOZJo8+IsWGGVHVW4AUAXGyR7JNz6XC4ww9i0DJ5rWUEabg3n8jk3BDYXYUFCZc3THAM5hZzJk
orCcy9jNYqWQ1GQEeQr+2YARyvdymxMOUhkO5y0os1y+wiVgFoVz1PU3F/k/c+nwb6yUSg6J+sx+
rp43Vw3KhkgZWPdqFDdptFQe7O6a13gEmDzZRrxFacgxoVL4oV4tHQBmaklw5f6B9Yr8aeO+d+K+
UbUTx/SCrE3rtjSuK4KIZaR5fde97Lq9teXMw8aW2y6N1/MXVzOD1mHtDa5XJKpmlo6wGPZtnQtX
AsjOdsFkBfThF6bzk4EwKN6sNYMDAkqBqlzumBvBz3t5L/wYRucshrz746Qgmb+jlp8SKmUN+48J
xVFsDOznme+ML4mIHz7DetK7w4vF/H71gxlOPjBz897O2Wd1i7teJUFUtY9XTelRaJ2Bs0+JBIA0
xOCm7FTh2aw+kD2GDC3HQ/d74HVv+j+BP8sbdE5eFBPVeMZObzr9lQKsIyCglzWlM8oo42PchQ+a
oFOeCGPMSd83DDkmDGm4R3WIlAuiJIXtk8ZKaPtt022DSK5FllRBa7G7P+G1zuDqnipnCIdU7VbU
G/y/hBcotpLNUi8zEsg2n6uLBXNATq5DsJ1PcsCHd619zHj6rRyZuO2K5bWAyKMoLFf75MOVBmsn
tx+nLn0zrJ4raRlfiJJNm7ne/2izbls2EB9QToRQpuLG2vUpj4XqjLwjLyooL0AD/W/iPP5XFYc9
8oBtSOAwUERWLhnHL86J353SNlPgIchXhg2bCzrllEJD4uhdc2kSLZTu/b+6ShyjQlpDDsB8poQ1
04zEWg26jMno8jKvp8cQ4QcZZU7sLvAQ4a8ImvE2h4mGphT/ZMhN2u1/+DXEX00BakT+gQCbDZWY
g/e4Y1wf+pvFWOScRSchkSgAJIi48wmwDB5+bTZOJm+jk+mdtO/0AXvZHUgPmEoMJ9lW7lQJtg3b
tjSJpp3ZkZvaHIncJ8rwyn6yU3GcpgskXuhTmBLLbu1Bd0NrQCwTG0ElQiruT2jj9AlmZchfnY9R
meeac2iNmvL4L/2YneeEmanq2BUTI+wVwvttnbWzEyHyAU6vtBxrSGo1QQ7L4Dmr1nkkDH0nOlcQ
A5d1LcmSf97YVRWRzdyOLXHQGM7bf17xgtSCB3TeX0cWUWmkNmMdppI7/gkVp8tFlY0VA06hMh18
MKq6meTTF0kRRsiR+deA7UCkqbK3X5NCgVRlGW1Wfc1Bdh1iKYQIpXnHIqlsXUhNsd3u9Y/VMeFT
/xGpKGHze7Lj6UBm1di9RLj5S2Kl5FzVsdwIcg6LBirY/n+ZHVzJko5UZMyEWpHwnEa9bLQYV/Cx
yKcn4ExlUTDaGWDgAlRjrQK6BaHy2EtW2KRmvUOj6Vy8lMYguR+WH7PPaKS3Poe8ZqICAzuIVF2t
Qe1G1VibYNu2HyvosXYLYO1TJYc470ZDlyrSJJoi+0G7eDCHM7OD3PTHYHnYAsNAk8/G8oseTCfj
KkmhbyJcWSqzsyII2PTypPbdwbhAxyov+IMj8w5q16y2LWFxwTX52utrIlWcy2lJXuoV172TcbAH
3ZCt+wwC1ICtsZBqhwTJpOMX81pVo7p3q7/QP7uMIqmQZN87uloYOsPWYIlKQC4Goi41+KMdeyTC
34olTIzsTWN6plmfRT58yn0gCw+MqitaUZjGNQiDa9cOSqyh6dIgUPTRQLn4gtau/HatEGeTyXKV
0DNxL77+Hi9VBRsr/ehHMPJd94pJ3vi0IchPtv3YvAR0E5no1uAku+6lpXVXcuwS9DoFvZM3SrYz
9aqqhR6MimKvFzD7/0/ndhI7TsVse0Nz/nmYK4eBOGGSRFRHQut0ycDZek4VtFZ0s76lRsShH7FF
Uc6kkULPlrIpMg5XyMD2y24tuUCAYJQnDg7CIznbWGcsIQVUKIfJABLjXWuIrnMxgyiK2V0xf+rs
Kqn1/PQZMphYejwjs75zu7DgUO3Gv+wmu1V3cy6Xffnp93faPo5oCnitmU2S4amCI9lA/dp/s4c8
KDcaHjr/6AoH3tow198Zb0aHyPf1o+rn77G4IdVVd5vuSBTyGdqh3O2fl69dTEEdoBmuStzyHDl+
R87lOpJGAvFTpt40RqeDKhYnSh7T0njFaQc5iim59VtyOc4zogaHpewju9BBvTmEKqdGeKLYHrUH
mi9ffDHWobCso4w2QJmDrlEN/bJfXH0qYEtFQ4l6DL/BwNxU1Ysg33XpApqeiiUD/3qo6CI73i2M
wJgqgEmDReslrqW2OV+g12BujwnyB2nb0teLZlJKMyBeE/w3JMykxHjpOT9AwMQjXZpvnbOxGn6D
v7xdSAAXOXjBgXvLipe8MFUSX/S0DDDNM28+Zqeenj9KPeZBTomO+iHqe2ZrLxz5uAaVdwtN1gjN
9zz1rFhg6XBDRVn9j07rv6Ep0BeebVkK585E8nkJ1uQfEeMPb9ZhsWMdOSK9jKyWBSxHIVIC5//n
w52BeW3gOQ+4gS2gw5ZUV1T1bjAm0ycbvlrBtD/9s6M8WHZ9VNYOZHgxCl7bn0DKZq1jae8fr4b7
Ax4K6yMyC7sJP1KyVXWmV+G2gZRg8xBaOr/F9zgbO9e8E2arRIvMdJi1yvGwqE/rXvwq8r2nKzX6
HYBykEaqTzpf1YQ9/rGEHhZByi73ekJAC+ePKBoJSVL9CNNzM450PPgCb7lo/WqVKlZDQOHVLKXQ
xMeO0AKDqXz0o67pqukiCnMxl5/LElP9yuhynjT2kzq02muXIbMz6dSgFlZDHeVFTehiQnKTr9Y3
IOS6HAfISQvcruzPjHJv4+pdKMtzWfBdrl2nAgJ7VuXYHwRjk5j1/PyoN4cW3xQ265RnaVFSBMzx
NsdfI2ZqYo8cEM0E9816aEXbBC3WxNlEGUwrjtI+xCcWihcXC8eICMzX0eFmsV8moc0NYqTM4AFt
X26ddtokUilCfCWTiyBo6kTg/r0QfGyCp4MYEvR2p9vbTqU5bLt3L5Dl/o+4cTC2ODO4aYNaBw5R
CrN2XnMJO/vE6hAVyTXjFKpeoGyEpjvAZmva/CLYziuKd8CkxveJAEv5eYOhcIBvejbX3Yj2QyG3
Q5x1/N0pbq/W88Vqsi22XnnedRUNA4tWqOWruxdFPXGWNQz8IJV/CKJObDLIvsLR/mHdOUXzvaVH
g6CRl7Q443w1ElaH0/pAOcNTObwxNUc5qU8KKTFeliHr70V0kRYT6Tefy82O7kuqVuYPb6JLfgwf
NyK9f8OHufFhdotB62BVW3MvOdzpCd2vaxzVvmG5zDhBzNfiYq+RDBY7Z1hXHFN7E+UcDuZFBxwK
HIa+7tg6oZgwrZYMZE6b593lKU+PDJ5Wa78lO1XqIjklKWL8+yQXhyFFA2Bl1XVdAiMVpKD6h3zL
4tqt1KFykoMbHZs8PhQppqyGcJ0rzw2BYDzpU48GA8M654wE9pqpx5P3f5/d7cK75ViTzCneIXR1
ROfAkRIhlSEunmYgXeW3dVNQzHVfSa31eqRSd8fl3AjsOmHOc6Z98TR69i0DuqwnyzLnElgeU5ue
f6zZe4p6NR8V5uMjlOwm+OpnxgP635LISmSljzaeYAHOYwLqO1XjPXKYZ+rq4WEhxK3SPkdFDJCF
3R8iqwo3bhbXjalqUqCmfdfUNJI9GrlnMLBewPes8EhfHOvJHEaEpkkXKgoAFLPmy0XCWaJ4hzmW
T7gh/PywqDwKbQDM9Yn0IoGoXYXpoQAEZw8Z2IDgphuoB8/gkXGXzbnPJwaN8JSnd/6ejSLWSXkx
lEx755xrj7va3zcmMhP3G9/2MPs65O+hdflw9ZeP9U4Df1yDYe3DdcCHeOb/yyAcUkuHq2W+bdEp
98Vtx7yH4MdjIQ/p7+Uj76VQN1rkdmhaWWWnx7g6ydCKbJSLCdiPLwr9dBbMLBBpnxDE5ExWLBqb
9XFxdvBPcMwtG7LY39tbWpg5Y9/0sD94WTilQHY1uYfldxyOprWDhhomhEAxanryStjAUNXr+mg9
W1+SQMDsHDr9Oc7SwFJVK4+x5Z8aTKCKPW/8SqmBunxxHGU/A245l4q18AGK5wNZPEk30oq48D3F
3SRLSkwcMFRlJWZG55iQHxlhV5FOCQCNt+/tW/qjJihI22GYakj+a32bQ+wI8SQsq6HwegUDnpcb
fsRm89HigeBytUS/lMLzwUNjypnv3yXr6oM6U39GouVPbfro+xDBbbfnnH7B6YsUA8EVtBd3tBA9
vRwiQZYCoSi90+JE4uN595uPthFnObdExJKnceLUdGyF7Gn/3ZXoK/g0T2qGTuNHHwkqT+awH6oY
8XyRnIMbQQP+sgnvx0L5/DYXf2UvlgnGcOd4JSORx0FltFAhinv4u7FnPmyswDA8B3TdsMIqPHLV
XWOAfVKbDBX6CV6cJo+1NeImlrDiiM05AWooyE6BK9foRulYbc66BJ3orQHtx+xgCBv/lN5F+EHF
PhljhwzUP1sPYoXEaWjcHy/GRk8PFyn1j2caWfSaCVbqBhU5jOijYsUuRsq7zohNu47XzAvhba1D
JYkNMXi2IogAml5fYJhicc5EDXzFvgIzcOP1Oczf6FFFLL8U+76uv3RTT17N+NHURbEU8J6Iul9n
RDgE5ExOjjAxp/nYVRZO50jyaoUN5Nvi9+MAHkLb/DyuKGlvzEz3pNUINjN39H42OOwOgNvuBMVg
O++UjqnbHe89jOTAiAXYZqbGJ/5jt997K4qvvwtK87pIPzMHKQzDDhv0ouN/RbkylDzFxOBcl9h9
wcitBkrffqjSnliogO8JuS4Z8v+o9GZpuo18KqxeIvljJTRH0+43f4hOeGvTfyu15vEPPsAlHqsz
8mNLRMeVnoJ9qfTo+qYgmNdcgHGRWcnQSv3sGnbxYxZIj+0ONf5m4vHPs0w35RlczdwnbNYGgqZC
wAxPpIcXu0uIqD5WZCeVgfvPW0Z2I6q2eqemrAGJ2ab1dmMcaVRtSOH6QPzLWTQ3gwItaJdVvCYD
ITYCHpgu48cr5yNZxEEQKrec0QJheMzKKVrJCFxxCC859BifVwDcHs87M5DzcSd9ONnyg2eyyFB6
aAqFFTfNOgrn5TMSaMsmBH0G3stPa28XZ3S4AyYr5suG5qw6lhJMij2yYsGGXraD40U8Ouy9iSkK
21yz3OBvGiv1sOH2t7cQ2e6fWgZ6dDPiszQc91lpNf1wo/jPRW7hsYkvcy5gm3/uXJwM4KRAkAMh
M+H5TbeZxVuz6f3VCkyZu5uR2ZCmefhXEX9yHedoEKrQWcS/gnd44AkYXr0Dhg1xqT+G5whnFKVJ
gKtl4duSqY6OwGzkIPCDbhJTWkyX1KhF/eS14lOuproGbQeW+BVy+Jw6rKkBI5atXmC60QRFt3/l
4BT+UQ6nCmBy4FyJYpRO5AYNUl8JjuTaQXHd5hixxzsfZvHLTbOKYQIpT6W464S9GfgpR0c32wt+
BL9UEl4wEtCtFVovxReGmRRiVlPcQrAIdHgCvf7WsKZULpDG3Ftga4IW+4X4NlHy0rnp2iQlxaAl
fbtKShyYSOf96sVUmzGwQUpQoEHFc8eT9rIgAA+THI2RfYdjHIJ4DggrmqkJPCvFeTqRZU1FIPrn
wpJWcFTBYTNZ5H0GkBhzVN9k4AJvluCZjFByChMb2is/SrmV+sszEvUCGBoi2Lz+5+f3Hw4q4X7t
XSyo9wpHtJa1naOcDCinfIsHoF9kZWxeKa6p5hMLoMPLvj7W5D3ULHie+BHK+XLPRMpNGC8uRCdn
PVJZZZ74XLjWv9RRREN2bNM37Jl2UirsL4Cibl0M/ufyqpIzb2XdurBYo9LDwPArfkeKn3XYaP68
VhQDUtVdVU84Cesq7CyBSU3B/Gdh++0w+ImZuFPd8cQ5aw1osxrnUFv0eiE9dWtv5WKhbyHJfzIs
u8KiFCelWODrdxBX4Vj6ggN+v6F+zFnGh69jkb8H4Vxax/PXwN8SFy63mJO0Jo7kxuy7zvsJByGY
ZSE/nUvF/Jz0H/vs9qU6MIEMDENuqrCqMlnVx88W/7YOhT9bIIpFCRSnOQNgV3HOg+a1jB8pDBJ5
/GU8VjteTHIP34DK7/AFYspr+0HV/R8zwp7A4/L9Oi7xiZs9bgYnwp3IZrToWc7mmLMvtuxsOj5/
Qj6DF3AFfasG9w0aJpR3Al2RdmuXYBYIHM7l0uVebyDdlVKS2ZHj3yHjQOS/BEpkwfyH5MuBOlM9
nJGllOrsZ/8PkyMMLZyI+hYQ5YjzldG6SQFkt3ddARSewMbo4Ih9piZ16U3SySIS0zg9qWtaJQYL
dASNhiJtHoiNNfALljn5KXzhZcfFMQZOsFs4Dcw5QX29J7iZD2FAe47BSnNP7s/jJXfwYZo9sp2d
G4MCLT3J3hVHeHrewMQ0MYRzLs+1tTx+RHYyPVU2jgnVABLXoIVynmjYX3+3aY0PDr/G7omWGfF9
lwL+bcYcANTzd3C97S1RA/4OzKUkwe9qroMR17dDNFklaqrPtPc+GID2ExdqDWGmpsniS0TKNTPi
aqTEHerQwlram3/VzsRLdwJUrMxZ+O5Ddlv6TqmI+qWYcBgVOXRxRCaaNWCyByZshTG6YZzCb6Pq
otl//w5HWCij/JU+/CxVcsEGubWwPxtG78+x/EQ85abokcQoRrqA35tbtKmEvspHU0LQO0+u3ycE
6wCj9OUkljY1lkvZ6D4FqEusx2PC6H1tOcDdPgrsKHkBP1KjQBNEmo7CT+yYvSZYQxJjuiLK3q9+
lt4iO+YCiJFTlyTcVyhzFlqKhR6OcyHA734UTlfvI6E98xnRnyulHUlHTvb4YTqF+l2ezAi6ahCj
oXhLr1XDm0xjyNQAT4J/jJz4wB3fLVpIdoWxArpcxj6akWIuXdDT+HYmNTF931b6gDFZ+VLEit0c
2wFnAj4QuBPD0nUQNqHOhUcPOh+DEw20mpZmWxfHSzn33WNVOoNJxVEJ/gd3cdclmBPzMO4/hMbd
mbL5zmsTnHeoyHMlvdxEG5PSqkyqLZp3NvramK7sjUpVaTSwEnRA3gi/DneyNTD3YaeXstqpfqgO
2ig1jtID2X96Aw495q+7Q6CGhKvrT6RA7oHx4AUodvfB4cIuXfgPnRN/9Ey37VZY97L4CdNGKu6a
riNCcs582MCav0ZqxrMNc+O/Uk2t3mk/Va+WEX56xn7jGdCffIMclp3QbzjSKZ9RcC0hGBzdAfDm
mvh7JXjBP8ULcZlQnzvGKaa5LbNeVASQRXVZfhWcgRamqZqHnxbS1xXUnfKXKucqcPQzcmkkFFgN
a1frbohfUwn5nTIZ3cInzdg1tartX93+JeSlsBrLMRqLKECoB2qq9KnXxAWFLSBJOTI0GaifwCid
DXArWKCJi8WsIdJsnIc5ENyhmozDTtbPH7BPotoG0T4CQZ/RrYD2GN6wJNukHkH4mitmBEet+P6Y
g6r5GjMtuTD1WYLtfCCW2D1llrr3RYB+hGWFTlSzNqeILDxmCyAajx9eP+0YYuxDX/9RS5Iic4wK
wAlqEzPc4iXblQUGq6Lf0kB8YXXu/7YgsP4QFWoqnPK38vz2GsLdIhX2R21KQJfrbw/s8AqLIF2A
ZuMY2vuOKpH+Ze8+dJl45dYjtzv9Yckjyl5RtBMsoQKOc2FKyofQjK2LOS++Pdo3X/a6gXtoXayw
zazdmoCz9Rtslj2vB/VcKxNiwxqqWSXMjoRqj17y+IgiQWCr9ZHo9aTJiQrQbr3BKVaKFd1hfFDk
Em/XB4xAwzuBe6jJ3lTkntmoEfd7HR/6cYFFrJRelgcz6U3+1L9qkDOO2AZBSkVEIbYffonOwFdi
iJgKgIPnQoKQ1rEziW80kRQ65FTak/bi71jO0OodvyjNtamcsQEwLL/0PAuZizdv19cGgAc5JOVa
Mk1ibD4xc5+Zc6KN3uCX51rIB3QZlJ8O7hOvVYXN/S8ENtfnFl7t5U9IzFqBTrFkcHwRK0hHBhNo
Vm2F+Lvf3AjIlNuD5ofWM3bhzi2Yj3u59qmupU+y52nRqkWTNK79ISgNO3MBCD1RjuP9y717cZF9
tUQQYi9sXLdbWfaALErjKZMLVGKIGlwCFvuxqOBU9iy6o4Ro3G+YqWqSnQ3/pLIufFSx/b7BQlsF
rNnaCD6eMxmQpQpw45+wYeOgORmbz/aDP9XF8j1fobBUwQfAa/BbehxwF+EQKGPcP7pfiy+vn5i5
tcu3mWFg3QazaVm0N8zKPca14tTHdTMEo82mYt4JNpAzMq8fTyNXLSeY3+vJIEEkQNpyomPQlILJ
p9lqafrPsUa9U5pjZU9LhekADAqnzZbXe46CNEmwPHYjXqwpSh08zTWH5R+P6d0Ajza8gcPFRSqK
8LWoyXJWYGpdZzLFBURbl6ZFM+zlKiVvfyP00E1d2WPMywIXYwZU2zcFBHicRLa9xM+R4c/IQEbY
eO+QqBTTGrI/c1OOSlgw4QNJv6HW687xuxUkf+XpaAAcWXwREyLIKS8z0GiTbXt+x64aSzv6Bb/k
aK4MKF3R0oLNIpy6a5s4wTmsb8R5yMaMOHe/ookFskQKJIlmXrqBEidb/FEVMNdxphtQ0+/x6yGt
Ky+ZFsylh7OtpX1mfVbe9LrvqZR+glsjYzKsHosDGCmH1Hng2td2/JeBS+YEj+sQTp/J3pRNlHr1
vScghasTdURShrJ5UY7+B9ZmMrrDqIcC2dl8ytATkjwcGC1XAdkr//bXVdtrztkOz4mu2DFWPlh1
BXAE3vKmE1HYAzXhDZR5QmHt9rywyuczgdI6F3jJbj08PpnQ/dNqLdUZULfnS67BCvrTx4vywUNf
ud9nRr+ckNzZRvzxwaGTCJEea+bN4k0kteoJPzaIs+JvY5TKGhWTNaZk2T8Xe48NsqNKeshssA2Z
nHbIC8vGzlNw/46xLibZUZKhT9tQ3fMmIbrpJ8+hS09dC1j7Qkjn4k0+BkOEEwykdYLc8rRTy/gm
LQKXoMS9JE4FiBcscxLJ6mpSWQmZanP5GAufFGC2xRzLHJhlu8ZQQa/eZMeaX8RjxhOxuJfsqLhO
Xa9CRrsX5eLq3BIgKHodvdhWrM/2vYI2/nwVu5rutgjnSE9BRnI8OLmLzYk6bmWyOj54IRpHKnAq
IY6Tt4h2mAyUx6W00zwrDduI1OQdsEBYbusR98NEpx5f2xFRFYbO6fIhap0NRsIqDqMJYG36xxIc
fIT1NeLjpmgFJKV+2xiqpXPENSd6vf1m5nqUaAsR6r0lVt3hyV1kXDNRkb+wj6zyLwySAnhhD0Gd
xJdtEi0m0zEalTplhBwYK7bDF9/dQa8kh5MxClTjo47eHmQU5pLe8VAxt1SqjNVxGCW0rzJ7WnqF
MA3RkIyH99Gk5oYjaJa501xrnao0/qnw4YsLdmKSZTMIpFVqBd4/tcmJ3dKil4oErvmIRtMiOThQ
xBWDSJuogXPL7h6Uw3naQ8+HWvlVMqyVE5jwGH1kd+Zl96Ny1sfAEDatxXL+3dR7eEnHWgb4O97u
4MWV2QU32xf+AU9e78ntj3ucjLqOThcFvddUTzdmWNgQ53xrunds8Da4217NqnY8OEQMJrVokiif
KXfcMtLQzW9kUsv2i69XGpoDoesxiD742JyxgVbR1OGtyby9auusRptvFs7ZwMTeuCxiwFUheG+u
kDfwywBDbTr0UXqTfLVXq0GOEEuzXv50zYzXSOJgndgQD3lhMbFi1H9MjLqQaXynhWiBBzafYqyt
Keo1J4j7pqJWbKwbxlgx3mTMJ211VnUTge0IF6tzrAJ3DftziGqkBUyzPAuWYHZsywDxNjN0rPgI
oQMEfy/L/G5W3MZxZvPklkcpWREilC3bTpQVG+hWTVJ3vqLRcwH4ItUJRE5+LQLdcgL49mrLj5ER
d07cVgvE7SqV8kl4cYjy1p4dhESs1rQLXiyzOpoLFQKT3Eaq/BYuBUvE1DS95LpJOp7np1KJgYty
fKJ2141pDUx1c9cli3XdXqJSebRVbbDZvQBizInjXsxsyThME5k1bBJQTibl8LZpLHrrq7Era0Mo
m7CZIARgki2YSAcSjZHbUs8M2pXZiTWPLLWyezWLe0PSPz4TjByl0JaqKUUO/72+sT+LBUuTNgFJ
Np8KF08DWgOws7YeDCWbJ42tjrgnWarjJ/doJZhocoUScv0/xF+jpP2c5BharHF69ybo9MpfDk1y
HnwGUDcVAcFDmSub8EXA6W7wlw7fbXY/NfqnuDMZYLjjWlINlrf/PjOwi9MnHSM0/6xaiFPE9XJj
LwmgLlwtyk7Ct+otYbocYZSNh9WP/f+TBGUJ0S4AX/G1BEfY7pZ3PoOW7zcRJq01g/Eu8b8fNbOs
6SjPu0h13wQtwvt4gy+L5o+rSuYv/cEHKjoeo+Xx+IQEvxFxlaC9ZM01YaXJ8p7KP5Z3QUBaPHN8
gKtY39amkPnOC8sMr/jezdz+wTarX9ZiUqcp+PM1Rrc/XR4+vS5ZGvPzMaHWKt3kRPkiGJ4PCj8J
t7pL5KuNu3KQB1IbWZIKkjhqxUR6LHVrBlZvbQCiBg8AHjQaAGf+GysHshOCGbDeJIJ5gtc4hT73
d6CvdMIZ/rHD3m64jyumwri1u7+ibSkXbF6ko6vTV2XRiHcJins6iVGPlY8Mzs+12hBqVa6G6a24
m5j44T65HjsPPFd/nkhb4HFaoKR95w2BEqTKvDQ5IMjkl9QemKW8Eh+VfGcQpmqZpKVMiC7PLfkH
Vxi5PJKkGOdiskDvHtPom5vwy08jc92v0HUQwiizzkeZPApadyWaJD9GBzHlNVdZIq1shGyf/uxp
7aec4kmE7usa8WC9ai+40fTSZeMTIsvN633UpnJ2CVknEWBP0/vyNc7QgKAj3vDC0hM6+CNKbcoi
URt4lg7LG7THb3UgWYGo5u/KB2/bUdRLIeXx9RRqwBHRaOenu3wlutRaeZ9MK7bKQAMeJlj9LdPM
AkMUC3Mow1vrR8pmgd4v9cPsS2QIaA9IN7Y2EDC8ooicEKdpArE3J2/wsXAMgDzW70dJWf1cK99i
9kvCrlPvFSxp8pmSZUt9lmnkK8j8IU7H8QE9kqg/SM5aZL+WWBvg0PCqlnw5MuSWDDK6/P9EYst/
XXWECZeeoed4lI0IAmt1RfD580qTgCyxVxuVaVGKfX/M/5NQNWXuFVxWVo2lejchsoXDzwfvNi/E
eTfmhjViA7aNDvKt1qOiDExXy/+vGzoQF7s1cgo6x7thxUK7fqPH0NLpvYagj94YZfdln/CLcnt8
NokU1hFESyjIoC2vRskmxXY5v5THFbRnFspSWOiYM71iG2WZaLdihX5N5GO4tmfMSHnVJZgfuAif
62b03VY2ybjG6v7+hlhxkfKrXqK0xQiqfPqILXhExShT7fqiwRCushBb65g53v/WimkuuerVs237
THnPrVc9hg7L5WL8u9CxD+mnahrOLyHAt65ErvL1TqexKOV4Xr8x3gfQth8WA9BHjZWA1CWu7PVc
K0KnMH0uJ/GdRI0BKcqQDtsUkTBokuYh0MfQlHa3sYN6oxQAdeZpcHZ99vDFoW85Ki8ojf+zXbXy
W57vj0/RRVoA8GItxEEEn3zvfPr7kBy8sTBrzL2lsgb0Xo3dabV7glwipVrqbqPPhwBPOk3J+TMT
XYoywfDZeSX3Nx/awXq1N2oUap7SEZJ25hXa1dD0Be70JSnJbtQWVUwgZtqGYSHHveWjx6HNv51m
laIXPlV4daAyNnszyXwanj9p8nLSA3dKWEqqjMr9MdPJ2qQ0eyJaGSg7E6/wTXuMusUZKjNmbaNc
eZ3MvtEIGzhVbpUYyeKa24TslAyxojOxMprqlXPhsgsC2afMdbAdC1ra9y9qnE9PGauAUNUlVxZp
Q54PUfWHNgPqaaZpGz3gbOAiRpVOBy17Pd85ZSrofOJ2kXrPuxDRKKj0i1CSSXsrI8nZ+Eg7Jdrg
TjEgl1x7CMCVnlQQGkM06OnF7aH3Kt8evkkOWRgocNgcGTT6yQ2sq809TwLMaIihYK2Fz/vg59Gb
jDarpA/APYnJm4AMVF36spheaFaSHLW1x68tFKFy91SIlzDVLLgE1GygC6yM8HiGruxycl8kn2Gj
VCU0s9c1bAl6OsNy5ngsfUdnJeUaI++JloyUZpW73Ybwbz91vRCEHgm9KHmp2jxSo4BU5+3c9CmK
kNx/AHJOyAqjFlMcoGSg/XnAY1gnKjtpAis1E7JSiZb/MclIdNukKUXsTXRBoEiV7AVRByWtc3ND
5ifwzsTHVbV/qGFoyfYsPAn11bao0tmgOi1zO7da9R3lXjN6HGvaSQGJqp81OMhXJ3qVTi50tVhK
TDGyRuH2xPdfk18nAtU4yNz1+gD9ex5syxnEaRxZd6fn8Ku3EIi3WbqUthjVFY/M7PyJoKl+HTtR
l+v76luUdlrR5MpHXCBCr13ILzwvyxnKjI5LvS9AD2P8WyyD0JSlM68rhgwUq3rfAwKoi79cy406
xG1tFvv2Jra0jjrp6C1rYY2aDbpz8f//Rhiejkj/8pQTdfs9j4FLMSrHs62vncrOtPFPwR7K+xbx
huKFGbtJXQokOZh4KE/xqv+zPJxteQdA/ZIzHiCsy3p6WmoHf/gO9EGn2DPB3MQkEKeojIsv8Pkn
vAyD/KH3kO1s7mJ5uHKzfPM0bpjly3MyEqiaJT/b4UoKTH+qQL/LTzcfyv5NzVwNCR7S/AJAkxXB
uExbYer6OSoGHhWfYRFUBa25XTpJhwPIMFMgF1wWrUEYjN6fDclyycTnQRKWjPnlFS4XlPN2sUge
uGUC0CBK344sY7AQ15jQWGnKIYZQi8NQwWkisr+l179kx2ChS3+EyG+fv5S1xJQunLC+Wg+kEHme
aSImJvI7lpBkwt4skHWJAa/3Vy2l19MCw34d+YkhcPruvFNZHOES1uIsuO9SNjCvjcpzUC6E+My6
EAK/VdiA4nRIQMyta80oHYLrn7NQpjKEGXI9BZ4wfUzFVpALNqT7U4XVlyk01Q7YAeZXIHFV2keF
I4duKRvgFlGZL7xceDx6Bqui1wd52XKe/hgwnfWhYWtpwgUCprviPsuXmRqnv2sSjMvWSffAz8PV
Q0tBA2FrznGisJCsCIb3WwUPvxqt6V2Tqu8X0SaLUuL7H5JXuSuV9EL2tKT0pCiNw9C1oRffW2Ds
cbNOrWwNSMDBZ608UFO3dzofFRvlKTfKrdTFctjTT/ZjsCttPnhZ3Exrox5BjmRRmVA2ifHq5zUv
rUMpsS9omGAZvWJIVQREBBdV0hNJVQ1Bsly03XxegOU7u2uhaic+hbD9Xu3E695WcDL3rbARHn/D
bF7swtyvMG1xfGyB2rfR0za5eiV5/JOEQeVptIEExyx6swfG4uszMVQxwXt0OErUvk+xKufdmzOF
OgUTdFYr749B1r5MoJbd1GzjlEfxgAwTWZch8JpbRkwUrXXx6RvoRuxcwnHm5ywLIsXK7SZm1gTP
NqoKkrMaIbcbE6Z1kLLxHEHkgS8ZVhSx3Ll4m3zwMHMiQ5TJf2Z0EVU2hXB2iQUGPqvEsCPgJZ/A
eRqWDS7R/FLbLLnjvl4zERZvtKmGmx2xptF00R9WOqrezo72rKPZdJ/udKH/7kBFJdTGCzPyCtp9
u6Of7R9fmPO76ZRRfyIGoNgui0xQT5R8x1RxcGxiI+1UapZrQpQxZ6QHiurVsDCcrbk/fmZboHgQ
JGukrgBnG8kUmaaPJmhbT9oEdA9DjSW+HyAwN8ZcJytU7N0qUELTJnyerxeS6+deOPXyMwx92Wxx
rAYCf8ybLnJUVYoop2sYMY5p/WhwmdUGPNMPI+HicprQx/6b6K2HlGT58w7X0OxCEGXrvrFg85kP
e1qLhFcq+mB2bIXiCtUUt9RMTUxeMQnO5LcdeZA1BmUo4OR7+PozsACwXMp1JRCmCvq55fJ72+Ph
8WQ5ROF5e1xQQd5oElSr1NIeWpm01lBlPS/xxA4hWDJou1uEHMi5+C0O5diU8SCsfuFAC3t2rJkY
Bur4NP6yC9LNcQvlH+C3hU0grDVj8w8bLlnO0NFwm1D14hn53A+cSLD9RjiSLp1etwsaZgIT38kb
UZsttBsgsgXEiBDOxR2iC7pyiFxLsnNgkmPc6Ss68CD5D1kzgPIh6qnNbSJhntW/hjnknWl5WvJl
+0WOI0zlxmqre8NNarXHDJPCa4w5IBVX6IdqTBasHxmONeGWLOKMGlaw0dZumaMrayeqm1aAWjlO
cltcoFMkK/qOBFo2FtdIIXHH0mCCcK4HTRCoeDFJNjX45ThS7upcIjCJw2OHbbSDdr1bmQNH9rXX
7Gtbvw5PKduInX3XNvf276ahs94Po3tHpgkuG4QlY7u6k/UU5MEXed9FRJSlD3p6Xe0CoDWaIT0e
yPV8+3d8p7l+GF5lJfqAbrWkyW/9/dv1qVizqOYCoH4kuYNZZmuNwFGpEOVkWeHIvYkbY5iiGFfY
sNau/qcTHV1R9hnYjmw+ALF98Gv6vQHixrcktJqvc7Ac0lNabghGAKvLkwdQO/AGSiGFJOeWvU7N
DaV99eJuOAJZRT/iNX3arN/UPjuzXe9yu23MZvyUcSUAiw3ANn8CkBX/ufxPRNga4PcbDfjTvoLG
0mRn7+qH51YEworPuQNMSgWCKTu5QoDOZC711hH2Pj1eshHn71XPWlp6lvAei0JMtK4SbWi8bTiS
rZTOpYkz44pRNIXj19QGjWJ1GqIyhNvQqZ5WEMpc9eqUaxzkTDfWbmTptjXkqcIokE0hT/2z0QkM
NSePiA+L1E73OzC0XUK47YsaUkqygi4MmuuWbGtdtPNuJT4U7Y57o+FLZaL0mPpPhs6Zbz8VKvL9
qLZcie2EfKtot92TqNCuCA+McWBAVJeD8MF0hEigK8304AzMfaxgHg1WhxgE2B/ZOr63RJlFb+h0
ZckrhL9dtUUNDHwW+kFdF0yZOJ1L2Ldewjf5Z7nX59OSC0nhEpSy3HKM/aEElOVvQkGYqs/t35+m
mnwCYUVkgSPYu3i6pwWv5FHwrh/c0GTlcT14vMxnBT/LQCN2fqrnHHBwJZEO6CqlCQqP5H9trWzy
8zs8QmTiP1cBobAd92JDIO88vUL+GeB6zLje9fYMG2f8QjoQoyhScsz+ViYIyzyJOV6c07lWfPAd
GESvIN5o0v4EBknSwghXo2eurs2gd6n2cscgy+O8mVaVJR9AqURspAK8J24A63dlYKkBoUcZS0ZZ
l6UUz1INwkpOCoqlahv4ycE0+0mOAwAbG7Yk7E/AJW5bW6HW0zjOIRl3ZwQGfoEmOCLtNXbdCEh1
cSA9n0RcaJujRcGo7JCBGnY8q52C/gldkTXIK4cm6h63ethZzXKqrSCgsbhfAX/s9Tcm+ICdvR7B
KbjrIPQOBm9iWzsNL0+k/5ieDiI9tJSV2oYvaFoG3KEIAa6Ejhfa4k5q+/jRfPSUv6OzdEBghuYa
Myyb8Vejw/qlVcRVoyLmEyAZ9RQ5DEjBroZ8qvVpK8+VxEXT1cKGc45SwFIivHc4zzaMOqUOKu01
/GT7bYzTUX+7Sj6jWnnT10elMZ82PGCxBSlmJwsCno/HrrkzHWO0zGfLKJccCLAL435ix6WYYXAh
QJhlqpTLIxdoEZdORCIoFZtxQPeWddOEDUAQ7Q0Lj8tB0ggyqehCvT7HKOV6H2IX8TNQSXfF7WPh
fVpWKud4hkkTVN9Oen60JQXDPp7LveBaTqbkEgRSuBMycb39S4aL+W34/4EvQkTOyLS2FuB+8GkQ
V+MjtYP1SIVFMCLfKJyUlQNl39k5cxYTSUV2qT1V32x/1HVmhDZEsT09qJcLLbNQxYPfwhwuFkES
xGE8VJmHUgQAn/052cNlE17DEpqTBM71Abl5CUlu8CW3q1T2vr62Z7TTiMag8Slsz+9E7KHLGfMN
jrhkibcxqYv3ozY3bTTZb7av9vfK44xzfeLERplpG/KUSr8xG2NdeFx2/nCXDmQ2+dC6u6ubPj03
Mrcy8FJui99D2IsCh0bpa6DOR9zIFPCKC37ge7rEd9W3tqoqcq2FBxJR7u5/fxA3NzBThz75fVFQ
KWVhgXRy8IKV4iwJY42aRVeKmS+lZ0yaBcaf5SNmo+5lyzCmk5UJuOpOJUHbDkGMeN4oG0+fQQSS
CCutE59gi+Up2y8Lr78A1DdGrttiTCdTGFF2ojrYXAXppgbBddZ5rfnZ/Dp0tcv0qHsdcttmuDci
YOpraKTTzEtpvAP8Sddci+e+CHBg4u8j8sEl6I6RxlPlmZ5KcWhUyQHYYBrF1bU7QeSzy6elCzPo
BAqAN2xXCqnlZG6r5a8vQpmCj0Ys7ICNFvLHpFlVhir0A/V5kbIoHmBDgVFB4g7pYPcxTLFUdej+
onk6c0RviIhyyWYg0oWpmX67TtAYmQp1mWr8Lba7ZP/7axT6YtbbAM240DgJ+rS5xExKGGlK/J2T
23XUdSLnWep2JXCq0RjnLeo3lvr7rAZtQSsUHgnJgeU1wrGnYUo4HMbVOx02107chJJ8EnRZ8tg9
MjjGEeL2tFeFohxIWvWY/4hcIOmw7k4jdz3Xi6WDbGcXSiJLt2dqBllco3VZKkPD4OB4StkQrXrj
l3K5LzOeFLP6sq/QvNj8rVT99g99zYkWL6DKHgesvYE5YNIpJLeXnBVW6Kxq7zR3lK8iLJkyKMax
zTwQWc/UXCh0JSlILoTRWTP2T12skDsbQrYColAvdDpqiRcgs2DBC5V9mjph75Y4ogO5L0VitcSa
COsaI/9jSqakZNqR19teoDi6YKuvJ7RPXgCeoIJzcEe6MXnOEL/9JZ4OLh9JwwXvOk/D3oQeDiJ+
NwICnn5xDxfWtGWKsGXNhQxQnYRvPv41f+kQARBhwK6CgfCslzbzuzj0reF3Pn3QnGdFaAJUDEhe
pjJLRxfumpEcQI3apm89/CDwwcjILZtp1TUgAFXbjntE8Obbm7I7QbVtVIPaRgVRw2Blb1zAibRm
4Q7Ign2LHzXIcTeVtP/HoWYRTGZh2sClIHWz0cA+lD288+75uOfDgSRfga0tVNZIUZHuL/R6HlP+
UfedNCSdC847J4efTyfeJJr+GqKX8lmJ4OKKZvbHs5o1ClO0jv7PoKR3HSiKBB0nmRCU1OLw8hNc
4//TVVkXA4sBlFWjMLm4L1fgdlgsxY8mB0WBpUZMC+NAfsp/QfkGWa+VQApY+j6Gj7xO7aoakmJy
6ugsdWgINtutKpvUCYpp3v8laOGcwKfAmlCeymddU2sd79GHbxWB4mcT8/fwpyM5EmeWzmgusW3H
c5pimPp1hNFPEv8p7r5d50CYhcH8y14IYzGJkN9lWivJU5juEwGJMCq+AepVBwDUy7VT9v5S74ce
VzaaYXs0tMMJ2bG9xkCWGG4w29V9k8sJ1J5w9ylE4SOP6UEnN1jsnS8xqF7TMp8hXNjodBIB822a
+miMLV7+FWMNohioHp34AxSAR689FKdrlecLHVJYQnZeJkHYRCXuASTv1qy+9GSNwkVlGhgi4xMm
3m+ZazwC58JLBknqpVlm7e7XIi6DDOPjH4UiY92hf7TDqjb81cPLthL2FGExPY1JlEk81zT9PFhM
xbon4dEaxESslImxu9CddXJEYgZ/Cq7YThVGQr4+dsm1J0oy+P7Hkve398fGtrONZKMtn/yXniYf
LTklpGe0k84yJ3LySpeChBqI2bOJKSOkjLl0FXYCNdTTYmLZLWC5FhbdTAJlSu3GGxwSmHX5fiq9
nlzgSPr4K48sfa/v/FWMVYblmaWU6ZKCDg1/WV3dC2L841mIzb4X8TVsQSSrQHFdz9pdbM2zDY7O
/Xqg7t4/y38XA9zv1GBOUcA7eooqBeNNCboV9G0kyoYmHMf0btSaInVNQQKRGs/6BcQ6dix/oq/L
P6o97UWOGDKN5D+QAEH/ZI4a+gF0zlLXgbLj8mdMW2dLylvQRY0wfVUlCOeDvqYpShCl/jB329Ij
GZwzgICjHhfP+wsSHWDMF6QD/9H8MyGXjPvES236PHd0j6K0Lq6uPLQ6VStolzmRRb9F3VY28rAl
lluN+e822WnaQSaiFBaTTjMrY4D0lpegaMcnJEPf4eKNb4HzvOgNPRTvCAWanGhLlATDcR5iXtq2
/ikUsQBYDKTa+pb3KEdZnElKqtUXiP5U1e9Xxxu8n0NWdsfYYM8IeAoTfW/WCMkhsBOllQMqQ1w/
wBgzEwDFPH7TLLbJD+JPfT6TzK8wQ7ZRuQx1uA4TRCHcV4JvVawD/dMtTJzT5o8cMtT6M/gJPdXI
E/CyUdpATtxlCo2YgPbhSHuH3AsvgIm5rr32H/IDvNdLVEmRRtDP0qoigFQv5qU8xS0shY0iTwGW
JTOP4npVSNEwey0qCwiIfL+J19BCA4Z1ka2bYbJk+VoImSZT/dkrt4P87OnhEmEl6a5sOq3n+dpg
HF62BqOaqHbgHnUWrR0Odic7WOJeIiRAd/alpHTJNs8KYQcLy2ozgZmKTNNrR4lOBPdgm30JisJk
0c4N4jqqgyv15q5wK3VweMT5WRIypqGTgXXX/YZUG3IX65S4EH9I5ftI6Ob0tQtPRsoKdy+ThlBA
hTG5uMv3kDkgNNE+H7QpWLjcioM6n+SkfGxoEzbrkvtxbcQX6YJ9vJN5X0Mc9ERCZ5IVnp2X4K5f
LZICAEFkuW5P23U7YxiOCEX8F61yYXVhAv4S1W+3ROZL5tEPjExiNp6yygNaIbpAkw8gRrEU7BbB
aIFWOcBO1PyOidtgVqznVzyPXj29jm4cSwohs4vqB6t7wFvLuP3XhnG9HEITzY4bYJEMm55dwAD3
g5MI/XXWSEAiHbaS3GzK3ANxf+gH0BY4PzH5wD+keMkb6+kGVIMNTeEWPak9cUuya6lV9bp8fWuQ
++moIGjmR+CRxxFvbYINZWtQzLJskU8rHic7S1P8ipQ67xAJbCapJYdtugEHoHTOmW9qTgRCpmEb
t8ocCLt+x+//Ek28+LAu3OI84adYHcEBqkaozMSBSEB8jQftZTph7y0ljhnFkvTiqJ7o2P1JhZHy
/kivZW2m5fQXerJacPtRI9pV6tiklQT5lM70fiqYS5HeebhBg80I2rmqW/Yk4k5JYr1R0ntYIAlQ
CfcqQ+z9RQfNv5A80NxxRcbXy/mvmkyN3Azbny1PHzbqz+klESXtef0baLTSUQBVQF6ZG4Eur/Jl
gIIBlKbn9wYhzbJlPa1COIvUKhySRkCmUZJDN6gZzLc8hFXM6KYXdMfPR1sClIjtNMMkb398j1Kq
hMolbxfPfqbQU1CqmcMQEiPf4+5OEIUfSHgtgPH2h/xqW9B1ASRfNb5cRlr4XsAQYcI5kUbwi3CP
EGCBEn/snXwGRO1wKGVetK03WRoFjDUGGE2vC/NYFSKPAO1jMIBTIGm5ACHh4Z0Vs3D0ivUrPtYi
kr3l9du8P7LRi0VpK9bykRNzR857hV6DAG5uCTVN1HYSYET1L3eAgB2miE5UXm7lZS6gcV0ToVDa
f748doJVrIP9G0qR6lRv+Wvi9mZQyvL3DD7eHtBZLVJCImlSWF7B6Z10dTs8OjpmHcCzWyfZK0Dx
8tFt/mFebdMYVpyvzZGJvomKFGtxLL2XJDM/S6QOdOIsas+jHbIx/8c8B01dSPvQR5sTXuvqKOYK
mQ2E+QEIzvlUkqHQk1U+/V2iHHpSHTc/vGvGNtXDxIPaaXKqoXGWBw/fGna7hpV5AXl8MJo1PmHR
kUFGsOrzkuJVRwMC+U98nHJMfd8Uj2quRMM4cEFo2Lm5fydvQDb1q5nCKiw52Itf5h7plvqiMrYN
3MihWD5bYodBr74MC+Orh0EU0Igp9UWX88pEqknbbxy/tfYTBoCUPFnmWILYIxt5sW/dGtMn7N5w
GtiVoWuzMtisGQ7Inm2yPZAKY66agQZeHykw/1juwr010YgomvMvamq3RtsYmZcSvEiy1eh0hd9d
MoKs9ij7mFigdHXXu+oDn+sgI+djHibBGYWiv5mFqITE0HfEiUKH+WdHtkmBwPMGOK8JFAkFs0ZV
5R7Rgqyyjb73aPc7UEEDa8hPD1pfKWPoz/xjlzohBb4hSZzb6JTMd0gfU0WOCVIRHykf+Zd9w8Uy
8RNIULVD8RFZ4puaLDfV8tRp+U51yYBEQa3yrJgp7WR2sAxY8QkNAl+SGzvyR8Yz5lpFVk+8Ra/e
Xo40WSX2n97SImKka4mSLyAE8bFFsdXOjpHm+bU1m8j1eQugB+KVMBDzu98saK8mlO/1ozWnHd+8
AbQ6WfC3Cf23pIeYWK7Tp9rkSa4aX8i6Mvb3yYDeXBqgJjQN0pMMkuOs3Ht8GFhj8ZYCeh6jz8NO
7zvXbCGjRPFwhPViwHfD616mbuEbCpIxFOf1i3tuvGSw4s3ZFFNTFgJXsRp4ERvuv2nw1gHF1C2J
h49ATkLDlB4Bjp85BIXVjdBbTJECIGM/gSn+vAhq02uJPSMSCHxEgjlK6YHIxwPdg4R6B109Xk75
nIh0BF3QRY1yt/UVti6lMGrHrtoEj2r69uYjOEh/8QZqsG69PncqBv5SE/oMIqUGDXbB3D0QmsgU
IP3WM1Ok2XgIg3zCll3tQB8mTIv3mY8T6bTiwUcY1XFPjJWwY3pa8gOgsTNSJe2JsnKky8/wOCmh
4k1AWXphoGv5M7K3WCobqUkIRJ253prG5ruz1WkwWhx2+NZE5UEKV/8+3YV/kzmD9etSsfFWFFkv
XjTqfHo44seR/gDmKyYCvD97lc49jQ5MssWHJ+MM7bGu7fxhVsBhSPDu2a4VaRJlXeVM9uLwLEkH
cxSYKpNhO22NJll2ZBeJ4ZJyhyJR35jCr/SjnLFVFTUL5rnwc2zH9lHhUBQn6JU4RRN5eWAYzOLd
qdG/68YCwzUn/XfIIjiM7WBkfRxMD06b+F6Y0cRVlGXkhstKnrjD645pUAQu7hu15R5C8E0+ZpQ3
jpw6ou6KkVsyKVBgDNJAM7ZXidn/dKKeuJCm72fu8enRfWS7W+X6UpfEQNiwCNDhQKkR+NIlExKj
xAIW5T5Cqh9CZ8tnCSmZF27dbT1lnoOozRclv05rQfI3sQTL4jR6sMKsmU1OXCZwvjhaVdS9FAOO
N9EZQs3Fvrp9Gw9En8VJPN2QSEgGuydEYlSWXfBQk/7VP/YUf9tSbwJKHqUc4qZc9AygxxaPwauQ
Xrm7KxJUWwGxV0iF/pbMrT2YJFL1UDlCVoUsOBdj36unA8f0MZQHek7hdyJFJuweZrez3hK9+YT1
69meFZagAoHDKPZGgcJUPMcoPBuvvZx4i2twvWSycBI3H2DtavkET41K1fPmT3gh9AMLUoy4UMZs
5zSgRxkDzT9GlsqiVvOOpQzHWkQgm/xpU+BZFbc1cRaeNTYyvOsMBlwEktIw5OhOH/Y42xj3WBhH
4p/mYVN3GmDS5dR1B2j0A2u2wdlJy8OAnu8XU9i7dhyBncgk0xza6DBbkAxxVJqeEobl7lTHqShQ
HDSmkao45Via77oSVlFddCErXprm2blrO+d8cTDvjT3Vh4Gc8HtcmyjE2v6NWHDPdPvZIOwYhU5t
kwKOp28/mE5eNMeNHz7jGcJC/hj4ZROQYCrcgKLJEa0UNF85UvTFe1oTB1v+yonA3qrgwOXqS3nd
Ocn00iVSuq1hTNlIj/Yr+SKKRb8fSFlNm8rtDX+Ar2CKgMdQdxjTKk+Calikd48jEw/3VIgMeORN
dv1pqs+MB+eRIikG1kF0JBrjXtan5K9f7gPzdwVCBEMdVaLrrN3Re7yoTrVJw5FWRI0Y+ar3fELl
ApH3PdJ2rOUF9avwwPRYFBxHc4JmtpL2vlD/BERbqSlnLefLU5Uoa32mHAizcM1fzj/shvG4stGi
OVjMG55tZAcY75kZqfQZVlUh1ubbOni525oYldFuH+/V9uFOE+qk/qFdCnfBpJu5Wkaa1G2g676w
0nQDU1o9ThfKtixvW9CSVdz3Rpu09DNnxv91EY7+lihQant7ip3JzI+E/T8apx/+6xpaVzLWelDI
MaG4j6VVUAmYiSW1RkAGT+rWceJm5QZJ2I+8FcMH856sTKRa7k5AkgmpJVWN4DvrviazBCO7t5zb
kDRam30jxsUiG0kErOB8OWuMjmgZv1LtwaRdo80dsuqZeRsR5mSOG5kNz/b19lWq86Lj5UkcEYA4
QnuUKU9ED9xhpJhPoihPpKZnzYhG7Y5G/vRrtcGGWNnoAx4U4aSTjQRk0tKwgUrEMFTtdooj0xrR
65FPXdzjdoM/ornAnME5lAq9SFdTKvxRofhF85fo0PdWgfRzfdeVzyqk9bTplZnm5VW2NE1hF3lb
AoqDwTZjqAUZHDPhcVbKkMjAU77kfYqwrOfafHHxWU6Kj8dWVgBmvzA63HkEpwsvdoR1SmYI6Juj
KDWyDEjqdKP5XPSFFNnQ1vXxCQpinVj+wIWVJjC8qykDPfWmRghv2MuS5FAFN6C459Lf3Ly27+fC
+8mbf5d8oRIfrLzAUamsPFKtH/8pE6pj1vio+Kk2CMlmmGjMuDOhS5Tw9BDeLITBLYTq1jzjTCJf
JpdnB/6eVmSGPHrgw/BlS/2sLebMmvHu8yt3rVzg9GvCAK/2MXAeIjCwV5ay4au3kJ3gnjkv6JHo
/JUOtRjzyKFh9yd9vW8D6gCAeqPh1ciYTkVNsrx4INgvHbWk2rC6W8Hlx5Khlr6z3+F0dsoDSgo1
tSEwoIzp1/mYeXWQuhYaRudgpNlB+cgBGSkp/UgeY8RCx6d1uPkkgTO3+7C33mxg2JHFNohpLHm8
kvON5SeCE97lU8e/6fx3IH13Zl+JH/A7oHoLZc5lknBf5zNpEo1bnb2yJ9L+H9fV2IPbg+AHZq+8
bta7zfesatuOvllG0G/PtDqm65/cKtJblJPatJ/lLA51/dB7QO07+mMLke9M1/C1SzK+yBNX9QHy
XfFTJuOOT+/t/PqPZtNjXVF6nFEKXySY/m+2nuxYFypO1vtCGg71mOl8FZJdVPAmmRBCjptPYHDf
eAjzD/RkRENQTZ1z6zaD8LoIjw89It2wEdrxkCwy64Mal/DLTSajgYVlMacv3Aal2IiN9fzlzLuc
nt2CYOFx2V0SL9OuEF5XqgjhmvL3PXnlH5LD8J2+U+V7Uo++LELCuuSyCIf5Buh7RbPpf5N6hxy3
c5In3ZpL22EBXUNCvDjUyfUOffxeJLdd5qWZ5KRh4PVDUDOWD3dNpRszgXyZDLGja+jckPNFN+u1
0ja8gBgrcO5JUrRAju2mbD8nRTR8f+b61NifzV/AZxubU+gkbLM/id0tYb1M5NzMzW3sSFjk1fej
v9BCHgKGHgjbvWDOOuHH03TcCD4Ir3uCDYPeGx0xC7KDVAR6WwKfoNoStWMEMVoeFH8J6uofKqi/
ggFspMoYKpYD5pyo/rqwSl4ACf8A1WkAQnYltW7qEX/HXUtwcF53T9WSYh6ybXIGVVl7x8GX48Yg
fzn87vMrIestfpFRTSan9u7eXOeSotRkjxvyKna722v7/nrUCllTXtnYtOdDOngqu6YUFEG9HkCZ
Rb0eo6XxPuCK0aDr9hKa6i7mLfom/NFXMMY2H1ErCZ2dxARHwuIAqq/CnefpMMWdeyOuiWA2RZnM
hWaZnfNM+074mTNjXR9k8HRSqE3AGSD46Vb13xJY+rESIsArp8ZTBv+OY6IbOmh/Wp4Iylj6/jbw
g8qvRhly2uvhBqj2GYgPW8FmmXn4FJ0T8qy7L3UjNZWgB8XqRvk3IdAiHrMorpZMe7h3RqliW5jL
Inu6s3nxl/EOYogFGIHG6k9bPv5Oll3z56A5DKL3fXaz/8pQhRQ8jlr3BokgD0An0EGHg0zeDxF2
vvxMJMaUIDblgWAErdIV0TYwxS0AtATJS6re3c4NbxpeGCbCQ7vkjK1BHHjsJ2M5MPYXr6VPPHYx
fuFnAlMh3BY3p49TFOF8F45qsLmOsaMOYIJrGjiKJZ8RfUvz4xRIbxt7nPXuL4zKvzttx9+XZ3pC
inwAiGx++LqaRcJ0eMxJA2wCW2IUuQBdloF5CDUE6NoLBUlmQHpwYQdil++ZYjKAfBHZbQWRXm1B
WbyUurk8BVtn8NVNmrScbbxzIntrXUfgMVN1nQKQcpEotdH9rMhA5PKvf1my2EcA+9iNilmWZWFO
ygOybJE3et+OIpVxv6V5DzsjozTDBqZFwdR/yBLfRWb9U7dDrKaaOjo5nolq7ag4rNBmYwj1XDfq
rCG6BvU233/ik0WaBW2wxOmO+q6ce7Y7HIIYmklQ1eZFtfLtN4+gJHsr4X527aJUips+ANbAqa4U
3pVTYhABmxEEjV5qPUMVLe7uz5x6jJFFiI6hYBeGZECraQnnhnlASWrnUWHdNu7Xt+NTs9sE71eJ
Kf9PxldyZtAlIKqHdAzqfcfKRsaell96p7qxV/JeTol5w8KxIKZVeBDvErc0R5yBaMnnuZU0RgSV
zletIu1N1Du/SxuFgrG4rqH3awysW8/4TDnxZpu0O0cToChA002kEPKLMgdZ7g68C/dy0tPKwVCk
DSF4KfIM1uz2J5x3+FbzQLThNTqL8NBJkadK1mXm+E9+CUrqQGHjqPuHRN4xZnbwYsOau6YswXcN
kzFdfYt9620FmdmeVz4MW/Ovo1k+oOuLmX0PFDn+JREcBAvsIvDch1TLph6JafALsjRZotTGKR4P
XqnTJzncLN+APG5SFeTHIEgMBSaEi2A0ynAkvfpgylgCriBzhKpWE41Fo13WYX9fUkt4g4E9/f7g
Ys6x+44K8aDpXYd6c2SX7k5VVIncbzP3Dw/Pswep30b0RmJ1fwpC+B3S9wmjPCrrGq9NaGusd8tz
M4BVTJm5x+7yuOJ3mocBWO91HcJp+y5cWTDXkCGd4yYVZB1UtKDVYyyuCIP1ajU3J9WCkVHnu5wN
3RjVrFuYfmF8gIoOy0lb7vmpe4WPm8dZecldqwmdkU/bWr7E2a4TjZslEHwq6igPCESTpYP/AREO
0P6sL0YTJ8kdC3Jt/8lxJe8OCvB0n01BtLCDYTg9lSBo71sDIM/B6Yuq0fD19AkkxZo6wyC5VwaG
fDlFHeC9hVAqPN4rF9eocAFC4aC7ggicXM/pEYLxx5sOpgavgMfketAwgyCKgqFfOf2gktP/WmCU
IP+pDRCBIUV/BLtwNNiLki+emQyGJfp0K/iE5+SBPCMuQHd3x5U3elo8ab7N2/IFeQ3qcceggZPq
x6VBEuRvmsYsXiJTntQM1pZBiCAD63oB3eGXJEJhRENIRiSkk5RfsdsmKpMwCwEQr990vGWxVUkZ
/SDoeP+Uay+R26qDtC71S+d2CUeImWg8PHo3k20HcGxKuIBsURivHaw4wPuROLCQLhCE1wmw9LBy
/ScnHg8ss3SGOuzcpEr5zXcg+3l+bzvOPysUmTzEKoEXatcM1gQXQMzvSQFBz655qlJWbeTIGWLu
HphRZsA+oCUoY6ne2wNamL+vebzRkHW28I1gphNuXgg2usdxUTZIQgyE2anxlNZL8QvZQU9306Zv
6TSgqfZskMK2m3V+iJuh0T0royd/oY07SXyqjjUxeRSMMY1UV9SEJI4lakS93yphlGvVVSWqUAD2
YH9OboVrmxszGvB51YcrHRLW9mNCL+bkHPSPyqledDik15ldOeqZPAZLmMyUfWFWfV4+wL5q0eBE
uNc0irY8Zx4IizZI7CxmRumFk8Ag8HbcnIp2bGsdkZM8Bpno3DlC6d2L0G6jXpp8cxVxDLzsOLzZ
dbEveqAnCFJnJuVkBsorOWxLEfjAzdQGUVuN7OCKZenldqq2Hhaik7QRu8+V7pk2eGHiENK6xNKn
4/00R/2dJy94kKWWKkBfu7OUP3FfMavcqKv2ry1G9qIZ7uzmA4wnpdo3h/SBbXuPUq2Vb7A8uaLf
mLAgPkbqTnOAUGtul0vX8m8acwXYMQTBAjmjPN31vq36rFyoibpGys/T38mTiBrOvfC6O0H7lMxR
Vql/ykLxCWZo9bkUamDqd/Bgmk5HnSw+dU6zor0XWYbP4YNdIUaVVrMqzClYf6xyV5ouj+tZ1VFb
JKZV0STVs8hIT8gvjGq+ui3TIZMsFYn86w2CZEvizCc+CFRi/cZ5Am377ibYMDM1Mvq+WdxbEGau
P/uRDQ7bK8Mlc1mAEPAD8CxARO9UJNv0eZvm7HMUzm3p/zye8iyXUWAbGNCnZC6zhz7GjevTiGga
CNjlnKSdxP0xas2KiT+iYYmFvRcLFJCQ8Q5qLrDmxnIZzXYa9oIqKibh0rL6n50wJi1Do7ukMu5i
TJAkdUBKKj56Tk53cQ9ET3z590MxgsVFT0/C8j9zWvBh/Pl/GEEopnmIOciS+KyAs8ZeSPLS2M1A
bteJ/b9TRNFGWa3VbwCuGSU+/yAeSj1sRWEvg1KXIRsh+nxZnPBxYDnU6o9RufP/WbZrQ0oaGv4L
IrRvGLRCoG+MrufC2mrrPvJkj7GKbWsDmzaJkdh5YI3ldbXUC5MudfMtK54GL/pVRz398/KGqU5H
bgmxc8c21Btyxt1jfsu/ddfy4cV9IgoABvf4RyNUuD2nCCJuWbCbQ4aPouRppsPs0XLjCqhEjdFP
04pbUOFva/kbk43FOAASqAxQIRjMF52vJMy+siImgNtyL5t5Daw65b7EwRdUjPHW8duNkMNQjTBf
ssB80/xDFHsBYorwGU7ANElaQeQBLA2rQfh1z4SBAAyAZ+ogXSfR5bRg+/EYV1JUQrjoJGJ7S//g
aa4WYSmtdvn6eWrEBn0rikVLJT8QRqd24dnJk4ZKJCjaN5AFel8r+ypXuNtDpPYMFsDHpJB/UGMy
XCrP2eR6duAkD0fSSfyq2bO2thdBUU/4QLqz+nR68Aa0CTLv7A90s9FpErDP7l4TvtT9pv1mq1Di
hrNF7mbTtrcVCGo5pl1c2eWfKppP0AEyb3/zxFrFLpXC235TRtVh+PeOagARdyAQUn3DhtYNjO+3
fL1Mr1R3HM1gKQHA1Cuj7ZUsKya0upjE2YaqtEtCd21MrlQcHobPqN61BvgNRUZc5dTjg8qJDd5T
QccczxqiXt2lmi1nktPezpbYZ5ACP0Ds/UsO79kZ6y5eJV6JisEsglOxmh6i4jBe+fZP8HO+Y0pi
eQudteftwuC7clyDFAEt8ZhPdkx9c2qAddjkw8UEcG2gqzJQdw+VmTGZNfzGM0rnLV2ZiggW2M74
F1XnQQmB7gMnN54X0Tdt110CeizgFA8ugzjszSGCiFKyihOB9/XwJPEY5HGQzScurHYJ/tA3bydi
SxWFJXnOHL6CWbfZUR7YUJ7XSSberSjVtIw2BC0IEDajefGgkAnFWI0jMXPagOuqAStpKIklNZJT
fcGBAO/ESdCr9hB7ykL6XaQiSfk8n3QYujLmokSGho1kInHGvyrYdBSPdjv0RZoBbSm8NN295IFu
/QlI05C+pMUHRALrYafbzQFnYzokrwUO4YuBUY7mtTZIOYpS96iqOqBsmP4vDmF8v29gwM3g6oUp
jUnRycr8vBFP64jiwbT+bGczgIaDpvV03fh0hWW+Wm8XbdfIxoY/6gPiakrtYjBX5uIhQEMvSgo+
sUTwLLouw5A2vLqYxuA91N8BQ9VN91GSgSCPdtNRbvQMTDQTVXaC2XCX3TuXJAqqkghhLPdxAs0T
bYuILwxyQe2fzU9jLC67aMf3CSmfnyfZWnzNAWhUM3zXpOgGVSNJYD64ZnkNej6edZBF1qXj0+V9
BXYTZy0skn7KfNWxhKDO6hqRpgS1746hqazKovtGZxO0muZkKxUZq+mpvpI1193THGdheXvw8gX3
bMUndh/vm784dFIhiIbgdSgaSqPfuAM8soiiusYnE5CqAcmKEQcarzVkQOqtdycbhr2VpBB53EJU
txMAfzB0BWm/eQQAYJwO7F8C7wVnajv6vhUPuaghShZiyERFePqunh52d0Xq+xCu2nbBFMTmoVZn
iK0urO7eLLpCPYyYaO4iRBVem6xM0DbQpgVJdAYH2IFS5rmE5d+MOvRlXkdTJ3NzOFUOkzZ8COa9
fE3Xndh6Duc1mLSCVCXAEWg6N301H1JhWsP92RKq7sZswecE35XZORX3YZrXPh+ssdS7wtfbUAX4
FXHAAS4netVHsBMSSsgbJ9zNKjtQq7Wkk6oqLGWMuqjkVZM+96Sk5f1Mxg1DHXf5f7ZioFE7F3Pq
mgdcJTLR4U/pgqWe6nzK7CvdPfEdXFO3b+P5PSvnX3f1j96fNMUGS+mEXZBGk0Y/fTHInUPM6cRr
X7rAwwBSHAcD07CaFK6NDlw+k4MxbsEnFIWMrOkedFqZarXMMqilxq6mLAdxid4IclvReo9T0QIQ
BKD4AjG1WkXBTVj+YODpjGvrCwt0NrHbC42sdaJjZ6xA2CPtknc6eKz+th3j5AtevmInCUmhg3qK
f1cev6te2kX4KAuKjMhvHDZjQJiSNeDlOzR9E3iq6q8i0ERIbORvrhLrxEPmpqoRuTn5H6QO2fy1
Q4ZacgaFRlQ4voEzBZDKUU2/oFawwRXBd1tPG96Ql1uL12uwJQwAF3neJVpmcovSjvaweTZGpSMe
+HCa4EtYZL0IhpVWLxyZXwDVbVMCK2Vh9bgk/lcuu6UaZWVm2ZJ/lVTlklneliKrSXGbvDnZjZ7H
BTLDvYMWQyB9WjE6+ZUUmvzROqscoFlL8k6iSbuTQ3Gbc3KdslPJAHcF+/LoXYnlxMBFj5rqwUIS
RmjIKv3z0hidz49YOu84pTpCHFTY7m6pWC4iTr3D5Gzkorj325AFY6lqdzjsd4JztFiD0f1aXlLk
NmNdyPIOuQvZzO0qFJRdGFG/oKHaFdNBh3MNGzngA420sBVPFR+qXXRWzVFhhE4+1X7Le/frYQ0a
ZORBD97yrOJrOhG0gMrjg7xQcc3fBsNnKsPO0ZFNg8wHB+rrF7B5UNa3CA3RNgNxOmh5pDELLZdY
GRkR/24g1uR4pT9mit5C4rDhzDdZ9uE4HYJvoTM4mInqVWWAsXmknuxmPqVbcX5nm7BEwuBVnzlM
fFzGemfzpNWcxJzRAqHB4zzDXD/MhN+MUQceFmyT7oZPQ3+/B10QtZeCmeNKEehXnDAjIYClLdZ/
ZxNxU7Q2muPaWdBpT8OAGxj/vPNskx6XQV6rD4rxMSSN1LLTMq+5+PTZ/5ZxT9SvP7bqNrwmnwlc
f8E2Y9EfgSTNNP2wHBLiXLtlAgG/m/Zc1fwS88sZ7+iOy20iUNpmUziaMl4eHLHdixav1qjSzroW
L35P5YvZvTh6ZecJUh4HscZRPthw3B1ikZ1YkgrZnG9Y5dtitcf7TOiQFNlIZ3210BKIhqAUpHx6
97ESaXeSY8IR4zq172/ADgBUg69waMZi2fNjovzMCy2gqc83TfUDqc8GaVkqNbYlg8NY5LhRuKq9
hhOCPKXmIVFLEqMckKN4B/3yFT7c2u8b0m1mZz0quLlk0iH+AJO0l9m1+qDmu0bTT3psgZGOJN8I
3M3Z/1q8sXWXHxdS7Oi79U25mobIf+C6PMBEhssrph/7NG9e7B3h9D5VcIlcaR8/ZaodTELKKRzw
auosyqkGv4HLUC8JFBWzuA6z9ctiIzNZhwDGeRYdM4hEFter48sVOHqBffGxbbVhMkHE/t26tkSr
g2rQiY4++3nMB/5FVgC3PrHHnwG20dH1/kFOwUqUO65K0yzMLZK98hER8u5hGDQNoLsMaK9o/4Ah
LUpfTJpxF+dIe7nTomsNAteFjp1+8JCYPHI+hTHuos8+AaXLNrzOtyw1B6/etaveQIC6EIPR4y8+
yk2aPHHPUc3yCJywXfM3FnUU33DmZPn3d/1YUtfGXH7iHLXyzI+wCvzNk46Je12Yaoav3ijCoty7
PQPVKu/W6zR2j2PXED7jAr0z7vvKT3rJNrby1a3rSz2c3Zhl6OnAR6FRd13FMbcHDxdE3wpSVoeu
OYhjuVZNLslIGPra83JZ7rfvTyqDyTLg7pvcN+Dg7wk/BDXa+yBpBwnuMHvpyOdCoSuO2R/oVhgp
cEYep3IYKc+zRN9m4eMXHdI2ufFV/rAFCe/j1YxqP/Et9SWWuevKuNL74BfundxhEMA3OBiXbDQT
8QmQmm9fjf3n6EgRlrTRHgPynfFdfFZCcIU4Waj567v180KVWIcvJMU9wfNWWF6b3nGAA4A5Yy7G
Ly57lkgn+OQTWwEK2dlojPURpH3EJlfi68SV7Um2WlQqInyBR53w/b7XKMcAcjXInZh7XAWwakHi
fIHsOhMbD7/kvSpgzAyoEytFvu7Er0g0zpUqYh8qhuJCqffw3IdZBXqDHJl6vcrtL9B5ixhkSj2r
CyD+4r8pGug2A/kU6Uwo4sqc23wBunUqemp3O6uo0BR9Q8s8SdZYpl8OWkt3JOQ3clVJQIFDMOX/
a7G5CiwkSmvfzNGGuyIw8vzE+D4dKEHIc5is573M+xWpzXYF0+yodv8E75opFqN7JtUA3vfFrCNo
TkVdnmmfGRzDWT5Mb9ZcKR0XMxWaFy96dOKmxltYKUzp43by+YYlKemqiueSMl4SUW+bFWZqgz53
q1mvPnQG+b70YtaLqchcQHBHJejnIV0MVsVHEik17I4c/Xt5bL6lC7lMsUpMUZ6h2DkFKbg3rt6X
DGhS1HUVj/xNenFegr9wMPYL2Y4FazO30OMf9wYK9IVh7Ia53TqAgH04ywhUEoNdjcKJyzc6UWal
xp7obBUamd3H4KHFLgs5pDmL2DLisvapMHXWHhwcixAKogv5snH4qlyLzag0mHoUsA/YoFUKAXAV
BFar4wpt+AuIihvo553D+wnj9hoIMEKCi4I840kGrvnj3AB9Q/mMPh3XKowua5MwhU2F7XKNMuSQ
NFqDLJDOyEvruOe74ZGGfIQFM3ih2cVA/02Sl/KhMtqi4gBSZ2QlI3AY08QjFCSZyJZQh1nfhlCz
pcRueWQ1fY5sX+RLE1SIKrQpxoi1CURf3W/WOfK+Vyik/1CgfiuRwF/QFe6RgoV5bkd5V0cDLFjD
8gcTrAtIGyhnj6lRXNRAMCjXlP8FstCH3tT5fBEZSSflOyDh6ewCiT5dbUKe7utRQnkH5ELB+yiM
QZsZjZU77cNA58HsiFfHJBySSS5WnfcHuIT2vERDbfheG8NmrCtJSElckmb6Tj9X7HzVsMYRTD/X
e/NCe2LwijoI/x9rvX7mBxqG5TYRit4jHMxwJ9BxsSV8nTSUGdGhnDZoQVZJVPjpXSIZBIDex/PZ
4up1Ufh07MMqRkW2gwoJfVkrF6Ev/dw0AgJZ3IchOSa3G+juQVwsgTygx2opFhQNol5YFe/HDPha
KxiSCUBlXysM2zAx5iW02CLtbAV6FjfAke5dmciXvk2V9Djso5wr1EoUVppQXb3f/N1he/hK2yBR
UdJzS0Ccnoebtte4GhhePymDC5fZJUXB+5slMBWtNUMBDKSJQObWJnqEUHptsDFRjqMrl1anmZWx
sSUQ/4OIGgUuE/d32gfEpb6aiAW1fFpi5i7WlwvhsVLgqPnHuQyG9eHLreOO120QJOMHYdDC60KM
v8+m9iNtFKb3DM5L7DR4vDlkjEzWZrBhD7UqbC772dpcPtktD9EvL33511DYm7XQMkgBF0rnxuG8
6Y09OJQLYoezjpy0u84L0TxA4pByR5shiPzHYmAW1qPvD8PT7hFnEqvbjcKfhKMO/DccPO1Dmzja
ugDWmcx0+hvfVcTTRmt4Dfa5lZs7/dtqy+WddNZvt1pSD+ifdQRAS4NgzmM1KgJrWF7Z0NWpb3Qm
DoRwY3UVB++sgZdzWP7hj6QPIVpPpAIAXiRg9DtaxxRMqOY6FmVSbWY2wUJXD4GfnM1mejGeeR6M
oKLf1VFRw1hkWlrNdqnhjRTO2FkgHvVocmfz0OM+sTTS+E0v0I0gBBS0zpYyGz9BOwj+KuF9G7qp
G4Jsd2qUsqbWPqZ+PhSV8+gafCAeBXvh0VC1zjwJrysPWLPh4XrjG7CmdoGJ+lG0e4mNQUFEMj67
ej8cMhRxMpCo+gFehIw1jtO1HDUe4qrBOM2B6Cb8fizNPSv2kBkwFBP0hLxd6bQG8D4meB87CS/m
9LZ+BI00PKOiEoOSB54z8BgBcmX1AyAM9750TV7xo5pYbFvLdRhMIZ8/a+xg8lCiOrQLmEM6LDoZ
I0BkKLaxGfobOlncPiWYjSTQcUEnKt9F2i6Vp12AeDjPvGE/rtXiyR06W887m5xL6CGQXXfNVKtZ
j0w0CTVrkmrjh0U7/riLd9CxtjhjmlbmdLv0EkBmKsSowpZE1HG5z9LVHZ6Rk36bVHXNOKhvD/SS
5Oj6rN8SnsfCleEsybGfbw6AbfKTQNuMZkB11wGiDEuLpSpv6W7zKf5aCiDKr0Gc9eigeXm93pXB
Bv+MmR6xlGnyKm6GaPkpFNqLVd4F3bS3OX2T6RtD2ErZfVXQ45kvvPYv0XRv7EMkqPCbAXhgclUi
DbBzzNFdV8alUaudhsTN7NNNPob/5TzWzhQV+2PVlrGOjSI6F8Pd7WUzuEvILotVnb7KxD7jlKGZ
+pC3DxKRrHTL+pK27W+Ilgp6oLmXy6uZi3uqfy5h+KQWrZe8E15FDVMAP7vJK20SQ4z/nvcjIqbE
mXEh7ddIJMOSemKxAZk59FsMk8/t6CPQKSIV4PGevxnv7W0/GsdCJLAcpaEi8cfGTfQEWep1esDk
HZ9/hjTuntYY/8R0pjUzegXDF/CF4zAgWWe+s9SMgJPYTYTeg6BXZUZl+eVgHtKFx0ke4dSyN2bK
JXkmy13UYFk4AWbpvnybpXmTnS0mHPT3djWq/8uTcnJcvjTJN0oBmMkSXzj1msPdoAxo1cHiTpBD
fBcPrQZIF1vwGmNqp+20a/8utcBwcEQhKPVpKKl9LFrJmvZd6jzc/sI1oC0HEAi/UkaZprFPYChJ
kXo/anhuVP1Y+m0bA5Nv3T2Mz7xH97a5U5X8DlkJPPdBditbmkSFiFO9aWqHV1u83GRIIEatcxk1
XJrh9fArdAILMlDcbQuenmngBwuh6sU8tFgrR4kvvsNJty4GRtVd3nseGwce9lKpj+l5G/Y5Ezf8
TrAwqeeXsnsviuGWAnTuLKGMYVpwR2ws9VeW7o2vy/KHTg8IogqQ/kkiA1Kdlb/m5sO0IwIJ0WSC
/BT2TpD2jJ6+K/E9WOeM/e+n3YA3x1B4H/YPLAr72LojEzGbr2ojND9PdVVa1jn7Vw6fajfuqF5m
3+T8cf4mXpAjy6xcqFSESdpSDhRC26cNpxhdNeoLFQhdLcKdB5Bqr7wK+ba2I/N3tO3gvbspiwty
9i0Kl3CJzT+pQWPv/YnvsggOypsI2dj3XW1Rvshx7dFQ4jAN/yI83E8E0BVSDZ9+5Zh8loGLtw6M
O5PXbtMLqppuBslwys8Rm0CoSee8dEmF0aDWIPXc3Dj9CmW+PuUn2DBTuoo5sOAIKsKwaq4g+6KL
6ObY5pGFB4P2hvaraFDUG/QD4kGVpSJHaoFBAFEIrMpLJc3rH34zGHmiqA5p9igNBfTX/79+I5h5
5KFNut1JQuQEM60EFmEw/fzEw7DrpqjnWrnHq4uP749nxiIqhtucfuGr1p4TSfW/LHKzBZ2nOI80
nTHLhVpYl8JYnBBPlnO1zO0JOE4qlbIbSWZzIcE5yYlyQTuG64f89Zs2t+P4/D/Ct9i00twDfU3f
jWIjkImR+LHSo61ko2k2wxv68/+FNY+AoenuT+9D44T/izoJVWFeE76YqKteD44RcKqrUQO6u00A
sRkY9VdjQHPpW8Pz125SVa/hLE6Ik9DybILOir+dvP0aSTt0+2zTPI1zh3fXok+SnzPzkyC/9mee
iYYYiveed7Bf4CgGTpieJPiRRLOu7faUVBKl9Em3AV7v2ihlY21SFQGQ9RWUQmATHv4AdMpNrCEk
K31iWaE9zxWf08tQZoo6gpblvN+WEveKWZuHHMsyaCOxsLUl1NXdo4S/YK85mPKeGAEUixdXKFns
yDgfpnXFayorOYy+FtrregY0KEpi2eK3nX3pPmqY66C8PV+5lClbJ40L4xu7n8ofRK9SrtZzGSiz
GRVGfJATQbLWPxhmfW0MPqfU74d7TysvMspaSOm56NjliAy1JQh0v5jf3z3HZI3v290rolqSSQSi
k3OI34UsfRJjtLadvr0DxCveSsC9P7JYE8dlFoOhSFErH7ohHoid0OU+AAfs0o5uZRUGeEo5lFFd
OhSDD4o6NLZecyAuKJr+y16hCjuutjgVGDbFcRK74ufl88U/9E3qeSHLbluhRW9g3zPID3Gb9LUa
x4xo/in5JH1VpjT2Qe3EEI+e6RhNtkhW4gMvME4K8GN4osfBgD8ntyw5mj16Z9wID42or8EB0yZr
LQpCo6tRR7T1VGDFMwWx786bNb8NDXX9nFMdWKKKUxdmuV8dxER2HYDg6AFhYM8BiV05RXUGDIOH
I2MJlnwnUtrlFqnjeRbCcgu6tPMvtJcBa50Kp5cdZaZpegoAUik/sAZoCQZrPIcYsx2leWMBSRIL
JvTAW6eLIBln5KC7cWfX8zqn+h5EsPisAd6pw2Ni6WDaXN3yygsS+4hyKDz6x244gh5Zbse3CBHX
SwZuHMLyzC8RsKdFJ9qwAWDiks/sh36Vt8UnMgTxkGuxWVNigYtwItaG6vleBSpcNmU8d2/8grRJ
GlSOHd896+PGVj9qEVILkjOu5K6XOOeojzA00dmL9fc4iyX103e5UHEkpSun3XSAM4Wa9sA7Ud20
W+C6/IgRJR9RAijO/LjoIvFqgKS2oWOt1IuEoTWqgjNyq1bc8YNpx6YvoIL6NcgX9J5m50/xpoU7
Gve+vTENAmr6gyy0fF1AW+IaRgFavDyoW5Pqs3BGL+0OBvHLv8XawDTYBqF/zk++d1tqzwwf47rQ
ZDU3fMBBo3fVVonVl5oN0denfOj+zswNmwtRQb1gf/qzbwbmTRr1fx12YgMEdZiMpsjCL/imueSZ
pu+VDvWyJ7oKr8mf4vMoggVIHY8ivy9wqOpWS/FXN21mcHuNXBRlqaeZzEMgl315iR5/0NaknkHh
bvXyjiMTfkwFTNg6PFf2rGlqv/c08geM1W/p0b89PmLGcTrNcaFWcbmzP8y7AXuEJcbB7dVRHJUn
AUicjb9pvMBwYOaWDgqxPuNDgxsv8vNBprmrazlBuw3wd5+tno8nJj/SvzJFPKNUkigiTh27d3Xk
jNxBNkUxqoEO7ZhRDdBMPvNnw+QgyqhBYrq9INeobX/2SGCoyEBcjcAkPZZTcBLxFdHGisTZpmrd
NP6GJqxvamsKksKALWBQWTHvnuoT53gmENn38DHE9BNCDU3qrigtVkLKG2izIe9IC1vJwRhJEM7K
MOgLTJOfMtYZdZZKv/WxOeF+G89Qm91+UkAe7Wb7Sc3LgATysbvdDpX1fkabZtKBEVFbxo/tqg9v
caEatR9dm0IWw5NCfMN58V6zDKLcir+U+5xyu7Q5Mb3TQguqJm8K/KEGIM5Xqlrx6IvtcHW52H7k
Vc5MhG28bq+koC7dJ2udfLSzqjeMAw0knxbPDaCPZMzJrEJA7wuP1wpfFRKZW0KSrh0jgIRhcSpZ
8eVz8LR3zkSNXilUYh0icFOEwjwCNDsqmP1NEOLBPOjcz14YklK2tneSVs8nrvgI/KVu1Wyk9s/x
STWTdls7svVUMbQkTeCeyFzj541Y0QxNHNyIB+f0f57DpF9cAabqXoHhgf71hD+x9n9uOSb1lPpM
MV5aG0Cr7FLUgsAZxR2qD5yBcibULylhgcRMg/Ue1JRINLwD6rCHtEINdd33GVZe6R6JLwVn3prR
pM9CawsrHuaEYhKvUNp/raXi/fv/EfwevPoE0U+J9jVEJkUX5yHUaPimt2gEo81GsSNMcoJAhURA
PNloHn1G2ubCFD3jNCdc+VegaYCfQdB6c/uwyvsHvdsGzYEuh1DJNQOACfbrNRpxtXJ/IEezUU2c
r9mJIegtPioOd2iP6bT8kOX7oCLSZPGwIgPq4EO/OhyU8n7E9pqgGd/XjqT7pSqZSPO5duzVIpKc
XpkDiAB3mlnuNotTDNmdyq6zMxHmbEJzWLS1AlBz+IzmhWgtq6O8zTtsaQeCz+SbMAMiIjWt4Wpc
2oO9xpy0qEYNc/BKZRFpo5RM8e0L/d4i5WBUn9nHlRiBCXelBjBxEuLlr/89n2eEBjDZYHsLKSKU
Nr1uDLzKWwJyacykCvT5Q6UkfLk2GLWCN8/CCKOi0+bGorJGkQKqttclHgzBoTUC8a6B9zxtcu83
o5CKPx3apOr6gNmndLGwv8ARn7NF8oFJCzi8Jf6bbdZ1GMtjDq9fdG9kWa4sduwCLfBMZUEofSzR
2pxvkW75YrUKIgru+ERgVoa32aI2p0UUrYdPwjUIGT+cN+q4izE+DOpwSBZNrtKE8+lFw73szlqp
ntSofz1taJ3Zp/9UzIe+g5XxQKjmV1auCr4ZEaCkv91+I8imbF/G27fxnYDtfkoySt9OaNj4EVL4
6jo0mjU2es1kEvwcOJ38/haecBaO38GGqrfLyPP/BU6eN198vhF4bj62BafZZQ/fKANlfJnVgV+v
vzuBgvDnohnb5fkedqk7JfhZy4+rgyxp+Ad+exby3VbxzRA1Or8L/tykC71Z7YsVxG35lIZaMhwt
LS52rJ/W0LVj/VeHG0mnyCQiY04xwde0d7mXwApLGOn1j7oJA/t//yzcYjpPMFmOUKv83k58mIvD
WUtskptC+11ODfIYAPng/qmNMFHT69hkvw5rVgZRr3Xhfeb0s+lf+tBOZ3gysHEYJOBQAzKuMIZ0
FEIEqM7Mex+kghtajK0QfwmBeE2hctlCHD5V8Xjhj61dz7wpYvZMT067Wk3D1H80BixwuQNtjOsV
hAhSSnuF2ExeMf1IGWik68AsWXJp6uhmHwylcXUsa3vPGZ1z18f2Sa0LC59ygHn+2IhoZGlExqr0
HXVTNK+d2ZhZsiwtmaqTMvKGKl1NkrU2Yhj4wT4Fe1CaiM9elWe9jHhE4mCQKZhQ03jNi/SjPh1z
X4EEVFlNvBHEY13NI57ivuos6OXi5J+cdtfebNIU7S9HwbeGPqum/iThaFv2wKKbUzAc+mTb3+NR
tq9QIMtQtkFaqU++JP6bgBNA5m8ACrlC8NhBXQ3nDe7f/RmzhN/TeEd/hE8pbJ1cVt/FFdFFxaPo
LX+LAgMygc8gfGyFGY3vrHoKMSNQDgBdKKdALWiSxUi0kLLe6+Rfq1yf4XDLLRvnbpBDPQ+Ibgvb
irVBuKkJHeHm+Rjfuxrw9TuQjpdY1ngg9kQuWGFqqQYJtQguNAC5eHDMdydGJ4arXspl6abXQgEJ
pzUoMImluVCBtFpJ/Vzg8gDrjfUm8O2OeqXzcOctdD7BOVtZwvDW42mh9Gd7c77J7gdLko8FJ2Wy
NhI4QHZV8SRRDqRfXdoijTrFxNN3TXJoyE+2pUTGHyJCFPB/iFlYRNnR1nnoz0C56iMyqVB2t12M
WaswaE2nhlxNrXI7Llpc4rsYYcl+HqWhpk+AYq2nUFQ4PRDRPOIcodp2j8DurTRiFhyyFQptzZed
ILFyNGjnF7Gys3rpIDSjsdX9I1ONGIbsPuIQG62DyVlpnPxrkM6wh/mQv6+amCIf/BwbQJiSVal/
vWNiBuROmrAiJo27h2o7ORgy4PgvCpWMA3VHXOJ2AS4+BMVd9GJTjWVV8d2rm1UKUIZGfV2VO71d
dfy+wXtepHkuYDjruJ2WEvvZgcc7qcfz2rDeYEb85A5EG9pCXFeAgENWFtPagAVVYjU6j8FQsIpg
LYaVkZH9NtQInOttN/eU/z69QZIRtEg1CLohi0+7iWooHB1kk1cOAhOEM2fQ2POeyz7EAN8l1Tpk
/T6a6MbZ2Z/edES24Ou+ZEI4Qf1e+UmCwSPsnOQVA7xOR2RNXarfyXHNIrLcdp4P91LEdkaEtJJA
v0nRpXNZRGrzFiEbtJQPzD/S/uULteIEJIbDWFdBfc2oBJhDV2txUUTRTc5LPrcc68NQhiB6Hcas
g9hC92uQHZ2pCYY6Jtx8xUzQDtuTgE4wS+EXU5KVwsmkds88KOFOiRF+lR1UOnZtMiwRPb77rr8F
JU/4tPSv4xy+Y+xU/YTmgsQqcf75zImzVUsQRhKVTlmWNyLN6QvzDune3jImzrGQpfwA7ChAWwhl
8/aRQeyT/DdaxmUrunxN0vsFNQHDLlBamXQ4zFY0zZuAfYNEnfY4Lcykw9C3bILVeTrY5CkPaiWM
YjW0WDmAncR5WIh0iGuJSrPm10det/ny5qnTuBoXxxUapi9R0ZxcmP8OJM0lAxiarEK8Q8eItgeS
zSCPfnTv/WxupKtrBzcwB+zEgVbCSnTvSVs4KjneLyYinXSFlXuY37yk4vYf46RStjVIfmMNaGlo
We6OLCHMIVIIdtaU2R/6ZSNRCZvOmRTNg3AkrbneibI6owsV2nAOc/oM2cYyagphW6DOyuhM7dIq
P+sp9c51t518Yz0nWEZAUFw8K6hIa1DAzDf6id27D5iBkp4Ct/M9Url5SdJnDWznzJWFHIweltov
Z7btT7atL9vHWTSjY+7czMhBBkXCeEX55mOZQv5NDDsbjbsSacNlyaFkP4o7A8pT9xj6q6ciGS9p
KXx2eHvCfrFB1zeGLNgcfNbCrqb583TtN+9FZlH/unlQMWtJhy2M50SThwjePgivK5O7cs0ay4KW
hvGFfM0t/atNRf6to8Fms5JL80dSYEwL0sBIXDerT8CS2ERw6r2Uf3opoIhkl/GY008WBnl5R/YU
eBgyJjTju7p489z3XTxJr8+knzWF9xmxRVlI0V2vVzBYLdKLFohiD3vPfITHd4BaWm2KfIc2+6uA
HRCDZ+SHJ4bB4W4kABgD775ISk9ll/A6NzximOMSnqPb0Jn3M6qeH1tjM5agBSsplp8Eqe1m9uMH
GELDeVUJu5B6AyitSohHkD78Ks7BQJ3acjtPjcH+2ejMikpbX7BJnvU4KHHxAaY1KVtCQLfqTs9W
V2b9rnJPse4GqbSiUocNqKnC8dpAiGWmhXezfI0kX0MxjVRr+n5l6A/c1uCA1muCI1JWabCtNHGJ
NzNAoYnoglWQfUYzlZ+QXOrQdbxT/TXY0LhJKOcuYFq1G323HnaeXfFlBJ3VIo62HbLRW4h+zIVD
4BW097cSTmI9ulGCR1q4ZPIhyUERT5DO82LUuuiZOFZm+Td6htxkbmAB78TOVMZ9a6o+TLE+DQED
h9FpG5zM9rOn2B+SjbTnSoUetmR8GzKQNXm2AqnZfaIb9boXxBuKsQxYI+dKwceexqd9VatAyeOw
ojgkbZ8e6J/tTqz1vj2EbMkSdmJifRKxOPazRKjqw0n3/jlNgRs+pEiyUIK4uKJCZYKollAlS6EV
EgLJCiszUvaTawF/h4ggsDL7dulKk5m//iz5sNnIgfqDL9ZEQeiyog+i9s383QD7PkKVjNDa+45q
ClxTFmGTCXeOGoixbSzVebmg6X4nIOPi8KiiHXueTrXiOElyUnDb8wdoUtH0cOZdDV6BBw5mN0HZ
S0fr8wV4EyWf+kXdvm6LS4g6+s/iR5lBhQfmDMd2k7mHz4NsAO4xN8v+DVdKZS9ygs2Y+AH6aPEd
4bz8KT8a11+tgYS7cLdATdZRycVP2itucz246+5n4dNxa7gpw8i4oMWvG24ya1IgDv+pkBHFPXvn
YRqu9EEPMhiD4uw4c7du4phOTooAS8cqW6BU7rfWdr/FYBsz/iJy8x8XxGbu0odeE8nx78ToLJHT
IeISNTuvaksVemvAIOT7zwyokPjEfSvsA+0be9xzpJjsLbtnd5aT7PRq0sVgdr7F6a1r9smzjN9I
OzL1bEtMkY0kj7/wgD5o3RihEqGufeDBg/4zyQ/a7wnMh9++vo/zDuXChnf2PbMo1xK3gqRDSJoK
rWGrYvGWeXllO8sBKy4yZ4SiB0xLYmpmeKJ3tW3GYIi87vR1YASTLuxgYUjceJr2jeaBhcefhdBX
bXwlFdyD/Eik+Pqj0NSEVMGzrGL9MkmQCjmWr3OQ0cnWwnsXSuKbQNZtm6Tw948dMpCAYwm++cZP
VSLynXc56V+g+t8Vt9KvdyaAaAwF1jSmkOSPZ68psc0Yos7lquSPHzybb1t5Kcoz6Y9+aFjb0M8M
uNgp98frwnHrS6XRpp8QpFlnv3nAo93ET0uMsYCh9IYBB7E5Ag8EXrO030I8i0e50Gvbm/zBDmGE
geX75GIJhop3hl/emfZRffOatpeAaYpxwkRSB1t5+qog47qzQ49k0FctpnJCvV4alBwZLyGUG4fq
mWCCJwSXz6VZNwD6r2wsFPjiUd6MlqjI4lD+7sSGQ5n8gFqItEAhhxNZk8Xh+RkpYfvwF7Rv19wZ
p+zEMGWyI8pUzSbHvVATIbUNbgh8AIyw16E8u6yCEK29HPUN8XsynBWOY/CvUVEdy8Xii5JsCisk
jwbvXmHdM+u8ii2/2HfhRyfcwctOx3DNW0ETlgBo/PSdINLFUBympFw6KlKnzscN4yLNC6Rn/zJ0
bb5RtWxsjud3klpKcNJE4W4oZe06NmvIZ5gHj5FCS/MjCD1AcC6vTg6oo5Xokashx9K2NaGkRvX5
HZ6X3xC7WqAQdhoOEZi6vz1OnnMjjJ6PlHCMw2AK4IjXt3eomeUOcggN41mW0Zq4YjZ97I0AwDyJ
PfAGREnyB+PbG2Srr3K19sCuwZ8jd2EH7QXWykkx23rKRWv3Dh/TgN9ZhHQV2wzet7JPEkyNZa2d
t6BXOQj9TqE15PwZG5k78cdrpatbYfDXqZ+uibtJSyHoNi+A+NYACnMGe2qujmMhoSW5slaWG4Nt
bubqT/bAkJI0GZgYl2nS8DxiJILmR2LMJlA5PJawEkmf0YpsCYj5+IN8tFG+hp3gZhMm/z6Z6PGa
n2d8dKY3gBvaHc1LNbI4vd0G2hdjXJXeBjYnfRQlfkgbYMQCaRMlQa9Had0e4VbGvdBb+tFhVuq6
nTKll2CQ1PxZMNrrJz8ecRYP6SyNGRsQZ8hvZKRrAkPnqC6WAOjthsYwviBcQ4VDpAIqml3ywGlQ
tW100AsR2niB3FprU7Mdj/DCW5Vzatb0+eILycF7npK/QmTvAvQktfCCMEbkcEumJ03s+5xvGpSB
A4hyB1+g2dPAgSHgz/48HDNT/NvVxM1nxKdg74jODZ3EX2RwMB55xHCyV5RqVZ31c2c+Kp1eLAFU
Z8tV/lErArgNZN9zlS4dXxZBMqPIv0YtCUAbhhgnQ6dLAbKNMchdIAbJscXMuDYOus9UW2y4AOxR
ir60/R1ivHGhLSutHey1txhC4hV25ZkbOLT99Ofzk91HQQ1wPBY6otfUXcjFDYg4P8lMz8+xWp+P
+9BMRIxhmXfVyH9uyao+99J5+m3aQ+/aXQ9piRDp6Xsd5XHt46kqxgYrbPgucGY1+97a2u2rDHPo
qGf3gb3ZV9XLYvVLvAqaQzFA4SCzSblS9S8WIKY36zqQAQiT9PMtXBNUzSwqmqN+stScGO5dnz1r
N02a6OTq6I0yTckOZ8cj+pIYGmEhVTEc78VEoezNaDmjJKopSAbigummOivEvvH93cOZbe5BPu1l
ZS+TPK0/es5cDDXvsgob3usZoTHvWpYbSDe/mjbFevzSvFaqhp4pIQ5RRGdU9oarxmHovWgAJytH
ole8qtuQlnVA/5BHO1h9NLmhJb7GGeVJylH02vJPrcNX99oBR3GdMVYPWAXY5dFfYNQXUlP2GSUX
Ya9g1PdFxvTxilTq6Y0l0DeHGzTlLU2d1Y1sRspA/krIwELMJDUb84kq6KVxA61e5fvJfrRWPcdw
dF2NA7B7/2Huh55CSwo6cCmo6WqSz55SRfIibInIBPpVeWuD25ir4VR+ctAUZi/OiG4446U0hFou
iKVHr2qLQfjG1acuvDKFpQTRtZeV9fRJDMKFIbHGGXUGn397b6oWr6GNpSQ2H0m0BJbaTVdwcUc1
hdE4BZapxJF+tWLwfaslRj3sahF7fLdNbl6yuuWNzGqJK1Ssn9SwmZpo9XI79MBfbyk9OMApwP72
8fgK2PAspTiEKj+Odq3o4q27Kz+gcHbGyoQstvmOKSt1bHB9zOzs03oy6/hfGszo5RG0c25ZJBlf
pzobqetisyFcT7uTcOSqpIie9JVb52oeFHXPRLxs4bLVqgNnVs5C0ZdyF4Ra4f2KHNc10X+DTQQV
+tmTQki0BDo0ilvRPxYX76J7ljbISiRtahHaR8K+sHiUmR63/gHgU2QJfeHAQQ9v7bEOMwMTaGDf
jUPt6K0r9rtJResa4MycMVT/rH6CCqgYbLddjUgxFxTvm5aoMapBsZAgZCYvcdvkSdC2WpWTlyJR
dBOQHCxlBhkhwshvl/+mk2nDFrnlu6jAi3xo5DP4KYEwSuifiqrgkp4/+SqffEePNuCL0TJiB6U1
gUunPQPFA/OkP3pYaolpAmfrSJNqVGM7gxP4Ov7dAXKx9WdOlgfm+I6oveWJWeD/+2hblYW1k2pK
WXBS4RYKRgnZ16HkwsOrgBmfNsioGPikK12+cSlUw9hCIvrWufq/tgXF5qyUq6pY/4X9gdPGucTn
rsVh6MS87HmZXUzKLuo88TQiGiiDuRFPw6TShK+N+G8/WjB/u0PmRelVkcrHSHBJ1sRO3kL/yjPe
O96j2mkgOokICm4eKDL0RKosO5TVdYrJ/Yv6TYXTViJsoCWfc/Gq43M/JZKiANdtO7HsWRALHbaK
wv+PWqUwwXAdgt32ej70Y6CSngUZBeQNlit4gD1ESbF6GUrG60/eqI5wDHrMy4U+U3Pyl7wASnEq
wzUqj6yoBq0h69CgNB5BaligkufWaUJM+PzOjgZf6OQb8j4KysmHOVefthRCD2B2/W9QfLG9Qcpw
XFU+aHNgSrrRtCyjW40SUoZIo6qUIezdfADiBn3wz6c5YYPBsTtvd2o2Omhhoz2R7mI0aY4GTjlX
P/RWqsY0FflgB6HNOumkooTsdYmXP/ySfamog1ovMe9UEGYMGfLD2d068JZlvvIDYEez6LbRwWoB
ASHdgW6V7dMUKA/9XpZOIV5JH28Fc6GEv0fOojdInTuHrLBDBXF2j6UgWRgp4y5p5fGBJWO+MLCX
XciqVmXnAZ+N/gUY99YFyS+Q5zAlgHGa4XTqL78Iixhb/pnpzDygKH6xkmn0cgzBhdm/DPbm6OaN
W01/yIK2mSc44QAFKx4er7VomnC26B/11363bCjdweZCe0NUTj0B9sWtC6F+y+OJAsDQOITtovUc
xWHZCwxHewkuM+klSr4BMAFkDne44qVNeGtSBzS9mBBuXRV302ha4PVz/HMQc9xsyg2hX6TCmToU
D570MYJc+OxJ2Y8LYD6mqguopEuMPCJosT0xS6nDNr5a7hvceeDvENQ+VxwaDXWungzlSA+vDpej
Z0qJp3G9OCrvsqp/3fzqsjmQK3OsZNqhrSpq0vDGE6XWNKJOrGi2g/Tqmj9T2atRvrLKmc/q3OBH
Vwoh/rhGQF9fjn+W3W59HYVktK/tBK5A6Qu0qMEXuRd+mUQJ07P/729MW9aBxbuB9i825k4i8TT2
pSN3kCOr3IzVFYJfJCDtjFeuHXJtpgNhKaQRSIK/neP9+1nicbxG3Bj74nAUoe8OlcM9yd2zvY8G
E5b143i8wEwI2g7ZrsRRQTsNWykK9PmTy5fo7VDlg8q8y3F0w0V9tG2jl6CjUhiOxmnQPxvvNiFw
DO92+xB+PCS1+f6redqjFfQlrSoXUBknaSXpABUqOxgHbYiBPCF2mbjWnZKBGRJvMIDgOGmdanLN
FhRBgqOwmA9xcH++ivgH33CqIkHGYSNfzfdDy0cjgkL/ZZCG5LMP3l5fByhGuhDwzRQOny+4Viee
XMG9fEAhipcj2Al0TguoPnguDwasczlk5qNvaaPk4HXHp0z3B2VMqqEiMMOiZzVyaO/JGUF65QVo
ndh30GIK/ZVTjcoS9Hp9RrIbdwhp62TP+6vg3zovKOAFGCx27wsk/xrufcgZjd2q3ocXUw3huiVS
RLzqz1GpojErwFOTXZ9wDAAkTiEuOU/YUfc11EYr9aP4vguwahuC/FyPhUXbn9r3+UPEjCsbyMG/
tDilE9cvfjwX2izKZNo0WAPxtDoqCt79rnUBdkkmuOAdJb1IuHubMpJRrSgJJu68U0UummTkSvwy
xWPiFHPMBq88+guX8nxGqu5GZP+fMkBAs+YGN3il5vLytDc7L/bifbonOKxdWGIlvLohiUY8uI41
fvySfAYfKXmEHgGm/Ni/6SE933esv1VBEPXduuS5WaeHY8JFJCBYwLwHf8+DkdseWiAGcUXQA6fC
wMboO/Rccwncv4DFi9yD4FpjjLwOBQ6r49VO05cbyCAf6EVujgtDhhVnPjSPJ4/xwgG39m5u9IfK
sz8Ql/eX1Fw8CFUvCO86H4n5kyywVaeHWRkeDmiFFAayN35TKug8C1pX4Ka3D8NvQR7suMDlEDr8
wR7sszvQmffxyKJwoMPe8dWFCMovMwqmGeMK18DqLczcUyvFz56CX/rUvbvAXd4HiGYdZpDgNPsW
RVyXAJf/fqJr2A07O4AkvOaZdqQjS8Docq0yUD65v7muzDyXzPjLhfnbdQTAO3oQcTF+Cafa4nlm
M1cZtLnlCxxGrK/7eyKlMeACVlWsmM7m9FBeLMQJe4IwVyAQxuReQkZFZZTJbAvB3FhqgoHL9vh6
QT0J+apkFMPg1COOowWmWbOflKEhNhHNP+tzvYu6SszxKR/4JDHfTBxP2wMWEIf5IM9xqlw9qfEF
54lFybhDoeKXo/31j9HL5de1fNSqfxZ9LvimKQhviRHdb0kI9RGZ6Xs7AVbRq/i7mY+kk17dIpMC
v3M9cv5ieZHTm0qeQ4+v0YVJN3rYHmaC/UNl0yzk3c4fTOF5lihLqrn8jDhzp69QJAcnLfh2TXkt
qQO6CAw5DRbGOUP6zsnTHLoOq7n60wVaOh31JotevD51BvR9WTltRjEVCf9fcAYfHe7fn8b/Fvpf
FQxguoC2oluKBe+NORxRARc17oxrZvFa8hNYkWKUjnWPae53eqbO89GocujVHscgBBVsw3BsNoCG
j0z5GegXHwh7ZUzz9wN5AM21gocedslRI7pcgfShH9Q/8c1ObpMZrufdmyVQV+4K4ArG5Q7K+8Ck
PCkPlnW/aP7ArihIePWNg4AM4s/OrhCnvVyL6SMLDuO44NTPjKCdMdskFLQQvSpcnUhxUKac+W83
mfy5zhVtov4w7Bakm4zp3OQW49/nPl9mmGjfeXIXQOC/NezLLQp8S/cyiL0CJcSRcP/mPfXHV1gr
PN3zqkagQOOnXszbGioTP6DpJULYM9zUMTpLt+UGS8u+GjATTBhDw3zfWbkB+RMY+KZI6UINBF7z
2EZyseqdxvFV376CLMApwpBiDIaXF2Rfs9+7zbAjaSyYcDT7fq42HyJThpW2DKmsFtVlJ4cZyqF2
70NcpdvU1mwBi/LnL8aCJDYFS86idMkLVWVme033niO5bZOtAREXRcse+cxBy4ExYE44/FIicjbF
E4j3zTD1QLDfqTx5eM1/pF75wMZOIEFeRiT+S3lI/Z6H7no2BygXOn4BoMpmlnaVT0F/LEgp+91N
wxunq4KaKu1IHvSGFsGL0HU5wUzYXvjuKkfKK1zN+ARem9cWIw6/B8i+Fk3GcfGV9o43hfVj/zvE
wCT+bRLoSzADjEjZTUW98sxiVA6x8Dy1ljU/Sk7UyDrMqzRZNuil7HEdHS+vmho+lOaw2Vw+vFmS
gbVLofhbYlb3aNnxOvGOvL28TD8gBfMv0pl6NnYaJ9gU4Nwo+bQGQCkJuoYqcCxU0xfVbS3EbjFr
xVc2kla4X7+kiHRa8dSpO6xP+FvxaEULN4kB21VKL473FHudKoPGX0oee1g0eeH4mtd+Uv4MDpMe
TA1Yn6EYX5WnM3TTxrMfubvUQyxACPhzhz9+2D9k0nO8d/6LqEMREMdC3bjnJaduOl69ofPXwQxZ
VcHYmDPepCrkV0jQ87d58obIYjVSCz79hkHyoXpbkbiW/j8DPzv43pFGcYbSZEYi92JXBIMbEszi
exrMGjbNgnjTwE+Ind3Jdw5Hpb45Ospjp7XT/arZtTXtUhj9IK+EneQb4P97g/rx7Q/gswd49oxi
zm85mDn0RTbCeF5BxQhDhPXBXcaIRk88CAfGaoZhN4wFeCRjiYTyZaU/g6n9oO2xIqw7+ZpfIemB
SPL9dQ+rEfBRKMd3PISJvu9iDTVH3fPEwqR2KUMhmRPvE84lbzSSZSjurthoyPILwBdyWOWipgLZ
eUtIB3/InI5uSjEE4Zm8sDDILzmznyQGAgs6yXGZZivODUfKZBzhxaTBEiLSaZch9LMxwr4wUaJU
TkA+1CBSpDdpYPX/YspIfKwcBYSZsIp8ODvLF2oxETwRr3T70S5X8o25/0R9mnaa6/EQw3Gb29f7
S0lcQiNUA2QB/hxmF/ZZlH1r13n8lgun8vk3FOCbPpTGZRvBgJClsFdDx1j/x69LQIbJHRgGPC32
jkMVWE8eQkHUSW2kpsS5ghOTVxMKcZMUxBI9wyJKJ76LSCcg6WyL0LtCBknxLRUg9YKzh7pSMPbv
lnWjnh0a/Fa36llWLF0ztpYwU9GedaGuO1P5EtLvGAT8QoNqlRx8tQKWwk45e0gGf25KyRVfQU+t
NpQWx47Kd2KepcWy0a8u4w+LwZpF+Iy9g7paVtYju7PrjLn3wsrWbDv9fpOITcBX8mhl8NtM7B45
qa4IZ480z6lE1wLb5cwvreZxFoKSV482BglbJpjJWHUxRCLzeqScu0hFWq5k+w3kyWEn+bql/qYZ
zvOr02+b4m+xMGPK7QK5Oj85KuTuLhurjPytgNfxjk4GsY5k3gSVmHn6GXqfIKZHibwyyr1itNxa
1FoDra9GGtTjBmaStezDP1Y7bKlv4g4z/D5tDLJoTJEX1bozdnA+mL0PUgjKYTr1ZA5BPdVoPJAQ
wMg/gbb2CaRf1J71jHgdXOmQmV3ZLN7G7DOJmpF0uyK8MS58QJmBA+peWiVnqEIsYc0/ULtHyJnD
kk1gbBzi6waNwP0glW3SNRtekjhjEZCkcy1OTouYH+q4luqP75Bm7/ZEhVTdJkiNTR+Qg+AsABG6
ev+iC6xj7/Pa/+iEl1Vk37uYxnXLm9TitedoWYWshJ/Zy5CY9fHYRQohCLGxuaeHnZp8AKIm7SqO
VTHc7S9bGhVeWj+Hx1KIEYPhv7nDBIHFYixywXoepPfw8hgeMtki9Ixtr1yWqraA/H3XGaJ0F7Bl
4oh647gIlnpT6ZHaY7opK48yK9ERFsfAcrnH0Hinkl/CzDaKnu0yMuNWk+A+bx2RgMupKuyfOwBZ
CyrUVrX5QmSgwTiLPJsKxCP5x4ZjFfW3torGq/FBjXpViiSKkeEtYX4aNs6ERxqE6xn8zO8Rguwi
jsRwePYmLa0t2gTQzG0RYstTJ3Yjx7jDcl+jaoRrVvhxsBqV5FAhg8i7nWEOwbuOmlLUGsMh2doV
QY5mR6H1AtiSQRqm/DmLGHLowFZLH67y3CTDdslamDGZKdBfSe6Y+JWMe5x0yuCzakBz6fCjaqcZ
74wOfo34qbFMyXU+XpYgO/SMNEfi0x/6CcOups44AVCib+mbzS5mhvPJg9JciK+z+hdpQBey3hfm
z3vHUMWqmc4O2Y1MvnlmtAI03Tb5zUjFOJY6UyLMLclITYQ3y+2Yv16z1nRCOslGdKhvQgOUJGg8
K7MdgtbbisK3zxFULpuqjSwQOdGhXyp8d5fvnugnD3cQRmbFkoKkYqfR4BP6jzRHpg5PVCjNbfTk
ueWJQOiY/E/kICkk8P3pRHxOkHVTegSxFWewo133ZdpI8rt2fqoabXeR3ylWTV98QJlorxvCfUuW
zX5bN7FMtkAjqTsmWLlvD0plROQMTlU3Zx2xZDpRxRaRlA0CU0/3p0n7VbCx/nlIJ5Mo7LoWOza8
PIpcHTdsbdMbQXsLgIX9ONyJV52Fb6p6LDwv19ohHCSO/VJ0QIs/WZhLCZjshB1vjnJ8y6CUuaVM
0OpXotHzXVxqyQ0+2f4DippQxtRa0ApfGuOg/6zlmkWw6vcwMPL62S47/q49vNnOK8/DP+8ruj6P
/hUM1Lrpu4X3q7mHuiZZCVahUnpcBzM/WgcmnntXbkmNKAU4421xG8hIbLZpzoHThKd1hG7eTwxc
rUN4Lz4O7A341CC6jslywIl7HDSyCyl5uEXxQEwn4PVfyxR8oDJY3nPqw6q204muBGPRhV+dsHhe
L2MdKISTAm2cbiWvEkysVC6luynwTYLpGCoNARoBkt2Agu0IanJxf4kotrUAeg0X3SWfLntB9pQo
CGwLbAqG8JSX7IyCHOdNj2p9HZ4hOuahLaXB9GZduVXk2wjzdxRBij9QRIvPmjWbS1hxWh7V90fu
advWjjaOUqaclqefuCRgEN+ZFJuj4JmVioPUikjN0bUJx9+Yl+4L6d8hMVfumyCAiwvXIMPY1EcP
GKwrTGWxtgoCudK/EvLNAjeo+FOjH4pDyMt0Sm24WH9CDSossX27PBQT5zQYCZpKRPDDl+KqjfGt
gZ3rm3LyyVnaHFRs72eV4PvbAiphdhO00c1oq3JtCzkzpDLqbFxbQpASg8O0TydFX6EgeglmXWsO
60fDI9rCuSUOkWMke8zm0A7cndrD42ujXxKWmVNpUFI1j4T4xpb82NovI2/u8xWJHPmKzW5E7LQx
/kLRGjBKXA71bLlegttQHCoeZVasVn/Oypxn2pfed7gUDGEy1ajiRVXzYERxWG/B/2Aci7fsFtZb
PMFAThtW6SkZGO0KiZXanUsqaW7ONHK0r6IGztZ69fuocS1LbzGXqmi2vsRQ1qVufN1fgGnGClui
WOO6MBhmpOovFY5i+vHXSr8Y+3VgIVJpaUdf/dq5WWTwxlMH+vKtGqaWQ3GXCDNEaTXzGtEMTaAC
dr8PeS+kI0KZU83zEBrztoKjnRmDg4sbQ1VCo6ci3n8vG3t/H8eHiptKEHxfc6gggPVcksi5bNEx
jYWJY967evmzqK2A88yn39XOT+Wsdo2fsc1gUT8BeuLl2lu8QSY1HFi0U+yoPn6MBaZ+aDtXj5aY
Gi4GTLDJ9hxPQKGffTKqK4CPgnd5Skv00yWPrqxr0iu2XLMCjictpgUnmhPc0hmridfwGXZwXC4E
N1MxGJmeY0RwXGX234YgqkG6L0Sk63KIL/IETDAHEfaipy1M5WARl6s+Igzbnag66kiFbA5I8RCz
gbSRdJ3Y0VVe+0m/4KrClb8ORj3QPc6CG/x8BMsWOZ5OEAMjhkaN2BqSQYJP9zhcY43jTPEQftPg
iAYw+FVT75V7PBdXGTN5ixAi3aEc+rcTLWBzngU7WoDz7Ozkn7a2cwRjCRD8QWrVa8S0zEAjh/GA
iWLa+7wvPm6XBv7Q+U4eytKfmPUkprN6Ze3zV/Vfuzhqc9XEfgD/dDKBRILPVyobSM8uLw+8xZye
u3ACmdF3tDZU2XEKDWFw3t9DeEZ+isaKjcxigDztgxA8P0YnCBR2I7GkbPxCunbIJDKicR3wRC/g
3e7zYbQec7uMqFP6kJao2DeZgwOPb6ILkXNt9PEoO+RIgoWWaJwAI2u6QcqqI9ivt7e92Y6Y8pzq
hWPDdQwJ3gdBnb4r5pTyyT2IVk0Mvfw8/6bEDpZADQAlNf9hrb+OQZ7NVOqiGE/hqQntWE0qHwlE
kpniZii9T6pbuhfKECWIQhlh3Rs/kioDAE0jj87uAygIwiPsAWx+9MGDJeMmBS+kBVdj99YnC9AS
LSOFqvPKd1DJON2qo0kwb8HOcFhYDwLRTL13bT1VJoK3sMHIWR5IKCc0jzDXwCJ4VAt13VbHyiqS
LMCagdk997gObDv8/8jVV3exXHdokEz0+9VztRDH06vz+uhdfKMrJgpBH0sxjc+V3FkneyGORfIc
IX5REQP+3ncQZH/SoeRS18pEZ82XtBXeNzxl+Ivi3S08Z4lY2tU5/XHbTb4joKhZYyVm8z9S0TfP
TzwtW3iJsqgSc6FxRlTnZUukr+kpzb9SEHyVrFiykyokZ7L7rpSW9ZES5ZY99qN/bwFsFkzXPGk9
ZnVJZ9wB9hTeyPe60WdhAfX+zQIco27QuiMrJAM78TpFELCHCIoKsnAh1dbSYtZbjzXzR0VVQLao
SBDk6d005qYGeJaW7fOJNzosT1KkNj/U/9zk+G8WwDQrhsik2ddQZK8oVft0fTsA8b0D4N2pVFcn
4k7d5/9+N+kay1v8K4rGGCHIo48teiHbt8PSPqcnEQ3cAaXqj+IJzfOL4tJddkeA+MatIOJXj7t9
e+fdoATmZ7WfS/1avuw8LKxDeJqjDLORM1hwhE7kNdXyugxffg0F3qBH/yDoMciYFwX3KIOWSQCK
POcmDmqhh5o7aPFiijS/pn7fiWW6FVq9FTiYMrXuCYUVey5Yve2ToNdb6p2G5Hi3hgbE5kPOAHKc
l54v3pMhOoYD0AQis9mIMn787SSRijVA9Zo4+KnwVclDrhDbgn0zc12hdTfMfr1wJgWUbQ6cKRxK
jbKCFh5B/m2LG14ElIivi9P9FoTMeIGJIrauyyyLzp/8i/94moyS7QhOyPPvHmB1ZNWiaZlFcKqz
09gtf3T4QkgASi26xm47oBHzGLgFmpN5gUIfp/1OqLIC/q+N+zzIPVy/nfFx+cwNE8cK6WE3T8RM
fPoli9aJWaKIEnOWLwJU7pl7nnnxl+bsvel/mMp5OZK6KwO0BuJeR9/psyAqtYVbjO1cFGhxOf/D
MbQwJ8nDzD6WlWmilQVj+0D/E8nGerSoTDzSuyMJvw00zFHw5hHlffv8mefLG+6yf2NJUbAGE97c
YSIxYslpLOF+z2fksxFJmt4dIzTtpCIIQQbKHpek9oFnU+jqXDwSp4Rxw6K+J1v6Lkg2DSQ+FZ3F
Tn2cJkLkqpQazNayAvf3dRR+pBr2vlEI6TMcqJ5kd37wVrZPRnn9SW6tu1hl07gqFAtOE0XPfXJ6
iEaa9YrTZpyFM+lAdTGk1SijaqT1OCrZTuB6yLqr0zbfMcL5XnxymEmVBmWRrpGG5tkh9BKrxM9C
rGheqYXEoDRL0WzMLZrZlA6btRdlcnt+KoQ585y42DhJaa7fSWIv2X0Ii/7Ve3DmLIyHDEWipVEV
hHDKLwoSq02S3NUaQi8gB/FByjcNdaN2AOmZwRejAK6AqHOeVUlUHnAFCWHLVPBTq3vRfuZPESxg
DINoOIEXnRiuuHOuBWir6vh84Q0mhNRqRPZCP2BDk3smmhv0Aqz0LGXo22uJgXP3fJVn6hBWg64w
CCcd7+co7CHxVVV0Tvxmby3eGJQLRoUP6Dn0BJfdzWeQpEVA+3Sx45ZHN7DAun6atXXUZ80C/zCh
Tex//cg3jIZ+jTMTa8UEtz2v2QhiIDVGJeYK/kkUjWOtxOOkIzr3pyG+/jzqOZA6JDrL6IUHhNSX
4Dr6DMa6Wu6CNMcnG5QZl3WQFST5LjXlef1WOOM2HBsAQL0K54b1SGssWqkhfXHGo71lnsmUoa/y
9X1eVujYC+HEVo5LXn/ixL+rx9mSgkLJN/bO0zfpw02ma5wls0NpXL2XHPnRQj2dTpUXTsAU/SaY
tUI9dN05FDc+kM0710g6l2J3YRZEOWE+6fbVXgJ9kLvVWRcjd/SuGntJiuAYsRIjcSWXHURM14/g
sS/1oCbW2nKNHCLEi2mzQ086rGw1yJZCmNl+TZQeZhcEg4dHvxVodt2486lvwpeVErxCAbPcK11B
GgA6fkHnin0oNIK9hHtGQEbBBALKBoDyEFpHdvWRl22frNUjCwvJk/ktpSREXfEamw/NvzzI9FtO
CK4QPIK0VlotsK09/vcNUylXjaPgbjn4XQmJT3eQNOoXL/CDlSV1bAvswxX55wUJwOCHQ4HG0tyr
9aZTSPAOej+nYa6I5kVaGDMdVeD4kGjXZcyULXvTBqF7Zga7y1Cu4FKOKFFfJBqpCTflBIBILNNX
462nNnkiyMWG9u+tQpwPzxv7lVvSBELL/9sJLUA7ZJ8tWvkqPbeCMqxY/1kZupifs+F5sperawIb
dmZhL9nMNx5COt3U5Q4CC1V7+frxhpIp13etlS0d/1yUGUXjygxP1JpYlVPLhA685JQMhNl0BvCa
qeSGypFSAcY082YxUP0NnVkzIstrcO49X7PDLDfBSk6faRFBxQSM/0ojRj+pfkDAUCKiqtalu2kw
DKNPxt7Rn3/wgPLaUnEfbgk6k11GR3Esu40qNnrdokenVulgd6nvYo3zC252OVKJzKv/NMi9j6qx
p+stjH7o+ENrcQZQ4cSe0sPMXPot+EQI8ibRbu2wQAMF/Kymt8Sq942VKpx0ELtf/GvK+wHNyF5U
EGmcXkSFSrD8t9MgmHvVoB9suDPGghOLEgk/LKJbGFeCoOe/t90bKetK3FKuoj401NATCrtqXWo1
SvQpW+xrIb/0Sj/Tdc9FR0uf5dwQn/8agmQgD7vxmMstq209+wrrl4tJfrdm309yr21A9WU9VebS
IPRiDoR0UV4UYmM3iYv+8Q9Xu8W+lign1OP6LE1L33XVqJ+Hjq4Tyw9pfgBVM4E0yxxp//dqEXwS
AuK1e4agTHf0oUl6Vzi/Jw/RJmh7XmpQG230ceN45kZ2p6ncWHMT5yDFbYUjHtGCHDDPrrI08UZJ
iA5GNp1v50aSEnaqkQb4X+CnXhlEs6YfXz4DEhYFN332ZKuWEXyqXpwG5DXoJcC/DWZ1Ej2CBN4v
1MiFZyS6MMsFo7LDWVgVueos9gclJUuuuYwKbp41pc0ZL8J9dxTEkgyHpcMXqZjv7ra0WzVL8M5j
MnUmHQE1ufE8sZVqpXVo7gxMpdImkZ6H/yykh2V0hFSckhgydm+nIinSkgZtVKkoYDSjdR2KUd4b
eIR4EVW7SHj9OZQOYsMrWlw6sxzDgapd/ICDOg1ZdzVrmeQYSTZqBtJhlsxVCzzTQLyj/1/GWDjO
kmsNFIGgS/GEs/adfUlxuKJkPJj3D3nCxAvc/FSDJEn/DcClJssW1AeEv7NvtE6wjfhB3t4ZHeAC
6vvj3pAHSCQ0jiwlwCyKj6eJ84n6WXF4qtNV+akV23PP5zLUsHXKb7xzmeCpJSanVXfyqEWpCLjE
MZzOlD5tVxeS6IGvN3LiO54mucJk4pXWv8UUTemSHLkXAs5xzmQim6SpR2W8O2RKyi62OjIYxgwI
KLd5jso1sfIInx9UMgVo3jXV/cw41uXKgvHtIN9hXdcy9mPQaDUtCAlMqjCYPr4ywCQJw9nYbioY
Td0QpmdkKUzfZBRzI6zOZ/LV433We0RH6rKhoxlTVAHti2Jz/wMeDRu+VCa+49WH7OuP7341ICH+
yvEL0gNXYVakZLxyivBU0VBwyGN3pIL8EyeLkp3j56OFORtQ2OIbEx8HP4l7nVpPlfJxDaog9Q2J
adzqH+cJzirgRMilWwQTAi+PTZytBXvn0pU8mWHFjXlJ6OgmQ1tlX0YZR1msY6ZIZ9yHqw8iYDYk
0LMC5XdijMhjgVTAtEKLIZ/b8N2zwNI4Q53e+Qchhfg9AJzrPz8gmLNhQuPfQP+WPmLtOir1yeh3
UiZR30Ko+fqiL16Tf7E6+kFZWuOJQCQ27qqRGxMBlRVGJitd1Jk0w2lFwDBbfzM7Y+qVVkKe9sE/
HlooHOnshghlJ1tLLu6QwqnJsaIuS2x8aIIkKIznmCFQeTzeOhei5U74xULdjZA0gzho4FiLOgTZ
56vzVtlkcW4Mv8gAWOOAg+suBCadNTdYbf2vBnkRNgT4f7IlVW3uAtOION9DroeIB/I521dO10zH
K2V+MWqP/louVc6GTZ31DdKaMADNpB0xvXRWTGAW73frGPNE0N2al0I1/6ipsKhx0SEtjAjiCXrd
AUzeFY1LKt/ozPwkyghpRdBDVr8Gc7bn0VgKmL1hVCSLakdBq301PalczC2roI/tBqJSITxtmXUt
r/4F/iA3sie5T+vFunHc57UDt9vrlGyhq/7rnIil21E/88wV0MR7fhD91JhqvKTFL5rnfpKuHzSN
W60uTGvp7++qG92c7jiM93Rphhd/4MLnqtw4KQjQTyvNjQRr3YSbvRYXGCsTjrSwzyHLz4ERJtyg
ItfDBnpjAut8MdWgw8Ho14lF9GgY2yvpomH3YapRnDs4i7EztnXeXbl80Vm5hvpwhA7WqTJ8aiKR
cT0gVu3DYfamxpgyrscT0AGJeQndb/pFrszBMbzmUPP8B/gQZWEQFYToA2Kt2EqKTlT3ZthQxscU
+AbZccG0TF+yQe1qQslnWzPgV8Ii+61tT7KySyy122i/ZIgEc/aon11meM1Y5kWTtH2EwBhqe3e3
wE8G3Lh/8PAmK47jWJKS/swEMQM8GT2VfTke/tZ+NesN+tI1dHDcuGvn1JRhHjSXbvfWbVMfi217
Qz2S8aAOaRhlKoubEybZkUOsqCddlBAyI1wqdPJRSE7f5JBfe7I69Iy8I4EVQbJPcVkNzYRQjtq0
OciyB1DALl/pr9TPaH0HFMl8SQ9tx4Gi9CdjKS1nmtzjgAjymZmTKXD5B9uxO4idgkQkRNc6Nw6u
mzLbrTC5z0gLzd/gytZq5PbkyL+Q7JM6G7HgP5uQlxCuM70PnS9P3moRVpPg+wdjCuXnlOyQXAXh
JoWnhhdx0i7zq9CZTsmIn8zH2yGqfO0+zmE9rwiKR/Fav3Kn2rP4a7/CrAUSKyZLqHgls9LU5eV9
B2vZwa5M/KrYNAWg3zznOqniYfvOcL8XIorEGp7xd41L9c6wHjNuDN2edXPg+xKrtW8Pk//9b+3c
9j1GzgTgLJ0sB4Q7YisBF0wBSNi/bAv6lq2HRR8t1x861stq3kjOKHqFOVBJtWz8U8XrnHEoZsQO
xf6pcYMwO+JJfBd+X/RP/kgKuhVu7D8hOPV8V/Jtk7ujxg05jf0vQyXGmKAGpMJBGMeTTRh5jHSh
W8w1mdGri9c6jEcy0SCj80NyYAcOFzWj024SW3AD8FvjYkuBFz9MNYu7aKiPCSnrtxuo3HCEAKeW
sJnESxdGm+0uaTqN0wOPTux6iy/bWqxLPvlgyTM4D7/8KRZbYsYkS0R6u5N/E5/ZckcO47IW87r8
/CJlBUKKTcHuVHWbrRRXSbiUknjfmEs49+ROkQqmEJPV8p7YoVFWQ03+P69llLCLMdKHIt42cwjr
q24xYM6fGzN7/tbUS5V9FbdIbbWaTLAu0vbesJId/pm3yAztshRmjO8QIVDqpmFoMpKvP2ivaJpe
rBv2+F12YfnwJO6YlweuX/Er69/AAf1c5OUDZzq7Ogxyw/0HTO0CpZUGLXOHYeNLpPfYC6QAEK8J
TwgZHHxPRWDvpt1+pX5AAhrCLIk9ji/BaxYbpp7cqSkqNseTeMzJukXu0nufGd6BuP9O1INVGXeZ
y6FF4SRYLb+Rg0m74RN7BNyS1Q9/3hUhKJI5mubDZBp/7ci4yWhcUdZIOmvjK2/ysGb+H69SdNPK
9YLFmDYD/3H10ZAv6YNyCMyWhRzXhymI/BIqLmXSffZfBkwW8j2Vkz9MhgONSUOYvJohqAFsd3wz
Js4w5UDByVHfkHbQg8QnoYvRIFunwGHpXWfA5bsh4/Erz8462e6+dGtp51rlQDRJwBXnSVy2cIAx
DSCUr4cBVGl5YROL1zdl6IqSBDCKGSEETM6lKUod/H6SiTA0i8E3CvDqbxrM9PQLYhaW1kZSgqqH
ml60OcmgRHkGXv8X3ryEGJMGltlZOWwCIVESR4E/EqnlXevZyjSDwJYKUuuoLDmASmHt5uNljRn2
setfqEWcRihARl1jro/4RQSYTHrMcUH0q3LEeW373DkYg8hxbkdKxJvBNHLu2P9g732YtUEAHxwG
863jYSBU1lzzR4lL5xDLHjtB5HZO9Rst5Cihrcr9Fcpj98hWshprqu4sm72O1VkN5IRXRRUc4ejJ
eKcxtzN/KsE7Ss8h5I4uVmoeQvD6pEIisuFsNGSIOqgGpaINMlg+pzyy2pWP+tdzWvcYUayoRoWF
QnU1iRTHrPJOf6TaW1NBSIX5CEz6EF0m2PVBBnkNbccoST4t1Fy1EfmgGoxR2opQHaQAXJq6uFFp
g/hlh2I+SBbLv6FA9kgkvTD+AQkJZWN8/1Y4/08qb9yr3avAEhqEBQF35/FzbYdR59eyBUxfECx6
FNuxIu31XmrUOwLMR2hhm3/3E8TmaxdfvbNm6Yr7Kshm2IkwIyeQAI2YaPX0PjYlJC6bPkp7Ou1l
PnXBF841AOQf7wiXYaoiR5UpP9D8/aUnGQ+8FyUrgevqxjnF9cA7qzbjR5OTrDXy4WI1AdGuYbYC
qQ8Z2AoV8OBmQbrZw1uPYU+CvESt7AkD2eyxTQU1uIM95Y8Vz7pQnMDmUNGnV/tEykxFQnwTgUpc
h5/2BoJ/scyIjxafPA94m8vJZd1knxMnY4fGMnO91zvnESdKeeMzqLgXLoYDpSZM3VFfycqNLu6z
JhjWFswwWXFAW4MR+rRQ7OfF5nozJok140BwJY09HHKpev7owCdLCF2tUwDkTKVtjhvqrWghG6Na
B/0vuG2PPoGtvObLejV9+A3rJePghis98eNXpVEjEsHfz9YjVSPigyXHK8dAudlHtJVFKaffX/DC
QeezrKiwkxLqq2zzJ7DSa4u2tN1+Jtxi2aJgTpmhkNcYmE+s+017gJmMMLKQ8pFoE+CAfVmrnBKJ
KTRFP0nJdXkytJIqYiX2X7U70sKHOdyRCHw2GWeKtBwWZxTVl+LLTJiYPQZYgtjxMSEHmOY0yDRB
jyIYJwAUrANm5E/X8OR5YhYcD74GVs7E9w/DV4vcWxuuDPRygxHfwICwbf4WbGUVgi2p5lZR0bJe
nWUdqVEyAjTyErXzX5qiU3rK8lrMhKPQg8je5xu79xSuPMZpohPooqsjZP4PjlGLJlYl9W64wLhh
gu03O5A3/nLOEyf+EPxoQkcO3c3zyw3NbKPT1uv6ggFLUNHcQ5K+pY1WofXO7WO1S9oegrE9b7Z2
LpeS9dXeELWZZvB9NSwFfAZLbCyodE/dlFsPO3DaqL/V5rsLNFbOb9CEZupRucPWB9OAbLCDPgcL
ci8PQPDuSoldpU23f3aEA5XSbe4fe6q/nzRhVrhVfWMGvNlzcz5HyGGG04a1jk88br7Smuhd7L1q
FRUqW97FE2G7HkgRTb5Chsv6/pJRVN70s7eXHCpEVJKg6yEV5LYyuvPBeFU6NNF1KZx0nbRsh/qB
qwpg3GrXT+HVD9tdJ3VOqjx2C+79pobH/8Rnc+sZPs9RpaepSnX45i6NWei8AkxrLQL16Pm8djGp
HPkf1A/Jj6rjaCZNhlu+WzTggSqgIqQGFP2ObEaOcvaCa7esu7SqgJutsrXwCxE3MlcOIw5SElkj
Jsyzmk2bwJXTSct8ld+5f2wNLbUQdI+mzlISimrbtBweAp+zZfbFNOkqppHYBYKEco+iCQzS7AHS
7KDzmgnFNuGL5Nb5QQ18czrhN6wd02wqSCWy8hSWRNDwL0787V9MJU/rCgfpyKco2rSHUAxvzbUr
vG+5PC2YrBBZF/+ti2oY2caI74kVBNs7AaQq4fHL/WQzRASwg6nsuqIh8Re6yBqIR0/nbchwTc6i
jb8P2jSEEPFMs//O6QY9pCcUHKMA0M/cwRfSsE5m/wK8Do+wjwWmfXHjwJJy1D4cWnVCPLnEbLei
+N9EW4PVYxUYdWwxE8RLRFseAZ7+U5wNGlTUsxNIdgKgcZeW4uTFr/sAsx6wUDsTjVg2+8QHWLK7
GCA1+a+DUzWbut4IfmeOm0ro+SVSm6E05b9BLH44c7Yv0aEojBS85F6WWM5eQcXX94JDAeW5b08B
CdaXfIqMDYgtZOjXaaCOmwlJxCuzGp1DHmkLWVJhWFo+CsnKkZ5Eolz/eKmS7zPsvkHC2pMM3gC2
lIM+C07a5xxfLfySVGkjCECx5f330Zfi7CMX65Dx39DLygoYw2/IMJ/Hbj+aOj+/2I1yh3uyXPXJ
PLlkbgcc4ozsHkOBBKvj2qoYUBu4RiR6FD4R70qaCTygeXmqI0GsA0C42emeJOYT7YPQUk1TiKrS
MylS6vfA8wQZWtd4nDEb3DYbNgJzH30IB5tYdNZF9PvaZWjPchcD+KlqYAMHwpeo/3668zLTnjYQ
aTwuhJBXvBlEgoiU2Dr7kaaeZ7CjWDq0RC3MWf10OYAZgO+bIqxgApJTe2qmQ+MXwIMH0MHeNs6J
HktOnIbKBsSms6oijWbAC9HXVuN8+UYpeL3syTEsDJKjq2z0VMOHRGzYnT9xCs2Gsn1DTUNEKeoA
bpuBYlgSY8QMcihlYvllUZTx/dD0WzW5bnuNEx427hd870AJzYTOyyJdXJ9faIfXEcY9f2C6eoaO
ekzSEHF7mmiZQXEQNCSx0L7AdvV3z3DpDjUY6SaT8MrgxCQDJLC+PFEtAeVLbmDG4yFDj8kwwI8M
0AtcPkE3eaVT447AIeapG9kIPk8FC9sephlxzwwA+D4bcOYwGi7yG0nV85wy1wrjLTtvwMIK4YBr
KKnuh+7ew8Qm+rkIiQbQbDyRedga6bpizDvo8S8xuSpDj/et45PxoTrRfV2kGVW3kQRsamFRRniE
GMGT85eiEbBAAvYeXVEBV04BXFpbomBOZfnnUbBbGqsuEYm7MrWsI/Gabu9j51hpRHBY7fcKIVwZ
VzUUW6qKtVUGn+RPmOyrINe29g+JGDEgMv3xitsdwda248hI5Oo6oBVGSK+XeCo8HdScQXBS7aY1
EwMCVZoXohzJnaJTRCkkO2YJgcvqJIUKZ1JxaVYM6Akp5+nqsIk7tP4cCYSKXonDWM+otwYv+ZX0
jshnkPWfi/gwAx01J63HUgi9GlsVqBOhKrDf7B4H8GZAGJFxO8zQzE7++e5MfR2yClLBDeI+ZgD4
OVvSJnjRckxTJ6E8iDak2/TxIFDaSQnfrC0MDFNGsgVdzeWi2G/nyn4L2wUESM04l+bIk81hTBGH
Ld9qQktHknmM1PhbKpFf/qXJwCggKx1z3DF3lakyEaQ+crFzt5/TQ6c8hd81GyDOB1cZx8tDJCh9
GMO+MUlZVF20AitviL/n3uqxysglpCg9TKwprh38ia4XWkFbxANqfU2PMm8ua110A1xU1CQ/YPjR
SQsIwSGX1hHPJek/6409weeZ0lotuB6kzOAtjiYqqciFcewqakZ1CRCLuEUumvl4enk2v+xlOgKu
D6rnm8Bgqfhr++ZdF0ya7lBkxN1Sc5mf7lmbllJtQwhIF1p9c0oSIABKMZQLJ/5xBd4W69sUkNJ7
NdA0sdtF4RMYrU+aSlhOAOv4DWgmVqUZ3IJhTpTBXpJALcQaG38atRHNgGGTN9WJTdmTReaCFFmd
rU+yFkGDaf9V+jq15Cv2GESrvHtI4Ir6Ib0tfYXTX6R/KIwgoXaO5Ch7QZDPjkQ0sb1KbtRtp1Yw
ds81rCExZzQrZot4+ytQfPF2fpibNYrjFvH6FPvuWXOYUbvJHPRcff5fRL6GUgKk0Sfx7oc8L7Rk
09qcVpmaP73qKFQar/610LvTm1N/yb45+dbq+RR5chozSCG4l2V/IarRWmHoLCV++ZE/5QjM701C
oW8mjId43RQ9N7uER3awvnQ7zaWR8sG/0xaKc8MTEM/Wsq8PrW/pMWEQtuZ8fLsL5+1nPvhoGxMF
yRfu6u84kSjYq5h9z0ZX1couJ6ErM/TlwYJ95Q/2MCGjnXmroIM6RRis2PfiiPzVmXh5z/GkwYUC
I82tYmobR9EdERKiWK9M6nfXEfTSCb2M9/4tR3uF6REPhTWCX9iGLYzKKAFsxd8XUJ/xelF5t1XX
p9Nv3ACmRkEHxbdDQwCdJtdWIP8gAeKhI0UmjLvSG0rj4Z07qIgnEARQYea+f2nrw3OFzhMVecjl
eb1mIsZUP07h/YqIa3uSzdmbjUSG++wngB9/ZIcsSRkc734pCNj21kntFJ8EwT/BNn9rYkvXHI5U
qhuGvAHurnbBqADNQ0hXc/uAiUQXyhOqAVcCXeB9lKvUFQmIY1tTcjNahFipj7e7QZfA1Jjqltw5
xZFMBMLsKJ9E2PAE0zwmvOd1jcf74p0TBUvvWZe7KfMLHt0baoKGjYpRx9S/bCCPdVvskh9bid3/
wtVvcGZ6i1lpRCx/bG5t6k6PsdvDVIisEPRTb7mvXsOGucmbQ2OE3FzSmVLF7gS/m8aa8s0Dyo12
TLrH4sQx/Q4jzlOT6KUeasc7LY9dlM/R618835oo/Q96ZLkfqxg0bh7Y9hAfoDhEku+xZmRQXtHM
d6P/Mbk4sijjfRykU/Pe9ocazWOP1vMQBUCJIxbhG19YPGeLwidBQ0MrXrMkAUCEey40j1L/DYLJ
8xM0qW5XqYTr2cpFvvaUbR55uM1MQBvqSKfNtwAOfe6QIxPiEBChXqtUXez83BquqiIwTpv+4gLe
50KFSEkNEjpQiQU8WxmR0VlL1Pshq7G+u0Lj/t6KT125dF8lN0ApUVjw/47TPX5C6Ar5Ix98qd65
OxQjPV+X6BvW/1XkL1mfMxHFz6ZNLfcasdbzM2EwqUC3jWDN4YFx2BZmazxJUqYncE6kwWf3GSfs
WvupvvDSvUNxS0QvUSsdxe1hJVZ9asmRkVo3iPVNGiUpjYcwst7QhsUGeraJXmUx5no5KFjs3x60
LRSpX/g2FmaMCVAjhnENcfH+9/QSEfahFXrmphcqA1uMxJUCKFo5sLUv+1fEZxBhIHz3QpUgydsp
7NKqRuPPQi25N0m/F6kJjz6GYO920ksd9tOucev8Vg87wck5bW8OU/L0lGISBZWmuZXccBQIIIsD
sfWdJA9FmOF60JMF/9oOPkoIHA3JsmsYBsIYdbAO1d+IGrfVbMj3gnStgq4ahUjKuDgBgoqk1wEy
iOgCAK/3VC7OoWMoiv+kNsYrYIL6ZrAwTLJcuRusFKYaNDH8byoz9xhOj8mPpbcmc90rj7CPI2Q6
HTXF7wQk9j74G2cyYmF2GrB5ajSPA6rcxZVuQgVmpsBpxoF61bSaxGPqy3hDvsz+qRgbL0o35lMz
16C37P6cSUII1Yd0TV5iAyg7Y+P3w2DpvNM9SAAAoAGCkYqD9AUA0LraNV5rmJdDyh/bwSWTpiK+
1A0PGVBdBIUBskUtGvpVjki+n6StnpnWheQm19tEGu2zlpSxTSF2OArnA01z6K0JPa9FLC9f7csq
xWhxZVyeHfteLSVXevQC57Fopnv9VYRmnOIwT4/t4yr2xVLNMJsiPpuGyRZ5AV/WyhQuFuCdn2E3
HGVUoIlO2D4ZRd/BiuU2toTzh6pIwvRtyy0hK6ble1EOq1/9yfOD4N73GAezGT9Er6/AY1PMaqVu
Br+GSEv4NvYBbjnHEXiuyty0Ol3EbWA4hCMdmm/sCcRDZ4l+P37XQMnOHbqnyKcpldS6m3dTB5Tu
nLmDpcNg14/jRFy1+Q0Rv7UI9NNJcQ30z0whQgKizUry9zVugtBhnjLULe1VLr7oZXFCM5FU+ijk
9A41/sKqNmxo9r8DApVXHC6HFcgDsPKIdNnvDqyU2Id+XEf6SEOVJakb94EygvfB543HiHSa1PEk
2xH1gS+2E9GVFxWyr+ffVeegnuyQjiVzcyZJ2Py0W6dGl30GT1RP4G2PahrlYhvFuDqpkk0DDLWL
KQXO5quumSmitynmvQd9mEnNOFH6y5oTGxQVWr1s1yffwTfdr6SOopgaGgmhOcGozDtSIFYdDg/I
mqbo1nAekAZL4zvRoUqa9iHU++d92o64yu90fydcy+qLlR11CUnY8b5OMOgeroYde3vmWTmLdECR
uHi7gNA5QWDguGm43j1IkE3l5h8xo9soGRFFI170Zy3q11UXn0kggWJHO5zvGeEFtDjHLxWfv32r
Srb7BKh0yKHxeE8K1Dr0q+ZP1Lq8LfWhbC8CPTBhnmG6TJM5VlD8krOoP+YyKvV7nApvP9Ase61m
qcyc96lTy5wsiVfn0TlGhry195i0Qpy9kvOScGYs8gLcj+Q6qJXXNoylnuXJ27CHJC8/k3ID3Qiw
nua3PaHXxrbCIWCf1hQfl1Im1EqiqCDK16jSJV/84uQMRiU2htcZtpUoiZQNWmcHAUMbGyscnaGe
NsQK2B0RFt4OyNZcnDqOokTqJbV0RRZ9Ak588WOmShvyZkqfzLWuqtaLyQ22lTWPgivBDxjU8eum
lzQr/sdOoOqI2taUX7TOXQt8FR5K+5pSy8nVlHF43D1Ub6LnP1Ee/7r9qu02vu5/QXuOqKWdy0sb
tL6faEyO3fJH3BYl6MyxH+LD54X54t1X56kudcCTgLgA3qmM6lo4lX7i4NzAY2SvwgbJjl7ZcQyO
7Pojk4UceAax/dioryToqNeEZbOvDh77qIAn1NsjnbNeQeBaiiPE3GhCCMte3NaFVIEOVIispi7C
TYKOkUC4TJIa92KqRIkthYhswoOxfBkNTJhmXX1YqgciNJKZkHMCAEPa5rZNI+pAG738iXyy+bgO
OvDSLSIaQNUnWOlb8GHYzI9iVwPnQOwnO09EymfoOG516OYODCNek5leB11BY6755W7qdP3PLlpO
SavwAstzc5U/vAoBExHSZlA7x3/9aHwlYtISLTkqqs9P6ZdtwY12tGN/OrleWLlz1+VrWBaukm8G
a7GVktRax/3ICIo1Yz2ldvBABdWV32qoYPw1KfYETmBZ4OWwvcBlrCIYMKWkib+6ESG/cUtSWhi3
mURfN0kOdr2DsSHBiJ0CKBZu701iXiQesETeHFHXAhKZS/2+2+SvS6VCFgHsEFB+j241NGsipx3W
XgOIlvDhLkUORgqeW2Y1YuvdVG78gSlry0LmWKtWVeDU1qtvdFpAyyOkdpCkClGCJaZA+67i4HEa
3W5k9ax9lXTF2gbQ3XDNZVEXf44UD/JT+E0XiqjOK5Pn3zUFaUH5uVkkzzgAq5NrPMijkqy+tWqy
fvlzL6rLdrgMsEdU5jFSacsoy9jhINLq08t7Dv/hsa6tJ8/pKN4+gaJcbo4B2YYbMrxIktLrISjU
mauHdRNOG4Rs2rVIxzkPRnIqnrkDqyaG1rua3kENBM5h+5+aDjGoJP0BFiWCwOqpUWL84dEy9x58
mYFpnYogjRbctECKnxGfFNA4b5a9PgjL6K2/z+6PTZCAUiz1KhHzjpV8b7G0IlIkOHoCChS3JotV
CMZT23MygJKPvW5kjY3jIJ/6v8nXl7s2kamzj0elGB/3BXnlkpn3R2vae7jIrvnpN0kP3HqCNdYu
UYnzwmj5Lo86Lu4xgQpMZPAOPJv1PyE7VGU1P8Xj5InkiQlnlE58zD78//XH6004CTLGvzvIR2ii
M/19SzIbz58Zmitwftku1nZ8Yq7YmmN7dOcGyFuWYIZIsAwf668qMzEyVtZdg/BQg+02dR3t7yJB
bWUfaynaCLGxHZTiDOLXbJwAkFbZzs/BMbWCUSqzBP+tvNdn5cxBp8NDHlMVWbYJ9DUKDMWn9qPO
jkvtDtwAnFRV+/2q8g/X5OAb+VWX7M7h5SZys40RXbs9lfAOPcVkBWNuNegs6eBtA3Fxvyj+pXeN
tywUaIsXQJ1EJWIaV/rBKKgSvcDKkC00NvKyyNGaRoZ3T3TFh3mGt2mVUQIJdBgHvZRB3G8h0pUI
Fn9Fzk1ZyN2y40d+5e+0HPJEzDv2ngonln9TcO3s0oxQk/rtHFKMHSVbtEVihkcMYtTuNB0vlBW3
XtKk0Mmnihkg7nXfbagKQudzg+gU4C7gaPsQJkzc39OSeyiVuNi6D3DLuU5+N1fNBEzjanjJsNQB
943KYKw5UteP1qpKPgwJqr3jidqyYPEhoNgDA5xapPsFIxyJjetgqXv6Nc6uYCRgH8dpaVLA0W5s
7DYtgQwhjaVdwOZjQl68dx8YKtP/lEFVFDcdg0oEsHIv0jC2MWvMdzIHNDx3r+9XNbiilvy0Aq0C
abVYABmTGGiXKDZStTSm4V8XcHC4Xs/oq8oDRX6c4mqWM9ma8DLW0NIU4FSkdrAvS8qNmjbwrQz4
Oud1KrEtlx6Vmzy0DEoP3W/5fLDb8qeUhYBS9v3Pz2F3mvhwynLU3nSaitsFEfgK5YqNwj8Vjsm5
NuL5EU9khdT58E2NYQ9sPyr050++Dp/YgyuujDvi91RARuaRP4rFhEVN0MZLXxSFppgSFaPiw+13
sy6RRTWDOOAGiOLOKuZSKiCS86+6HqFNDgv6E9FPJh+kpvf7mhYxfbRakN//RbZ/OTh8DCETvd1b
BKKWDLw1ti6T75BHNLqSVVN93w1Uu2EewTqy2WuIeYkoOFkLBWPgwtIHqBKPKoy1ZxH6oapIiNZC
b7Ebn5es1CDQ/XG9PZrULa9qYvEtAMSGRai3zmjuzrQ854Fi+FWWSkNq/QW5qvqTeYOhHvwJ1+U9
iZnZ0SXz+PjNd+BNoLaYcqV6+RvG707DCj6XyXMFfvai8FN39vfiitUXsexuzxBwbu0S2M6rb62K
wrlBgOskLfmjrP7mtNta6A5BMea+D5yLVXZ8FWenW8hNiO0GEPdc9Y7Jkh12nP7FFQQMcNF7QjY+
tJewLJq6sHPv3B55ZRL3+oV2hqE9BnNOQ3XlVzyrI5+fldP1piuho2SnH32KU3HoIOqiJ1PlzZAE
v7LIcAWI62JUw3tWqqVM9oCcaWVqu5xVwfTfdcO8hRjUtT3EMoR4cK4Q1rE+ET0HKZpJVGt6Wq3Y
ICA2Ro71C6nOP43bwmp6e+OYYh9AdB3u1Jbaq58JDEaNA1xY9CvyiFPNYzIqbm+0JCCcZjDu9ffb
ABBXJaxUCsLYtti/fEPxsyQY45v0MWrYeMwxrfNls+/uaS94lOdWJXGILlKsTYY3skgPCKj9fV+7
OSu6SIEDhdofYOjnmQQbwsr050arv+k3cNlvNH6SMkgtZohsq0/XubXiHaOSSHx0U/qp9N7CpFRZ
QVTgO/7L+hj1XasZ/BG9soTySnpgru9uLzkhD27e9quu+8ZC5vOKuB8YWBBvX+hgaaxJGVYCVCyo
zMT9rDiovSbPgv274K++5KgpU+QfN0uQY8vHiQ32+SX4OQwI0pafFu0H7z3oKUHp58RChFi9E2wO
keCQd+nyL8AKqKEIpVtsds27zD2zWZgQMosiOk5P8QaBzVKf4y5rQz2Nl6DxNAr8oRWbghd+bLbK
TmKHn6jJv17ESnbU1RhHYjZoNVQ68qTkMrV2BLCee+zyd33zyNNLohXPlfUX+z7OwJNBHP3UDzES
dYfpmghj92GP/B2CsXHCtU3c4ueZnRYixeLrubT54w5btJNsiNUKisz+J3QAaBRnWbQhmz4lLSXX
4Wnxx4uxkupdzcottVUHtCBIRLDiuXmVp0XWs9lH7PaY5tVzc9dZOXcFVwMu0UOv3DdbIlGwYnkq
xptJNyhav1+ODUjJ8eTOgAO2lW6E9A/2eiDztvWOdHn76YhQj/AXZY+yqhgEcZQjqNvxJiJGzqnN
FKlQCuDPtfov6ejbROeSEVmwBicS/nPxQ6bQK/R+cWCOQ2bfPuFfvhEZeVDQoxLEXyDtPCml4IG5
rcK0KMWmS/ZkwRuvQUJ55k5bmZhUKh7pSQrPhWxbUWY3GzPlNTcOXFogspCziWpW6cyf5Wz2+XIM
r+kkQIK1gDCSu4n7x0t0UH7QaVrnwM7RXjrypZfWtPa6S3+SINaGB7nq8OiGmb8Zv+4OmInQ8pZf
zN1gMW2eVW1uFeV6l4RIy2SGTNJhX7WV9oA+PcnrUPsb58Rlno52tkHQhP1Vx8ouNg+LYiPIxgpr
zhB7MOQeaQzZiayBR/7FKWqpYw6bdL/WaZTsSe6VzH3p7b3mX7u0LSL4G4DHr2ofewYNn/Dsvmay
/IhZIND5VEcUTbBHNg4gTeA2Cufg0eaXVJ8ag1dmQ/CHzp1tSHxNOvowemDtw12bBCt6xKnVBXRj
WcqnZNF35X5cNufOCvrYhyj1bAL1o8jJkI4q9kh4ZZWUt7ZOvcVfVXwJk1CBuK3//K9XGy8axuow
+nGDdpKOghkFafojj8WY2Uizfw7U81QHEY/Ymb/cgCucDQja1LaLSiYD+eHQ1u75q6Nj/J+0hqmf
hQL3200qG1jrip9cZ6VzDSuGZxdmsGQeSyG9PqtUhDrz+1oqB5JZGPEI7AftQlTZo+F9Amp7Ycq/
bcf7lAhAm/MWbcDMKWSTTEBe5V1W5KtNknA36HM32BZOkzietVBsRgvWNKyWEyTpv6vrKE4vx/ZK
FCD8B7zRwqjnXAYV+WG0okXsChAht1vv5i+VlfPogS/+qzHZ5Fvmg2sx5qab/x9wpGn3D5lLlvh4
hW0W1TykV5xfQIVyiZTxz9h1Bb8Zn2qnUqgbn55SCFqvNApg9Jft8jVwAmpY1xiAAzJJIlX5klN1
wAaHxElfcjH6sFVJQX3knIMMBY92Erw3qQz6JUP/un6P+G0ja5Hd233PNPafZSuPs5HKWEYyJiby
55y0sPpyVfgc5REwO8M52AQYOboubjFILV3yaXGCgFdU9XSbMSn5AKEvOvYKOMC8jmXL7P43k26C
BCRvwbxD5srSvxgU1HA4v4B/rjC4GWP3NVZ+lEAvoIAfQ0Nz66RvY4crdqGc0Jbeqm7j0YXXD9aF
P/EkhrZudcchIP90rPPQcVc8bhZXMWs30GfvBUhXmn2lM56A9ou91YgNKI6jxphW32qxKX5vtedv
BOAnpvjZgUnSiq0zc40qgJkb4COBl8VsueRRzFavdYGkOO1j3OXM0MKMgbGqpmWDU9UF1JHYM+yh
129EqcPRdTR9uxpCkHnTVwmzJy0uP1pvutIRH7TQHLIvpIvtfIDq9XeLoBQO8xYI/RufRWJmWUBQ
ykGFlEXBSt3ra2zxLvuYXNcrVmrkHUs1vwbSg5LeKH8qMcT56vpKwHdXjc8duBGYGwzWr3Xp8SXv
9Fsci5qgguypDMWOVGKEk9wfTXIHg+AOBYz2RPlunuVtqngVqHYqoxa/g7qG2mK4WsC7TQFrhCXJ
HEtV8esFhox4ATZ+AyjDLo7T3fqB4OHs4bibj54lRspBDsvuNkNy6H8lFRjEqYyKg71VVDPNMc1+
wMaBDKJzUFZg15r1SM35fPNAcBITf1Cgv64DH8b+LtY1dMAU8s8de2kmAdXaqWmw7ulHQe6LCHpB
h9iIKw2Et3EMP5d7NfEBFmH8sj3Rkh2kOgG1aZNP/RKZtLXvLPuRBvJfBwIHH/yPYi3dMjCJisP4
9zFVtGxvLDCKlikSdIccqC8915tYTDg0pWGddrgtCk+Ra34DOy0wraSXuITugTi5/orxNbBj4L5W
1F+MOPWAnII7tQQ17iRw0mJ24hr3QyC2aSJdChwP3bLJiWUMxFdh9JTjEaGik61L33HyIs2HHVDL
Kuqdhxtx9oJaM5Az3mzHMiUHOZI9spIBXmnP+EqJtToipyvZgwZYe6nSBKKzi4EiMpWtTIAyiE1n
xN2IPGbLVIoBfieM6Rac9UX1h9TQUa2YoQT3Ai3ReBhCmIz9lrzxjTOnsL26qLS70xDS61i/ScUy
6jxT3H3itvUPxTCyjIUtp6ipeLjJ0Rb3687CpM98MyA+a5uNiiQikXkMd8478+KAi1U+8fF1Ow3U
+ns/G1p+EFFnCuY1r8RiGsc3co4mAwCZma0wXj6J7BfVV07DrODNRhZ+xyxd4cQapj7sM48qRPyw
jKz4bGkq5nGx2uOQhks7+3Pnhy+JjJdiVMqNSeX0U98OrC1ppiL5XlRl8jR6AGuYHTpJGXPbE1eu
Cgu1B50cb7HB++kYOAgf7ikfiTGC8btnkQUTxrZ6gOyfft35rTYDocO3B4DvK/raQhxj7ZA9kk5Y
kL6Ac81MHm3lscgBKMgIa8z0QoFdwiJKBH7t6JiyZCyNbpHyG/oMFCM9XA0KIDSOU9FJ7bwkg5LQ
btBDlRZvMoCjcpnBkzkp1ve3u4z3AAe/To7xoxmBrtqIPsTTNpZitqsOYmFqVj/feiq/IjxGl7nX
/YXeAgkbjsN+WicJjL1zzzxX9SOzRhIYr0x3i+mrA21Q6fV5uz0Nu9B16r5SN+qRAkoV+yvKbcFc
qZbMa2Jzs+YjWvGDxR0OWC596LoZCKCmMsLItPT33n0T0w2phpvBtMzcNvIMFq6OELu1OSNjUiBI
ZUNmCCapObdw77Vs3MGQfe4zseb6Bbq3Vh6eRz6PH1GCKCfQUCxt8/Ys1JJP/2zHPdlL+fGzwfQ3
PkcBM19vKLzAB0TymF+EGXS0yrnsqcDtZ0b9zwNfv5r+raFIMTOd6ZBuZ8lRu7u/GM3ymp7+lpem
Vvfc+x06ci2rYwu2aCgoEyxb2OvDl49shlaNG43Vya9kDiYyBbe3OcZwhMQxayrpodnkSJl2Uy9Y
GUoKHPy3GWZzmJz1hqGzHNonO0Tqbv4ZBVH13xP6kVO60R+hhliRSGOcQa1MXPAhTxCJlsE0AaLS
4Pxwp6aBJ5RP/K/9mejMu4ED4Q8QYQFL/owaf0hShx3VoTkUpwTh5bX4KsmL+j1IMwUdzSFtS9wX
spC58ZzJWtu1KOAghc6CTDASSczcYwcpDpHCjGzBRSNCb3UhLAib0eXynt2+/KRLM+uAIFDV2NH0
IwFEGJg33+I0Z9LwjXewj+CxtslqeGpVUp4aYeqtVdkxfU2CaHXQ879nSmxC4OFCqUWQBsgPQHBj
GDasVck1IdnTWj+0CKUwY8AZzy+4h7H4y9Qf1w946BJpneOw65PhqIGR9DqNYeyX+YKiWCr4mG61
VzVIO+Qj92ongagEjG4yzoqg6j/jDBxgVoBv488KSJCZWx/BVE2UA3X4WKuh9O4tkPZEvbw0Z9pO
2xPQ0JHbK/7fRdmaT1prRR+LazYR8FwCE+Rw3hAVoa7zzrT5WmyRWlV6J5sQRG5zL/X6VglGI25k
5ge0rXK0TDzWWqI+lQAyLTt7bpJNdp3SjB/wcnwBDEccX9S+pcT+4C30ei7AVyiAK/Je81SiKXnc
/7Ut6ch+aO+vj+YP2HmgEOyTmRNSC4QNoKtA/TOL36ZJ3NbYbpcM5vyTwSxxjXAepzn2LBOt6vQh
430Hbz8G0QpKP1lioqacqcvMw5ZLV6AgLqv94GSwoafBhjDz3Xk8KESvDN+AeQR/P+oIKKSIkX2U
naM1lq8PxiT1sT1dTeYf7sZVkh1vC1tv8DHZpC/saHvX4ExiTfjZR4Rby8k1g5Nnnso0ehJgpqAl
28LTlOmZYNkDpFxD/Eud1YzQSHHbx39vsqkrZ0sf8RfmQ8Q646bC/6fakABFUQ55psMnrScJARKp
FkiNmNykxsbYpH/FyHyZW/FR5EbY1BGe/3JaamEQTUcy5r4S/OyjQELqUDIsC2qolDMKLHgmlJRw
dsZijABVPuZu7xQ1S0FcfepWZ3HwIoYHu/nbqNwEP6JusP3nabOeW8Z3R+MsLaGT83rBYghj6F8d
cCkfvx/omE/oqjXHt71NL1w+IfrzLnnTIk2k/MNIxF3n+0KMkUV/MHBxHSt8l4gEQ8e162AeEa7y
65rV81BZcRD64GjKcUpRUlkN0pscmFv8zGSwijKak79zv/6Rvg9IG9iJnETPnf2rNZwxDUvpfFJF
6mkGX5TXvUrxXoxkl5NOcOU9ZVzXgmaMKcRUkRMzHx/A5kZrC7XWhusndefQbgIpoakgl3/dIX4Q
fpmBRK9PZlUbNHqFWelfznQETXGkZjcfh1Rn8rhJxkd/znLvgaC3jQ6u38irvJ1rT6/4RY1lhPA8
iNbHlz2iRRzSTUU0QS3BW/woIn367z3TEWApbIoXsaX4v7GD6w0AxlWFSrJb1jQeQAbUI6a2oOYd
rQ2oUPd1Iw9a36boQpPBVGmTG78TuMezI3UtZEgv3+7lRcpeUa1xuqPnFE0fwfoMNqdzJ/9Lw+VX
PXdrCdg45pA6EvHJbLp55STdxTyMKfKMXj+CRl2VrPNvso8hhxqJAs+KCYFezFw3XAZTCuZaGHW6
vA8SWq2pn6lFczaUmzBoYtFJZN3JMEq9nV9WjNGzYiPHvcSUwPL8NvjW3Z/SabrcFjqc5N38kML2
wXDtM09+9khW48xwIgLzFOTB6AtcQK634QjkxNZE4Vsn/d3jYP0++olptoVqXYRkIB+XQHLBsaUN
M5IxSxfK83FHmDmd6r40R0ZyOTgoK8Bx3SWmYqzdGvjipOTJV8tlDuQkureKOieD2LewEUpaEaYj
eKCQHGfChaL3tmq0ouaEFN/28LmLOiJ7Xe2B6xbp2ybO04tgWB/1QZiHqgox/EOwnpnzJGJq0Dlt
/Ov1wHjkRgbJ6yR8TueUrs7y1HTkaAzXU+dJRf6v6c5CU6wcQoQNd4tQbWbyiDYiU0dG7f7tAQmf
mR5Lli7kl/01YnU5yZi+kLbXvy6FVNDFfnWZCgAib0P/OjICd53WrOdBSAtTnO5KTceoBYuQT7Vp
feh9tVwPzdMjRiI36BNC2JTAKPkl7XZEn6HhJ75ws4CIAfBb7DwZN1590hA8QatR9gjegiVZLq2H
CyYP262Cj2KHZk6bb3POEc5BktUySHZ1L3UmCaPRT07gyEJab7Kn1KrZba2NFsLPRH/TTYHDUK2B
1Pi6ca7Tm4k+RFpi4jXZZ7UYQ05CJSrtBc9Sq1/DCY69CHCnkgxy7aBR1GJjbvNLKMyyb5qLUX2d
XTuDle4W6urDywtPlgAfLLeZWfGNR4oFZeabWVoeT9DRT5rUK2Hb7RvdfM1Nv66SK/NwdMIwhXqA
N3UjMeo4WF/8FOpXjAwKTSa2GJYE74LvO8EiHKB5irDviF8APT4dAC/qg53Rlt3rSrdRqY6E6Ck8
nn3IvCQ9/DgpiF6gD7H6tzrw8+19AUJfe+gEOW6frVmor0qPp0sWkDjMrAbiQe+Bb/96tlRUNt2T
90LfBiZ/kolzcI9+WyVKG0JsZwzOWRZnTAwVnVJgk5gnhWd0RqgP92oFHUS9G2HGfEXEnM3NUaP9
DIOinWaIbU/AcwVpDdzEnj3UR4IozSwXf2Fi0YwFnEDE6WgNZfjHOSxhOoNPDG3qBm33LLLyFl6k
RnuQ+tiDR9lXf1VaccATJwlO/gPoKKCWiZL+/ZdveydUI3I/mpita083mm+iahEjnCfS0KYQLUqR
SMUDW1AcUxRmgGxzDi/icX2ep8sgkX1gsvimJiNh/gUWLlImom/Mc51cnO9S60QBbBRIzn0H9XuN
fzfpWSqbRD00rue8Vavgdm9UT321Go9cR21hTEh/KTTp0DeMdW3v1VJ/KFX7zLXahb1eKcmEmSZY
dGhEOsjBmNyOVmOivCgoMfnTqhHvSjY6EfByAg6mNI3ykPVxfzqIVhmKaqaDTw1K2jADek6tsBw+
XISWXLUNkYyAj3C4Z5troePvYZ26iVF2+44R/70AwUHnoelkBfTBOuJsozkFWkSa9CBeBbgvS1Gp
7H2FK8bJQWvI+1PS5ljyrGnJ4k3IWINmfPeWuAUbfWhBxs8Z2k2UO/nQTZ4ro1jPs1/GMjDMvsFt
gdcqlTXuoo+ktaFciqQ6HNWLHzmxtkn4yq3Oa5qlRmDEtiO8thU9OlVzO9eJE6z4A9OUh6hG1PKa
Q6FzSHLtAy9JOKB/GI1PwmoY2080uEt8oMudAYwAaSTrh1c5et+/18dtp4hd4Z+4IvJgkkljQwzr
s1NaJxDyZjYbO6zLEFr2R2pXTxEQuD5DgVy77YPZmM6aJVRnV6RlqSioWPqwWQtxByGzbCAexnKP
I8hRgSzhoZ/SZOigtwcglyiR+KcwcY3pbQZBGzEqhZBVQZdc0052bDj2hsFOgL3svkskIVYXVz1m
c5gEn9H6R5BFMas/PZ2OiksIbiY2ZPe9o89i0l/GiVHBaFQV+VmgdYaIiL8TSonNj1U1rtOFe0Ne
vv4hV/CURkXbecBA+utut1ybvJBt4RaqROwWm2/KgSUKtUiN/mvGJwux1XdgWTwrC2c1D+2uBzqM
04g6a48Q3u5ojdP/LZN4yKRU7N1k/iROIR2jiO2DY2yWkkjiwOA0gHM39yi1GTd0WoEX9CDse6Ee
7mTy4YGr+PjKbwq4mpFbaEMZGak6c9Bt2wfNrZQz1LWLYTRVQgHHyxpVOi2W7/FRsmN8XYMmPywo
52LOBN/bXLkKq7zAG+gxVBBuJxQCBJtpSeB2B/sndMSg+VRwL0M0jUz3x8jDi78t3R504L8I81xb
Cr5FDnw2sxtmJLjtOrZ1cLJfhdmzFkwpOkyxbTwKYDl5GdX4++Al78fkrlV3q2AbJbcNlTL6hYeu
PpFPJf2c4JKcOd4Tw+n24k+a5NFtgJc//iClk9sMtegUVAJ2EgU+xu8AGWHV7hU5sR7UZ6aV2uWx
Cl4nJvsZAwAHKxnnOc2Pcc7PKYgruzW780xfiqqzXBCC1AJW+FbbRV7lydJgczHl5cV1xRnheGLR
HPt9T/tpQi2mOGJwKoVdlxRVdJe0J0g3yYTxyEAUCDp1F0G8+hLx9CT80dcu9CPWXc35bZ4mtqNc
i01jY0ZamKn6nYuAYWZjwlbFUy03EGZ0Y8X+Chm8aMT/1LgyqDuzaL0qr8OeOnLMN7/KkK1rdMCH
UCRYV2kpn/fJjuPEw/LuMgxLh4yunQ8kjq3QaXR6XG26e03y9Zv/n/eVp24+xB7a+1SQUBo3r9I5
Zkm/Aavo+VYi0YPcGfz1QrYKVMBelap3bMWN1KNw7Tc+OUex/NxxCfhJkN6t3iRh1fm0yyCn9wFI
7U8scOyC4MZxXpItwrGT9AWsy0p1q7HUYcTfjzCWICFwOg9zZXtZsShoPqsb4z+7BURRMmnw6p2c
eB0bIIrUuh97rZUCTpcHM9L5gbjhhQWkg8tbiJkeVyx7cbdIse8opjhvjl6ul3NAPtRiTB8Q87sV
aFuYAluLztQvhvWcG/XLAwQ/PvNqF4EwzVpfKrz2xEE3iDGO8Ps/jr3VSwiIxGrPyFhDKMrJr0tZ
4RE/PVDJ4PG+vqj2kdxIYiSLQBVGE4UJ74g7xip0e9fk+tnx7WicebYRqqPLIcPrUKrhj+Hz0U7w
p+yhBpHGxnwewuCdD9pE+FejtCZaOLhB4HU8btXFNQrnBmI3cGCn30dTUXEUNsxYoC7NcLavGOk6
d8GO71cDKcURaNI0UHtsIyYA9Y/y+WJ316D9zDIEW1F4ZfcMZwOWk3YJ29V2CKbJg2kBYteGOQMb
xH5sR4hJSgUP9DJnDjhAmRHnnmRmPKB48yNli+AlZgiMsrzEl9nno+HGdrpUW8xPyIzmWVoefuf8
trKr5GAwsJXB/QqZcAW6IpPNQGSc2tnenlj8A51bQiGoVsdlyP0TqY5GuMSKXGcS8f23+/H56uB6
WujHYV+sOOxKFL0vid/IXmSv1VyPFKGIwkwWOqSBmH8/aNd6X67cQAPYqyAWgld5HpHYxu/N+hql
SMUpuvxW6IuvkEzYzguMmv5gwbXefqewSPSDe+PWChVdmg+j4ZdXGvLtO2cEdIW9KJ6CR/NNSuMK
N7MzwfFkWQzNhxzSCgUC0+FJ8kozZGo7tseoM0FFAwXibP52oRBVMDpUOuiZzRIyQt9uig4zlwfz
daJ6u0BXf06V+jGND3Ou5a0WjCQ1qSCU8ZjOwV2mHcUQNLfdJqtqX7kzy8SZJJ1ZDjPWlJK/HPFX
vWHor2dmZ3iIfoAuJemV256XkAP5d6H7PfDsq/97mJvEBLE3LWE/s67M56QJlLpAqUoneacJhWlq
YFV0fTojyc99cmFt8oLbV59d4WM1wCWCZy71nSI4NcUF1UuFLBqjgaue8pOAifxnp3ySxWLF65nt
OPxr8KisklyNokQRtpTKfe8exFC8piHkmIkZge8pcFlSm34OUmR+sFElMUwb5uFhPPSJzHd/e4JR
SWd/+y/8dr9lNOGweUzHimwNcp2ZPrARHZIpEadsYWqUUal3lvFGF0jGDPH6U+9vPsKIPVF4WAQ4
1k2aMkKJTXC9aZsVNGsIbJtfq1/BXJXLLJU9bYInzPhSdEZ3bvbTXNqFFOwI61FEmBzGNxgfB5lH
+aBNDQJd4Bu0ZmOE4yymasUX5T+b+os6yHru7tNbuXKqHlbbrDAL4kNvM6N5hYmBjxnSToupJi+H
GoKnC90pUCEUZHSg9rWnN/tcCBHKK7TRnrton9KZzlfFSawMW21wSkVGpY5DZUe8oEXCeqopcGjp
qUxuT137/LgT9NbsuudkKmI5OzxVvaaaqCzDRpwSnngau50esTBGototvh575WtdmpGYRG3a9GgB
/FVeSiZcIyuPCEFRz7sVf6wizQS7f6PxFhophRDCC01Jap/ltalwcS8powJf1dMC1KM9LL3Jb9Qt
ithjxyn3V3EIuE6ITT7RU74o4NMNvOrWidw6jjaBGCsV6yX624UZizqaznwLBjdCiuKfmn5ONKMd
Vxgt2N9R+SJ47dDqYotKAUtMAGkAD8h4jqZN7ze2WiiCeATDu2vg8sZuhWy7bj9gfF3V3200wNUr
1C7aF0ql14KG45jOtP9Mr7zTkTWp4CFB6xkAgVtpIhSNyD+j25c/AhxF7EZ31pQqUWMVnQNiphXD
j90n8q9WIKuBDl/eI0WTsVY2PQ/I2eQ/edkaj0d6MhHv9q3b6rlnESXal0y+07El7bT9CAqt4PnW
LtFTh+yN0xicehuaKsbWmzq/JR95bsgFhbkuHOXyqyxX+MMuY0fZ4MN37BsRvfFRhUbRYQS4KqxC
eFX8U1uYmCLJHHqGIl0YcNNisLsHknuu+eJiwWleY/oDfCwNxWW7eOiYO0RSK4xRZvGeJoIv16UB
SEltoFU/W4SY/cPkbEUsHHhTYTIv+TsWuD535CNdNRlgkIgLD+pKIgiF5iErgpnNfyaXkZ0LGWap
GE87+7cTvolcVB6W48tmU9LGCJO6ftfzNpOWCM/BTmoM7M+fDtw2fsZwV/X+hXGJf3kqYPrD/qyA
Rj4tCb4OZ9vScovsN6jZY0K6gz5Sa6raHJBDkukTweMY3Q1PpvfM+WiaKXQMJJ3SPJgdc6S1yAnR
lFt+QuPQ6ODPFl3k3dyOEDy+xl5OLGAmStfm1gOj7R+jRJ49almqvvYuqHxtcirC8k1L8ndbnuWI
VpegeYb4DgrcIlojV6AJWjlrCHg9Z1YIXWnb8CFgvLRhXKAW1qP7NnP6VHomeVqKnDErv+V/tao9
2cMLB1RE43iCp1xnFh0vYMoGgHtwXPGYB6qRN0uHY5zrDvd0dXko8L4rkTCv+CypWT2jBP3jyFGH
A0YvQ0XcG3t3xEEj7pwtO6liBMz1K8E1jqY/DywHwsNWeb4qVv8/fCpIu8v1Mzjyythj99Fh8wmX
HVurUOL9mPYNSv9S1CQypCmQ5GtSAHQKXpBOV4mf6pIb075OV2SrC1txkSMwqnGb+AWybDERIQ+r
JUNOe3tefmi6FD/bxJZ5cLJx9PA7H2/iRNjOOTuqD9LH8vJcYmMKLsXhMT6kD6EAFt1qTEh+qi4e
IWtAlGfdv2cFLUy0gOITBitOmddI1VOK9838wcd3Q+kaIr57xh9K+k5QhIGOubbzPHJjbZ9LE9Vc
uBOSQK7QNwP4CWANzyQ2D7a6aIWzzc/wdFv6TiICwq8+IFDILXUF5Tho05S8JNMA6c7U44eYQywA
fsgYUfRH+Ze5o9QZCrWS2knhtRnxQC/kIJt7vlQQFBCoNr6Pko/WdQV4ySUeKEBeX0R3vfbkS7IA
muueRy8FpiObofccXoDmC3XTX90IMFiwew6CVPhJe7uTb2xEntJbhHJab8zQObt5gEKzfjkI7n0y
HIVdR0ECWlEqyJ/5m/488ZdkuvwhPBp8WVa+VxMR6EmHl6SayFs0hfH4MoMDy9WC1ijVk4gRZT85
uIMea0OppjxFFZfnX1npOn0Cn2nhCgjxMEeDbaR4OVY+pEkekYWJaeMquz/Hp8O0/0MHF9LmmuJM
qegb1VEwnIxhGUmAAfx9Q9ZztMuIQMEHjLrUsWf8WpX9dkAe6HC9MGM3/vogirn5JvEA3N9DzOnx
OoWhpNnm1q0v9fFL7oqQx2UUwE1jF3u+HNhIVW33DzGI44cNnTJsrujBNGdqXzCPJjkMcX6wEnkf
EZUxM50YgfDTTvCRXbAmw/OPjU+hzsBAFv6IRcH5B3Q8+R9anX9Tc35rQlyEEjIBSko5fhpHvEa6
dwtziTmVGFXAUjY1IxR8MOiPcACmQgAmCnS+xEOM+aISLasL61CmMCvNYfaHhHPwQrrnvgZygUJ2
AZ52remIQGu8VuhQ2Y4/v/uwpJ1MAm/1vGy22ZMf1zwoeim6R3M2iEnPKiAOJEqDL35ojyRKO4EJ
GztbifX0TtIobSS73F/B5JKDhblnB8R/H64cElMY39HjtPetwVzjllxJlZF0VB/r4x3qO9Fah54S
1X32Faq+5//oZ6OumFV6nqrKu3ITRZ74cAONNKbom1lDU7U8+spmf6oaipdUSzbXKyaGDb9rXHGt
ZeE0ejBx7szyHbk+K+yhDhEiPaYUr+YMjlSAY285dpN4St8LdD2Y5DFQ5O4bGIuwIx75gYA9yksd
HltMtfge68EZs6JlsyZbHWqBLeXx24/+QAQcMYdFcCCpuhmpvwoXbilSDUOd8jg7P2R9cCdpgMh9
WXMS2QmLdXzeWzq6M2zOYa5sQStryl9Zyjr+AuZTbc+wmk0z0iLRtTEvwm59VfSOT0sgFVUiHfdV
3ZGemdSSMvwqkCbPFWa/cyGgZg3WjkfW9L/o4zcfYiClAfclBnvRcN/RrvYKUC/QOwGWw+XoUvaa
77f44RPoEGb+17l2kte4+NalHkV3A1NoCUIWE+xAn3gfF7PtakbGFBtQHDqoE+vnpG39riCv1f8m
7fPpMhBvgM7rq8x+yfTPa9eJ+rnQFQuerGUNlVL+S+c+zfurSN7chTBoOmip+ll4tGJnw1G6g16f
/09tJdr93LWsU65+K5mQ77ID6lgFRynI6/Cguc/0CFEGch/8TOaOaMOUzuzzgk05MCD6E8fI6Puh
Xub2LlAjXDPfzN3e2Tf9P7ZfzdRabSxj+wGkKddo2nO4X6ZeM4Y60k/uHYOi2jgM0tIQUkJFcJhB
+Q9usqP/LHz+Yzd4UGukt+AH1uLyOERdeFUAvdsd3XC90Gq2J0HxDqP2nLd0vXIowblpTpgd1olD
xP1Uqk+ZKl304an1Ipc6m+wm42ro1GA6EXpzyx4q8gS5LXzet0vlSIFFmplF4mADzs5Lmd1qwx5O
rClQqHuTm6M9uDOXD4MSAtnQYiGsoo0nrPNfAJ+3tDDFf8rudUR8crS4h9CLYH8di5LihIqZNtt8
xwkfFwaf6IPgAnnuEfVOsPZ0bNKBbH8SL2chn8g4cpgVdkl0MP/xNCasRgoTpOnL8VuB6ePLHMG6
/FIt9xnvMOxxLC/IBv8NwTsa03CGg/Ejia7/8kFdJLUKhZziLWxluUGWmvNrd865IBsGEhElr8B7
TbMrjCEHzqOri2TaN+F++T4tgQLMPLunsb+Ns2ujyx3v3x6hZdIOLS08RRiKBqpdTW7v4wGGkg1N
44QaJVfgyfj2EyZ0jix69uQ2ZqxQWpn7pYYtCii6ELNBUwpY7rBnH0KdKI0WT1qkGTnKcDKhAbWW
n5cN+Ulu5RbjYYCA+iF6PsM0AaSoRpY3/FkY6wXgS8lqC9+F8T1hh+13l3+LNZav4ShFNbtZhS/6
X9ZXDAS86tab17hDN/WjS5xhUUg2kHnQCWWQyIgMc2EqoFxxTIhnCjKN1OHxz2mocyC15nmZUO7N
qsHWs4u1D1gctLsnQeiBjVRlP0VnyhGrMiOKrxnM5n1r6B1PYB7rsShI1QvAHCtjf2EPvVi6xO1S
5d/arkfvUC4rEtZaennyxENcsAaV7WSAsTOxe/QhprnlJ+ZuZxdKltOH+ELaE1JkiMQbK4bw3Jy+
OhGyqsDLBuxr1Rj3ZnQ/dV34DSwOYcUG+TqZrYWSN10gJPEs1W+2FKAohSOmTYmiTdZqZEqKCBf8
rMEp4zyrENzccOpRs5pqoHPzPeCKnBqq00hXFZCpIKAKDeArpC3gyMk07JCCNL0WxGUGqhkKBeWZ
E1YQBsXBs0JAfoGl6eXAjiPSKn8Nu4itePG8zSpwuLnwqlPB6yc5Xhr2NXixmcJm5Z8oum2X0hvD
MY2XOuN9Fcq3tyMPQv4UcjpJU76PjnVraXthEHdpilkDyuhqNb0dRMKi5t/saL/+JSwf3mpHgqLO
tOzceqVc+kbeCXId8IJzApA429vG/pYPjwf+KUcfsxvrPlovepG/kWlp0oGD57zCaQmz1bXYzdlw
MNYY56AHsjfvdmDq8P99cqbNhzuSI6tAnR8awuTWYkMp+KGdOweZaNvTVdW2wwcsdAwwIIh6FjeF
6WFYPEzjSFnKpTk9jXHHMN1/SadukgSncHtWNYSDYLSIKU5pkXiOStAMQELfegGj4eJrMG+7vpEm
tX1Fbfhq6nCiL8VIrmGf5GtW9ZECVfyYfiL+99+4XjG6qGZMfIcbF/MY7sDZNUU1b92S/rRA26w4
Pzw3RVXIQ3ud6tf5eSbD/saaA49Ppga8mWqGGUbsaLyFr8+SA2iQ2GBqCwxdfBoTds4E/WvaTT5t
Pmt4lc1eJpUqMYlX35YQ0khVEILztn3rzPLrlK3L1sqqE6iLF+BIF75Cyx+ch14Urc8YDavBuqQW
xKvSVgwInYy+QvF2Ckhq/Fi1CRuD3zyxvuqxils4y5kvMVSSamhOH5X/VC/FTzmxlpe8Nl1QvuX2
3TjHc+ysUP5OlmXnDvbXQlJtgP2Ewj3SU+Ap9UiY+aoN5WMiKDLkBM8REorwQ8YjWp9OywFVcYaj
E9TIuD6o4z4AyleMyaLSVsu0O7fCt0MioFS0/sDpWMh1qW5EyTTGKGezkPr3oR/kRGLdZ2Eulxt6
SI4ouU+5Pzqq6OUMEXrgPA7zjZthQtVFG6xmH/kNtZpz7TnPwx35Fszms3+x28rM7uMA7PvtOHi4
+Ca+CH1IdsBwBW8yMLDCtEPB92ja7tVfjim5hBBrfNs5fJgIHygG9GlNvM53Ov31sRXvmcBZ2/H7
dE17lPJD3ADQCZq3mgaqWJ6e5DjiH7OwDvGdBgfjLIGQrxzb8y/W9IKFHw5JtJWkb/VMm596fNgB
om0MNZCR13EkwclHriwRCHWns809s66pqwKwy4Glj5qaY3PKXTI58W6F6wL2v/FkpM1uuN5aFzhK
pNbjwCX84MRHWXWMPssVpVEBY1MMtWhrm3Bi0fUovO7obujTkqZg+kXLwSPr+VQ2lt8tbtSS85NB
g03dIKO21QXqd4Fa2UE6EDI9Co6nzJRADU1v+Lmxi5IHzgxnw5fKFjUGMnSBs/pQMHIFyhjy5wig
hGElp5dBZ3XJ4p1W+VfrbuKupUiUxDe89gE26Cx9GC22mhKa2y7yVnG8rT4t6UqU+iDPawIYvmQr
XJIsm88dFJ3oSEiC3q6/b16g8Khv+tJGLXXJG2zP1ifzt9sGpKOk8tzH+igTOSfti8qFJ0A8lbUO
Ff5h/wiVUOLC8rIm2iVg1S4MXPmMXIdo9zupdYT05lukUkxPvKblUxYVTjIa7zykPYH1eMQMK7Xk
l+4Soc2c/UXrDVI/CPWMilzJqFoRpdOT2anFEW62a66NLvYi4OCoTEdVsQ1wWAw1eDLSxwpnNXMS
SJGce4dd+SChjq6/o8dBFm7jy4KAjoK1Q6lv+F0KlIIBzV1/RX7Fi6QnL5ELLTvSa9zAED14gmOp
i+nbAIdxjZZSNTmGmeEcWNcyB27yqQILdQB83U8MsJGyNHZ1AQvdaHJCsF/uIUOARA0/9jdodKFL
dfPcUVcdgHhwpYMxDBOqBuPO6MaeZanJ6d8ibHwjyo0XHIBDKqYpdnuZP2dp49ta5v8b8SHXsRnx
tCVkAj7h3tj/g6kB+EIcxn8ETl6kO7l5O2kV02K2F87S0Qxlv7VDAy7xBQakIWVEatfQ/GDuAIIi
ykm7YiRdOMXIgDrDIde9IdvtiUbFTJSzHV1WUesmJZ55sOy70/c6w+6Gg5wnLpbsAJ3wDEbDaoJm
IoIM6fhBnXb2BU2+VutnUT6xGXK2g/Ma6BmTuhgtfcdVgwd0OpkqcLQcLH22iCDPwo73AiGcGa6i
x7cHx1SjdawHBbZMwi/WXTRn6lUHEBlJb104SQiad6hLjjaavY4PI5Q4BoWUzujmbW4Cyb2LNgGO
UNe74a0ORJh0lt6vmavF5gE8d0bMDfwdtksgAusX2TyzFlpDULA+nb91ubeUF0o2jzrKsgmvEvqf
j2/yhnnbwRdDC4q+aUNITqGzoS231fesKAlbL0bV9XfMSY0FMQ/bK0Xh5X4SIzXSgK7CAO6wHwyY
xWPtE4C7kWnmk8Ov8nwHDsDZ38/ek2biunpIsmm5qPN3kWOYAtgdfMEtifZUC+M9qslMnEcYJPFt
uMBuRQdrmHH9W2MHBexPsvDZdUQfM/LLSTAF/Se0CdbANdgHhOZhArhlwAaMre0DYfobfJviMLdF
QufFTJpxohuubUeBFB+bYeq8ccTsLbq0Fmxeh2yMW8bc4rDvH6Ya+fTspc1zKmWdrz7CjR2jaezn
hUiqZfQOYkcT3bNwl6suyTAtV7EuKMGHd6xwDpXkJst3MYwCKlRer0LxoiWxv3YnDBqbogdseHSw
4J6lNSgS4neFLM4+t+g6/pSm5HVRUk1v8LKmjkFdYDfJaRKgbuN0+uvM25k9akSOgoUlXQSjD3Sw
cL+mHTvODZNz1EFATf/OhYtEDM0OJBsd7nBNT46kU2gYZO1fp/4ITRlkDlYYy/C655p9eAtfHet4
R7td8oHgOfF3xX/AZuvY4lUMnp+Ses3du07uwCkWX7gXi4+DO6a2ucHq4mVx9QR6SQjNy3AtP9yZ
IqT/2Wml66LbyhMcjdxhBkXGQNVIIQC5AuFzWS9fsL5XzI3YgckXSgjghApagN6HpQOtVohbPTil
vpwyO0vu7GK8XB0e/3pOA/QeYDrKPhLr1O1fRk1rvyIR//3xHO94UFdStcKg5Sv8WJ7Z3jMfnBZQ
319vXwQm5qcCX2gtQXAbTfhslGW1/fDBgUK7+StRDH7h2/crSrliqTltm7CdmVXxjUvYac9MeQ3H
6o16TuXPB4ek28n3bhQXlFyV8xJSLmCMQLzWoExTII1Ch3OJLY091BnszWiET4UuOGqafyaJWw0W
2K1UFw1DoE7pLzFaV7swlwSRH6lmd5GFTlo0VxbwieunDt4JU3Hg/y90lz4hohE80OryM2RtAdAv
qKJkcWi2PfaIUI2VryeU93X2z9QewCrboHww91tIQyGgi4piIl1cLDHmIpGQJg64P6NrhZ+HW9ro
bBAcX/B3Rv/5GS8PaefLICeE14mCshqhHBK5BfadYwSQfVX0C+eEHI8NG3Kx2dfRNyTKg3SqQ0Kb
22wQxDyqmxdNWT2WOTBl0GNDLENtvYuWWLTWm3yrlnjXIp9hV9mT60hscloXdkEvGUTAQLnTshkV
YFyq1XVBGgI4RFpO/1pPlu6SB+3OZ0yOn9PSLcI4oWrPiL5UJYUmR9auJiuqS4NzmMGs5NGSLFso
wvGaBInkpylAjYeIOsz9+9iCnwXJXrwkv75KNhFQuL/kH0uQ93ecV6iYuhBaWfV/kqC1S/JVwVu7
kCYJa8mnHQgM2Yjho5+37Q3SJSeJLuGDEe9TaM9KdW4whdxYySoQk0ird1PDmCdArEzBRKviskVq
yKWUIAKRyn01CdXlDlzYEg8gM2qaItXoKOSc1Gjenl/RM493rw5aY4WwHPBm1joW9WxKZBD+EKaN
LKORjSGu8DU7XrTWdPZHDz/S0osT1fpdj+7kybXceNtLiRhSzG7uQiMhyXUzhTOXlGcxGw3IYrVx
t3Vx0DoAFNyy4hg8huPjxNR+L1lWSaXwYyD0QphQO+Vsj2ndF1+Xiee1kvg4/RcRhbe/ShMBxnZk
pTWO94ZiYTneCQGMiAvZBlahmAYdFxideGqKo0+PuOnmttm7wmdIlW0qIUz5HqKbqa1MdCt3DPGj
gPOFUD+a1tNoxRF34SuDeqKKjkHKUX2OAwwzLaUhhuoG7n9EbLbJ1i1VlaODknCdBqwK3c90UbS8
6YtKcTtAodBsYFxcRG0MyRLhuGDE8RvapcgBruUPBQxc3iLrLubl0zk9CR9y4Kz/Sqw1RGO/rIkn
mXKunJIMW4eUt9WaWR60ylVQt/nYJzblOZY1XBbNmpDeywu+8jz+UemsYBI+2uqHLSUtKuvozuaz
LYT5lQE079/0HmcWjRKH0Mj3NpwA8Yqpo97bm3GOHE176zPflEL9wOFre5y4/PCDG20x8BT696LE
Iqy5kM7EbaagXGjf8zJdU6LZiTYQq4q87gweb9Pm8t9RuAinujY5K/nUH4ScJ4PwtXdYC3Hf5EQL
OkV9EX3zCcwgmJfZ5I8XhxLZ8XN0ybIUz6JOvncM0Bmi4PoFm6a0VQ2EOe+yGz6Vw0zZshKA3gDx
D3jPuiBjvAJIarYVVnM/FwZ2IpwjQULtT0OtDBszslwpgpY5aWTiFns+TZqeflOo13F+AZlcI4o1
/lDKrUJARBQnCi6JY4PV7J4qWpiTMlFqRCHjZ84qV+KUz3DL+uyfLYMgftbiZIZqw0WcA6gSPq8o
6xQQT1IxeF8z3x7kQv9zokeUbd41rFwhx728L62WsbYIOgpcnYEvuhM8kfcb3HRWtfKWcywvtnI6
Uqb3S6UOtFX2PoUOEr0/B23iCXK9ctu5j2DYvwt+xGUcym84JecUnMOiQ8/t45CbUfZJ7JJ7dm72
sGlzbLd95D3RlaHFYD85qmL4StODCuMAxIZwYpDoQ47hqsne+eU21q2LT7CyFO3IQQgrtWHVwC3o
JLCs9CJ2CLuKpVVcqGVX5oeq66c7se2OkP+aiehoHQx3nQkD2yG2juoYLQ0AxpE9tJFx0MjTQg4n
bY+ajIyYn5enkDkj0hYEaL9+ECLwL6ThXpjuLXm51hPDSW4BMv++yqGAFIrmFejhxq3smtnAkmGP
Eet3mK95BhYjvbX4pGRYQ8bH/gwrbjgaI83y43rcCaenU6sNgmuhBfMyPpCOZqe1v68u+cQ9TJjh
5MnfUxNMtFfBZNAH0NQ8dGeJo9W1cyWCztClSQg3KiNjDXN1UOgNMi32397qNreNphbjDtHXMWIN
NiwNYAtGMczu3fxGVTlQxvYuLwFI7TTNfVq6BjXpVB/wsuxEz0vT0SXAQ3NgRrfjZ72GHkrBn7Ml
VX+gR5g4oN19QI2FNjnfaNem3TU7KIm/4b3bJFOUcN47iuvMv2WqbrowpDpZIGAPqreLjLVNRSSu
BbK1eUobXAfVrJYbf/PSp5NZY3EYK3/QPMjIU49cxo1iDFomBB/Gy/blmP53WUqI9myuDlbHFwpk
6LfCYs9MeKN1tz9guLo+wT8fDWD6Ulrg7krZf4zR/pDVVg6dAkIMuwUyY73VGWoWvqTkIJKLfDRT
Bygd+mXwIJz6wu1r/9mHi7rqvfOFnAOd48Su73ifQHzi1UFBWNbBborujPQGHD+3JFC/hALQnNhG
xZhORFQWi/WYhad3OMlLPljlxiEVJQ2JkvSIVTr3SMYnF2UgtGVAKeSCU/J0BXLx3leZV+G9GQ6m
7O2j/LV5U2ZFGAiDHjWIXzYqHZNZSFjWvXt08NnrwkqcPlvTbTe2Fi6Gbc3V71G6LaynL46SlvXk
DrCz13animKNVX5jzdwXPrRjmLO9iQeNZwOY2N0fm0ItoztnRes9bBIPd2j//cs2IIg/Qc0xgqkZ
Uwnz++7xz05yLavMiEA2SggY8WlqDeEs80EYlwGgk8BgDEy+j28TmcBWhGDt8ZrdDOibNVk3fZPe
PVvJp02s7MO+sxjPeZxn/vYqi9+J9wh37GG/UKxldN6tFYVSYWwLkcJxYxbYFxvoikOdx95ODtwl
Q/xqFI9v8OOM6HW11xKHCotOYD9bE6IO2osV++D2LVdU1obmfewLNySfdg2D5qyuN657K/40rnvx
rjGbnwNb+eTHS/WjWon3RoJagfh1yuFMKVKoxwPhQCso2Ml0oYjU6ZWl1AI1yHzMrl7EuU+Dm7L3
CIc9w++MV89NDtN1mSutyai/RzwicXSukCs7CD91iJyE/Hg9D0KPfVYsIMXMlXh2OdDkS6/Q/63N
EDtnt/ZBzmy8NmoaWzxXA9WeiYxgQaLNdnNhW7pvgXbALQj77+N9d2xevnCwqggVg1QiQ71XJiuh
1QBHtA4OVEq204yK9/tzZ2auDOAxDiwE6bnVHzKiVDpSINAxJoQlAUrU2WOobkQlZt0BGBY+cvl9
jN2HsrcOdGnQ+8d3E3Xv3cBNpa2zlIssI54K0iT+9Hwwt7BClZ/DweVN1PDOY5k9dLHahTiGwREC
ZRrSdFCwP9WSgi6iCNP0Okz1pRPwP0SlokTFNNZB6yr718ckf2rAIUxHiMGXvr5tTh/WWcLNsfrX
WlkcYpaT1TNw2KOJvP/doCQ+H9L4yXgNiSbDglBTJII10+FkLGTVafnB/VWT8qtAL5nmJT1anQhl
XW7fXZNdiQb3Td5B+kguO+pv81cNbtpckpKl0rHkLlXXgJfRki8s3QYl+F9x5EkTGp6/YJmLbhRz
aEx63HmlS4xOxDDEjbLm6A+GHvQ+MwN0l2BgCnk8oDB/yOVFXUkiC9Bcrke2QNOw5pqfpk9cWokm
LfUgKWaHEHoXdysUo3KtklEqthS6Vqz8Kmk2XfXCD4ucXumXgzhqABnnRabNq5DrNnojCfTtGdHo
XOZWuGKevs0qvk3fCw9FLUggRriehP1vXhn8utbwddbdhyHsogv/o4p/fsac8eYP4D9dq/HW307T
NooNwa5zAmPMES3voVaRAkhFuh34nuFozeQMwd6/J/ctmm/c0p1lVYDTYhDfscb8HcF+5sih5EUP
c+hb+D+E5l0T5I+6QfK0h7tpGn0iuxkYwRXV28rg+D1z8N5dlMDrKVmZhdWlzy3gFQ+hIXNfKgtz
UPLIguDqMdsyVRmdjRyvATjfs2b0gbVLtTpCZPVaQKGMUoPcjunOEj9mmQmjX/52CqHovwF6m8j5
Z0QGljmrVtN3fhxIPIezwhmsVkoEhbvX4i/fTMpl5LrC9bhh0ztkL7+XRbGz89OMX6izRJVYQgrM
yIXZvcjqqzyqSDnvaqQAlu+sHKVh10ofLO7IJC2SEEQsRbuV/vikiMWxb1jZXPHx0tTGXQAx1nRI
1Lfi2r5kX3ZMceiBPJD2jGZPZhS79MHAnZR2+N2DcBOWLVhSHc8JMZ9boBq7LwfA1JrhyRuEwPSi
DGm0mKqjTIidrtxquYLxjrW8k56BmZ9uGVYbP7WOqnyNllc0hTsN9OpAMcFW0p3/E1LHeo9AJAoe
35pHasNVpWIQFmzG3XkvCCpr1C/SZghl1bMr03DNXwUdZGDjOvdeHtFN3g2a5wDjaqmowCH/D4l6
9c8Gs/gE7BpEiUUam2NwLyG422qBumHgWmQopmSOKblCDNL6ApJfuYeDfcLunbmznJjj/oisasS5
ZHd6wcMfOHsxwBGIY9XrBSCjMkpdwjynb0zUYgs2f4Jwn19H3zLwCHdf1UKcKjmI7+4DVOQAeOBr
9+SjIs6B51qVFuYvMw++nngkbAS5Ddy+7XUREICEemkMXoytFKsbdHbk97lmj42qD3/KZiiDDLBo
Xku8AXbcsZCEQuM6hcm5nBBC6YFfoeFtNgLRaF68BpT/tfp63g2Zv34wCym4bSPu5bZfAx84tknm
QLNbCAW9V1OAP/70qxD52B+D2BJhhLcTh1+SP6Ul6V9e2wFVNZ18iU64JcshT+67oozOz252NEjf
SyhKkgGQvgjxS5NhrCMOmFMu7P02JZBLpfhH3TDsDbReSkV5axCY9gauJp77Vf9ogHd4QxBgP+PL
JGut2e96NoRcZpRqvNDlJoJfBuwGcH2WZrKHCObENf0JDqxCGU/gxxvp02rv9c5h+QTCVGxrix45
AxNfjcJmaXTjJVNdEwk8OoL0eCo8+OVYdXxiaxB/V+eniOIR6ChZA712klxo3BRzwsJww7JKP2Bt
/nJAk8T8kmCED51k3PIzRCm6eJL+oqxZDeUwginwsc21tAOkVo1IEtuCO3YAtEVmk2YqmrXFpRZO
nohJidKOuS7/JQxHUt+MNtaNYcZ7EcXy8QhizoPhf5nG3+2lmgSrSXWrRzL0odDDbCoQoM7qSFQO
RjEwFBx9UPxWNRxwAeMjNeX9niSj8sWmTKRrYHb33ZR7PYowxn7MrYEEuUDOfdA8e7UOCU3uBdQB
+bTJmwNnOtkA1L+plgDR7dU0lBbdy9os/CR18kW9OPmWCAFVRnQ6VxYiWkPvkGyiF80wjDoCmXoq
dpYBFDNnGIVfh9J7onfbre0AIQqNV9hNYAkcM/fYp8GuPtnSXrtI9oj8KDs3ErbBE4qAaS+Vcacq
l5ofwcM2cpGdU/ZhBY1QRktvkkI6CyNfYUWeLr34Zl+kh0BovSxkZoGmVcWr86/DYWFCACXWqy2t
YBwMyBOGZIjDdpjCzCQfcZdEU122269VF8BvrCFFB2xzyhkdztvSD4pv7XR6Q1o1sD2FJO19ny78
rXeacjCMykOwyPHSx1D8xzzzCDupU5TBzMLmEAPT57RXyD0it3wJhbXy3v2U5Tq64rJb19+dYz94
FycgNt5I26u30dWL+ceJtMySNy8SI8FIx/62U3q2eLJj0qWVLa3i89roCftZoyA8HQXOnN/xifAP
5INWFjP4rv123v2LjWgZfowIwBkDoGOVDoWXgtfBo0mbaUZuvPaSJPbVQ0o3KjTj4KWwoquzbym8
eeQXaE9zP/VPea0YQ7OpvBionMOCkd66bE+s3tSM4bMDQTWjip5SNHEWvCszY6C5LKyrK7j65aAX
xXTY9xV2bRpdpRRw+ThVuQcoTLmI360luSa36R6KXlJPEU63MFhTYMRDA7U90AQ4z7t4VSnSwPxU
h0JBBKp6fP0ocDh/Ia+lkSgAcWTiMNL7wxmsO2KncbN7yJ2gbR2gDpzUPsJC/UXcFTod8BVia/hN
rH0QK8FPjPPznTu2w+fIDgkSy1ZqVD2gmiJ8ksjInL9hwagaTMdc9eH0H135XZU1WdoZyglaOfgx
zH7S3mIVt7+FgCG3MAOzRRUisVlzEMAMhik3XxWGocyEdyKriYgTdBdJk+BgDglqJts3fIgzC2Qp
jHx3/PfECty3PecU9/ign5mAmSik8UuXFZHsWYh59o2I18QUtKQnEk4nNWTY4MMsw7OLvISKynqO
xrb23ze/hDoex/SJRnQMR6+ku/sZcW/2HX3j7IdOllsyDFNRtKb6W87gqo377E/Ru5DKA5aS5OBz
EjMsatrUy6bHJWRBu2IDFkhzAZ+Gf2ThTSEdwWoOm8Dd14v+5snAoHH0xX0LrAnbNpThumkIeaba
l54vqZaAs+ELC07dUQcP0+LcDW+SJarEkwc1ScfplPXvCQS/2bgGlx1oYS0A7yD513l2ZTUQaB8Z
f8hQq8TBxLiE2BRofQsbelqg1lbDfWpDM+31zld+ZCzve/EHbxuwpApRjlc5mQ7SEYAGnrqary1G
uuOL0uIFRsSUBTvFXZnictWkuknRLmwN4sTymNf9Qlh7y1XuSzmwDPBOPgUtEtXH3fCrzdS2oHAL
GyIx1mX4TpQB65kJWBZoHb147fpR51KutOUVcpwXHh+GIXUmaFyAlNSjeMtWIysKFihteMDsyMjK
pQPuqBsjJM1ZkWZN21w7jviRErqHoPWPv/9KARXZ0kJDE29C1ecem8P0QtG7Nd4W4Nm9fbBJIJUQ
bf/Dw3Q0ONKMG1V2lpz7vjs6fDe3d7MAw5GWU/BlvB22ZY9NEp4Q2w7ZoDMx9R8LzbNXxgEpnjio
hVJ8CyfZ3mY9wfSZQrEgRt1ZKpymnvJpEDRE4W3d/UUZoQFOs0SyX34Wdm+60hn5YnLfsHyPo+Dq
HCL0iA3KtceUc+5XAzWWmZmPAO1ozX0Tgi3/bLGf1oyY3NsnAAj/rZFN4HMDEmbabBl2lvGlr4QO
ZhlRMim6uVcOL6ZItfnjVMiL8bkX2VbcoAS1JVAJkpOGypJIc5OEaHZLp6izpz9JdkiPvTKzE4mW
12utLdpwW04dFXURxyz7BkwMXbLOMuDN/37AFsqjKNYYbkaDSFwNB0ogBbEW6Xe5QZLJgtnOjQok
d2DDYtPIqXtQjUDdxB1wvNVONLL30C17nRLCd+0O8xaYT0BWX36p7iVWKPZLej1CZrY+9RJJA5jY
QBsDYq6aWfgyTY+3jOfA8TwKYckcjD9iaEwAK/fuEK/rFvHbnFTJ4p9GUIua0OOL6U2p4gUQ6RfP
6AtZNwhhKaGuCqJ+ZjOtOKqb1FfFZolZW5wVBM39EHoaQrFqdcbGHW3P/rTdYtfFF5azkb10y2jK
wcpcRj8cwefwerjfelO5xhz8UQw/4zaM67kapJB0eEjOkoOOgN73OZWymB4esL83VOEDmUqjF3mu
nSJOFkSjGsfnvCI541dXxCKmfpkh9ks4RSRNAzjMv547OCLZFPM8V5vAXJQFXFyrTsWC/dpytoWo
ImVNHUXHvfYF58NpFTnQmgiZP3GIisewyuWmt8E++J0BIkFSeSCHOxfAlvfiaX5dNoLp57XBYErJ
0GQ2W/MAp94jpRWYCQxp93iNyKhM7ib3Csswo8zd6Don84ITtW0kR5BupCylDrAdupqqjNoM0SjY
PV8Q26TAjt3erAl4FOzmy9gnaR2sAOaLm7UBhDMpE1+jbbDNEBEc683IERiQ2gJqkzn0uepMcyE2
N8qkyIS9NH0rta2gBWy2gxkhrzlb5cwthHlhUoWviaLU58knGQ2nS2f3iUsEEJS1PUwaNXmpKdJT
Yn6oUJJMqRnECd/8eClBWXcAdBraDG7/p1AhT7LeACsYsap94D5tm6Oiglf+02VafrFvYSEk05S3
Ex5K5qZXhYowNScfkRN4GuSAMIYL34Gh4qQVacJ6jsT23ZXl/RXUBumyMhAB1ad1i2mRLu2pZTPD
fTtqJyCg7dh7nBFDoZe+x7vEYEWK8p4I8VKHuYuECieC0f1C4RYjkfj2EtnyQb4BHosul5naCfuZ
UtHQiFy6jNgsPsP2XiQvJ/q5loK8ncPD9NvFAw1a2z13Yh9GZUO2l9BWKEwW3Q14NedgkFhakUIW
v7Gttt1Mqs5ix5/zoQJzXz386UzKwXSwZ5PZ83Xj3WdgfYwtSn8SAhb2opO1w11FEsT1b8bp30q1
YqZQ/ldETEQB3ddwycu1P972JdrRKHDdvB8c8XoXCfCIIW+79DXaxcVnDywIVeDevwpgRYMI1o5F
Qwx6pswjNdw3JJ3F9Dtc6tdo8tjDgdbKm2JPVcxNyadOrRU5DHepna/SIgw6qwB5Yps4zME9qhZ0
1JAArNLrFT+5112it0hmtmQFpx86dmniwHPyg+LbTKtmlgb1joCaWLHZN9BdXIfINTJnXYIAZYpQ
4je4rMZKWCpVy/fUtdw5w5/UAC7a8D83zdE43AKYQVQD61mCRGLpHZtk+ChLT/HJouds8y7xfGZq
e2nxkVpU7gqL46Gt4aIzqa4d6MmCgLHXXeL/pRglxyhseaqwBurE1tXo+NrTzXXSJiTSX26yzhZ2
Zu2gVhtWMEKe4QalLqhodn00uqaAxx7iPnTPtm/JZnkXgvjkamLpc4ov7SK+S3+QtooLlsEsWrHl
cctIHX43C4F9pNd9V1VQTmRBBwrawZq37/UBH9oDDlCpYqGXIpRKufKZQBDqvzns/L8/GBnQLAMY
vQiveRsyFwKMkuutp5AHWxGJgzPfbAXp+MiXW52fGNDSvp0V/ffbkf3SR4i71jFgt+1nHOd1Olqo
ob45EqqvdsUUy8iyYtryXjByV7lvgJqXCP1mNdJMWZktkH9nuZGSbWCcDjXkUG3S287DQSdpXd9/
foU4PbCx22T6SqhpKQk3P6tlhHEdm5C8j06UyvX7ADjii9/FeR+eCIM4StoOG8NdZjmHQEDup1UZ
/NWL6CmpQ03JtAJLe3WbasYp2t+WT9IyrRQNKmklElMGlfe8Vsu1oeDa1IS+t8afFPI+LbBP2Pti
jAO+i+LjFLv93AXWV8tsn5mWxVBMw7YPwDhUzgW9KTe9CqeBJgoPI8LLKRz6PDLncZt5b7IC8F7P
mESacs626qsCFxGodZ8fm/hUIbE/XRduQ+FZKIgOI2+EpG8S9FQVQZ5y6vCWlYQBKN+D2FkdmW/T
Bi0V2veghvC7DGQuG1M2b62cGVXd1vyPB7KXZmcY297Ue6pMo0x5yhtSOgM1xu4RiU1f/u+D3vqo
ytZqOvR7BL3qiq/1UogzJkqiStGC+iAvNXBGk/DlzWS9S25v84ssfWUVrNO4hI/Ec+zZYoPEp+M/
BfJ6qFVDXP2qUlTdUe8JAgFgDjApIUO2Mo9T/Z4w2l/cMfR7e4/57LHQZoCDZm1/hM/5mtyT/3Cx
buAvq0OLeRiIgziHBYpYHdgzOqwyKfLBI77EClnDYmQTj636DmsmfGPVye+IMUU1696Sahu8Y0r6
lGa9nX4EJY1hH7K3ToYGkuGs0jqIMXbQzGvg+ZGfObtaWgzafqsJPVXcBNoMs2Nz6hXGE3Ah/Ip4
YqTTsBlsFGXrhAJnL7GHMumFb38fqXj/DThcUY4nhPeFkY3ESwVkDzQ4mbTZCj6ON0WTjbpmDzeN
15oA97/hhRfGd4+dO2sE8MHZHo0ePBnbqnd1mCjLPHiyOx0qN6MDibG10TkYUgXV0Sy+xWNLPeC/
Jz38bfExQPRaH8ZcVpzU55svfRA949Rxw1WF3uoIUQCYPsbECFhCqVeEy3HxhD0+MsD3aqyh8p+q
VXR9vgauIifx1zMcxcq1ka6i4B8tvKbE49v4WkLtBkHlN7iVB4HuKquHbvb/IoZCnkNBwp9GyOpv
Pr1Hx4tMsRBik5L3CFX377dTvqiGNvkB3DAMeVO73j0XWJ+2L91UiAgRe1uW/atsMzXYXU93I/qr
PPSjqySUJ0t5CHXYZN+3hSZ8hCyfrR6PHQp58x0CPiqtifq/QAIxoh6lv8DZnquR4+vDO88l39C5
McfaLJnp7dJni+MC1PkfHLQKleeyjjuWvBli27sHXf7GMjoiZ89Rg2CAWbhdYHJcvIHJVUCCPamN
rDbEYzuQsoN3OX8hgP7ERWspHwYQUghzEdxbPGoRzvpbJkqKFAkkW26sZfz29t9601F/8Wdqt3mh
GzXJXa0ljwX3AT0rlGGOnVZjUhPufUGhDH0OX8htWX4zoUj2imcT/RDghHab5rWUbRK7Qa2Vn9Vq
Ru5Lkf2zShB+3jL2fM7WMEQQAk5QSWk5fuGJH5qjI3qBtgJ3i1xFIdrPa4EbguMVoEE5VOBnGqV4
N6+fKjDc9l4l9vgTab0illqdEINlnZ8SHBz8RmDvxOflo1n3ZGR6E2gJBkevkxpHz5dAqP0SXz+0
9ttqNOfMWpZhKXJwCOlSz79eNfhO0uKj9alwoE+sWvhulv4GPqFOXXu1UPIRtUj1gBmmfZzms37y
ayjJKKxwp/JfdTGbPB6o9e6PBZ4XSWH5Qac6M0kv1tSg6N4DCg1NkI7vi0dDz/ZxayzoAMUNkt4u
wqm+YwxDkLszRI97mw6QQH1auGM4j2k6CsDPN+TArYHlDxbd59KXLlATJyCS5h2DTKuFvSw1RtSc
OiZsArheTERx71Yleu4+x9WnDAH3QzLC0st86El/lls9E5MPipx5zgfsacCj94s+r+qF0EzV/etf
SgWqOjyOfNHNnEAGt4H2jt470JyCv7o/fQTXPSCxad4uHe2+8hiUhXbFc1IJ74fTh+omO8CT0bqn
p61/w4W+SLSSt4km2sBd14s4pxbb3tdStZqJ8UdrQBzZ08HQ3naCTwt/OoF/kMFsKC/4H8q3KDk7
doVgBkW7SirpQf0liEqqbvAQVl3p8cozVKaCLFoav0pmx1OVmQVD6yyeA3LfS1+iOPzcrdq+f9lZ
tjj6mYKiN4k7q83fxxVnIs7vJQNK4WL81A2iLrIgMnioYjqOkg4Rh9VYyWwh5GYT1wMVZSoK/2Vc
V/bolrDaXuLhOM7k0BTkwK5ZkRIkOvyZtvE/NprIE1lAd3E8c36es/UoqApxKf6hSpvELVRXPbWc
hj5YTbGsXswpC+i0B/VRsSOBA09kesV7TRu5HssklrIezHPZN3iDXGFaaT/EgTJi99WygSwmICja
AR0SSM6yPptaxh04+qZaVFH1Ho6evzDNLZOlhNy14MDItHYQvX/LQWXAH/IqfCa+YPw9wGdF1306
1F/TBTJIfghDPNiuXY8Ova0V960aieVdmbjgHMZ7/XR8i+iQPfxh9rNXusyB39mVAF0ZMbi2B/WN
c4BFSQE7ub9pNGsgSVQ9iDJUP7RGhUcwaUKLbFAot07TmNesA0O/o0OxoKCRKafFlSKLrbBuQ2o8
6nf/4bX/9mbHaBIBwS6LZBIkCLcBGOAXxNkDiJbx+GpiAGGiyrdSww3ExzG7NaRU0FkorGdqKtpv
3GDq4fTwqMPHQOr5YQmPhclJxDJ/q+QyJlQbCNxH3WKRMorUIsDTN0PTDDkcOTBl0/Oeh9waMtdw
IDehWO4SrLuRyb+yPtf5EzzMawpPoL6BPB+uKgDZaW/Fr3brU33jd9pOH/GJt/pQWWojUVDc6+7s
tWhKwHnQ/dfDLfY6FpC9OIlYnNsg3t2DY0vCL5laAl6/pWegkco2Gkkjd22brUZMWxNoqlZvaN/j
Kq/TcowvD+QlbfH/yvULrqlgSIjfJRL+lokUSmZ2Z+7yndvPiXb1xms6zgUUU6cs3RwUgdBHu8co
tP2CjTInvLBdI6LRZCcFANNncKTk5QG5f9cbeyW3QyPceJzjBkUtXjPW4sS2GGcPAqIhtrU/vcyH
KZu9if92AagHtBpw/TjnBRLuMKDNMA+r89lGsUIRioq4VM2Kx7lMfjiA2cQRXhnN6MYLaOkPG+7X
thgaHfwISS+sAWGMbtMNTWVyzl88lNNvGLPExvpa5t9+HrDpcEPizMO1IAqjSavphrzdFEAsgCf4
9E5pCxzq3I9Z4mXwIcEHv/d+KbaDCCr2srZ5bJzHuJrgpob60gOKCeNTIupwxQqhi1woBTYerU5E
k3k56SJFUteVmd4FOMHLz7U+c9xbX2EGqK7U1j3WHerju9alkI3kkvtCCrqiZNZYpwFe03gC+6pL
TnQqdWqiLzgedtR+slx4NtivRUHGnGFLhoDc5zuDM3Ad6Zn75c1ZKMHhevrXTrHAw0YPRbXfOmab
4OwyB4pg8C6y1rOEZEvMDNTv9pCqL5tAmChz8NNQehg30z5BIvua72tLlbNoogmX7SqoijwuojXD
STR1HzIxhPVB4Qt2aGVFSMBEOgXaW1yDA5u/lSpgy0lnTuWHpu3XMTj8J/unSshIMAy1fyltNNYe
dldEpz2ysGl6Yv0NnbIrgMQTLEH/hl1XZT1vgledMdO7/C/SKDKe7sYfqf3RCHh1oGYYNkuzF1aP
QdwNec6wLYxc5LS6ohkHwL777+PQcXaiVidhfjJRKIZht+r5jMPe3O2BcbvynwzV5om64WlmJyVx
y2zQkClJS1pZDBkgWA1T8AFjG+qge3W56G9m+cSbyh5iO5azM9oxdzZhFE35XViBmcL0wq3IxdGK
4/98YDurMB0P20UekbCpyMZPCgOcV1OgEi+pvPyrSzLVDAroJWniCZmymn6hP0yJ1Dv+JDNNhLrl
1inAf87dUjSk+tt2pdGUfvNw1I/vzHSGrIXewahJE3tMr9+SCrLwuG5wOH8RfldCc00u4M9kCRhv
LytZDkvqKIQ0ir5100iqm0eybayoYW00rYGZDekzVnwYdf8Av+3eqXUUVT0XzmT61KmUbe7zTf0/
7R4RwEv0RbydfEbFKWojMifvh2TxEMv4op8lolrd9VMcbrOq56gbuoYP4osbYc6Qq6nSdXy52/Vh
1DPNVESJaUyasOF5LOto0SYqGU0P8eYxOy1I28uKHjvZi9Ao1V/aB/mxhTjzG4MjPd9vqbUfot7v
mWD20YsxqmIFgf/XoJa7vRfYILR0Q/EvbmYAD23Pf8v+OAoJ9729gPWrtOmDGyRKnsjK0EgviYiA
Gpko19O1ug2DhNjnkL6ZqiNPdkyjsnaZmid3rfWw0LULp8Jnb7uVF8JwqrgtxSU3dG5OeO8vnOiu
NKrkvAjmMAxgOeCFfItwtHoZxOBwC7KJJv2d/OAxFsCXih+wLM6BY8ktMHukE4cyMPgejfL4aN5U
8v5kaJPiOzqpN1jDE44Jyn1tgDu16Ppa0Uj1n4x2sXQDV00yoORvUi64Sl1u02YvxTcaZmmItGr9
bZirZXwwtSA75eg3UNcb2kVscfCx2Ml2FN6YDATLCGWdHgw+L+70Za97KBdGlynoaIeW9CB0V/kc
EpWiRqWM0hMXT8VRpr3xHUGn8dZObBCX4aDwJh9naIzRm0wEtdbAL6Gjcv0YRAcLLfA220YVNIjG
XxpT+v2c8YsNP18RA5xOkvtIofYcEoQ1y9FXU7lU4z3fRT/Ru8ObVnEfIgmJz9TNPp+DMG86y0ZZ
Q7paK8Hz5lP5ZfveddRehH/Grp0ztF+FZy4fJaZh3A2hmpMAZW5LZhkfg28L7vNhtIOxF22viLl3
WzGpGY10ZU2pCcW9X2w3V8LPSixV6A2gsThKp86+eunS0f3aMmzLjNDKhKuYQRPIDXYR1a4K4rJj
/6WMI4tYUf6xOhoxayY2t6/3SLvX1jrzuokPNIraK9rQv1uD6XPfivyN2wzO3IhnaGg5DZoaH44E
tOhtZzJ2N23POxDOvX7VQFe9GwBFgNKqu/+tKIzlLLUljzW48zK9fTBxfaRht88bFoXi19OAQp0M
pAWOViwltTuxeF+DWtuCSfqN0C15m9MVC6qSgQ/YBPrgZaycv/upe/EmmPNYsCd7fWw2HtegYcNp
Zd+7kkldVj5r788Z6092lfV5y3g5XyvLyEmZWdt4vNjGSoggDjWNpO55PZXsG60mP5f/MYBjS9Cl
/6hNhS3EcmRjS6ioO0ecepzZd4IDdFpIIqRcdExv1MHznaXzb0k025gELjW9R9i9fsA2dHjYZHPS
vGunUSRu/bYpgvoq3kZixHKvaR5Lp2wqYiMHMIb/JSUSrLk2A3/WHvmpaWNkBUYuAac1EfCr9Pza
krda0dXVmQa7cj4Yq0dURJagxVNlLS57e5ZnLxtwS5f0p5iOeQjCtD5B+br7MMhJj0dTmDaBKWm7
5kYrY2xMJmzuwZ7HfwIpwfQ3arz5XZiKRgJ1AZ9nZJg8vBYOeUhBY6HFhxB9CojlkRxPh9m6xTPv
rE+Jo1LAZLY0roQ/LbAToDm2my37SLrwp+j7jL32x4Itqcrkz4iFtcIOWCso1LQnzjX+f3QTLHpv
rO7ncMX0qYPRVxgOjYIcSHyMNEAUSCml0kTUc3J3Ene/9DPepqR1jtrykt+tcMhNyez7tmFYDRbE
iQtst7P6rq/eBEcdnwzuB9AVa2GNkVJKhbYiwX82Y80Bh4i/nZxw+h0yUKxStpqyNnxLYWj3Wgto
iUqem9lBJ6MOIdm91sS/Rvx8bmsgILtVe5YBQNxqm4geJ4QnMwVmT/8KQzXb6+yZCX97dvmfjivy
eE1Y9HM+63HOCbsb8EiW93jhXMI7qpElnRZpwC2jQn8wpW8lfu2MHSIpxpihjfD9b6sWJ/C5c6y4
DWsi1o10HX/G+Ccre0U2uEYOyOOqoUXQHRjjv+zv/upD2LMhOmv3y8JT+4g3cDUC5iU+ZYeVBg0z
+A0CjQTLHz+JAONl4pqFbWt3lxqPlAkl7gTwiIL5i5aF6T9f6fkomCodJG62sFqF8ifS8yirivjD
4QMqu6Q2Imcxj+8FJRpfSxRK6fn0yvgw4p+GoC8jkRfG0g4uGQbSn+teopQYvzukc+QTwNgPQ7FR
JG6q2Z64ifMe/56M6gXPl+ZERdRfH1oB6t+nljFa9dm70s/TblT4NZTHDNtUvJgr0U0MjHFw/89c
N0VMxsW+MtzoaobWHPb2rXhmrE+DMbhslX6In/ZXWtTquwPR/6K0WXNZBirnsCN9QFSt/drAevsi
lWGEf5yFokI+lP1CeS5TN1YWRrlsPxJYiZRP8r8nSV5MGxzjDJV74V/SEGMeeTLOhFv1iheaNC1L
56QZc6OQQaHhKtQhKeEWkPbWupftzp13Y0RaEbUsI0Vpfwm+nxobtBRCmiUDOqoGVz8droVWd7HQ
ArrMzi1xt37JfFNQmos5nugmW3nlz7yDBmlaQUbNeMub2DUcWo3LMnb02Au+nEKDeOe82fq/2fIu
dtJQgGniaU1WFXrm1JUKBCRBPYjzCb5jsMmabzuLz2zNNkouEQYZjlnrL6+Sl7SlOqd7HAB2NNZv
iD4Z17fW065rSWmV8PVj52hvgouygTy3Rw+6CnHTm+vm6jtbdaDGL+OHIxAG2brOI45BMKyDLqlQ
yshJhhd0AEc+stlHCKwsjv7haaYVcH75jIguQpzoxRcg0uY35HjW+0ac01O5OYpWiCCxVtMdLLha
W0oftNEqKums0hSUbRJ6PM2lx0xrpwl5QDSPxksxhMX5we7vMXQvGFA98h0GE5V5UzYZ1GaUAJzv
bmRo+VK9SHudJnJ7NGsj5PCMB8TAkyI9+QXg2LbUjbyfsUBxJNFt1U3+lcAHbpJI6OeXkiP8uC34
CEGh/wpp/sm+XWAyriY6bC1yJkQs+i9HbWmLDDaT6lDyceBZLNxx67Sfmq66upcusQ9OXa3/dkUS
63pUMjagZQd648P7AZgHGISeZ3UjMWp1hgLZKxhKb2UOmDIC7Lnb+oSIdyC702mmChpiOHqKbJPd
UQynHCFQLDl2kLuCm5xHrIrhIGxRwdnrye7Da9UCRj2nCvZ46Z4R/ZTRz3OVfvvZZ+wngflP6ciI
1k5dimxc7vxGUgiKIDz2FMaNaOkR91sKgsB9FCw30GQequhI3/ER9cfIcziikePIZoluXoRB9a/f
Og82P9e38AAE9CExYHKZEM6VQHOCqscGG/GvGEtn904Qz10Ds2m/C6lKwiRtL/Zq+XPonOfQXsvI
mre94smdLeE/UOHaaFEYOr/fEIaGukQvW07PPOZoW7Pp60HeWrSLJC7q9EEvry+xpz5h2LXfGOaX
AyXpYcaKy+OnA4dn32yOxCAilWOdAmRqLlxJ7dOw8aZIeeW+fV8uvDEGsA/dIWdNerg+pY1W10pQ
YVtQc+Gn8d2+PtSTWbmMAPB2HqwXIXWWX9/Rlb6UyxajyKSXFD6LVpSymZnmG7Xa9h/sfYqFf/Qs
4Rp/EyjsucN6HjaspRQ0dNLzxAEspil8MrI9HR58WgfBK6+zTxone/tU3ecoIVtJZm6EuKoZmTz2
JuTkv/oUUXs60QQaR2k42Cy3WvmCiaTafzS9Zgkv2RKJEs46z3gTRLIXPPWi7HA0cJhD9im8XgQV
lxO3kAeCsfsz1ddbrknQREyxtCbXWQN5dZEbfkAiPiajX9e44tPq/CzEgWnYKyErQczOPv3nWtoZ
bqGh4qHJgYWsfeAGoC0SRBLoUJSXR8EZ1fNUaE3WbA3l8iCFNjM4xrF4nVt0h3usT+6kWq+axsPp
70RDhUZmR+Ccz2GnWXHCQEQGtF+am2JjH2FD8TdJnL62JNpJryBc7Ky9GvOP7v3kdriFZekPpR3O
2NFzaHvBIhQdvWoaWB5Qb+bI5sPkZZZS2fHMmcU3TRdowgw8MOpy120Sr/BBqF9A6plelgTvaTPN
GgoqZCv9JpWA8oxF726eB+mEzEPlylU6QXJ6S04X/wz51sfINvXo8TY6JXOoFjGIqOeV8rcZg4kT
GrJnoBcKLX1576gjWfkIk89c5PTNDgia2AheWYxY9ccc5Y5fgk/N2MQP/VL1EGKezYKbufS9cBCr
Ku/4q5oY9NzzfiBjx5HaDsVoSaqqUXawoc6Rgm6Q89O2IUqVzNg+gV9nd/BhJoooDWlUFiY8WUf7
+77E9ytfwwYkEBEb/8VMLLKRydpajlu6a7B+d5zYtsVdY249gL8tfXNUyRN3LPDnfLhVBDwNmrPK
AGqP1mRkoT4kpnUIX8NQPE/eDGwUZQJWpu+mPy2DYJhvmca1w0fP+uL3roN4PooXDsjR9Qftl3+d
wELvVZ4uwaaM7nB5/y3LBvxqzY5tK7Ypu1FBNl7HRVnNstAhNrxnPLMEyzZxOiVuvdnkzbjuX2lY
DlF/komv7k0XFqx1WvpfPqI+lDYFUO3GlgA2oDCnLCFuSkjPUL6MFFdVWrfOI36sMiYJGnUqvoHp
7cXUdCXrLdCDKkzSsh9zVjftpQxKj7iezhB66rpXJ9R8wK7vRUpHmpOsaAN1QrFXzzbScG2UJroo
kKliXARKDAwb4Ed5vEHTR2sHzAIEuIda4r/KXWSZCIC5ztkfmRCZySMoxZs/RN0tR2kRdeRyV/8x
xLcJOl4jybqzdNNtnSuBdLpbVcs8L+Onjq4HyC1jKcA53caeEbjuZPbAQzf0L4rkjtHK/EwKb0aU
G4yqS/SasRQemvhAFFhPBok2Fhty36SNLT1zeRcZdp73A6t2hCekFjZRdRktoGRmicYYNMkeBZex
+IRLZQWLaLiC8sK4YktZLoyyZXDxdnpOD4Xx96idM8fPOBHgpZmCNN/Zf19LrQ/5gW7iC1iOAjlN
5fpZ9ax2FZEWQNbvNf9dOSg6l2U1zD3Iegz/A6uG4gW0DxCf1xw+iRrqviWv81HmNdPkLOnD/oj1
2+S9BpYK2qiDoG4gEhSQQno4q0dQiJ0264V6aAhrJHS6bfUcnEm9xQNDi85vTJ3yQHuMJMvuDaFL
gDS8k+VyZB+KUA8YjUnWxelmymI+tY2dluswfCccGtcLslsPl037Kc+O4R3bF6iPvpZlp/EVtuZw
wAGMODtOpX+mNahxAsvFtD8GO7E2IPQA66Ss4s/vXttfO3BuWERQZRTX+je9nF9yH5MVvf/fnrxT
8gdB2e3lNLW0DwLkMWdz1+sWKNr+FFMtMulgoXaudeB+sICUvyZxOzRkoORwBuasMlT3DzBqiJTS
W+oR9XQ4xkkEo22ZcrduwwX8RIcadbkoUNDVSUa0nctUVHveeK9Y+0tI47qEWX/SLs/5tnjX4rZW
lvyvZUYnlB5O7WUzyPx0t5OL8aTr2egyIIeFGXXK+epKsOnQwr7mGWP1hJ6a9w87t7QG1FX3aOa5
rgfIwileubNZQ/xbB28eXdF3OPKXyBZTk0a72L+uynAqZKOyELpnhv+vCC+IFCy9UobvJtq4y4dl
O9YfMqNRu0pECvZfSNGrqOIBqIGDO026XFsTR6NZDyPofmLNDm0TMXSikwHbSjlYcNrPc4amrbkR
b6gXl5CF5+hcCQx+h3gi9haxQyGDHLTH1iM7kfC6WTJ8rrtmEAjz7cuoPtr1ZBTQ0OMWkochsXZJ
R21FPl5I83eJ6jDuC2mF9PCrp5G4x+bcwrFdd4CViLZe7cWmqKhulFo2lDZAqVwx/0h7CCkNqO30
3KVjO3OByxznVEsnsckALdkjNcg66ZAPQlKwYvUKeVJUeaJGbzD5B/VSTVobgTJ9BSN7OPeVcyc+
wseZqAQGOgB3c3hciJAn5bR/yYiSoa1BTOW08k0+93aRpbjeH+I+KhCmlwRR/N8JrktntJKxNmDO
I7yUoiRqARTUVRBUknynHG7fbci2CPiGiAVInPIiYg7uIKESfBE+bmslLaf6T77/jbzD25FKCCFZ
1q3zyyM0Jaya9z02W+HNbluNmJgGCE0DdOp4i4sqoktMXbbXQ1deOsy1VPglKTKrGkOGiOAo4R67
BmHUQnSe6MDRrDCN119SP204uQyMuI3uh5ButClBp4hiIHFoIOkkfQN/XdLGVg6g8fUdlP6UjxIo
poShaCLjWF+Ci+zPEcARAdBlxdJKv+jJbOhjiQxPSkYNaAjkV/N0vEpKnXJZh7vco3IoVYXJEtDs
8SaTfOhU9vWAnKTX27lDrWuEQt41etFnUWTji5a5Prp5hi/BVo2mpZJqTpQPx9bF9XfexvODwvq5
rLUyWt1uLeK5Ga+mBzRvVBlL2Dv3eFaTj5LoBhKB94RTrHqSl0pjghgk+1Hyyx/ZGT1AxVNPDNJ1
0/z/Y25486qJhxiby9sQp2kDLRtmI6lgI2ZMccJm1TrBSIBLpBkAnZR0tAc/oDbKsx/PTtIbhZam
wYudJ2rWiCCrPPwBlB3ikYsqLiKZF6cz46+FTHijSQZxhNf24FB2ThzXgGnJYHp7xK+ydzXjE0EG
mYQ7Cp6QRiFDydg84cZ0GkMH9wGyctgTOsrno8oIB+R940MTi1jqp0vxTJze2g+iCIk4+0dEnjVf
QvcBQVidKrMI1mlPyHoVJI7XNgsbXzzl8BhHZHLMfWfGdsUvc74nUrWjSQMMemky5kn5m7XPlewf
hhNCGGI1i4Ds8bG5fMtRNgk2UZhWxdpdlIoxSN62X46VMY7tEtjZ7tyliFOm++QXNvGn5fjU8mpI
w9oBqYuhWnorxW48NICAgZCN+6GawI68H1otsLxVDDt2kvhCBH0bstfY45BsYuFGo1zFI6lC0Bml
uBALt+unGqmqtLC6sLPnxRRxZ3CGH83MP6nmrAHkkXkXpQfuKK8NRqEFC18gq+duTyoLExqKX+nt
5cC0WUc2Yu9OK2Buh2Wc6ehtZqAJ430MPppOavtzcsusA7+Lfrtob7BBV5xx8j59yi97U0OQon8f
kzSd8lc1eLPnj0LsTxh2jKdmJmbNorxYhQRe1ei2t3hEqOXQX9vUiZoA5elgNgHoOUmgAhsRo3UJ
Ay1Irbf+4nWz0d/cBF2ahAMu6oEc9zSpzXY5WX+biLGCYgXKuj7W57vJNzpeG62Y5XiQbRRqjrT1
QArqeyUJQ++vm3VMOv0ftIJIdb7wMc0vGocadoU8Y8HYpv71e+34PaisskUpvVdbWYuAabcibTf6
koLvSm222ZNlZUaQnLcLLriGy4SlkTqoTnHB66TSAFeAuuoenh2D1IdKw942p6hRjmyvMD/lrrOi
cm43XivXwEK3/rkAHHf2hoaMT1hFkVx9lGpflqNHmG+15/ZzgvHWpGDiGrEHrA+CKJbBWS9TDVHc
Fs0CiC8yFnuedPBG5UdMBDi0QuM/Y55wL5YBv1f7g7d7Ppg1tM+yLTijThfA5tA2JLHw0O6WdEjV
9HA/Ac/zYy73v6JWJrfPun9tOor1RssNueEiS+BLWq5mnC1XOGdFKIibhFNDhgowwSHlFBcPsW7S
9P0iEgubaNcdxh0MqQoyEQeKTXovFEauc3wnXsjawI1IAXMyaYa9eVZ/mhU37E7rcguSEKo2ZFG7
9/cIge9KXlLUX6UxV7mih3nSjqHnH3HpX8hv92UQCQ1p+ItUOOrKJEmqo21mL8NQefXhdroerfcg
L9sBVWY1HHQbaaeV0CdL6dy4znSwSa2jXPngcNiLGdSJaWw3hl5sMXm3R9sqJT3JfcdEF/sGyPU2
xEyrRQSuYHSdpcsl5oRM++NCsWsj1EHD3JjYxDkVV9gHACa5vm/zkRTFIG8pLOfMwcZXTl1KLFfj
SZeU6T/1NFlocRGcGM2hfTxAcG1G8FbHgOi0otrt6WcwaRAiXhJGcANOIH3WLzOHqwCZ4mbo65tD
rDRYl9FlFNAMwwkiPuvt1H6x5k4SxwrMuuf6QDgn2dqzQVfUX476wTjQ7rVwwWv5FX+vBRN4rtRW
mymsm0whJSunJ4+PuZyubjJpnOPMUs643CzA3mFwoxhA6MIJfa9Bv66mn+fTRlfpXTtTepqQ3sPE
2Ji95eRBjrpbLcJh9nonBsHlfLqmFi8KNj5cOWFtZI3dS6kh1KLGV8Y5rpy41F7bJVN+JLznlbYo
Uvh9Ktqmn8wyx73mnbELxACyy2ZRfu87D8MFPaUh+Gvg8cgpG89hf0A1DpaPsrSwnIsDSH1DRKTJ
ScTEqOskeORYIeo1oejf54nRXN4ND5sPfFX8Qm8TPO6nymEjniMQtiIwMJSirpQu36YSjkfeK/W2
yAYcyezHshVv6IUkSfX3hy5JOjO+sD9KODLZW5epkBjtle86GCYrKMmRdCuKZJpQ6FdGMlljVdW/
V4jTcLfzPbF0qDHd7w3O4E/po0oVIwC7qMDlwp0uD+ppe/OmZzi4iWpMfwranP8r9cgBaysdd+kw
kwmp4DqbY9BG6igoVJAL+4A6L7notNK+s10lFEFvLgKiLaLy+/vOyPsC5qU2TnSKkT+mlGjHj9xl
rC1BzqNYBNPvBE2+4kkznJPrb3GlEXeQ25mv4jFaglthVf0DIyOtqkSWUlvkfb6s9ZB0DfffS5Sr
WIiZQ1XlM62sgVyEV+EwIQSnr1sG8AhX6eDlzQIL1wQMuhXnbVwksVjaNqmVP/RiNx2U00Iq2cfh
Uv6xZKfbfODp1fm/jGgnthNLJIOna53kcAVp8ZS8kmQSJjTv/vr6sq1UFbjpCsUi0D6NsvkgwxIF
m6rIeZ1flYNJgAYSCuace4h6XOxmgTwzGoV214WHvL5BgB2fAWln8x7ZtOXQlkmmKPss4QWBcJdL
zDqcn3Gq8/mJ/r/UT2q8ZyPzmqLK6kKvuNKmtllkELBbI62woEBvWw1q5V6flLBJUaz6crhoDdzJ
31SF19l7UHqIX4pF+oJYMHbJEEOQXyE+iQbLvpnc35bYjnGYIBDl6z2IOoT63s5If62lUPHMzHJv
p14StKWVrf3iOxC7pmW5N6OaEXT0wM3EBnXiTQir0LA9WaVggCshRywQ6GkdZZQQPL58YYAkWyYB
T/INNjxs5ePx2hMPEEIlxydhtARCFEwmOIOmhHz3H4yEovp6XH7OmEiaa6fGZvpi0PoSEmYhLClZ
a7mCihv9BeU8dCsHFo9lSP0h6dJw5byt6Qej0iHcoQMo86f/u22pys5QscHpFnBcFveylAcV3x9y
KqLtRMlABt+EZV6sflhxrTjP0X2LSMOZZeQMeKprPXAfarh3zPw71EkD73ZtAdEzEMjOCU/9h9QX
PT1LC8HH8RISlWBreDrbW2zre6sAynkflaE1KXlivhMsnKUIx5YEmTDFbm4g6gSlhmElj0kRuVON
VeDnVYv3sDmmxnGi9QR+RzFfA14sjT7g9De2Awb7s7+TCoP0tGlpSOU85yzyMf1CwVGVU0giHJ51
zX/fEoowTD9kEH7qOYuzsZxUo2/mrSyXmrejKZLaAq9ilXX3k9YXQ18b7HthbJukUSG6+XBhEXK9
PovLC1jlBVDb1ToODXLX9UpwOQ2lf7XFibAmuLeKp4Bs5GSQUpY57VeQaw+ugXT3NrhFpil7Dfza
khMP5n69s22gizYr91VxnSrhMR+6VAMy27DQgARKcdOUCdjEcJNxQvN3fnJmkBZCNACwpQ9zI2dS
n5ghk8oM6/qZ5IFNi0dZ/hQterq6fOU39g2gskE8HBeR6gzqP7fHi96hrXjd8MeLWnsAa3S3K28A
cp8zzUu4VCW/iQr6X+F9qJIr1sefCRUcC2Gq1y14d4VbmNpcBgEHKeiiVWZ2PBaAdHVZi0OCc5ND
i/dUnd255aGUw3/35uahKzyBsGG1R9EY/KxEweEWVdrLbHER/0TUV2q9s8rDFUUsEdgXRWvebHoF
kJ0iI4nG2OE+qdcSHoMpWgF3OTBQxJQXcdbZna0NH0ITH7JF92IA92taEYGL6D6iuzkgQ86zmzho
VnxE67qBL3cw1prf5s71vVXKcHAB5HWT7W58z8DJtKB3mAbMqt81nliy52wppmjpBnOUwDdYCOHb
9+n4fuYnAXWdo/6Zaom502E8QT+5kV7TaDkB53sugbpD2x2pXs5Tjnf7KeXl75+pW64mwCp6G4BC
LHkHxMblaaVzc+2X0IC5YdwqgGqLaIlG/ysh0TjhcfYv2xx0ghE9TEGUAqMfy0m6+5xcExO5sY5o
eqWY89HyIS9BfM7buvUthH6kA2c/GUEGKD/2YGPzcaMc9MbuIVqRlc5UZBdgv+zIY8yIN5ZdWC4c
LElElUgBo+mNawW5MlqmckUy3V5bKZoER0BOB1BivINV1szKeFTpOdhqJgnZfAJnjafHJkt6WKqH
74LNWVhrK0VDqrJD6a//Jm3ngR0rFE4QRSXOwYgevGsqn3CP+/SWad7cJRVix8HfIag+fEkepYbx
hJ6zFHbZ/pn4nApJzq/l2YRkToHKs4KwgPEnLKbGmnyRApUKO273yPY5QPk4kPFAOjOpQu5Lc3WK
f8ijs4D/OFSNX0IGpzUfBpsJg0GeQN0YrSCo/8+Um2vIBschoe41ZdBLkAXYlDpDH6NNGjiPjuva
pne9px9VfJOT8swe6ckRbwVsjU9UwQvc5IpoSKpzNDG0bFmkpnBrNiuUbH6GUo8Xf0gEgx+IWLEb
9pgzQ+i9wXEgBe34yfyuWQ3TuvU4YI+U5Fa0g6zuz/EjOT/uSuVtrM8lG+BZOmHGcEwUyJ3Bgltq
KYDPQCrwfkrNaaxtlTwO5G4tf+VM+bJeI0mpf02FBmY7n+4J6gFXUlaUZWU/afNRMQGTxwtKxnZc
m/Pwuf1fJ8jFfDAmWOz2CxpRTz0DFH/CwilujcZ7MDenwzyt9xeU2EjL3b0TUAnC+d7wU2/iJueZ
U0yu6E216ezy3dWARHszE0qqpwQOhFTwk7rBYj5vx/9+nD690tEfW1rMwRgCSbVK1ReHlUB/2zu5
FnL64N3B7qmc8EgVYcsuI4w/qIXIVne9Z7tQawJIlOVjmu3a6o0MzERq7b+xwEygn1P2i8NnTHDL
jPQ+oWV7aR6WcyglkqYAUHoGtPXxy3P6IH434WbsbHS8Qo0AxIU5hNEnYWj3uxPTIQu9zXMqfGmP
Ox7m9qpnFHwxin+WJh0bm3EfJtrlmkCJHGR2mwBzAqdKoTnLK3TWdF+tx2rsU21wkHVzI1nV/BJW
HzAbKpIG0Ks2gCc+qoYybhLpXU7xv8Dlz27L7bPvjmS/uP7r53Bp8iWWaxepAbpwNKqRdtzKVDs+
/8GvziaJ7Pze2fYhmfcGqT3x9UfAXdK4RNYPH6Qc/+fvM8cJbF/vyDDfg0HcgYvTOBfvTdePCpT4
wMfUBorfWeVuaJuyZ0Fj9gyyFJL57Hh7TgNBCwcgsQHM2KYIBhXi/pKs45M5WCvrZpAATZv7h94X
09soVEecRp8B8DbkzXJqzaFv6aZNnA85/lSrT319zwgmzzTVasNxe6Ea5GBIqoK0fqnzf6yWBdN7
mbRA7VOKicgtlJ+w0I/6KxwCHNKOqlTsDoi/TG7JLVB6k6Ialdm+bs+OxoBx5CBdUZcpdn1mbTF5
fxubH30kpaUFZPrdda1sQe6M92NPoeyXIMCDeDkT+icFXiwFw0OmwHtxPv50lvmK4UyukqdqZy5d
rjVNfnpRl39qdl8tGoIodrQtVdA2KNHPBE9Gkzt+MMqj0VRfMMX8WnPcAE92Xp8hkEVpoko1QhOB
AmiIdMOuJWstkgnB4rtmTRem5HfqePwnO9Mh9aS2st/Tlc6eDqZca953O5HUZj4grQXXqxrg93HN
tlHZyOA+v8SNL+zdW+g6MgboRmfZqc24DVav4MIdW66avDfeQd/d3zumDLF2KvR2x2xTu9Hkig2e
QzqeoEdkZ3Bpu+TkdQ5War3cjKFF1RZwNMWqIR3dvq/TwMBVqMSlMDnn/E2ceNfBpPhAmuhg/KW9
y1BD4pCKx9/hBek3kTckW/+ieY7V9OHSNZZpqKSN02Ko42eXV6visjqhq4K0/DgH/IM0iUM0EJ+9
415nVU0RdT1vOOUbSy2T6hBhatyWTLMFHss9YLvoPU8M8Rdt17aNDHyMPKqPAuYouuxb32dyJMW1
aMfO+Vgw8K352c68SCNrC+XpUKrfRoh5pjbpVfOV+PwDWxvx6zU/hiFeSvulMGzOKK2pTUKZZOTB
r99ds/iW1y6kLTXHLquEW/S/bvTrm2gUAoMvddBite3U59QLisX1bPoTC/938KUOvySuq1U+MOfJ
Zv3ONHCmpsb7PUkkcIsVUPOEY/jWe5cRGPTN7Z7Gcrz0eVO+hWmZv8XmwZsWc/IrbW3IbQ4lCo3q
SYlNysOQ8nZqsBvMf7VeLETM22IvL0CY9iSQ+1IYP0h9+hP74gvv4A/nc1y00ipRGCUw4gxjyagr
sG6OBT5VWqljg4SpmsRatAbIF2HNdvcMWMY7ffxmX54D1G1u/rPdmQn/S0QPNqVFSfRXv5zGpgU4
gM4sYw935jKRoFcPJVOUEsbTyGjMDxvONjlWrYqgMr0UijT/EsXFKadnN/yfABr6xvhUCWFtn6B8
c/p/nFY6g/J//GdWwXx6VMqzokd8PAhXqgpPB0RjTP8z5/GimIqwkDvOB3DVPK7JDIGXOuQ3UYub
q2wS7kZs7KjJoJaOTVgZ9Lx6rFLHZ7DgXgvmXIzpgZd9GyTFl2m4/PZzgXQJdkDPIcK7Gmrhdit3
IJm1XXcXzRUkUfuIJ/xVjvfeNGLF+BKMCR39y576rosFUWPASxHPz/uxMfiv4jXJNDO6NaqpsJMu
AdjKO4ajaY3hLeO0NXrsXsTJHZDaodc+r0PJ88BeEWsE/kqHV5AonEBueIjUSIvJbemuBVPbRaES
wjKZ8Kze44i4vxyQXsN2x2OupFhC5n0HLXDG1Hiq+vCaeavOqjLkI4FOMK8jFboMtZNwUIh9q43D
Oy3NJ/Wf+SFihn4vMo9bgg/eEXk+CPVRLwp7lfv64mjhTPUNmSq+cM4WGKGVEu3T+6Rx59UcVKc/
tGQX14ufV8WpskIaTx/YMeUJ3+6aoOD+tDLDkPAL28/5kRWAH7zXjYfjrY18lZDuoBYMG22WfTrv
cQh4YywqHgCOrfvl6NsnxBQDybGjBT95jMsOxkZFdcGrkevS+k7kYysxO/Kg2HLjbnwpD28kOrxh
NhcwcnqdRtst3eZ7Vryxa1mlREOfLxk6XCJjUoII2My5+UAHKKxJLDXbvnlIsecNtPbfwKnm3ZKt
7oaQ5LVRZqDkxqLPndYcOqSUF60ypiLf9J7oUlFM2a4ZAUUDxv1G9my6qdnUs+uQf3GuFCjZID5F
z0aCHKVU3wRcxLzbIYFWHDsFWawIG1obeVMxZSODZev86ZyDAsK/JeVWqB3wi9Lg00iY6UJVoqh3
NvH2pRwR7n4Ey6SRtB1ua8cW3J3HlC400rlQg+ZLVsTXLVPjo6fgWR5mZcMyU0zZhAoXEMha+G9M
Ao6CcRJPMyzk61Q8nbS4aowcWvG1tfF+G3STzSV+9zIJs3YZDi+bg8fS2oqsxkmNwNBKUy2OXXan
KIK1vNyoRDa+/v7GjbNLoAwJyn6ucHt2zFqpkyoFQUlaWRX7Tfu1vz8bLdgHpPtObq8a2q68RyV8
kmebZPZPyf1qx9Az9pTAQgt8mWtIToSPOqnM04KHfE7tnT0J2pPkg5ljICIenxCxRTQ204Xc7aOf
7qhP+9aL8ysbYfpggG8np8GYNJIt1JzGYgn3wnJOnrgpt8jfg9KP4np7rs6DeMhvOdWc+eoRQuDs
Np9YrZUlRPAaxSlbrhLR/7Gny2vv9Fc4IBiPg80BFyCGEgGIesDv1Z1PFhLR/gVv0FIZPwS6ucEk
olG+0EA4nLvxCQzQ19oSDmfGI823w27mfJiw8v3iyglVbj69IheouJlkZOapmViJYFoAN9RK+Jgv
8CKiaoRcVSTaNE/Am68mWcueOsD7uQ6bo9LjN0VDyWndoTinR2Hnm85xZXrCrkqkQQj3Tl9HXKjt
6iMbFhv9wPRrzdmNXdxGrLPiUJVMqKTRQovahYSi47liY911bS5IYfZRXN/oqGKlECkLj/v+3iDY
Z5gW7Fh67Ti4r7GFOMvN/rL9kvex5ENgElv/4JKhRfaGklBCFq5ho+svTroMXBDCTonPcw+3MScq
71vXG/0Uj94ledwVPAVTImB6c+XSefv3gc0ugBvoryjLwcZwfU3jNVNi6Cy8/tBXcmnDQCiPIJj7
/7XO9zEKd1oKAxh0ppNbCS8Cu65DsOJ5FJL4Qfd+g/S5A1zc9Y7McQUVDoD4gD7+nbrFPbz35QC5
oPRXXH0HCSJXF8KG9IqeQURaPONmkde10tWx+axlFL+w2FwhXwTUjVzwPqDACZBNe1N8AUAbwjS2
koWgBn39NMQHuAi5l8HL1TcuQPv67ukuN1gqiPJC+Fx6cAGzWaYr0d8KUoNQXLipPjGCF5WKJAUC
u9bJy9ZvzxFfFVDC/hRxqUq7EXMnpqAmaWaFhU6vZt/vMcd9u34kcbkL3XymINaUVv4o/h0xAgPV
abxZq8waIIjLljWZL/7SiDmI1eAdcJyC2Zlff0tYtzwoLksQFnsNExKfrBLwxq18UrwTHd7DrXzz
8oiiMX0DfUweY/NkawJv/4Pf+rFa5Y19WiqOYYmS+9OG6Zv6SAU7We+0E5cbyEAaplZVxx8KzgYf
spyIPDvkV5cChlUyl/yPo+naalyl5b8WKbUkc18weaHCmwF9BTOzfrR6AMI7SZkpRFSv8/Kyd83T
AHeUoF1AWFaeGIj2ZEMSBUAjivxXNNbWKU5/E6qQMi+Akgjs2mBbRd0lSjO7Q+3h6XoeAN7cP6Li
oYRRRkE9QB9O6u0oG/oJIvSth8+lAAdNodRNXyMwCoX/Qb8tEQCSCmtjBfXnZ4YYYE7FNV61jsVW
fU6fm57jmlAfsw2GTjygOOuCDUQFu79EeZwaBs/CpZUK/fnWX5xLhqimYMG4n4c2Z62jFSjCZSpd
zUP22hHSZ+hwG7LZHsFy3oAxqPGvK6+IV10rSu3GhjWBLx1UF97/kZFd1p4V6aNegZb3zPCfa0Wx
YpCdClyE5RWpp8kNvdZWHbWoYGS1EXiJuVdrAIgt4GDzdwGlibwLwSGNJO1Mb0up5B0qLrZ49/DS
kSTDtBEg34WTvbXeubKuFktKedso7LRvjDXKs64zgknwsgD5lkwra/vbQP0aJyc2GvCxGEEnwa7r
iaHj6+S+QC0Yn9yuTXcT2qrbB8n80G3cdI85EZSytlmMVpDQZVoNdNRa+2vFQ5BCzVJIYlD8BEh7
rJwOd9a/2MVDiIGCCo9kHiJrcReT6XfLhT0FXDNNa0QcbZJQpdOoriJBi/3wclAQDYNnruyXOj/L
+rjTJqB8JSZ0SfnyY0i6bPxgjEcsZyyuzdCWuen93XNu5X7QwzHsaD5qG8WAG6w8KKPTvnNgJnT4
PACH+XjjbCe5GfueD/I6EtRDmv057O3N82JwWpu7bEzRDdFqwA8diNnVTBwKOYfV1Fz1u8wJe+xr
IKmx0N09w6nb0sEFrZQVqUwIz6Z+1MD+NJ9HOCRpmg6p21zfjW/tCmpk7TcuptjUZtBJi8iQg+ay
F8Ak4fnKOtuAWliG9sMSSB75qhTU6jn310KK0uWp6A8fULLVGv2wda1e+7N+0ACOXRi2WMGhsQ6C
JHoYbRtoMM/0nb6DuJb/+s/srwU8yp0uidICydvI0faXfvODpvH7Fmqt17TfzR/kgs+BpKhxHaUF
6AUbVFTrdFQX7wyikPO806lc66stI5MiGCZeb35u19NQnFEb3/HrojYh20MrnVmo+dV+jaCAS2q4
Ev1tswaCgukTyoIAtiBdTkULzST7eu+eFhXpFpH3BvbxgzECAphZLZe998qK7zjKNPZxptSeVIyt
gj7ZYsWBC7s4GLyhW+ghBvFAiNomnAd6e7EsbN8A/CnVIah0mH6bYl254siAfDCgGjfFZUEtVduC
KvymJ4whJnuVFYkO6n1UEWZy71yqXN9boifk3eYC9vd4Qvnq2L1X8Ozz3Zp07QGHiVkhc+GSdoaS
gJggeK6g5S62qcc2+AriP3L4Fwg7HNWC2fbPEwyc2aXQRCIcSJHU1M1lhI2gwKh13sH73WfDnup2
IvZe/IMLQEPwhJJxKn2hGx4Rq3ihZFaU2uncGXSe7Vd/30nk8N3JSETtIbqGa/pXZ0c8uty7ZEkH
aRKLWsTVVYbGySBksrLimizWApUGIEWod41l7rCNtxUfXWSvWC0QyzxAHht5n0hXwxB7hmvXicwP
KMoicuYlgpyyTNdUuQoAijKglGcjPC5GMe9HKQXUEdZkJIlqHkXKpblE2fJ9GhGDAtZzSdPMzZX1
lJK/Y/Vx0lHA9YqGUf2W5u5ou4Mzo9ffrknPwSZDOoDv6S5M0kQxTDXPymAQCh9Nbva8OgNXo5Cj
Xu0ehRqhaz7gntTjnBm8CEGbzCxOmkRkpwA4QjZdWmkC01PENJ2uP4Mhn+09A2MnFpbhEX2AlXeu
1/6KmOqm1UMmgQgoWxHp0WWNnHCD8saGcGRM/cYeAI/XwpC/IisBkMXxacstgP55l51bHzBRZCyI
aVWsKEmakFKqlvp5kyhVbCuhr5190aoSrWsiH7XKvCDwVOx9w/sVuv1mU8plqUy2RyOrgvK5ha7n
7SGceZvb5jyzasD2rJF33wrrYVC5y2Mwu31gMRPr2uLKwVffKvcteW6W0nwb/7XcIhMhnInlL2WE
o06288hJEONfKwnoBnL5jNR3qZZd1usHMLUZ4vtMizCh2TwWTnjFuYLm6IJTbbCw8rz/6iwi22X4
+gely55H0+2nUTRMrRe27OKCTXtbDdDNfPE6kKP4TEv5xmlRtItNczDCUzhHDgsWqVJLZW+3mBbU
h7h3SKV35biH2oV7JOr3pcHHNCoQRPDKmFJtZhnBDwIjzLNaM3i1D/DzrFkazaC7aKEnmj+3C6MO
Hab14nFu7itNFVRqLfRfyBqc/9NxjmauRMGt+iUujkT6pLWIJjW/CkH0bvWO0Q/4HYuqpfGw2wBR
rIVVhdxJIO1ym+Y1IqqPkV9sFPM+iUYq7bep43tugL9GIoYUFeg2LDAPKAORrpFKT895o6qZYDqo
9k8gVy0jfQ4vtuL4DvoCqqtL7b3o3rhQg+BP+zqg3U7O1YZ+zvP1ERQdBoQNJeWIiBg6xR9JMBPD
Sr6Kt74t97gICFrXyNrSBRG+jjfN8CyGuMoxFMAaa7NdQCDyq2rGbzV2XQ/p6CQj6vsIK6fWLP2q
2e9X926STh+LMWixMPpnUJjjDSVN0qLOCwc74djqM6xKLiUc6DtjbHYNQ2jhBXBLaFouGD2PLtqu
fhgtw7jgRyhz0bpTBZ0VQIOqQRKp+QEYx+vhMid1YncTDejf8TWz6ZBwX/gVrKp1qT1YWWpiiGT0
RDQ/yBQR7TMqX+cq9ID/wE08OnwHarOP/6OxRDekkjDO6UjdA83ajNEJyTVOEXrZqfPVhVqJUuE+
fltzJB1eVR0Ed/ji7MinK29n18c7r/F2DpT0V7a2bS797GiSWGX1+e75qm1ePUNTjr6U4jlY8PSZ
c4qbAXXa/T4BIkAhspRe1r4RF1N9PQCo5u5L11ZJAqnYqT+gGolnh1xjAKSjGAx2LRyJLzfEMAQD
wauWZ7To9hx4s7hD9ztxvUq4VvVud/ujhB1dh1hO0iBrrlACAEH19ImdX0t+M0jX2RviXxsKihJM
JF8SwEljAndSA0aH7hQt6Vj8zUMkplRdM6J2kGie9lAUdj3Jc1lE4J+Dz8h+qyrUvsMARk9E6whG
oNKSoDphbNG/SIa/26LrOlaaRW7KwFiTxwmQzZGbfneBLqB0tmKdZ26UWABaWRToR6241uPjacZV
JHCmqg3p0dqSze6EwXGwOm9dImgcGctjU/h0CyZ7PP3Il7127MQFMDwYGycBakvAG1LPeb8aev8s
T+KjpaMaEye4TFvJdj33WQ6lwa/j8I3Q3bnRg31Ai/bobFJ77f+pXkuzpnYe5qDv3pJJZG2nHlNI
CvaikTsnkm747kpQNeWglKjZBuAAqaimeV5A6YS4pwSC+7BhG5IZNMcHOsQb9cuGwjld50uhKKCe
YH0i7BCFJpc6pzBrZ0/+7ObCbM0k03Gn/2ut6qejW54c0ZcnDE3ED4WDo6vQvvm4EODOoPhX9Zvy
A57P2U2bctDElSXLHj7Jh56iC1vU+lOIhZC9dayavvJ+sY3Z3crrOIy9oWwen403xn1PK7Ts9HTB
X5YnA5wvQCz4UOIR8UO6qlI5IWQaX8Y2Cr8y/fOXyFTOp4gMSfOZMDUkgGd/k0ZXcH6en32rstc3
yyv+IHVu3uNoduXPq5yEpEuvKp0smsTblYxvf3Gb575eGpMp1CLA20lOSJ34NswRZQLReDM82eWH
9l0l80LtVZRsEXBfUHueda0MLfUQN3+EqAbvfKKH3XAoKD4lCj1DqKzoHtuEwktD5b3aSF0aDl9s
LGd4lVKJn1SkHaqCMSua+HDJj+m0QJ679DL5M6X3R6y+drWP29W2SIaD9vO/yMmi7cM1Sdt4KrsS
XFiz1vY+c3XJwVgjEhLYOoXg4Xg4Al5ujmc8f4UJ9N8KJTzab3NRLTKa0UOi1JRZUTkysku0TfFp
PnjMip9VzZQx3CwK84+r1nmsTYz59tjaXcAzGRQUNxZhqv74IInEfQjp9qMtbQAwwtZ2idecuh2k
diZ7VK2WQeQi+YK3vb2HEXnOLzznjpfIHFQ7cBKfKfCjSGuxOF7iP2BGPJQGLY19AxnWaqcdY7I1
ZriHWAEgkDQL36f7i8CRh2IRspcbgy+1sQ3zb9p48iCru0ZXUJBp1b6DFIIVpV/tY4sf2hQ/vd4e
nsqyXTQPWWByl4S/P26gxMGk+lAywC0um6IXFIBELcGdmhcQ8QL/NUVOaDvPRDY/h8bs5aBzuDD+
xQ5YW6NmLm5jBUaiDRm3T4b+EzlI7yZWv2il+q097pEciqMatsEQpGkpcwKuQ8wtGM7jtAbhKmsO
YF5fP8i26kQk8FgQhfwNFQG3Zm5z8PBCg/n2evVurYzfkn5Wg7TGJM/slcC7ULq/htMdGGAk9kOz
duA9iPGTOy6UQRM/Wq86xM/RVdARjRvdAxkIWG72mtZrFsif35Tt6LUgs/tMtvSJRREWnLq83FEV
6EWN/dCBxRps+RXCe5QnY807MZcN2b++DQTeARuzVp28GQ2XpJVDgy4PZTlQgA2IFVl3R+j4YHmh
CzyDuqXgSMaG7Q1skoALswiU//efr0x6GigORFMThRVN0ftT5hpS6u6UzKqBK11eLroXoCdKptI5
GNRD5xlmGjKaXi3IsSA7d6o8eVodSiLYwXTmo35jQuiq809HdFbW+nhCRmuEw+Lc2MGC2x42OpST
ZmM2CIGd6s4H5EwRlluU46GZ0WvQBb68TULxYsznS58updZw8FFDzrckb/3hjY5QV2we+T6T1gnb
eVJizxWEJqFtAwjS0JBHxFWOZQbPHnsgE0EPGPjS5yooC6R+sTqHShhRP7ZHXXI47aRRHA8vacdZ
Jd5hrHNoknzQk+5rQvJDCFFRK1WfX3xB8S8G0fcubR97WY4WfVLCiBpUl4sZr7OYC73wBF6BjS+4
CyMcJIu3ionLiJWj0G+a0c6KZTR2Nxkisq7WxVkGKaEpyktKA3n6MLrLvBtHx4zGHt/3GBvHz1jv
45ZFt/S4glTJlHJxpllTkBQ6ZVOqe+geZgFzKigxfNloLX5seOOQiAMnjK0m7p/ljobw6/2cz5bD
dkkZkdXd33HBO2+iX1ExZkiR9DqeEj+W9pSpxBRCRIE0qUl6p4HdYjyEuEFxc+6363DKyUCBD8ZG
LbWIJEtJ2ldVrGP34UlNZtyK820whZsEriFuMPmXVvTsS6uTx9i7w7wYj0Wt19JxQUIJh0GPB85o
UG4UU7Brf+1m6w6IolXBkiOlyHk5xaqMbAaZbJEx0nbhEvNF2pS9DeQNpKdGFqIu5YNJ64xT3IYC
38TlECVG3EgDn4ptIoERYe748mioea2x9Xc0BvWSs6EDcUgeZyiKmMutzdF46gR8o3r46nRHUSlI
IlwUrxN2aFgVTXKJkvinlQJqs8h+2xg8kC1PkvhtVUN5CRPElPkCtIgf9yMMwaudgJZZYqzou77P
n23ZVfMC/oNrjM7dCIBsPSO7RcvvowkXX5hpp4ueYxH3ro4qz7dh97b3i+93RemR3kDiqtG6+0EF
caAj4kgUf9syPiUpQw98WbgC2A+p6aAYzjGW04ZSo9P60bxqMfMGkNJgGi1THL2hjhXCk4h/ftBm
XBWu612C3Ue6wnSl69tAKo7goq1ZcODWNdXoiVJJDA7+ZgITdrwn1pvXeZlPjPBb1nWioswhJh74
7DzE3fdAZd7OOony6q/DfenKHnxJ6hsHb2+4mCLTJWvy/VlYwfS2Yx8528VWU4/sKfACl+R7kTS9
QAOFCqkYj9bEId5gBQF7zmTThlEFTbUgu7RV7erwaXmKoPIvtlKTWcE1CI1B0GRv2IdKknkjchRc
XJ6lfddvuoM32keiihhFVk6obLopRErLAGdVog1CdG2Rlxruan5+1100axtE/p7bS1xltLuxcep0
2+Tyeyac3fqWssMO4kjmqIhPY0frk2kMLSnKDm5Z7qWNz8jZuKGAtZNRI7Zdfse7nOyBTdsaBg2c
IVUriNEz7kn5UYFuA3VWer8ZTib8wMzFkWqXq6e8tuO3pQDJ7XLv9BQXDoT5uBUXm6fN6a39OUl7
EX4/si4MNByzskpnL6AS/6n757u0H7RlQ+e07E6sv7Mv3NsDBvtgCwhUkLnPgQyjVI1fExOGyMZX
cM67b2CuMxmZ3izfqKj63JIeNR3PLBnrs01qa4Vh++WaDu15VXIUuKL+gJx1YLN6F8abxdwnAJId
yFGyGxRkO4NDTJ3p50RaIkH3lhSfr4PwNLTRNHh95Bqlm7oNENCcVyJodCcwV9UT8HlXo35UQ26l
3852c0mUy+h4hVYyMZmqzpYAX/4xyA8+aCAv87dzVqdA0V3OxoK7bXfGUlvdsyUYBCVOUU4rMgSG
L7sxknHXBxo012HfEl207+kT4sEQdzwg7A7cx5MjEe78ytSmAzZUapkw7MQW+pMVEDckyfXv1kq1
wzvcSlfjjPI2wLu1FdZ8midkUYx8WN1ikbV1A0R28NqQtaQMZVidk/wTWbG5/p8VsJefd+YPphX6
uaSks130qEYR/cqo+6aRe8OMFZgQtEL/Ch/8uv6tE6Aj9Yl4qe+ZTkY0RnEGv0fXqtwGGB9G6mCa
H+Oss9WCofqvsH4nOXAEkVORNQMgMU4fXJPTpVWtmHr9fBCehST7nxUD35yS76qZeBrSwSJMLDCh
71xkMMJrNsKSi2ZtXa6g0zUM723T+DmGCPApaE/1XJWi9bBvoIze6xUZkeEIgnUGIUvKhW/5mBvF
z2Nh8Xc+eNlNJG1FkHaETo+f6p81V7UxKLI9qAzK6hCLppHG2gMb40xYqUa2NDVxrV8QbeSh4vQF
ZrPvNBtxsQ2PysIEutHtSw/Y6V1v607I7ONUSTAs5qSl+yZGo4Ugr2/fMgpv8IT41B257tp67vqk
k9UhM913fUJvPX7+se48z1wn0SBvB545+MPUDvnhbJtfCLgSyFt6SO+O7yJLiDmFRW+Hxa4ZtvZr
mHrjgFMoi64mZzsa2xlgNH8JE5phiFNuJGCfi2WXnw8AdlxxKg4KirVOtMwGxSt1qPXgmX/I9XF5
W5XooNTgSCybXMGxdF7COOX4RPL00e4bqXNMY+IRuRvYyhzHsfgP9ZTIULEAdtDo9QgKwGX5Ntor
2PHYa7bEbJbX/T7/dfcD+5EebXRJUyHoeyeB8kGl3NyT4lf3tsCSMnNw09MVh33oc68/Tihmk34h
0Fm2tGgNexEUBuwqGk1QNkqbufR/JcZ0/DPM30lJPPZ8kuWRmeSDN0lRY9FsE80SmEQVgTC1d3oo
aqulIaJrZnZHiwsmlMvkCiazJkRW3VctWHlF0axO0myNhCYVlUQnxAuXwAKtdWEWptlP1ru58xvT
tismcUH9U1I9X+mJWzbTGREy1/YJksl1iyOEh2cibPeo9XOrZ5Bcuzn64XLDjv38Yj6YFI4QwDZt
UQ2u2uxvibGf1R4Coaf2LgvuUPLKbhsFHV2pCgvgkAbJgqtX4YN67GrCJisytbb9N+zY+oILGvgy
H9LaIvAn7/3IgjDbydWllYyahXBkSrJyhcY9pEtCOQ8zeOMbfxmInIQdYv2hfRRu/JkmriyfBSMi
XMmN/9LUw8FTNvJzgb5sZapqrE61dBDAKWT10mBa5RbbNIzmwuBSR9yBUrJQ50w0cZ1xZpDP9m6K
pp+N2/yli+OfIVWGFHW8UxeaCWL7mluVU6DwA4HXA1n7oPr9xqJM5X/cVwp10QqNb0ouy+cFLoOj
gBvqNp2E6XMdqN7rH2Ml+6RdY20YbRGieJMMcy9VUy6vlSWvo/y6XBBTJNVhlLPO5OR4SulpBAzq
WCu6226h0n+fC/H990ixnT3jBU7XGU0ZkJXtAcw09QQEsM3vqJ8Keeh8td1ndogCf60Pkb4oAX4d
Q7vttbXMF0YHJSwhYy5gVnEHXm7OXETSu9/IfM3f/RhIEJwUfNgAAqlDhBuiTxEwtAemsYTP4hL7
J4+1MB2Mo2zkV8pW8WsxH1UUHA+BhvTTAY0dMbZq2BKivTJdmhfC2g3R6SVEBHVV3Y694UF4r15S
LUe/z9/zwJt3rcL8lVR5U372f4X0Bt/xbsc6e1FHuIUbRJRdtrEe8hf+wxVnfTl/lCZmAdCVlVPy
J0C236KbiEDLjA3mKUTS3dComOdPOAnYGMlA/PwdtMuhQXhAI3lPCcqn8rypBVmYV7NMyPcnhDR7
l6SmE09Yv6SqxEI0ndHxl8PmshW3yFFk8gM2c5bcqZM3YvjwlHVDFOV63ZQwqrO7VBGGkONFPVTv
66Rzl+5ugJC5+9zBmiJ9f2h9/KkkYMETU/9SvlmT6m7uD/TqhQfAFlYfacxe1O3ImODXExJGeQWP
TsuYO7Y8gPZ8IeOzemKkIJYDpU873LTFHLJoebCO8JJOFeMwtJ7aRBXmL/Za4otB/5d7IMQdd3TZ
TqVp1h+Pnr1fkoYfOv1hz1ZYuOyx2ooZPSVgW0I31bijng9N8dyb1s0uZ/dMl8Oo5HZIRPMVA818
1qJWc0uGHZazQa1Ql27CW8tI8qhiOv9MLt5OAKV8ekRxdCKzNMRtWtNo2H8MoKNDSlmmB74/zPMS
6CZJNwtmeyBn4juLejyCH9C9uWyf+8DJLje7XRCy2RVt6y+LFQqqdSk1M1EAJaiPNZjqVtydsJFt
JHqYAAVUtRQzj6cCuP1DKbk344XgP0mreQukCOVO/0esDZIayhP2G9vaWg4Ck+jXWDgcSCWVTmJ4
/BUfAssCty6qokeQpxAVCexUXTbqYP6yI6Rgt6bn2slMZtQApc4JvusLBZR9PsxwyzWo0F7H9Wem
egNwq5D0cdYWu5TLRVDqVCM4/wGw02lA2zx+kRQ1o3GxU3UMCr3g7xzx3S7rYlwc4P6eJP+KPwL7
GIpFSgi4ppb68C6r73TbaTgHJRbkH9NB09h3zcbSUmboaGjCfNzzP5+m7JyrJb6P+Q7Eec/G97Tp
aM8y8aFWQ1YK/lzy7XriQqua+/48Eu2BEYqbdnO/LKamwbTuCbqzDWweTuKuvUQChi45OMCcU4M2
Sk1jXtXY3TR+a3O1VR/SewwKt2oIJWcl4J6g4f52gDTgSNYiL/3BVjJIdM8CBlMGnuBOstPoyka8
hf5hlqJKkxZE/5D1ffTLP5Uhps+vTYZrnkfIDxnclS4Fz9NsilnW+o7BNUZ8PMKV5kXbH5QTBGB2
CqhRk1lBaXq8pzMTSyXcm3/6el366F/v7EFITWIeVIFOSGn/VcHxI+wDWkZCNxODUZuHwSV6hfKu
LcLAQdz1VrmSzdB8C0IqJpKC/D5b0MQUan/Ya6+niPn93VOqMJwH4niwSx6vfvgXg9yKyBItkgxX
AXfoBpO+N6R/n2OMgvuyx96kinWweguX7YBABu/h9VKba7NOaEVNENnPmep8GwCQvaffUWW9TAjv
8ApWSg26i6ceWxzAtS+uUAJ3EBhXtpQw2HDOpWqPQmiuo9k3rZIAvmdV4iEWWH+5eiJ1GH9uSUjl
+KiAgp46eJnECJa2eHmYtKqD1USJYIM2sjMQfhc4cajclErAF7lxss9KxTWOpcjSj3nfSsWb0c5f
Qh4DBNzfCEISQvINZBlavgcSMibghG8jH1wJAfxNh3koAauwteujaWImztTP4JSVTtFGUBe+oIL9
+jerSOKcVrvMqlhnN22RoIIhQWtHSlk0Ndk8ulDRxucPPW/04M7kSeL7Icoev4G8IdJRTtkab0EW
hD8trr/JKszMbSReJ1XciGR/ZQ7OfVhL+dXkrisZz3T5p+j/k2bWR10VK9dw5erCzthG6y/xvH2R
BKDvKmLhn8uMaeIw1BIG5L3upcJ3NDY00L5YyQ0szbclsVAS4sFLBVMYmklyqucDVrrrkjk9DdYU
cQbSciqgO4SavVZlebkTCQ+PxhyXlqmLAMrHFl7hKRm2ZlvH3m8rPH3z2nPYuHH13Z/mKlauC2Zp
+de2uASs2lBaiDUp5NETwioqG9D+mjFXP4uH9WQcgOiG8RX2CHXm9EU2MFS23Ylf+14B1GxUgv/j
oJh+wwqOwvb1mkncC8Lt1ROYUJ9vt0GmyPTij0m0XgcArlUL1SNxLYaGXLdRV4LnZrHc6/hijcrk
V7s1HAZ4/7f7ifd7hZ5Snw5vZPycKOUUh3QDTm9IRrUFUmqVTgpg9dOIlMBuGKxWhKoxIEodYOM0
f1FGNTGjTDlLa+fyCU0QDDdMOWaft598+pjzZdsqT7EDzcMSSFZiHX40yDuIYTrnHg/PqRB7dzwQ
Caw2m/TdA6Hh2mw1nBmfMo8uTEW3nhd/KG81adp7q1sEpPSuJGvWVjEZGof0FWjslJc4s7Hs31KM
7po0tF269+owJfsSEUQh68GIjnJPbIZRaAsc0jKkVLmBNmFvSGT6j5hpUC9t5IYoPhTv8fA7FD4y
7rtrpwy1IceJ5/PUaJSCWAbUdUZ/gVqTmRlYlb1chqRLKzLTsz/XdavbQpPXpCrDEoT5IIQGI4qO
1pPlVXaCmcs+68sFAGkaxEoPzxxT6Rd6wTPIjL13T61oUTmDvVhw4BHIzd9dZYJH4qgzlQELNw5X
8EIuIi2GK3G3w9gH4bKVvo+Vm1v32iba6fBRMpFdKMIv21MgF5KZq+0x6RKQ0jkhfxZmaxJpky/h
yaIt5zzlH0ICZMu1IHlhoiZYrtZyAopBK9mcxxWywWhQI290S3jG+icyD6yVXI/0kTO6V8GajvaS
z2pnk9C0AcW/TXTpWcV8NS1QuVh6HfjMaaEOOjyci51tDEVj2R8Zu/e6r3XUA6NNZhPGxcjsFFKR
mv1f4ZYxhrujbXlOGEJe0py6USjdaILW8uatbmninn7BCDS+Iy3eNkLursO1EW9+Shg50Cwi7BlH
110axVmEmx6A0XVbiP0pq0Tr+CYLEVHuiQ0qLQzm498Wjbr7S/zsgOkkIT9R5ndkZlv64Y6+jrui
hYrvZQAhXAaKrgV5QewfRI0MKTXki4t0ivlTJgbsmXxzHs0/pTUcnga2C2WfEU2ey3SLyFw+U2wG
7maqVR/yrUA6afJGxIKQfr0mHM7Ai15RuKz43z5YkAhIt9XTREQr8Cp6Z7nfFVL4Y1ceiitkg4xF
fLtiRY7zJNRC4mRlW+99mqE9C9qlVfxcp9X3tkHu1dg93Tgq4JyzblLd7Ucd7XyOx3AEEI+tvOdl
XvMdX80j53CWRN70XWczH0H5fTg9bUghct0FLytnz145HMfnNk5K1g0Curcr4U2a1swTnVNCEy2s
D1zJC1CbbLB1GuukIfl8Z2UiJQ5o6vG6I8AgGrW/HZFlxKabwsp07r1HVt1WuhuB43hmQr45NYiC
VA0a0PsdsAr1/HpLYwiqvR3VNnirNbiHshvTBuL0p24s1je5cC6F3cHcx1sd/eJj8xsSo1m5eoc8
N6WuBY5XCaCXtJzc1hHQbouxUK+ohGfPrp4KJFERircNNShsytBB2Tj9F0c9pC565OCs+uc9xt+i
rAriaI7JSivuXbj2Ff1xdjLw0jNhl2VOZ0m40g827KsgVbE4OGf99kLyUIeeZsnOuMRaPyjZUMre
ub3eSl4aeqztvsQSaJ8JgWqyZ9qnZ85I/Z1LuUaE4Lz3omxYOVW+06oPg6GmoXrHY99nZYAPyKs8
R3t0Cq1+Cy9lII8NUrUlf6pW2hdf0hNubVLFGRvizdAp/PWIHJOunF81HtP34i4VAYCAE97CcwEa
TjAX0jl/Bq7bYCvuNwDetag9/Dcsrnw/dXTeAHWWeDoiUN2YftNbd9p4CsOKIAfEH+8OexE6A+Ni
gLhbY7zE/IAON+pTqcPq3wzH3kZBWrHyhjozwJ7kkGV9I71YVcYjvhESaOn1NzfdTLmUaTWS/ccD
4lAzxO799T+CcHKn99HiXvdYrZQcCD/kuBd6S4vgnkeVmFWuOWNjbzIWntj8WgFZBJzaMMq1avRO
nuTHfvmmqA8bdSb7fk8Zup49MQfYB1g5i/WV2/PhPCW9ZWuWD4KtoVN4utDK09UY5jGIfZodTgPY
PKVN0beVZPn8lerh3D7xJzK337aaH9m7TcgahQChzRcr724x0Zh8kZ6Mo7sVeMT64d1MTjj7OotI
lu4Vd7AEmmcW2dmMGG8ymIrrwtwisAWbgUEuXz0VffmYXUvL8jexMZS5dPta68+IaXcf50ATeKP+
x39Lej2WN1+pbF0ODk3TYNW2jM+GYKSlWfgCit/UfM/zvXMsgiaZmrBoZq3PUjUfNNWF2rpSXJR4
CT6CW40RfKj3eNtj8dhKKqaBkG6h/hTnPgsYcV2T69BZ92LxMRTRU/I6qh2ddRjjOm09EB0fSC15
m3q9UanvxhKVkM3VAaysl43LUiW9rGugrSuPElQksiDpvmGQB3Jh2mHT7+eXFrg6pKb9EOQLRbjM
eFaLUpOd6u/FW9FlwhnOq/jJE2iaGjQOQoGypHQNv/ABns3FD1eUGcLUkW5sojGpbkTiftT7QiaM
e7PY2mqFe2ONqxg/lgTqjD2CWZuqYiNSmP3bOuR1Pa3MStmrT7XhxvistSurx9S072huBn35k2Iq
hi4ijeL9M/q3ej6Cj6AnSKVpOqQXP7hl9PNK2HzwP0h/IK33Wnjx0LjpD6raD2R21djgV82PVEzq
67elzA/7U3HUY6i5nH6Myna8wUK7sYw4f0gT2lchmQ/hjUepVIa3neH1H8A/Tt6lf9LFqPS66glf
y301x5iy/YbfjmjGjZPM8NcaA49Z20t5AOauDpOn7Ie38ENmTXsMtxLEnneAiXsTmoWTeoADSE3x
mOaQatmpiMMuv+0b/rfpaMEUlDXJoHm2dH6g0l8XaeRH1JsJmAvZ5cfqAr6qe2oRFHgc39C46RR1
bj2zfeFJpyLiggGf4IqYS2qWnsoRJyERlSfEZVjKDfZmXi5BZC6ZO+h1efr125fo8jcRPF2kTVZO
Ua5OV8hRPLr8CAKEAeglDt2WoknKm1BadbeWFMLOHbk+cqdkKTKKonPzV9SiNpK+2c3oLXge+M5C
H14dNCAcostvFzA3PHTA0OBdjii1eZDxk9R0yyXmsTqsHnywskMbwgkXg29B4bK3qOYp69UmA9W1
FAqWvHS555B/U8ZsU9DWCRz1UQw7m1xr/nT624Kiq6EAwLRqZp4w0t97ayqIMDg19l3YDC7nIHf3
tF4hKXAD8p73YK59NrEQLevcOzF4X6LMUkAQarE2pfyX8yflkCfF2avd3ZgrXdMY22q1F4eJvno3
/f7LbrOkxBvMEiEnFrWBdaWDu0/kJfQFpBVdCqgsnx+6P2Qtt5Bt2u0GtV7hxDtLBseGC50zPXPv
Tmzqx8I6LhPMucC+r5ZgjBHPPkL8q2XaYuKS3PxEvH513wMbiwkPD4DtLA+j7SOIh4KHdqNhRdWi
PR8SrBMLrpFEDemMKuAzF0K7zQw56L01vo32Oq9Gs09OooGSKFQn+w1EjGRN8AZwlld2bKv3yal/
eJWq+U9q+nocihtjaqbGA+AjzoDmP4BiarXg7TUoPMe0Dw6oJ2g5hv8RzE1COSViQOHea+BfqtBo
S6lpwXSPbaPgzCvHdR2PpJQZmXeLsIUgQr0p/gMjMJ3k1QaKpw6QB+fF57XyrlsLzoY9wL2fCjnz
L/ybN2tMfTPp+t+i215H6LIvdnf5XRnKnwTXm1ZnuqvNndmZFmdbIbrWVr/nu2t4FeRYniCt+YrW
1FxHqD8hjHFyTh1tz/o+RhxKGCvdY48k9oK22qEIjErQTUvWzgZ8R8OY87kSLWS1zbAiSq1DZlO1
zYj8sSKA0ttuiyHcV1+EQ+HINr8sJP+o6A9JM5K5EjAnzfM6NO99GvYurG7SYbGJKqb3WpPVxBR2
Q4vj23FEsiGhWf/5sJ0yoNiQ/sFy9QeqzwEUOYx8l3wuZ+rScKJdla2tRiqJR9Lrn+3MK3RMMAM9
SxyKuT8xKe5hkUG3I4jn1ntPT+s3sNqO53UD1I6AUtcvAxFL+sbpuKyulVZquyGPvR1FPUjC618f
zzYeyUYSrrm15oZPXg/CaiNuQh+RF7Gpq8WtDgNlPLnPy6RCAuJYcRNPy+9fwYUIUPyAQaj28Jkd
zcOJ1eDbQaIyY4JjtSeX3SQD4sjk4QObkLosZmUjAaaBryU/WMeSJsHketg2DIqLXU+lxY3KWsDA
0TGxzOTLM+E0tcy51BJiDMzNpJF7NqjObh6uu60jQDSe5PRwmnE0e2nSa08VL/aUJxX+aAnrRPjv
URi9QIT3PRnjolgzpbk8WP6scoXtibMxMeq7nSjdFdbE0a+48Hx9UxBSz4+2aB53ZPhnAUV66Ecd
dNRibTkfbCnAMivqGvFtgjKEo4Y/tedP4kQ4yJ2GQHo8UFv+k9mJNpGdgrwiO/1bETqgYO1jNSZ7
kvhOA3YbPGc1io31KqvG0NopU3SKL+qCeRbEoFjMXq3mep2scFtEInsyt34z6yrVb8vNIky0exlw
TF2o/vWhO7k6Vm5Gc0qpIekzDLq5Rmy8vGcKERngLhKH/aeWBOKYYqwMTUB4l0vaSzKYmsawd1DA
Ep3jZIr+cd2wVlBzbhspdFGwKtLs2aoHFMOQ0CJhD81dkj7aXXud/SWn7Dky+KAdEgYXWwF43EVs
8MjOKGqxDMZJc0JxqqNfSSUMH1nHrc4RzsPzxPxS5ucOxS3bKymeOAnP00Jl0UjljHcFjVTeFMpA
Zm/W2FypKFuPKvu0Nxigvy5WSrAt17+zcils8Qp7JQ45Sd1QoDu7N33sgDEzKT2c5pZwFmPq5zCd
eBfDbCa1MWEaXbGo+h1d0dTzGZhtzxphqNsPGq6pu76PDT7AgKQyH52iq65tjeazmlCnMtg8A7eq
5TzW5zfEqP5taTtZvOSjLQadkdlviFK44gYuJqFE37oUjoSwtvAs6SdSDszEypC49OFK8muq4XEn
QvPK1eVvUVl3M08f0f+BVyMpajk/xzkAptxIJ7KjtkWBwy6qsAm3wqNmX0GHdnwr1uq5dklCJte0
9oy8DgRsWlQqAgHmF6LEIgnlKtX7rOKgLPNH/zK7OlrSgDLe21fzOmOAlAR2khy3FJ7NsDclQ5fD
Imu53kjwwiVC9jGpJ+fZnBhGPaxLjBmwSuoW6BKvVmGZZ8JzwK2wpWr20QI9b+MmoBVnsgxeII5T
ChUGqcCG8QI+El9hQ0olsuiYIGNVn3+5RHZvO11eXwdhTIFW1HDrPfuJpUeNqwVjpEdmy19rIRtw
kaY1EIVfXdDnYlLQmObeq8/oi//Ycy1QOfIpwHKijOQRZWZQHYs2bM9QpVU7qyTQ/mLMf9awq/uS
d/mKBWFfCqL5KT9eizrjgmXxudD5trDKz1ZtjwshMyQb5nooqPmqZcIFZloRYDRYBLuLUgPDsS4y
tMyEuCvVXgsuGXAM9PpIYdzHlNJIsWqvl6TaQ/bg//hFJ96LcVOmn5W80byEOC0bLO7ixkfv0x+1
fLkFICfttuzSmHZcKIDC4idGrYSBk51tJkSk2fFjsF0TY5OjOhfjCC1cZCO3ArFRSMsO07ApHY7q
GqSpjqZb64HoPbfpiG15abryS2UZArRfzl3IJEAcLfQLSUE3E1rdEbYEwLolqHDUu9D2b3mNrQaR
769T1ou502or6hvJbGG9eIn3anv/f1wmo18+K8uPIC3N+z8VlB1FUxlOqzMmXPq0BcUtN/0IAhR7
7Wact/s7eUmaHfFsRaYdxpFcVvwpAjsmIcInlZsLI5534G1I1d026Vd3FKvyP9dDUGXq7UWxKwoV
bT96KU2FUJJSaQI4MRW7mP6S4x0aTaXYSkb7qC+GYhJg5cvsNcj/gqIm7zu+QcJZPRWH0YmCQH/J
pDmoSAARXHo0v5lhiiFkNrsgnJWWME7NgzNTPovhto0hrvfl4dQN9hgGg4C+i16GZRSF2VROepIX
Cq3Xs1TYzp5kP7oIgOct1Rns0JGg+pbATFcdMmAXGrRgpv8KCwWvrLP5IcH+49m+2bikUwfvbnbE
d/v9XeEptXc3Bl5jUF1tryI+Ot87mAJU44xgnMsiNTNm/9/ppJgJO13IkGCVH8M1EeuuF9TKTCAs
JrC/fKSafuF8GnVsK4zAYuqF2WyjngoLVzUnPEXfNuJsDSQ/IX9iZtYazEmRZEWjRAcW359eaFmj
dg/jupkoNvOx3+QiQ0t6GcZxON6TvdTqHdwxSkDlcF44zRiR7Tb1j5YfVlAZctgGJ1m2AKUR0xd6
2gGy4F/5qxN47Gzjwyj4z9opmUKec/JpIvRbXOyk1ECyrhlhU4rtay84WXoYPGJ38NZ5nP3Rg4jI
QajgP/87r+0Ci+1hh4EszB/sF81EovRiCSTUOF60e8sRyUhC5zCobrsUFlbzC/OyS3n6RIW9Ij8d
SE+HsYufkS8CJ7pbIvVU2z9G0vrJIlbCPYCnLv3rDUDXalni0yP55gowXoUInZ8Iv/E8gOw45L94
4BvYz2O1ooeObkyAQBjzRxd913IQxgPGpPRchpYZBgxZcL6wuRJ3HlwadflyxuJSiyXo5oag85ra
HmX/vm524BbyOfHtzpjueoO4yxTAiPuy4L7twDxd9RgyTCJwI+vFlsDemUYNp7ij/FjbA9ScUqka
ySfXGkH3osDJ+VQG5hm3w7gcoSxkBFrkbvVRPv5C0jaZvkC8ZINc9g0BIZBzVwZCLEf0fdI0TSya
7SivQXRU45dGXKNAsW+eOPmpB+IczkeMO0VNaV2Oh1QB4wbOCGg11i/UfMJpzPNM4WlAHoRogMN2
VO2HNXlNcuTAsMxNU5cx0qCVjkzbDKElbMJsvMTAmOwdYN/hR0Bi9+4qQWHLajlBKzLNL8cfenzV
NcGkawhkZPVsMBR/D+Tox5d3XyodGcRCKianzIJPQFCCEEJrNyVXHleSc3AKv5iTOCwGX/winsr/
vUgg8clNurUZD7Tq7MMQqSa5vfHhNit23pJa8ks+sS5t1BgMKlAPmkvaOX+CgXX27YOrm5Gzcig8
FWKe8nftBKpBZkgjYjB+qmcaH2oCIZ9j61lfNPf9+KlZtyb6klUAc7xtjWGuaT46lZFcvn5evTh/
Crb7iSs6dN0MRutxlqFiMC8acfgDJ+Gn2JIuAKGeGaiibB2Y12VJx8a/yUnHGoxCnJSCvpZ1gq+r
TIT8R4i99C3P6enkQODlMT8av8yLvShzPTVZnOsGT3Dt3FsX35V9J3I0GvjzVq53a0m8Fwt+bEq1
+7K+xW9obXrILkchHe1yjtwKtnK5ri+Bbap6LC2NyYxB9ob+WGw+tTxHA0zryphqLpO1H7njEX7w
8a8ULLfSjHb/J0qhhxomRF4tvsNcPRtN9PFJCklYxlUzqicob0Qu3eGa36XQGYm99acC/AwYgRaD
B+Z5hUCY99yi7thygEfP762ZfFo6pAVc7kDVXg6aTt57DtoWfkgUm1GmgJqezhbLZwqw5UkCJ7ZI
5OmwPcKjyiqId0UlOK5nvFuXfCpmnzJTul5Dt+DPwaLAT1fQHfsV7zxB2NMQ0ynWqB7trU/+AxzQ
RbfmNiWByCL3R+d42+4C9kRAVRrF0QjLmudeZGHQxksqtS/b+OpicEZFNqD+446Go8x24dX/aAi4
PSNyHbtvqUiqk6A4pejqyc3fnIdDIJi/ScGU1Eo7LS888AglXij0xoJewdQkiOSE15NEYAz14+kw
XMFlh73cW3R5UEUC+QHD4zDAdx+LyuhQdwVEUqDeHuVmqNtcvwFO65rift56j9MCka83BbGveFpg
PUBo672cvE4cTv2cSbyV91L/horLYs7nJC8nuyYSFmjb6WMa+wRnSvxZm86GARW8tnUxcbBEy9vX
TU9etLKOwlVEBdkuTHqb/ZmCJ2W3gzu3V6GJrvAlBiUcCz5514a1uv/JlZRZMCa6CsHjN0qH27ZI
REjvAn8FnB7aorJ7WcgCrNnVV7VLCcoyZOSkq6Ijn80xXw6YPTKtnXFP2BMkVvo/hXm80jqJKX3Q
q8mgSCZKbRwXTxx864hGLT0/NWX2EKFiJWqIudpoLybE9tajJmC8sAZgwn2xS+przfZOhsmg+2Kc
VdcyuQOiXEtZhYJ3z1DxLgszSi7G2gGJ0lh20Op9kWIMtcwtLB9lS0/IaoZmkhIMLJ99G4GMYScZ
HfTji2se8C7Xxd8Fz1l4v+DXr8dh7MzXnUpGBBUUdp4E3oDw9mnQP1ncCFYQa8CLcxeNTj1+NGBS
zkTnJVuryAECHEW9McVd6Z11liKnnfklI03GGABQ+NvzPStn3St/vJ9rMWbI8eeoN0owTIP2M/3M
r0In/uGzbK4JWfF546QM7x6flm6Vz6W3JDRR7xIfypn5sMdVXsE7iTkDpRr78vn1Sn73684We4uS
HHtAlUbGU/LhhAMZltdfKi33vC4iu3IoK9hRetqSReaHz8H+gzjHAiOk5NsHPrpfDTy5Rnb/3azJ
+lOU754wsSOZ8lFbfxjArKswhlEh3c5Bf4P54OthqDHJqpJSVx4kFgdDeCQ0qGRdAwiyFqS+OqoF
hxXLt3OyziAvL+DFWtJyNAFySYxxpChvSFYtcUyWlONTPw2o5aaTVyao3taxB/ulQJCtvCWje6YS
hCyaCUExZQYPqVXY8yRdrC87fdcllWG6LM2brR9X6cluW5NMmwCq6b5TbsXq8ps27kcbHbzqsdcA
7VZwKO5BzqygzRAdxhdYe7oLgicjXnYtP7agDBOb8VqO0WM+mQ5FriQqm/v15qiY92NrQi1MwAeU
68Wri/k4sqJskbiNKvqPTPD58wKkdUvkfFQ3cOp/aMsU0z+JmPlBshA/Cy4TSVKzJDCU2IFepZ3j
v4+C0o5ywOtFHmoTo1uSIyCbsBdc3sqPvQkf6wYspysv611wEpaeoAqIIZR3JgauN7fdRbCgDFOZ
AHRp8vVtiZEVHzY71qbVCBov7vxfSdcSBCxcnZTQ4nfYpqdrJ1OyRqmahMqpBxV5NP2hq6kf0Gpe
6NpJY4bY7vSn27QfAo0F9sp52OqYqQqFQ8wJJZX4JteYbsodxsv9ZUQPngwtignExn0sOFB7U9X6
3+YKx/NCq6NVEqHLQa3uwDgPn4xSKif1RGD8J0qkvCURIUDCZs4SJv7jwo39wICdemz4oOLK25Nb
hNm6qwIqwzvvDcAcaMzMF1H5EPbj/jEbrt5O6/uX8N49W/xidqpLdnslQCmz+dmmyVe8VglSASuU
VCIKFoPl/+2EtTV3T6NTeKSr5iTPSfTYoKZe/GVBNYvOx1wT1NGUIzLWSjd7xzBFSz9VrL91tQ7H
McgAb9sE4DhAB1Tpamvf52OXwe2SQt+K6AcHRb73ACQhFkVJTp6t5lh+0jnyQ+wvQKVDqdd8GGti
K6t9SRuZ5b6ApJJ7GDhYHWu/WlQsu0hOMtx0D9CquDMehMROGzk4CcH9VuaGFdJ1o/lmsEAJgz4k
yv2OuSejoWAfGrwEVgXaYwH8TmNQWbIDYddJeMbdr4BgAchmr6uWH8FYoEV2J17F/OjPWfH4MHx5
etUF1ZC/LEOjYzr8IG2oLdFkc/NK/atoNof26UePsEG63mAtMPwRC1hfIOGmCvBf9ZFi/6bY/omq
paxys9lNaLqSyDHIGvOwb2ce5annyKAEbWMKdUtYxmCZn1/XR7qdNx5jOjXd+QXBgBYvYGOxnWoA
FiDk0Kd7jhHXazpJ3GNx0EW70h40hrnNF2LU7VIoXX/c/xFST/hhU+1v1QgQNXakslTIyj8KK3rg
3RFvWY5BWBs4dRmKSEcazXMWA3/Gn2/1E84/OBpSRjJ4fJyOQCIOXrd83A9qqFk168VKQp5NJ8Gc
Ipui4KOP1J1hiMYDSzDyQaUD43s0WRJLBLNhgz2WSNQqRn87a1uUAishHxtRen2Ke79GaZFH+xE+
6Z9no3MRATHbgDmAUGTp6gCC5posuRhw7H7exBI2UeztQQa6zJH/xFSvBrdJg4WcZt8+C/Gmn7cM
cyVA0IHlUP0nyQDpGBx6hKr4+hpYWi3B8qndezzZktXblD44Oanx8REjcLFriqSBSwTYWnqhwBAl
r35rG6lRSnOGbSNw3MynZalh8O8h5ejIQAPJjekEd7vV2UCovv20Ys0+rdE7gqQ6giirebwhDhwv
4g371Zy1CMkLCQI+apQFc4HybdnYGNlAoM9O7Q/0cwoXgdeSl6TDER+0eKK4j/TcYHoV/awDffkg
iIukcWQSPKAPy2pLPh+xiroklN+WT4ksYkjpmaQHaPZOPoNqbXyhLDYSj7wjT2ElQnZ+pfZF7vvQ
xJYtcCTfIExRS+S/sQkBHPZPls2BRK4HulqGxsmTHbPBvKBuZahsngQb09S6+qVcQrxFHtEM9O/c
XuDorLki6Hdjoh13FlZqyO+G1mPMp11lI2b+3zvdMt+FWRmfa9BUJPpKBhEcHTwAqc1aU8WlDWre
sw/PnnS5C1JuVPVeuzBT+lLkbgWezB3KM6tvh83oJZD3WSSwObkgEQZe8c+m6BcFXtdec6eROigT
R51Orzqqpud/iGGXqmzaNtkXtArZZRhwr48/+8grSoQcjt4Hbx5NjG+aSJpQZKH986Vb1sKdnvtx
uEEH7E9zZdp/w9cFusg8yMWJn1su8G/8g9BehXyaUw1Z7cNC7HgWnB9Q9xxeXUMJ2ZFqIu79qs6w
1D1yhAYAVMR5mXQjvdEobztcDOb64mey25+gfdbh30GxurpTImntSr2MxPi3M6KdwccWVlQigex7
HXzVq9QcD1J3W/KUew+O+nIE/A5bF2GQNy7Dn0HSLATWB31KvegJdk91RSQ8aAQ/DDfAep7oLAUP
WMm0WK3xJ33SDeZjHOg1vqoNcsCbWTVS4bN3iDdJSZFRisv8Kb/qU0hD5C1aMGNbkpG0jIZkbLB4
tzez2nByXwLmHZip0DbHsw1okiInnygcZclyE8fKh2RB5KYfG0lfQfxduyXR5Auz1tQHU3spjJft
iLz/7sDkmFIfFykvz5NxgFLbfEX5VlwUAHkiJHy7sw6Lphk5nB9S85/RSI9rWH5gqng+F/L9+JGS
VmJOqytnj+avwK16r0nUsYBT41wDjR+EKn0RZdg9EpVlteYEOjKXaFakwUrlNpJWhKM3ZrP+gVmw
774RsWD6cA0/rq8150kRH+scyoe9fV9UT4R8gvZ1Y5McVGH+9w7asRW4//dJQ0E3diM2jCcEZenk
/r35xlreW8Kljfs9wM0A+U4O8b/4KWcHuhEBCr3lw0wdnbe8qxNqRxX8eTzudYQ+NNPjvvrft8AV
kaxWoHJldYUMObxGxi5RrAiLnMTph6/GBCmIT0V02VPq2ewkfPYcBVq+FOOprS+9VnWbinyoAu1+
m5U/DaxyXpre0nNF1ZqmKUud0HJ0FhJPSpZTzPvA+zrMzRmW3axKkOOirkaK/rQxs8VKGy7cYvHo
vkOjrsSkMBUfBH+6mY3tiDz77+qRhsTPYurBiPygYYl3cDWDzb7Y4TA7F+5FXvyRhXJOmWxCLilq
T7gDEVwCdcQmyJLTkTjrvLqwDGfdI8xirEXGYNrYcra2QqP6KEo0YJIcr0q6IrruSMFgxUD7dSeN
hQ6F0ZQtuYE4PQV73LncExPWnXiKiYb1UF6mVpKDtc2MB4vlu24nIiV7ZZ5e+tE4U71XdsTAiEi9
gwMyTVzYu3uXVUFVzNObJTg6RoIOLXHjBjL+OaElyWXE3koJS9nOMU1w6XWqGgyVGDQIAJFDUGoR
+KLH/JHpXrkEebEKfiOYYqr5Eq2kIsSSZ+HVGd+dArN7JyRULUfo2uY3Iu7gUEyCoP36sX8GivcY
mn57XBiVtw6FnQ6qeReN0ghYFBwCLVirVzYWRXuPU0f5V9y4oHQVmOD5yws9HnkwkkKkO/kZihXp
ZwVn11TYzmTtIXzfDV5F0hcoRJjlxEf6qTzwaGygi9v1ggjI2Ii4l9N+wYJQyvmyhlLZDBpXn6nS
aCyz5Po5yVxrFBVWSJ/jW3XwxYOFVtorUVHnEL2VVR0PC4ItEItZQJpCfWWUSr41bIkMM6ms0BLo
3aaBffyecQRD/i68qv8BThIcakWvVZ0RivDCisROmIlrudllTFMGWtAmoU2zn9BzU1UvCHDEGBy0
hk9NFdrKU5iZqnqSfDX4HOOZ7WAkXN0Mju8Tgs91j469WHcCi/T1nCxGaRxWpSd2PHE0kFGuO95x
aHyRvcIdhpPyD266johyyUCN2n4g7ezyc0Kj0+xXykjBGTt3L5zIijyo61ETs798T2ECYAP5CBdj
DUMKjQ1p6k1i5mNU/Zr0r4XqDhuAyg3HiGXazlVVz7UeLSmehhgKEE1EU0kSQ4fGhLJfpExUhIP7
tZWe9c3oxC4ApGFL1U02CCegHbF8Dpc/WlWRtFsQAKojLOH3f/7IHSOm0/h9lsH+GTBujjRdrB01
ril+GjweUYQH5UxCgCrD+OTS3DS3WZpBtOaaEZvLxL2IouZUbDnEuHivLhMY2Mq0hIfgeArS2jFj
hV/8r9ao6nj4h+a7Yg+vj6XIDliyX0DfQeExq2Ka7HV15Ht8PlOfVHgvGKDhGv4MYewV0533P0k5
6u1FnNGv78w0zAMnH6d8535EiC7+1JHnHGJcWuINwNnecEsJosDaPdz571mKr70H+RuOt22GteDi
HxkEJuua/FV/ns9uoH5HEeIUwxuRMTH6UgFXY1JrCcwBeN6lmJWcX+V8Utcl/s26f7lszHtOJ6Oc
SBF9iEQKy78aFAypqqwgA7Bz0J0Y+fFah2VRJl+SIKKOB3LiASUPDLlHWcRQZrmx/qXoiubUECA2
bH0APGQW1vKjlF9QfELM3r2KOHVHxjn3zsWIM32VCaVu4dpRbzd2PCUSic5RzPyhOdZpStjWDYSR
DczIooaJQzjvWazBEEUPA5o99IWUwFr0s1iG0l52JxZa3fbZEPmzGM442yD1oTd77Zl5lR5o5JsS
VEqlJpMIl2keLzSmlwfihKH/VsLdRWapN5ZNHsu0eoXE9dv540b0WWZo0NDv2LOCCsjvzr27zsFf
cxYQU4PkKFu+gaD5UUxcHNS/RTkgelpgSZOX3Ogqx8tjlT8Wfb6lR2C+F69V5Txrvv6FH5WmMGp2
E8YCvcx1dODp344YJ5Ee0o+S1SVAzUi9DmmtHCfxsL7fyFb9gCjCsC8OZCeoSaZL3xMkUkPVd3NG
bdcakVcsow+JJgXhybldSbRFbhCrLiC6oPeXlepNiYvTqZxBjUB29gKj8o9RHxShp2xXKJu0Lpmm
wxyqgPE8zcR++C3awC5gu8EyPWumwHpIW+AgjyJITBa7D8IyIxW7rmYGqzLRKCBduAqRbY3h2p02
GQGqsxeoIl2kszOVvI+aY3yF4ZMXOeiq3Pyv++Msy46GZ+XrRX5haAMkHyjqz6KwvraJZMTVccFK
+FSnEAJjKOWhQWdgYmlmJ5Lm2ZnRJfqXa+XDVaXCYbbtQA2a14GpCtOIINkHNkR5udUaogDDga0p
oZd4w3fb4l3Py1IRkFQrHXgNDB3hnzbAkCn8timO95t5dkZt1kFyzs52qj1QjO6w+0uxzHg/7aDb
fgPsDSXzMQmTVq/TcKE4SUmaSDbl6ROehXjvRMgiUwaMZPQACV32lu4QDFaWmykLpcmoUtL6mMrM
sB/14Udcn9GOnXquFBjCsy4/xuYSXsbZQbpvsu0iDCRz/i7C8STniXyZvRCSibaH3FAHfTYZhfNt
QKXW9bFCy61jpPjFvw1EIMJxL5RuGHeoKx6BV/AK2d2rmKxpUgb0HnYZ1dTO04/J9Bb5y/M1S/dp
SUkJm0/6FZ2Z2j1r9E/JyBqyQMvEcvsUfe3HunveHzuWX2OSUNBCWmFb6OOnEEic4RuqHp8aXLPN
X0tKfcZdSVuctrZ1A7wjQchI/vEZR+PCFnYUXAuD1/r4yF0qsSvdnkIdrii/m/bn72NnN3Ii+DOd
Pc/iPr4xwV20OMhMzQBaOJE/88BXD3duR65S/AdrGICI3pqH5CfrSkKiKJx1v42DBrR/jvqfQyP1
uevFAdILSFvPl1UmgM1+waiu/U5OzAXowfVGawgm7fhiwUobrUxA5TB+jQaV0DP2t1oOVTKwZd89
TlLvBuUoRHKSjZtx5o9dkBy/N/8D7o41ToihwIrdx+gcsId+4Wrwb+EVNBs0YF7d5+6qXvG3ddlR
IUKXvpBArYE4PPUf2RBYF2jEvCYvkrJdIjszIF3cMwsW96GM/IXzHJZJiBogvwbFaJ0VtOu43F23
fj7FRdtBXsBDne6h5EhkeO9PSFGTz2gcW6r2uO01KE11aYJJ0QBxPi2/D+yYVAzcXFgzIBMNF4wZ
+3hlAyhs22kvETugxyMtleP60KW2tu4jCVEcmYsvtD4Qc7iJhIwdfVgjdNV9J12mmZoHe1TvzrVg
VdaQ63GB80H9Zc1VrlEyPXg2iekm8w9m+z3vjZrXknIx9Vcbl/9cmeygRRCP1ahRnfKZRUI9xBre
3FIj5AcW4BeZrAZeGak/j8XIIc3BwhyJXX/ptGTfRIRgtXQD9zUb17VDN2GtfEoERmN3FEhhfwhz
6gKFFhw89sBMSnhVso4vGmWDgZ+BUlB9BoW1VUu+BqzvY5XDLyKx0NWBbO1CldF2gIMHdA4+ErmM
69mftwlSiRLKlrqi5vFRDtdkwu0YrGcHeX4+3osJdL0Io07/cTQEBCpII87FAVxwfOvmsmQUJhgr
t8/D4IP0dZR3yE8jQ2TRxV51R0SRrLKOCYKggOugde4mYaSokLVYUSIyvLvtdVPl196ZGUs7/zDn
s3XMvRRaoRrhkzwvHzgjcEeV9jTmdThayVjLkVvb90rwLP7McCLC95B/t9BYCUh5y28Yyk/KA39f
1vxZ90W6HAkQRKdczpuJxTGGNBQaBt4T/0XPY+11q4bDYk9ji/pgbD3OGxJKl6GEK+QSRCrwl/b2
ks7B5cGY550ZA3uo+XgG5XnZBwaULi41UYW4hZY1/JeY0J1e75HpcrP1ONoU1Abtf/luJA8IWvCi
/GOf9CDblhiT+rGOhrnTxW+H5Afn4mt35LkynEaQWzNeZUUH6fUPJP6UoFJJiu1MHEgojtX+u0Di
cbLREHtOVo4RYQwgaU0xDBDffIXTGEEZpOuDGXcy/Zph9cTJ8QB7Jp+pC47a6LlzQu2DPYuxPEvA
FoEpXh0EVXpU9VUhBAfyn9c7LfDE5Iz72Kz9bJyJVvvlVNaLFUODS9Og00L4ugMeXFLv1OE6Aspj
DQgYBBL2jWgFEF3mv8YsapG4cUzqnMN67X7SONUYgmvIwxNpO5bZM0/Qux5AUlMzqe4SE1er94y6
tApqJAWiLijduzTCgBOTWA4G4yW+w+vaBN3hc3yYuZE5xvVyuSI7fCdGZc/OTJjo/5f6dYfBFPNj
i2+QWVLTR7xNMLNhInPJH9KOtL3AUJSQMSeOCKt+IoWyHZvUBp7l9GkaXdqlswQdKvPh/RHxNWua
om2gdR5b28/vatAOhOANrrP0rOEXDu5oTxmNV+qXDu488BfMOLtjHwj3ju1/qwdffKqapHFtVEgP
paxOVW2M/tw4vTpwgT7fUWOw4TSJFfFGsvtUVEynHEcjN5AFoVi3gNB2oAchOFuKt3zVt8B4Date
uPPxdjuNTOzJ1bvzsUWoZsL6iirMiS4J/Y92C198H5qapvEe4P2zjF4MFi6zAasI+r3bgZI3u8SD
q3z2+sP9YNy9ickyWQKeads1pqPX3cYMeZcfH34H4b39UT5cIpztaP57udqhxehfgWiEHdeN3/gx
nxtAAQPtKaB7lhIubl2kIBakQW48EauXnGimF13EfgE/dV9ykihNgQZRfdI8kmlUzsBxmFJH8Z/Y
GxJf1R/zuTfJqnC4ImZDxp6UMFIDj8qnf5GNuuOW16bkdu7G+WgH3PkS4x8g8XeNIcPoVrMTHuTg
CPKoPBw/BzQ22ZyII8VJWUFnksXlUe0La/ryptBnKJFyI69vWAf3Xm+0fXrUiqnfxGeVgNWohtcr
XKXXhrpcGM5Ag6QV1DjUuLKp9jqtU7BmhGRdBXwPhG18cWbDDLj9scgdL+Gr2QTfpb0gBH51GSQG
Ln8YaFrtYLemA0rX51OSQS7LqPXckNKd4Jre7ZgQCnkIi8gsk2eUzWmTf10aN24o7o65OdYpxi2j
r6QNzAkyCPsL+F50HtkvcTUf5HjpPWtY3ODuEMoObAuvP2SItRrdukmoPVZ1YRPThhh49Idr7Dtg
PlzXaqK9Kq3UgWC1cfBi4M91VYUgPn4DSELbmQm4zxWwU/UVNQMJUxtZrAOEx7QW03W4MQ07XEZV
j3mPTfJoGn/MserMj1PLXreFkPlKFmblMxbsan94h9HyidRrZABXYsbObq1zx4Geq/q5LaE0gzPU
kfgNLXo1v/2z6nmkFHXnIpxtZyiCGyg4LAkTgr6meURIRa+u6LRbX5BASOhtwBZOq7KJZRT6yJZa
TJ5OZYA9Vsv/x+CaayNWeFolVqScH4J0XV4eMvQxpq08zBmkb3V4ez7Ac/VSiCO80Y3Wlp12IQrr
dn+WaSgTkBp3sKvfA+DGB+xF4DnCid7DrIuTVpAm/HI6cophtnNKb7Lrv+4gkAZu0P5FokwgOYqq
ckIYFEH+jTNFaI01ACaMAN1jEYe4b4hZeQCOYzDOLdX13N6LY63wFP6vIGusO7xZxX5v6EFA860z
qxr/ym7jEi1/bkouJbYq8Hfxby3VN2QVTWD9rml4wZOUxsNaOCuxgjrG5boAc4xse66ITwV9Bh8J
+76H5LhU3W0X1NbfbqqHeOlE/+oRd2sdJhAt+wtOucPZFlodnRARDRR+0+WjP8Rs0ecfZyG4WH4c
d90wVAtGr7b4jnSiQL+WB/ETLwKi008MhEdmDI9zt3gJJb7+zZkX4ZfyIYH+pP+ZDza5IcWNKVtI
HdyUdkZcbX0VZnWm5a6lAGuBo0tsjgJI8Uvqo9j0xrKR9ZEep03IaSOCiRY9rQH5jxCYNdw9xHiW
RiTPryTbGT+sdiJCRTIz0nl1KItpMkbXvBPCCLdTluLsthk6FL0Vh8sUPbe+ESHjk54KjJO3AAw9
MFwRrKL779RCvW/xiI803Uz2l3VyqUtyjY7/ikkHSken4d/SD0plHmltXmkEl3i6L29nmmCzyLht
d8y7LTh6xa0UBk/nr3emy11h7UfuCgriKtf3rxEft5EyU2XZ97yPVatEGjMCVWbxI3vRH4fPbMpl
orr8B4uXG/ivO3mGbEbEwKmeuqrrxEBORMWAMeq7r7Bs0MaVaHFdCF0SueYFhZlXxGp4hdYkiqc7
7y2GCmE+iqY8Ek6WSPZpASdHuAmFh+t7sXYfPs5mwgxYOpWOT3Qqa5N/lsddl1DPs0KTlQKHE9TE
9r2DB39esnG0vn4+IKp8U7fGW54g7bBH5e+NDh6LV/EWYAUDkM0UddP9mB8mMqGxcybq0RPD8fr0
ZTLaHxXbN87G1L3ssQ1/7qDse454D4Jp7xX4a71w0Ij9zuFNWqMMwzrKfNrspGG8HUJUHLlH6IVW
ckGE7QSjbGWqEwjUH/ymcgJnLssThNSlse8nCW02zb8bjL0LY6QmF46xjLrDV11qyzNoH+tRBdW6
M2+tBGTj57aygma0FS/rvYQVZ5i1ePLAdohh2bXhzn3+ypEiDt88sCcieU6jgq7qKM4Qtkg24Q64
ImCA1l5P+2sFb+6sOYOMbDfaGVpUo9sW96ijePNAFeBcofZP7/STnYtZpPtGBJMgEn0XFBS1wZ7d
DwLNlDU6CLsso1N/Xsjutqk02lWJviurBvKUYWcEWY7+fWbhUSe60tCVh6kJb8bBxGW4L10U+BcC
dCMbAOnWr+8D8BWiSjBIiDf/C2NOX8+LfbRqGcctUSVZfPhLrV7pqbO/3oFN1NdNp+W5EHzmJNEW
FMu7RDoAvgN7sBShCaXN8lV7FzNQaPZGfR2kLD++oCGu/j6jIdugOYtXiHgGjeroP1Y1IDPOtqfs
2NBzZexFotNK0od4Uf17OYmC0Bn8jkUL7EE1jlqjgm+d4l6AM/X1rKSZFyyjON3i0yueqX5g73xK
mDlmDoZza9rR3uMCikiD0Q/JEkZGr3gj9OHbhBvreGJsROB5ZSFxNaLe92GckS9Nyo8oZHar7174
j1adEVmV9zLJ74C5/HX52GGxyJv5bzggk7Tt172TlYFBl0tguZoFJKRGJB4qruZj1Au23Bhd43/A
GZK/1sZLZKQRtmHh0gVNDY1XiJwaZY3AGX4/uBPiuu+5Tkrj9o02SAezzI1QzwJIeYE/iuW1P4cw
+ir27oEPH9mLnlmZ591tgErOGf0YyyZl+yyZ0tNtgdVH84B771SH1ZzXzYXRakqMZlEtQeHlyFgy
YLi8zHEysX2foPZsexn5SW3GIU1JBttY407Mq/bHfREGn1BQgPuTA97vXWrmTIyoD4Pm7Nmj0ZqY
KqhzgySWD1FKVA+L3xmMMcpFKEC343wJRQ5SQCINP+rvw8RE9ehBWV8csFT/2UgPoHkIyT4mJZ7v
+N+I8bUlI7NIYta5rgW1J7PZytN0e8V2YVfvFtONXc24QbQlnamNTS0Q+6U/9cy356gDTJCEr1YM
Rt2XL5MBkEnC1ISa1cY+5MtKJSingNjzKVRYJWRRxbWLfDRrF/LyFMewPtQWsxsRk8K0payWFZVt
tf24GBhOkFXAQsE2r2OahPKI1imVIAVsFOoAeOdlzgxvjhaPTRJmWBEbs0jdWJ+WIXR87PFZLv/E
Xn5NPKa7uSWYZIGwvVhhqeTOivniJbdE+iUdCpZbuma/RfOl8QYN2BKmhwTviUqOQLaBVUty8Fv8
yeNsEmqC107fLihJ4clzzykiA0b5ebhjqOi4I5fGkbIS3DevkY8NzeIDfFfA3l09M0qJvD7l8/2Z
JmMCsjhZH6vrlfQm5jHu6xoBbkPbQ077L2P3frvYWwdXtg7MiPnBfGWJBELaHk9BRaZ1WNQ3DNK0
ouKp0NaceelA6Pzk64a+Azg5I82rRcE5K32OrFHUOI+z2v8be48eL+YTLu3OeXSjKzp8IykphfMf
hl6HTzCueydDwU8bbk8Ii7KT9lChLxuMz5JwNT/OLLMBOiKoTnshzmmW+m6Yg0hjrjsTcdeS1tqd
DtSSkVaBBkMvr/kfdDmdCi+oOaFfmbl5+EUu6KNQqnWM8ajPIbdM3at/Ln5zA6ZDhHRS7xvq1ZIU
HjphzDGfcpRpPDShiBO14Rl1D5m7ywjNOAuztDqwbPk7gZKgbymTK8W/46FMQ9FlLCJTUKF9Pady
UfsN6swNHLL/Or2bQZH6SCwGgj1c+FBB9kjx549AjVPUT/SgE+8kmdY9lMOgJRv7uc1MquXo63eF
l5U0sZlKKCnorDfTUtXmdkiYTV0HF5ZRPbCWCK9s6AH5C3b+j9hYaGcLt/M3jnDcvfb/u80HI/0H
Ocexnl95A00uW/MVyOCnTvx5FbbD21AqqxaW0MIBQ9ySDES2puueNjS/Rw/tQ2KHlhq4fp14EUaR
Wuw1qNVTYegFXdy7AlxdJ8WQroiwifeDc9/SuzFoOX1qQQel3r9v7EZTu9JVz+qi0oGUVL2xXRs3
54egUgyHcfH+UG5My3f1dJv/tn8hPZXLGN8xoxxL/SQYNgBTDE/6G3t7OvXLi8rwwaIJiPyG98GG
vkYvJwOrqEyRlB8EsxWtOpj8conQYEPSzmBc7sDTJSNDwe5Qb8/CTmiFRlbuY7xz4X4ecjoWuw6Z
mJnVasvFgYM65Kqe7WaJM/xkZ6sKqpImMbgTM62SrGCn0Z5Wcc5An6Ww3IVVfXnL03CAdck4Z7m2
uz5oErl8hEdIvEU0aIRD+T54m3RPHCIMgJWnNdkfrV5JQSb2Y5qcs06JGKtTBYhDPLWEOONsv+LK
DcdkCj6tR2nMjab/rkUL30RJeQl1cDugaHgXMJUU+5JWbKATrRp0lp37c9emq8M0FelirYDMiFrm
+nMB2q8HUzA/VD3R4DrKEAlVc0+thr/JfvPQz0Vrjvyp+JxnXsmqA0yPn5yjAN05WLXEKW4D2i9O
YLZVJxR5C+XP8XCGR1zoJn7IiPgQaOSVPe9HCp3YRGkx6mBIX1CrkPAGQLltQR4E3EGnVpMpVVla
qeIbMzuRdTci7VLJoahyU4X6Y2aDsbRUWlc0FVWLW0GypBdXr9wLphwuUFr1YX6a9A5h08dJ4RxU
7DQ5gRjZFLRrrkRe94joVzsnM2+P8ZMlEqvODKn+K6Q+23i+WO9IMpAhlW7e7mzdVTz3U8IHx9zj
jcHNcxnDYOJqhRFO2w+qaM6VuUQn7aqwiiGUzcaMA34Ldd4UuZdL4gURWidTbqHUP09psh+4NAH8
hDfb5a8lSOLtMs15hhCk5p4kC1/B1mGcCpuDEArDQxu8mV0zzuBJ45f9cgw6Ca2CF3wq/k37sp8c
Qidf8m6qJup8+LsFRIRfGnnvIby7FTiMPgWK7H7utbANoEdHK5TmxOVykLwEBamUMuDWwuyWddE7
TitFkKI2KrYww05y1YO+aCraJOuzUQl2MGE0AdPm9+lDFUWBgGD72RR1dFWaUtSquLNqLA0wb2V9
aqDdLxSxqdJGXUyDgtokQsePuFhISui5Jnfs3195ilFkm2oirJgpI54u8gRUqsGHee4MDNBTuLkJ
wZt5tgE7Y3WaCQ+ovQnlbfny5xYK6p2DPqPRrIYrmW2AfoWvyCzZsFLGaHO9UukamY5wvC0P0+/n
xVPWUbTTrdxDsGE4Q09pGHJ6tMwbAiBFe8/ng5Dr2DQtXloEYocCP4kZv0vAsiQj9jaO9EtaXg+o
MHZDmbrEG1R69QedX3ooX5k84rH4X/xuGL2jw9GvY4390oUBiOzZuDDO4xZSNWyG0Ax8OOUvTexi
ADBN9SlUldT5EH3CzQJgqEJt2KirXclD39J7601xmpytDxhcNA60sDJsDejweqKhX5qZTTgZRsP1
GNRWzvxpwF00M6M0R0E38vCzoW042jOYJic9GIwBd17vq5dTKFB4r4kjj9iFxWr3HWoFx+vpwniy
RwzrrWHny34kVsEf30wtRbxWN0WkKNqNMZ0Edbmxuz75Czl0zyIdJBMDF/tU/n3C2Ri/DBAbVhpq
rtYreg0u1ykos8AJhCXtd57zGdDqzSrJmjTiZhKIcwol4FoPnZXINeM3/xHuKCmAhXujyMF3lSWd
UQbxFGrwuBH1238ej0YUSDMfrMid9gfLNl6eIq8kMriXxmNamwmaYdAZok1py/7atpIwiAVSB6gk
UmBYYUgeDdSfAu5e8DPiB7jE1KpxGealfdN+xCrBJDS0OVMNUOBmgVqOPbfSZxN3mne+LFaI60GL
mj6WPWWyQ6ea1Gv8V+LQLN3fvQZPQahK5eamkD6qAIiPM+FwvghfKRHYuYv6CgC9zoL4e9a7scdn
MDT9wxc283P6JkM5O+LYUBJv6By193siu7lwLZxhNvKCwZMVeOO+2+7sJghU0O7Zv29+J5rcHIc3
4V9FODDs5xthhQhvKrPtyJJvuI9cl4xNiVq0yPUUjmApnIVN4C0xtOFthkuY99uLz+eMn/jvkQjI
aMXmszd0TKOyWskjDbTLM24EHy8TFlxnO69Q/2vcxf/bBC1atssag5gFrKMa3wr/GA5LYTUzjcUo
Fe/bm8RitU24iJriE4LIIEOETVxsnQ7ZeOF2WwztmXzZ7Cp17Rc1SYux19E29EFjvtrrwSUSOK+7
EuLbh0B0cJ8nSk/7E/UHlyuapp/A5MFaUxVkyuzFSw4EWHs/8VWlTmrAIjbKRJ4rbr58yEvgtAsd
QoDtKn0rx77pcIfAxlexowpAnjSJdWHz7Auq58B6W63c06OlbaFPGsrQ836vamkBCY4XzP67D2vR
AG6Z/xygB7oOVyLoD9fAdC9nuk5AjewLKE2uW8tZ9r6aIDm5QV2eJ1AAWv7j3wvDNobOyyBRT7uX
iPUR65vxWSRkek6ZD4oH4Rm8lLgffcLpEsAQxbZ46r2M2oX9yPGE7mosXz16/f6UXI9gXeylSPCm
KFD+Lmx9HDAXMxY08NwAnAn9KZHniQSNdRe8PEOOrjqv8M/kZCrOyEka29PpTs9xAuRWJX3hTQ18
X6Z3NzHm/TLcyuh232vA7zVnD3DtW0NKr8WyCcE3r9ZpKgdHnqQ6Aq5jcBm5Kguo6Ogg96g2B2fz
iwuBQ8DWNpNxU7h8BgFtdOkrTPhUtiyw3hpRlvTwk+n6I6tBX6xzmqy+FRyyxR3z9TfQIu8G2Y0c
gWsihMijTgUgqmoRY1cxXlFWfy94nbb/skNiL5Y7vZuhT9/OsZPaPdOu4xkLBT4+93/YAHgO/n4X
70zEiSyKg2+KpWh+YBmiWAEWqu9lWTBbT2vQ4RZz2ZoQahEoMKY+qo0Zo+QMhYlTKD4SrcvRHWgD
ikrnYYTtr2w1rgOIDbFIyvxcgGh1LY91PoUEfa79MOPFoW+X74vVZe3Cls6k51gPnAop7bXOpsPH
0WSAzlFYan7tjBXAU2QMem8pwwivCP/74DSMpsah8cia1kdyt6lkFhvveIFmJJuGpNzxyH4I0EN8
uaB4T5GsnfGCjcV3/I4gaYd0Ju2r0lT5bSu2dULYu9rjStCVQv1iZBFUowkVucci3u1Dj6/2yLLE
oCXgS63UEU5syshI4KV7phD/7ANkBBPqtah9pUhcM3uMnQcxtOApML4R8Pnj7IcjUkc/VeQg0c2P
2ihX8nLAF3NsWRndKs3FEB7BmGAG09DUm2JZ8+BQiw7AuQxedoPQ2e/e9PmyjI3QgVsjjq6XKrk8
F9ZkS7t5e/WZZPUo7lp6jMQN2sCb1QoOmDOSenpc4Yzo17rp1uE60UC3LJAlnvp9EuFLKvjc01iN
Ms+pdoMrsuNtEtRyPyUr1UsXGeAP9AY2fR6e+3gqbiU0lTlEVot7/0ueXWWiTy1q8eOmzV82qYUB
u9X3/qKq+aDKlrbRbq9yuZF7pNLonoib4In8QFdeQTjlcNpDbjyWOUPXVZQQAqrS9HkAp2/WETUo
wUB+mhdKJUoLXm2YuQinQp3eOT9PwzfAsDLZ3wHK4lnilpC/eKepYFh92GT+65M/BBLewd43afC4
N+kXNIH185Cp6ozVcbdZXvinS+0aBI/WmYN30dfYgGppw79F/D/f7CVD6dZIL2PIeA6Bt74qMggV
wzHv1A4S00HupsUuED6rGAPYaauTA+iFzSPZh/ycIhT3tEqjiVhQpdBhDwYGwMZcXQ0qJT+kv/CU
rOJ0g10Imzg9Dw3sxQlcihGUuXaDH6laN9e3s7OXw6i2fTDUIvpksqbWvMu6qqrGYT5jefFmxVLG
ReNDa14LvxBrVXWNuVU/vdqswVYgzpz8J0KnInOnGyFrHjhgQXEU9lL/ZljuPMp57DcMi5sXsETv
1L2tcgcljmdgjkpTHJtJsnhNFMkgJoJclygQ0xS7GhZsNTDy58ENLIV70fO73MgvTb6+O8E3GH7Y
CH4uPV6tmq5f7ZU51p3pae0UjQG+mFiLFDjgXqweYljRLjhzhyW+nR8dYZnq9VqXetDLMci/1rtd
GuSdRkt+R3RbWiL8PugBPcfLXM8M/QQdIxP9n3djqdNzc3+frwttl48fLysnZPwR3addWCucb4+b
9uha1NJ1gqLGVzgAi+mCOzVP1NrlrpwWQvwvGsuywXu2K6WOZHpUcfh25XGyhYCDjfe4x0Av4zOA
KbVot6H4twnMry7CDa5E6R1n//3lKEAh9zAPa8ls79u15TpanAVAd9wyJNTCmPvUofydCf5LuNYO
+tS2veNS42I7BYQ5R//ZJFq1masZNGxE+E3hjb0+hyeM06yQvDIqsRWvXSuZ/RPqPR9hPsJY03vB
WaJazcTYBhKAIXbO+EcDKj8wsASTUD/DlvSGM1KZkMallRXpgi8Gt+NJTP/VqoIXTruks9FNXQGH
4tc9f/FIW+PZIWQ6jgI/Ad+elVPvW99Aa67WtE/uFIpnOEXNEikdt5PkBYwRKgkSMXK5fwqj1bNc
yh/yufC/kf5+jO1mPtWd6yttnnb43hgem0cbKsWqK4eD0Rbmh7x3mOCO94aq9K0VCMkfTsTbl6ZY
CGXkDv1W3y3kx/hw7hpIJpabndAb1e4LvG1x+mnToU3dgEXj3iZDmW8OQVRvf9nMok7MSXPPF6wS
Y+CWRxvz1hp2kdzeU0fzlTbpP0fDEiworWLxWIqw0i//QQkgS0ncry/xM71PABuRUBU7IVvteitR
STJu1fii5ylLYayM6kgKha4pBVdqoN/aSIu1lXhaOIdfVjNJ0iigp8d3ClB8L99jr5HExI2Sx5Nk
P8iyGRLYB62wCCMY84Yj9uyDnUxWvaoBvFElj0gbWTezfizpUrMzc9FmcXb5GqM2m5wCxZRYwi6i
ZQX7w6FcFDEy9g4BHMvHTD6/R6u0i/CY6YOq6tPmvKWNoomnTGJZE0KirAFdNQywOiBCKT+dTqHD
Ji1ki8j7TLsbehqasoQMG9Hm8OUuGTrg1jlAuyQOmnqztGZAsk4NCMBthe0OoQ7qRkpMu5L3LQsN
ePAbGYzHP+UFk45aLT4xAx2Mqemes7r171b4cvt1EEhDB0Io+xC3D7K5zJL7SEX3A/23O+Cm5Fqo
mwDx7uOmzWfPEP2zOqATA6nGnBmiX8noOH7j5sZv4oE9PUPtArlxFM+vAkkwOyV3rqarUdZesYo8
F9wz4+H7ft27HsRhjgqndY+wV4yCL3G2v4b7szQ1g5k41GM8Ui9jq01n15JKxx+DXZn2T2Goa45c
SrpQL6H/ZLiIYQJ206Vd2Zs6WtI6OUOQ1pNJUuMlvP+D1xM+HXWldv5PJoFXD5Wa7LXuxfY1MA3l
aFouj+8r4vEqMaYCLRMCG7K11ywOyLc5AAmIZ+FQP9Mkkqvhkco0J+G8sCjnRHGK1ysLTp1iHFA6
cKLLpd+QfFtFH40C5X5CoKwlL+W4sI8Z6CP6BJq8V6M+xpRr5eITUSAPXf8Hvt8ON7EjvNqBN1B+
rwBmqcvACf5JKwbq2fmnpYCI5ybLUJxlrZgiGfzavxP5i50t4DPTs/OIO+f0mYLKHXD9dZ6RbU2y
kYQRRe8qBIm/coENezr+7CS0Y/mkmycn7dIaP6FoPS9YUzUemlKgjTwckO4/4yUTLCtyoR7ixLQc
0PQLqAviXu/vaaIeAoAGfQFKMCav+YwOELtEjrNje9lBeFHfZE46mAdM9xkZC8DCDieJRatISvaD
8LZzRqq5DfP5yGOUmYQofJ6CdGTFRq5m7Xh3wcgZlupczpWkggO40YwYtBIaQfxjiDBm0S/KFnRZ
ldFwnzXbjk+9r4+L/SjPvJIKIwA3URQoRVtWHGONWkJlK+BYNWlOGHxI+giAlbRQgFeblVYtKU1b
/6MOTdVD5/dq2yN750bVA+yqCoaagnafELTC23aBsK1WOJqqcnWLc+LvorMCpAW5ui7flxrgRlsm
QHusqI3VyU5BVv4ko4cbPprN9vGOZfHPob2XNTJ5iKHXUgKMqQ5KVQy2nQwISAkr8Igj6GmP5eBU
/QCfUoBydPkcfv5r7w23r2nI1y4kyP2uwPax4DXmRWKN4A/JIkZAXo4Sahb44QDuxcmOI8OrY+kX
zUxQ44PGaLZFo0SW91+MS3Z/3SzK/Cp5lA846Wg0Ium4DgjV52kHjCwqn9BbS38y6Dv/HdsGi3RE
mEaw+scGKPw5eb5/rL75MUXw9EpiQqTmeRKOcrBsaBX6UiWZS78K1GNckNModX4rMW4Seff+EhBL
yxznUgbS+7xgR5x9aDnlR2gs+N+oPGFM1KlfGqqduyijGZ9qJivRUikN7p5uS35k8eUoow5wNZzu
J1d01mfAFcFCJdvSqZgsZsUbO0VQYN8xUnHyyibKOScmtHlnBtcQLBM/kR+OQVkAW+/vXi6A0ge5
NASf2KEMT5UPziplQHMErWLcM+Jea1JbiBrkoWQKurvCjMa2mu3h3jT5ObMJTiIu17Qh3waGxtN9
cGoNiBj+vJXV451iWmIF5Y7J6xebhRceMHKDw/0zFZmDs276qLtI0ng5BZyFf8vsj3pn0D1E42J9
/NGOFhmzQwKxHjT9AgPpfuvLO8Xq956PU0pKGOrbqDXb+dMnyf0ZKroHD0vmmKU115NeIFubdINd
bL6+gXafccWWBEaNCq5/gqGR8WL7c/JGVc7lQtVDwF/V41Hc3g4c3s6NcTHwfE45XZqATMYpz8hq
14bMK3kNg0Qa5mqaQPxurYQkoXBemcMV/4UOf4FmD5emrkCgLjtpNR1bmXtVloMcT0WkpP5Ys1ao
y3xW6L4gItphFMWE/PJRblFdhOXYeyBXkfBLqqyw2migvMLbncq3YsC1eOJb76WlbI890uRaoJlj
EWrQyyfT3KOoY9SKC39DSFXfQ98pK3Xtz757y/aUNCmpWsaGnNGiRqyQCUvMsC08bgi1Op2sFvyA
6fZbsn36LFWxqBJLpXARYaeK2SoGleXjriukuv95lsigOvmwwSC6mGU5MFrYKZQxyqU24zTgUQig
mGUzjm7a9jqptpYLLJH029YgxAFC3uzTrT9tM7oFBHOW16DKHBSYtHz8PD9fXI8Q1hfNNfiIEWdY
TvO+8A83j0kpR+lWEGb2Soukz/oBUkAxCtnhFwE+D4pgAQnAZjK33ESQezVyrpzZLhZJRquQWsQv
vUgYd4D9X668UjqDAXc0hNyIx85BhsR6rnNAd4E6QJ1bybxrQGawNz+e4C6lDCM3BPbkvgQv/ckc
tdyi/dbR1W37HHpo50TZKBe5B7zcY6GuBPTLCjl9WYYF2Rl8bb2ak9bz2na9qCSQ6jk3aRTbDYR5
5EDA96Q7rN9dFmGWOgBN3kwr1l/0TR6ZGaiVr4QkySpeeXDEKxVTbI+x5JSmX9tBoi7OS+EcYHQD
qISPiEega0hmGZEZDa3vbRQkmvUxb37Axr9mSqUuxobdm4U6SZd3KKAdODFV9KhHt2sr9+Lpq/6V
yn7FIMVOaMj5YR6lXJdhKLPdOicnp0rcWagzvYbZxvg4MpvVIZ4UYHFDrYhHhzGvsPDcNExn5gDR
1yltbGc+gNn4DlgRDC8/ogMw6ZFx0LSgigYkJM8jYc06qouevH5XGS+KqLrDhIuBCSlKbB64SSly
jWLVZyO10VDsH3xKxQFcRioFtdEFaOSq6sKdcTzrsmX3nQT0pUEEwM1o01QCRcldZpGxgEfz/J++
MyM7CHDBzkMZcQpVSFJhR5uNkIvC7QWt0al45tYkk/s2+cDW07mArHufmC+jokLOk+QTkEvTeLYn
7H4ukdQGq1UTAk4w6Q5odAXrEFOIA4CpFfwfdvks+bBRo8zod9vJEgKq0+jBfCkWHqsoi8VTcAAO
zBOe5QQ5AlvG681j0sqj8xZj5VzP/cfaBhF6hnlVaX1wEnLywXgKwVmFsHtiBJfGgKuoipHi/3cO
FoR2O3KIvwcUM8a7D6iZ51FAxjrrAS9ok5LSBgO3S7MIH1iZ3J2RDzuPnpXr7W3h5YWKGFalTJsn
LDu+m3UveU43e767wy4Nk1aBNYpVBMzvn/adJLoyVROhVc0w96O0Q6Xsbcj81KbnH3xFMBcCtpxo
y3C2ZW5elt8Ppcg+o9KUJ9P9X/2eLtiX6TMLsfSzJGh66owv0VKTf+w7oOiim/sAW/wOq3DP8lw5
VCzSpB2H+1ab24bMLNC/pEtzjnEJF63DnvURMNBoA3yN+HBTRA9xjHv1E8PifQsxcrEOgGqjSDic
KCm5pBTx0PUnVrXlh09Z93ibx4dQmN/QOHzHfKh7/WBKSqDz2mSVoJDG232imwsfZqJCgMFGyZBo
cMwA0NpDk6CRsiluH751qyzPupDoUR9DOLsPfXhjywe0xjzNygWj0Aa4KXFbwEnF1vfuiZ+NF55t
loJ1tychFjzFW9FX3zAu2bkM3qO8M2SuSUWk6q3/TJUDfJVTsIRnEvayDB473Jdfc2WuofP/CNUW
l+GR4a/7zka/v7ril4GiB/2CRktDvZVPT/t3M0w5KycGDfqwuARo2IyBSGds582NVVMEsqCRuZvn
nmQcESUDQTKpZdCEFT44hOfyDJE9gBEzlGUy+7Q6t3I1NmX+oH+4bdD3g/6VUCB/s5D+londREhT
eR2bp9bb7UPydaL4EyFzZHF0RfqMUV1IVGS7NW5JolHSfQDQ2Edkb+UyWmKBRxtPep3DcwH8bF5S
zNYRmma7Fu/Db6CG9h6OyiNdpE8QwtRwtCsaLHgyjS2EkAHEBCXp7QRdW1GKCkN8k4trPIOVESnx
/K3TRXs9o2o3LvQzdRhAnIi1z3yQUfxtfn1ZIG5YQnJx6WzGIDXRkk8RjZ7uaHRT/mQ44Dbz1Idw
M+wiz3V+xABMCTp+BuKQjJ4t1M9EmkoUNn0kKx1/ypAfGf9v2Mq8AVcnCufsyBsuIAaleOF8Ttg/
1maHNtQtAo/98Enr5qui4wXV61EXSjFgBaQtLzWthbHjjmCtRRovLNeI+aXEshhbHdvkUGiCJr36
nbX19XvAM+p8Xb/TVCWLcQmDoLKCwsns/kYDRtZ2ZFLAZJ+TKv7uDvc5nA/xULCwpL4Gha2dXWfm
paisoqPWkyF7PtyXpQDvBOB0gAMMykWa+SQkSOaS1lBTxhBS6iwQLPKJrIaGIFGKEK4HkgUFk1af
slA6SHoa0mPkvHPyslLEFJ8fyth7WYQnCcbIEPEXgfc0vaS+Imic5YDvo6u7puJ8w+K4pebFi84U
AICP5DrNz6XWvoAFHOK0v9BB8Ay6jd/ar3gYt2+HcoZ8vLEXO89jivEgkNg2l4+bVr5W8eohQrdn
7XIm6JOLTTya/K1gYJWaMlilhfGbBGY3+9fPpyz/6OaHSGuLlGlLcWHrwjJTY3mSem8KUQ3s8jlr
u1P08Id52AL1M/u3inkHbKnSNg4mGqcF6QMUax4Sopo7KFJIFMHGxYaCMr13K4RtCp7rkvN+E9jM
sf0thG9ZCeyeWNPWAIm5Jxd4uaQToWh053ojosZto1xppKI5F7TUTzuhGKqYtjtWj7L04n9seft+
aO2GYUo2bD055FN000myp1ZUPTXgnsQZN0foSTYD6q4h5F8KCD3W1jH8lTENTf7DBI28tAs/Qul6
XHgvPoyGHL+1jyMfrG34HSA6L3ZhPZJAqNAgk4qgTdVJuWUrRXXfbRE9nSfu2W5r+eJ9/BtfT8hO
9U3ALlAeCSCGCOUq5iz/rCzpSFh23rWTGScuLpsxHR5W574J36bXza5s+e9D23iAhSFAcfCQFvH9
ZvsPN8/nDqwWw7UqZA5qvFjCLmE/Cih45uQ3sz07ju6RwRBK3Kuee/MYvGrp3ug7LM/CxU7EB380
qy21tuAPyOexDBie5XZohNSyinaMINlIb/eFt++50sgxG8eRahi1yDLml1WbTIO9wI/5KejVNuN7
VdpTdS1iGSsu1XqrbWeWBhvYUOjDa1gEXTXyZQ29TmdsAr6VJfx7+MjO+HOSnSH22SWxx7N8/+xZ
7zBcxvZVGq08yUfQG0Pa2j9zMUAYbKX7b8ls6M42i6p4elmn7FAPXo9OE94X6u5ZuEfV3UBhKKBU
G3f6x/cwL3QGwdLsavoIahJy5ATIxI3K+LwFa5q56MVSI34trgyBdjVtwlNJjn7UKH3WGGzj6FJy
/7ehe/a6sKhi7xiEFgzk4wI1EXQBl4EmHWkYKkOyFTQ0rP5l9aRHOgrKK5yQ+IY5qGomATzaXuzG
dxPHmCVqOJ5fesK1nue2k5vXBFZ9YE8Pbeazuig3wG4DOS7htJu6Cp+8p83LH7M1Xff6iOSbraOS
ZotDb+P9C+tlDLOE4eGP+Nyg/Kkz09idZS4ch/2+rWLAo7r3SkEXG4RLXhr0YUjM9rCGruG4PDAo
2vcnkt2YZVZOVig/OBoekilTLLXHL6m7Zt25+zac/W3WcOQOrJF51jpEpEpbJiUHtA972PmXlg6T
haPQJmAnur/SE9dP5IoQ7xuEAdkn914GtHuy7zmi7Bwy47I6li02br28Ap4p1fxJQC4z8XfJPlYa
gSseJW7tpOoU18M+URB1BTGJlaOp8Twe5m3uc9eL3nY851xMjnoAXexwb868E/XPL2U/TT0n4dQv
5XPoHF3eKd2f/0q5s/f4tUStuN7aW8sH1b7zcZbGWy4dbUxsZJvKSrTmUnsieWH2y+D7QGq/18xR
bZTImxpqo9QSkRNxYY41593ff5j8rJep4d1rY/Ha+t1rNBHUTRzdSh8flFjDDDecDYAC9G+lGSaJ
C8oA8IgIx1CZzAsd8KMRC37hTIiFMxT4jkJsodlFDGWXipp3ovCbtHrH4/j1EVZRqyqDjarQfuXz
NrYgH5TIHcmejMn1g1B/H6sf7m8yiRBCC4rUHE9l8UJb9JxTWguCiMj/b3U8KrqkSf0PcLGVpzSv
Tx3LGfoBPuWGi8Iu82W+buWNQ9cT7eWH2TgwgsKuXg7Qw25R4xgDjMme4A6isIFE2QTeAvP6M6hl
bDQZQnYe5r8axzC1xdzsBu2Q47nHOXlKZewctIvWcXamhtycyl1t4DiL8UnXPj2ujw2ttaEfb5YD
cK2fI12aB5xND4y+oYWkTqSLmBmJXZAXZvv40j0qrpa8hTP42KXhW1/J5nbMbLgaK9pHmtKhhnpK
fOjh8GEhb5Y0rQDqGeejdB3mN9iaFBCeT+qYFlev9qKTrlH/TJUxRjSYh9NXPosHhWmFnRloesKf
S2WNYSFdVR7/MecM8U2v0+S2sRedLb9yZErzJvOk4bps3+xTqT7gs7t916h5pifdeeY4FzkKlcIV
mVIuOfQ0vIRnxl6avO8LejWKw8lEM4mkIRiwvXtcDi21Hnhp35oSyjAq1E260z8zpZE6dNzvLm5u
eR1ObOpWzOiaGOOmcWLklI/xUsTn3YMc5QFP5F3P967dunVXTltJqPYn9kzD6d3c9t5KI+U/gaiX
bRsqGJUtAMpcX49OT2ZeW3XDXK5Mjt3M23+aK7xURnCNyT8b9sZS9hxZnJ+qkv1T///ald9uEh+7
Hh6iurEl+4SZvAg23ywJIwFRU35jamWmi+PoNO3k55jSTnkUQHiwHDaH0ms3P7JGN/1xXBCmCdYT
rQwf/Mbo3Ep3S1x5gPqldA/GaLx5wamN/kMJCIGglvTMJMh44zQ1yYf/X59+vM7ossMjitSiape5
L6MlWMJNNGaxA0rMJF75kmOHD3gZbCV8vV1u8Wx9/hCmry8x1pJfy8LTJLk1Vi5el2O2inXG87hl
sJ4DsExBMqH+s6q1bCVuIMIEzzwEJP6cCs1w4BA/b/vt6Vog88kiT0sE4GYJBBgjNtw9j5n6tSMM
V17fYmpqDPGdxnmHyIcCXdj5mtiTpU/29IbJk/Y8geaetg8WO4ZKcOwrMMODZYs/76bd8PkXy3hM
eA3GQDT8xr1d7MQTq6vreQIFGlSYJG9Ic1VTMiFgxci+9fm/lrG//w849u/WCUWMGgdCocwS1J8Q
FD9Jo+pwD6LvZLZdi0iY7N0ySKlT9u4oUWYb4qBCf2C35ABqGMGkJy6rjB049xrnMAyvZPW51RBw
sZxccZAv/D6AY/EwScONbw0HkPuWyxdxCIZ4d6X30yzba0f6/l52Pqh7UGRaIR8B6BtexgN1QSMM
aUFDj+owDIlWbnA3qXf88wqvOV1c9Xz27kmi0sBixwTsuy1CouIAR1GA7J6ZmT6n8PWVUFpqlHaw
4WPQ21UtEqQw10WuA9t3k4H2gY7mD7CyxC1aID8qnUWxb+/3DOWf1R4CQc17b3NRV2s0hShYgVec
O6PGSdwwnGSTm2CLd4sZqFDoK2QXXeJmPbIYK/0zaJHYjiA2nJQiSAAfKpo3VugId+dolu72tu3W
UlIuEJnXWL+NDnmyGqjEg6XpkAZKVr8k6Vt7MVSyXOL8yLCGWCxtjcmBKNZcCPYej+FJehDALH2R
kPhG5KO/+sByjNdIMYggUCQ7+uVpHg2Ss5Il0CI0Q1s/YBoLXuuw0Km9D5Hkw1IDzW7Pln3jPd6E
/rcbWtZ93WDoHwAArsggQOCciGVO7X5F0lxMfR5xnoFcsHRgWzNcYGr8FOA/ayq0H2qNzlocaqm7
PsgQr4jh/yIR+RWD5FtzOtWOlVvTTD9Zv28btdHSEAz8Q7zNz4tBxnlmxYH0SX4RfXurmJtIvzk4
TjFIfH5Dj3GdYqxUaJcNdFjMGnILzKCKXUYWS9FBcmaD6rQjxqO5gxRIwfrdZLVnDBLlKo8MxdTl
3Onb7jTIXPUoUoG3qKZffLI2fQ6/uyGI8lQNvh+M8CT4VnTHfRFjSEp4xPsfG8LhyFRrVsuhYLff
VGaxXRxRy/j4KpD0juL+UEsR4h9EHKxjLsu1Um9ebXA3kWs/D5HTqkolkl8TSQ2JJFgE6CqmBicB
A7xWdNa3xXgmuGKReW+bxuxuZs1fl0HF2etbNIyNRB9YHy9reLC9dn2tpqOSbo6mdPbrkv9wE1ZX
tulK/n/Ug0CkF+0z3y3MpEDs/keuGYQ0CMWqgCSrDajr5msT7OJMASpLW+UPcVql0SUZfc80SDES
xfY8o5a0qGDHvTdnjZCpvGd/AXg/KH91uTrG2VtLzOUsu4gH+T8IcevT/EOumFe5CEEw0prqlfuJ
+c7xJdcEUPgQNE2Hf2yL3OTGIax+RVzrcOT3M+0XyNIOBegJhok4zbnkFBaOJZSqa3/bLE+9nRCS
ngUcpMes05rjl8O6xS/mO2Awc0PetAQdiPnUvU7WNsCEa2yRnop3c7UvB2k1wzxwePiHXB/QE4i3
4xEYLdIscmg0owvnCmoV6C0LReIEZwlcRF3aKer2nePyfeOsLsJTvtx7x/iGY4rne/xLA2oPDCLA
Yo/XuEDex9DuiyBn89rWlbe6y5bKU8tMcT1EkJIhQKbtrfnWLhdWrYP6TU1XjOSkNDuN7i2HA0R4
Q17KxwczrqHsxJmYEZor5sv/NQ7H1t/FXdFCpkwXZmQZ89pGto9jzBqrCjiIuMqBfgM0mtz4E8KS
MhR3I1D8iDYSYlJRuLTX4B/c5K6je6qHXLKZa9eK0mu8YU1MOi2QiH1+XJHzKBsXVKbpkoc4h2rM
3xHueHeNqvNydmwOy12m4wP37sgGNMyw0ShnfBzJQNOPdSV91LnZGpfGFPqFKt6UMhz1uuZy5UmE
kjN09uQLs4YUhZTXtTiKeJaYCAf4wPDpkg0asxogLbl7czuVdO9jWoDyDe2bk22i27FQlQ3BPNTg
S58tK9+8UKcGidc/DlA58FC4YTKW1Oum+/MSGPSWrnpumxUg55gJ6wwXMjrhmXSUFGcKRPUVY4L9
BotT/lmLOZTHTk2EnGv+cT1PcaBDA3OeXN49Gzl1gzWvCRDsIZUkQj57jRaDSH0eu/P/aSObZNJc
skaLIQATkQkgnao2UvcFlRpdjrQfKUILMnrX+I5uQpsw879BWtzOZdhcp8k30ajVXtG4tSFs+0uZ
KMOifEsoql/EifGUjDMCs9/J3SoEPGeS8PMSWYg43WurJZ46sTe9H7NkJWxjIf1l2QEsuTGRhStp
d/rYJ70HVf785NNgo3SQu6APLr40PtNHDvz2qahgHCXyTzjau2O7r8/EC8kjCc0fSqi3TqBQ9MxD
QjDpRj1VVxF3YRkfff8R3j/WaqQtc4WSIke/6KI2zLOBWRISmEOMaV2TQ6lEfIHH+AkD1CEouAJB
1x99+HjcyNpst4a8TH2yG+ryVhB0iaXK4hmdhi5v357fk1j3SSrmhtY6QjmeQvKOJ7AumEacTFnc
Uja2ns4GpFO+iR1mT6CsD0/eKYJuE+H41RD+A8GU8T0pZEa77ce3ddMGMyTO5ZdjcaX4JhHHIzlh
w516opipCtMuCjgACDcRilrsXPfllbMA5XSKuvcC/QCXiy4MXhojkB7FkgqpyNpwpEj+/UU9FuVD
amndeS9Hv9ZLKrs/2IDxFUvmSFc4vLXFcgokaKk4zcvubv+UgJIXyZTluEFzcKoLz8RH1Jk7BDE1
PonHVgSLzURd3ax0RBJVad75sfGo4u8rjNcH4upIE3GHcrRWz9N4wXcBl4OT3zXM+DLiRgMLGS8+
BKpJXgoAbUR7gfhlIk9/GTp7hX6VUYwJKg+QkNDYLTDm8qxm/kZSKxMAxv4EQpXH57Xn9g/YwWl6
iL5Bp6hTMjmz4OUmEEA6yS8AAozqgbssKGgLfV+LQbmU/bvUKFC6ugoCI844oWBhEi/14wMFBkTx
udxY7vTEYAcMew5UoTRX3m7S3wtG8kSuJZnmvIyKpKbBiN4tpK7Z7E6gcfOSeVYyh57IZzNm6LAy
dovZTdMr4gyl4HLWGwU4JbjU7BgA7aCJs1AVCUaeeYg/UxgED2hATeuTrdkJboQQUEws2v/S+kTg
xVrOHlyfkTsem87DC9qkqKJ5KebHN5UoPNHjMoTxM6ZiEo4ATeBtklt6CEu6UCEv6U6bQvAZrpNs
z1jJnBWkx+8beqvrnPZQlBfEFSybO7xFbwPqePmeLxHbqbGhpbOqUWHGikunol4izrKdcPbctD/e
B7X9b6hpcLVX+bL67qfif2w0QQw5pB9k7ByZz45LhL9Io+DqtG9Qda6+haCIEy6UyZP2kb5dVjOa
aoBfD+rrdeeY8+Kn/A+rpC7/taNLjj/Ho25vJ3wbDkHieHYs0FV7fisW/yc8NumOPsrmCVfXf/3z
G+hoR9BXMSW0eEDgG9N3eKuYHB6IL5znz6QVcsVc7aaYCzPco1D+xDPBPr9xmrUqC1wt/QDPAci7
5/4mAPh5TLbEcaiX8H43L1/3J1pJ/YajSMjLsE7x1lS5jHFjpta+AByBVula86yq8lDAhQQmnZ7I
SdGYi+8ZZdN1Zbh+PQjLAeNV+Ua1ozWSpXwTeTXJEKiW7GKwDcUWlhuz75O1lUbiyaTJ2hI3pTpC
9ZhP5sfRDuEraZil76u5ZrrnNceCnNpjFWQ/uA5H1YOLTfmBgLc17WTDdWBJSUtRWpDKPMh5dOss
FZ5lSQYFPr9s+A42TEpFQOy6/9QByA0cYQ/NTxhAzmX9deNIpMg9tIQnrQi2KZ0cXGTGh3kY3yVI
G4JmeNepG6iy2ZRol4XjlMc6JPTmmDgK2IVGaQ7jIouXrRyzgsq3RqsgO64h7BRPZnWTlwxtX+o/
tJIU48+O/a23rLuAONjNjbZqNtKBftrec5atZVlPRJIzc7vOmVIAssl+98eFM3vLe7SOvMkd9E0c
sfsNFHdSha2/yGEqFiNshBh0y6b94mqkf9nqIgZ7TQIf5+2Js4qE7sb/lUjFPgdLxPFHElsbcEAd
2tSg0qu+mSXpit4QCuEjF1uPLTiiTOHRT5rtvSF2vE0mQ2iPKWNzhXkU0EYcdNmzmRwT+LsufZHb
+TMb9dca3IoFD1GK9/tKXDHhhnbRhWLxT8MZHU40nUEpaXAnsn+XroTDu2x5uDqS9CU8mSGwg32O
SUtFowHJuKTRWQbVY34O0X2u/5zBkpwyrV9dkz7tvYDzvpdsLLp0M8azR6Lyy1ezskCxMN5Z7svI
UcSGa/xK227AakjkVjCmteD7lxAqNj+iraFfl5hwGvmVMRoXj8pk/9iSnpyDUvU3iOtJF69Z8CD9
qDrCCjsWSCcWf3iSE7dTT8p6V44RUZqIwfGHjflHn04DnUbRzlwdqStZeoXYyvUearujDJLH+lXz
gl3fmdv+2DZT4HPZINFMUOeT/kD9RPrDvQui5sTPF2eVlWHSpwSnowMAIl39QV8p+UvbIFgElGdp
/mRbqMeVV+rp1KhGSRc+ehHu2/bm0mLBSb0shjxY3HZO66w+y3Mgz7y7gbZtkoEDAEfVyceQGh72
i83NpNc24kZKRbbqRZeyHNiunUFD8db0jTGJempfEB5SLz0zG7DcXvBd0HWncOn+MyCBaSDqTcty
oUHHQiYbJIGnec4Des2b5MPGQLm2P/BMABlUYvVmoZQc9jTrpx1GR8aneYZzAZzjruCjLHZ48oNV
Jhrd2i2WNHuQak6KEhBPLxtee2N84A77NLLCBEJWk8slZ35kt/rFD6JWuHe0atpR2VHONUEqGIVU
nUuRquB5wevt0NKyGdvSEC5vsPTxHaG05FqIJdEtVw0SjWeGGgEbXgFRmPRQXaL3lUi9wqTTQviV
piJZQl62tb3ec+DUtVuQk3aD15IY0oDWuBzqnhwRBPLzL8YTRVtEFk4NcN1OjC61OxfW9T0WHroE
+KeINT6Z+XEQbQW9DvykBBpPXQcbH/746SnD+GkgsWVIbC8LFh9wOBg7DuCVpljEAxNv3/3kjAzt
uaPZli1/uICXni2L6VaKmW2Fux/pxeVjNc4c0EPyiG+GtXMbDtCbzEwy+v23juWyR4ZkSiuOf36d
FIJABZ60Qjz9DTdHCjqbGD7aHD1b4++p4hC+Oxc3nwE4BWoRs5LYFCYXkEYdw4n5zLc4HYXjhh3d
XZn+AUq8NYfsdgUFHsCDGGsR0Gl70lPj8LNcXaY7MUJxeRpK2J6GTXMOVqvkVHKG6Fd1PrRVp9a6
XsOM8FTVR5DFV2Z4LMUWif8dUg9Ibps+/TkpUVgzltGKNz5n4HlXgV0FrB7C/z2IHHnDLWowI48E
jSDXc5sGwWkHRpeeaKH8JqCrAjUxNAOhf45AVNzJwmtKlI9uB5RmeFb9Y0uZ1wkUM9o5V1asIwQM
s/95msWC/2oEY26Xa63oaCJATyJOWc0pwUL67MSKiPX4igt35B0U8zqq5+oDNpRRDtFXI+LdkHmT
C/5qRgDMrmm7QGcd8mcw3mVCzmkRD9iRQAQiBv6SSL+nCnppBH463eS7uN4jQhFTtgiBto43AihS
ubJHxD2sbo7tMRBrZx3mLbxpRuetY5nOXFkDGOgbdfyFZezrL6/TsS7/lAfFQDMUzH9iaPOf66D+
lK5s6Bni9eCVdZX+gRjUauQL3qdOBQRi0bB3ibn21SVcOXAxaEU7XgMhh5L9dJNpzPIiWERSnNlw
Yd6fZiD7tnw0jdforpC/l8Gzs2zVKrgd4D7tpQlP1fRTU1RCu6hodOkV9Hyt4Lrn+f2WvwmnYEqI
j/polOTkdZczgbkIp80TAvUr+IR2hEJ1iQsxTRJBtvnKEYgl5uldPMRgwqCM4MVY1ZI2eZZMuNaN
+61Qz9pKnOmQe+cuj67yAyZQw5Y5I6pFCzwX8esihgPBs3b3qxrJfPWEwOSscYNFtB7ufWwcGaE/
qgjtBmnEEpKMupjSpIkKD63tv78/p9Um1Y4HmvR2I9+WUPLma5iYGxXYabnY7OpE02l5BfokIDEk
ItiNERm4/j/iy4nW9VeJT3F/PTsmWo/CofLuMezV9BVFdTjLrea7P9q0NENQ52mLTOIqd0YiLdoq
3yAvz/3XlkXvZNk+BjfhlliGFg2nroq5g9spnhUG5J5W6vXW8TVec39cNVB2SQA3+gyJguba8Sbj
qW1yk1PsDhkm88RfVGt8mkAjx69boF1+1+MkTuxCuvo8D1PPCeBi3xR7wKMYQ5AWOrzOZu/VFmid
aF2V/vAkHwpqjBXZPhaz1GQAyso52WxPkURKPgQAWaV3sNMPWokkZPD23Y4qzlZdVuepxXNHpyqs
+qu7h1OK4l/Ip4ztKGcEnn/6U8HP7fIVARwQYRnMIOgIBBCKq6BTS18QmxBYF+7Yr9kfZf0Kvrhg
WUKNlZljjv5EOqVdgN3kYQZhnZfZve2Bw1EqvlHiwzwpQ7sql8+ycTpwHhzg0FMahOLJs4QLNkYM
GVdlkjMLYMA6/iFYvPapRPqnT69W+6MsCV6iXJT8Ozl+uQVuopQ7gyJwN4UtSwkI4hYLxHjEw4Vs
yCMpaX8yn8K1h9vP9EimHueuxqoWnnubrQ2B+dE+saeBVe50i5ZSfh+tYB/YinK96sC+oKvE5Css
DIaLcvoaKlmXM8YmvOEzW1Ummg0kEhj6CUjKllvrIkgrOZnS7lFhZFGSWwvDsJu2+W34xpuznfZT
d0rwu0YfUCN+meNK7vv+xeFs9djNH30pyq1KJhbCh7NhYeLa4+5G6QaA5TwkU4GtIneqH3xlBpw3
7lsb5kXxIbnPDQyQwbAldVtlIWxUjYGyzCK2zyoFsSp95bdDmXBsMBVIECpbf/iGD2u0HNeQIsm1
UQsnNZ4kIOchJB3TgB+1AzidEl3cRs8HpRhwSYFBy8Z3iFfQWOo6grCdcU4UlAJKw68rFLLOCr8U
DIIha5+X08iGZEbnBRMQhytu96oV2CDEaYGTQpSgr5GPmAs59FPpg1a5xY63X6hwMF0+xgKAFCl/
5ErJH4+0mkqdnQoROXuklFKFjBcrxtgN5VPdTvWbCljIVrgzkBE8TgOAzv+uFwaKYaBaw2ODqqU1
f3ir1IGoic6G3Xq+W9jMpAhmo+7u4g/jG22GyBr7qBY1ArpGX9MdJPv7Vs9mRO1d4+dqwJvA6hL7
t2ei76IdiDWypGr+vcIWAyXulWP+d8U1Ofezc179hyaTbMYX8kMRHS4l0hCYqoM1pXz+1qzydi6G
1g2s0iENh7Zuq3NLX0tzz2csvqv7RK6AixWViSkDvxF/iPOowlCeUyXNr274g9VVHrAwJYsFNX3e
W96AjvLj2bWgmkj8FjVNue4Rt74XdWhpawvjVRB8Fg0wrV7+v8GzkbeBLMZZB1Y4ZJTb4vEI0nca
gpBwO62mMyiNrjE11aBeqMeaauGdP2NCOV9Yt9ZRZNHHcVDRxlVlq3H/b1gOyTu2UiR1PIOqNu4j
gsat2R7PA01R1Xvm3pzCQ/zRagF9vVsGqBopBPlRTZStdipcIIkNKYOTMNKUvekUwHd99QdIKkKV
XwyVHyGgQDY0/AXuygPdinf2f8TAhwp91nIuqzPZdpAg2RLRcFQNwelLQANkSw2wezpZBPvn8bE/
nHADY3B/eiUCMY3UlFzFLadEZJUTFMEMGqhJEGAuIONTjw5V5ma2IDIQBekxhRgN+ykaxPiiogF0
KsiLzoqH6ssXyboLXuy18fWwAOvsai5E8/RTW3hOdlf6NozztVdX/9umMZ2lSMeKBAIBgZ730L54
w1p2xmPXrbcnaVRx9wvxUwD1Q+qndwAZMXic1a7MRY4kdVc37IrqVPa5FSuoVNhX4X8YkjAiVqGY
GGXddyF0yT1k4BntFdfoasfR9h331ro9+F7Jn14qwg8Xb+5sG1X7rY3bq7l1L0wU3tmjEkUbLoQd
q0yswnvreDkBCyNmyNwdkxfvw/cWUXYSR6DjWkSMqPkzkCbnfzCOhleAc8rWnXRgZbEj10NucJPz
T1hRBYLzWSsEqX8GnAtLFeDE5XrZjZiOzIlNtqKBSEfFZVzD/psKJx9/I+c/YIJo4ninci/LnQxe
696BOTWoIbsXTCx2ZuSzhliwHWM5UI6SlutOvlQKawSvPWqqAFbaruu+w9ZkidfK3WRDxVw0zg2Q
oA9SO/5aq2BIwWnctE+hQL6EaO8b3kTm+dfEwfvEikV0bPP4TbWNFTxnF4CNw8CmXgP8y/bsrh3t
BeLoJRCDoXyphisWja2RkerHl8rVk9SHEF/WHAGaE7MBixCWGKpZpqxAv1M3xstQ+SvftzFvskUZ
oKmt5FACPundv0yP7xjHI6IutvWP2yfhDmFeVEh/THVZDs1Hq990Q2eKA3L3o82KHBs8BsH9IJeC
ONW0Jmkjxm3iz1uzTuBsuXhuzFT7KEB7oPzE2DEhxMlt16wh5rCE3rE9cP2XQMAI+twb+wnBaWi2
U8IGV00dIMrG2D4uhlOCgt0bablbzP5UZf02m7P4/eGAjjSHbcP8JbKQXo8UodXHfB5J8r3C3e/o
5vW2Qw3PyEw5W5Y+a3i/qJjh2WHIwFkjNmcwHehusyyWQPYbDBgUgqKw+i/8svmzURk3N3Ncp4c1
ihNblSkIFGYParYPtuyJHn5xmygHj1b90yhv4znXFtGL95yucKHZ9i7Iblxd0xt43n3J8wm8DlOb
eilqP8V6xkbdze6h9NVDAryQqdfawEJxaTX2rt7EkFtcE9BWELyEMF6GkJBG9Fwl8w38FnpFtgMw
3S1ZkCqRkUuY05ZBWar6EZ1Setx+3379kAVsh3h2pUvLcsPd0lSG8+CVOdvk6JWHpj3e3I/MmS7L
tgVphWo+36Ywaansv8tgkHrSgqAsPAPgn3Z5++gO+Xy5B28jjp0nF7MuZUK9D80fbsNyJ8kR7Q3k
Wrdzouk1cnc0SISHE6FVVf2fFgOnvT4XkskTj+mElWpWil4ZnqiycG7I3StTEZMbXRbamOcYWgZk
qhBpRZfGGPQ04pwcLgqAjyZbgyD+XGf+FPr5cUGF+CiTWNtB9u1FUujIInEMe1aa0EBdJ7TWHOeN
SMTEhliSm6ZQBsHCm/qXXp1UChceUphOZa8s5CWbZTvDousV+3/0t4Ebk0vj4oAl9fie9xcMmm8I
2hWIaMC4Er8xXcq5v1ss2VxuWIov4v22DKbRzYJl1LEb1/ATSmhCA1TM1s4ZyMUNgtwHWCpwTtxe
aRMX5H8SRRyaur5xxhAXGfQmkh1fiYDLoanQHPWvNXXVYOfJ3jie8ySW0ucv0U1mUhnbqdcXhmIj
jBPIk6LvB7FqY4IGtiIrROZOrVPDoMkFvhit3RSt8aSe6jjK1IZ9DJC2YEIzzi1n/RwYQrsap/X+
aQyg7LURsbFx8RXKTTZxO3TpYV13TnxTVZbTNeKORPDtU3XtCJEJ4O3iuiIf5anBWqzVoqPb4Zqc
3HNWbHfqBngmCKpzh39LbwK6LXq2x4z3BsjEckRT9D+tWNCAZ1VI1kKpA54+fLQUcn6HA7qrMeRn
/GIsZWSZchxkjzg/BFfjuXmdZl65/OFS88YXTlSFEVxYV/NZaw3urzp+vI1hdznfVB3qVBzQXy76
qLSbAyvwHqf2QwIFB3HoDFk6dss3v0+pBcODHnm3eYTEOk7saDVGywRXqYKpr8C0uvSmOvM/Z8Iz
60Sch9NNDizCNmRhjXgNcFfmwHbeC9lAFHuNZEAOQizQoPLRc+YIukA0FRl7uV702PFCeOUiLKLG
SDyD20ScT8RTJnQmuPMQpEQ71xP+7wnOvLyX1GLLi79UXqjf7WuN32NKvxo/QRdmyNqAaJAVgO0H
Le3+wJ2kmQx79mY6czz5vtjiz73gmaxXoP9gQRSWybrnKAW3fNIMaA1IJiw/O0fxLOzo+RhE1dpf
hEdLnKojtaGpyjdROft42r9B2ThFm/qN3gDbsmWBTZKvzCuQHJXQ3/5RsAXc+DBwtBEKLCFJf5QB
ZdxmkyfbEt0hIv813olywqlRsDlctR5prmosjfmFN6HEqE55+UvsxmJevWj5VKR4uQkwW8YEYEWQ
jZe/FLOGIjvd7REtPhBcIBUPGEOdPYLiAGBbAiMS/9NPFd26WUHJjcHnafmA/UcvalPvakNZV8KS
VvpBvobGVOtIE6CvkfYh5GroBkyIQtEMbRrOgcDSOR+Xce0GX1v4ZKti/Yp7qTFBwikH7H/+yj6n
kD8iTvtNJNPIkXFpRetCUDRwtgNUCzN9TKZZ7rjKUut+yeAdVDkn0H0Pi4iBPuXdqcUulMZqmYaF
bAL/GP0BMOG+cLJCzzlkjOjQQ6+HF2SyOSn8ubz2KbjVJmNiZiIwzOaK6VlJoNUYxRpLW1GSYg0n
8rIcZOWH5/M8K6AAmzeBa6pHL9ThX1JGoWS73+5Yr43rm+CIv99UxR3J4NfYtsFQ+9H7z0TKoKOw
TY0QilfeJKRIhcOXn5xHnjWT0xF2vPjg4sWElW4sB8yq1D+QHNZjJYvS9ab9rwGA+zbWw4nhXEmm
g+3d4TQVwaUPtf3Oi8jFJVxaxQYVfGM3nnClfVguRx2j3btwz3Us66FmXVK2zAropWNfNN36kT4p
lnf2sNPLPOTcG4LcmZvZ9Jk8iO24G7BrZynOtXD4VxDucJs1mIoWfcjZWdqBk5ufNxxZ692bY8jQ
q7lKDlOFm8ty500T83ZFvAlVjI4s6wxciF6Ae2gI2CmIq6YVE+9CRtL6/bE9Q2epQOWuxXG4nsn/
9pr/7mjlcmJ3W9CfK26140czOR0/aiNYns3aKI0QpDZs9rLzs5+mz3j/ctRB+bzzpcfKOb1laiMX
+zDbZzuUjFEGNnDIXnu33aywlh0+netJAJhsbIRUhuNP9KmebjsVlQWTNZOM1oNfpbRb6td0Exhv
IxZQFo74i8aldUOcIZt4+SudnAU2KU1gZ4eXo0Z6Jevvax/cj6Ey5g1zRB6qVvld1i+sLSjBJr1G
fvnCp+KjBFJqN90IOf5qYBdfsBW592bUMRrPXas8pUVyHxg3fbRJC2Q81I0FD3NqtiSoeB8xv39z
hlHmx1rOwTcqJF8goGoMF3lNsWuED6qYu7k/CPQFg2+I4Y1HpdNcTezuSg+Own+QCyCt435TnmN6
WKJxbO9A9gtJGKwyV2+B2z+6nkn8i3lZk3X6biiYy7rh8B0sTvXSUvgYt/d68OKeU+o/pT8tU3V0
YAgoCesFLiHNi5zvzRcU8mcsVmw/53FwfJfWHnJX6JLx8q2UqVjZsOQAjj8ciJ8ZTeFKu90dr563
MEHPhprjHlsgo8/ELucktiGTMhkQZg4+8c7TMqLT2alAKFeqttkUyPSlNProf1GlUCB4wsAHHE1m
dGt9ELXTDLeiVgNS8IxLuV+Nt1zdBuKPA++FWXDK5yPS7Ycv+zZ7XKTTaU2A+daPpaK+/LtJZFO+
OEQose+/ml2lDRWV3QL9A/bYTF6LBWtDUqoxYh/YFat5MLlgfJpnIqoQKHrbrSFxhlLv6ETepxwz
U/FZjba7H3fNq3OBOUR79yx9oZ5DmMwToyCMxs8sxCCAIt2PrvqHs78cSL78e/NXKYDm7A9ARm2a
9IsDF+JVehXpBKbj27gopsqzVQ6eykBqI+pWtjYaohCS3jd0GRSCWxZ1qtJKu33Q8NAuRCY3oa71
CCDZQup9KJcAmTuohg2lDMvkoTrvuOikfG/uu5ESRH7GrtvEgF5LwaVhKiDWowHdpHE4T+bUhbyU
rF0+SkYFk0oQ5206gx9JGvLU3jnyNCkAvZwUpPS0DbM73pCb5fpKm8nE9mwY1K3423rlQ+lhnUBp
cv9/gPcFsNylDFcQlNEhC+krsKp6Wuzdd1TSAlSwnHhEelaj09tQG48fwHVW6iPgYLm5bXLGO1+M
Iu+C6djIArKgGhJ2ki3YM513R1YIkeuT2auGHJCYaYAZjbU15o6HfK+gYk1mdBIFiomyTSUXW4U7
F6YcG7IGhwoUv8XjHnG2GfQyyLp6paP1uhiffht1n6y1UXpuoxtIsOZ/xB8T590s7XIfU2NWIp8H
fTJV3BUR8MM1JWSWuEjJtnqkyem8pA640BJb2s/DiXbDnGRRMGvUo5dzBjHVXf49GkZF6DMfzPw6
oNitecuBWkXWB/3Yl571acEDHBpHpeO/TNhUle0O0ps7BptU4D2dU9oMe+ggqsLVjhyFwelPnKfx
LjPN/z8XpWt4fhsnJdmAWWMkLaUiC3Bg1Evi4w9A0SKZ8UaM6nllttNfR5jRjNYhZqcdh2Zco+/r
hUdXR3vHmUg1kPt2xHkreDSesdvrAzd8yb7R8ZhPERXaHEP4Nhd1j68FB6bH9MOC5NP3HK+jA7t8
cc/Y/gYBYFUHbrBFaTESQc9ahPNuYKFaXtOsqSbGkyaX0W/XxoEKJMPxYpni0zIRCwe4GAaWmDMG
Hia5qKFdttvbz/Ne7nD3bQcytJo6uOdvUDaFafu6MKI0jV/l87/EjMNXC1LsUloLIUvQjbdE4xJG
ExByVn/FcPQTaQvpbqJeGr4RMvObwfYYfG2h77WbDV0hKlAl7CMkvSTNgvZQ7B2ss6bnRfUSxprs
Y8xHWc5kWZr5YXf9gXUCuvGTwzgSZcmIHiGaDvKREXuKC3B4GBnzscSDtODjXHyHvIz2xXs+pgER
LcpzaccV0m/ZJyzFzR0Jw8hYbs/CoLa1WDCFuM9khW82zTdpFEpmFPImzAtJq7rdxJh1tGx9JiEd
yZuJcg7p8MCQt1qK7Td0j2Pefn/ebwiOK4OdwzVpJOvzDgY2+aZ59J3KVDs5DTptzX5EO/of8wOI
xoWp9koNZE5waoI3BajJn42T3pmXbh954ubapasicXAgkcmPdi5lAE+pGN9B3bPp0cUpnM/YAPem
va3m0PtjbvWbZyY0uVxWWYkePHnYOAACldwBSicq3C44+W838EzalLA4Z6dOpESuH7W4ZJBIOk0V
bidtSIdV9jPYNlWOxigzMw+/qsr00jyaorUMIkWS7LqC5C6htlaq3qrC4c3m7xwvjlVw9p7Z+y46
k2Cn9/BkFnPnlIgxATAAFZPjnKvVUTDB6eqgzMP3bv8Kma2OlgnZKZ+XZqtVboGv3S8GhpSmxgpp
d9ar0DWOw19gnr5f3XlRsh1awNSN2qKYaCfgEiKiU6LizmYi31WYHNCPqmCUU2gIWrl6OjscUp5Q
Gz64sadgyT6xFXPZXdU/xyBiHHrzHF5GATEQV+uOLVpK1UCvcBUh7APxzM99HfGZD8cP2/ud4rFe
jV1tYmr4EF02N3+j9iBcDG7+kUAZFoeNB8wrIsEjOKqaC6ZmJKRZdV4NKYrX6lbVHTvyJS1eSm4F
c8ttMpSlJhG8aidAkB0fE6iMEh0tBL+9kpTWs/d72ORFaho1uebc5RuLLoj7UzlzhMKk7ewVCCp3
ISHsD6nmSI3425+ds+fUE1iqZAExLlppXu5EYNv7Ojas++qHJ+ORGX4uNMu7zYb7hWck1evyWxrH
P4RhD2Wl89g+nbNBfhGy5+/qvKK9FlUCxtPUyRZGxAl41sZZDSRF0yqgDJfh3yMqQ41C61JPZiVz
+yUn3nabp3gkJvRamlhMT09xEAKb4vVgNTxNREixkMo5xTAMapBwITzHSPMek7YDIL1uuhrhm8+h
f0qdTc+hVz3ptNxx7oJ7Y4kAVcN1Av9pdQoVQdcu21D1po5pJ9uQWsmDzBx9vVloAg2uhZT5Ff0H
erM/YZL55NDMDmI7jkBFhowBzZxvCa3EfmzU/mAoy1AJYSoWG6McdxrapJgwB0IU7mXV2UT2yAvL
/n1FQHg7HO8Z0dLwzLnVy9X0FKX/l1entw3AJ8r1FdLtgpVeXsJ8yFv1SObEdRoPlNfzq7pPUa6H
vYkLxc3f0uTWZ11MlCJ15Ke1nHTlp24PEJ7eEtf9aH2bNrf3NQPch9ZKxvRpy+VuIAQAlRxdHDtB
iPv2xYISsQ0mEzCrFeIk8fxhfJYeiFruXpaKFKoU4nLcEicRBEH2Mt9iBwU46f9VO0TQ7UVHe5FH
Wb5sDbClpYtBfkrQQlJQ3O7SvyN3SlAI6aSTwOYy0wTvuLuV91P4Rd3tBI003tDjCHi0HlrBLC+q
rdJ6cUlahiUg+qQhJf03FjyHzYtwqsmdVrU8OcvI1PMReRWDIEb+9imO2X6NNtoz2kgUYBZAGhKs
KWaCAb7vjU4WIWnUApf5GuBJgRRiFQThecJ8NOIqOiMu3Lem2qG/SMf8ZTHz23a0RuJHjU+2tfcm
kFNDRamsnniPbzUxXma4mVtdkFOzW/fJINODsRHt1CTLO85QKP9KRRFxuBrxH3DUyH4hbl0wbYrQ
6I8QdY1WUgv5elfMGfNuTV/HXmwWh2bSQ+bOlyBIZOqL5VWZRnkmXdrInytZYvTubnf92oE+l+QY
zBmpYgTZ8uMGFSADcga9chLpYpf8Ey07i5S50ZBB6zG2efmBfjaSLjoF91Agxo31cfnVdqsqK+jO
rZWuwE6wwbew/SwQE3WgTgIE1b8k+fW7E0jdkkBF77KGvWw6ptG5ljlhcZ47sapFD9vAwWh7v6hJ
1UykK81byw1pLrUnY54Qz40bNIw10YXfdZRgMHYjmFlmxZcoq1TI3TXyMM41lotp36fS2HaoxySj
+qPJp0vPf0lpSTnhGAvTySco+1QfYrpO9V2iVtNUSgnalBMqlIM7y8aV53TJ8z8dCvCDsrRLnxaR
DDdVHTy2o9VzxZwotzuar0CRLh4i5ocTHUZXuWq8qWk52TuX5VNtnkeLYCjIhKitCDOveuYt5o3m
uTouTLqnqBKdoZ1cMDK3wcuuW/j1x55EwUhaH78FMne+i7pyfuyWR7JtRxJ6LpOTUXHnHH6z6gdo
NlsJl2N9PQvCXwOowVPFxl7w1razesj55THWRKS/yAzjWMUQJvr2WmVlgrF2H45ecj+8LcyEor2r
ABb1fOzvcfk9NuHWwda6YjR6UKLH/MtbJvtwxneM/rA5+G/H0JmmKuOsT1TEWZqvDn43UWb9cC4o
sqcqWgvoSJeoGd5eWp+WZ0llrvcJczkdiU+dIyEZewHA92D8YmlUav0flLp2DtCffvY/NUdJDmcn
JnrKhLIW4Vug/XCSbqK4vCR6befvnC0KxhG4W3VbMMmx8aiBaC7u/d5vyCkkHwTNdg+gbLOw8ymY
JHCgJKzKG1TczvL7pJyb+YfoK0dRNlU9PUa2+EJPhotwKKPAQBece2Bki2t1LKEqYpAHoJ6zHRSX
7PwSBSgNS8rDieAvqrTNmh8/iYEQ9sU6vVvFFOoPxjSk+xaOHTK3eg1blBxL5IOD5UXXCTaxEYHH
Bxj/geaUpaEwlS2nFi1Sm3l6WYPeAT0Gc/9Ck4AW5l0SOUuSeZVhWYJwv8m5hcQrrTJ7gUVC2I/5
A4EejgBTzKFMvt0X4b2P6zb7pDiT8Nc9NsJyiqvQG8/qvLYATco5NsQR598tF0P4t6Xkld0tm7Pa
46vSEa/PFjUxGnA1ZZK4WqM/DaARIz72eDQsTPWJ8qFy2MsW4CQhP/ZAYJYd3nyL+r6lT45BCWDY
bBkjrFN2Vr5cvMmfARVB+yyWzg49Mv5K9DgWMqHI/RDNTmIHXx5FnHBb79i59W81HZrlw27eeqEu
OSUMP6N5kQsqtI7SOYtROqu6sx5O/zk9nH6gxRO4kTSOc9lKU42b5QQHXlmR4TjpysIgzI5TniId
lnTrKjcAaYpHIJO1gOyby+/75UNOPmBhmtqVvu5uxSqtwdBvdU4c3mfuFGWJVgVtxJrc1zq4fMW9
NyzrCMkMORUq7tqIxg7WJi70wDTy7RIUxYv4flcCmj93JLHD0HcEZF3+m54XFDgKXYujdQ7jRoWr
s7A5EMyqyfzRsTZ6uWRlxpyOlbRBuW0exq2j3wPgTIc0KbowTSPlLuh2Czb1xhPQenweAPh6o6ny
GQKrLELJw2PesfE2TPl7IjyIAcFu0YUO5yAIU0E14W5kCCS+GCGQZiY9QC0WQxDaAFjtSHy+yU0T
FLyWYuEprdOQgajn9fFZGjsjUXjtW9e+EHwaJtXcuba7VPOi0MM+kySLJas7SwsOke05kE2B93zk
gAdG7cMHTa+arHVaiHBKXBucYAiGirVqPljg7CBdRI8eYKL7vkAnJQeZeIL3peCvrks9C02Nk0g0
DkZClDLRe9HVPrckURBSLEWAbsNAsbIxsJQBOq3h5mAgDWneWgrLc+0skAVVJvqyhMmPozctmmsN
2sRs6FT9hW221JEUjJ07DPCogktX9VD9IpAcRoSz/hWo9JQZ/R3Hx09Bnu3Ul5nMyjgr0MITsrwb
5T99ceYkr+Z/FEkS2aotV3RhnnUnq51HVB4AxjCb61fP8js7o2vPsD/xFYWER/nEmEOvwx82cEum
dX/2gMS0iwr2QwBWUetaba2F1SQ8csDjUw7TQw99yj/7dHJ3qLmmcAGUTPBifKArg6Ys3zEIbf+w
74k+go1T2DCZYHjAKJT+OMK3P2VHpLzeLxPPGWHkE+fK7Uj1QL5gbRVo/f25HCGcvREF7tK6kUTL
TEbrcswS8zcTOfO8nNiZEqwxBtgi4ObIS0jVOe0sEPAY/4c8uvncViWq3vtfbYYcKu9rVJtNs0WX
k1CS6LAG49vDuHoV49YRE1G/hEyGJ94r9QULqHiCUcTj9ceTZXw3MMCiHx2iTIxZjOPn9ffL1CE1
ZvN+/mTZEKy7xp5KYMcA9XuzS2oVnR+yazxNwdiTQ10BF7u3N/QDIXUcwapIlHVHYXcVD1nNA3tB
1s4ix9m90T1PaAptS9sOLW3ArELALEpS+B3cVuzUKDrWiy65vqz7vaLkhzLml7OEYpPIKM9PM7RD
xdz2kh6ibDV8M+zce5HuHk9rOmFcaOL34axvRBHXhMKUdzOie2eRACtTsqqSZ7J89eWJ685DHeAT
gZqlzqBDkCsnsQSqZ6xBcm1mtMuSbZzeooGYpJVmAuyNvK/oXXoj5u7G3zXnzLjqm2t/Nnb1rpQI
eEpR1mqG9fS0vdj2C57FapMK9TJF9VTBOK2btFdISciAJ6cE2mYLkVgaXdsWn25+E/cc+nOjja1A
5rXTdqTXU7z3Zl/eslMx95JWw29zXWe8n3kSEqn91V3aw12kdN8I0jv5N/8Gvl7PcrQ3StflwiWb
Jwf4QESiqRTvycKUEEI/3tPBKnizERJUu2B+XP/lJyEZeWcGWOrn7CvEGzIsGZ+cwrPj0V/Ymau5
ESXYQaRIDmI5v5rlkAXhXbAHbg4gSs8DEzpqxuibJGR85SGtK2TAePiHCHrfbyhWrZ2zQRN+K2ZV
mTudIFvuzGcuSTKbzDlw2ffsqljw0oEhAWjTlnVhXAmfTrtSOelKNpspABlXZakGmxxWc1c40ADT
0b97s2pggq7XVvpq213t5dD47dyI1qFcmhcVmOWKzA73VTuQVwiNqxGmVQQwj5cmtvsDCZF6v2d5
f3mvrm/K0AYGi/TIDib5E6eTCUop/+wo36CTIJJg1BR185d63UVCO+k4kdDLjrVhHrEPjLLnaVAS
zz8pnKlnI9rfcgpgRdb6LmvQGwSlbpGLeRFPQvODWLDjMaQnPto1eTW01dTomo2KH3NrIOw+mqIs
x8N8+b9uh53HoMM+VPE5M+f/fzmW4Q+sdzgHUae7vWoYpPVMXOaaK6JoJVgu4qAbUG0LWlYCN4cL
Fob4eOEPYGAbFMS6GT2PDnYUzSKx8/I6Xwt2VLZn8ACnskescoIyR2B+oaVs9bPe39bjzOTjRo9i
c81LRSaUZzPMqg/wP/xcoKLPy1qPZ2Lln9g4k5x04kGCJAzlpCxF+9u4ncFk1NrqJlEpT+BNrsuo
o1eBJthpWHFKkRgrXlFvvCBANz29VyRHhlbgKBnBxl/OFAPBFuZiLgtCq8y+/AXTLXq7xa2ntEAQ
ttEmPwrN4DEwFSFQSX22AevNP4BAaup/pCbBteMqSjjT32QXZTAJbjCGOK+w6JYyfmX1GLRtHTSM
OPvxOhByKr5mPValOLKdBm2G7tQVQYaZUv72OuzRTRCdXE2nVvtQmLMcBsVx8xTg4favakGwA/1A
eKU/x3sqVuDF85DkFpFZ/y5PmEjs6+9XixyeOaQYUkCOoDjh7AJPHO1e00qOdW+TQAVuhqwp/lrQ
G4dt+3bqrXGfIJu351cMF+8MUcvVA2B07nLv5Qv3fO/ymllxNBBM3wWOyxPPxrVPONb7U1D34i4u
+ZReIat9YjNCYHDRHKxPLyx2FGTDXpZPTnEkSJ0H9lUbS/OZ5O18URnmUJrmWLxF3I/F29QtHbUX
LmP8ykebWRAubabmBmd/P4TALj4PUyCkm4sjOPX0+ecM1DmdhlgSZhSdrsHAbAeaV6ZgIPYibYDh
DfU4/DRA+p30aNfq+bxrl6xfEFmIyGmhf2G2KOtMIeUNnTMa1EUu789ykN3eC7yZt+drSkJALKXt
/bYUXS9SmBdrQmWjnwKLX/wjMGgyKfnWltcyMirwd8EaigMd2ODukAId3Y1YdjX31cW4BhdTlsyM
92SsuwvzG9lrDalp7tAFpYqg6VKt6XPONTUh+P/qr4ayr9gnKttsSI5b++BNbqW/hwbtaa3ES+J9
LqNak7gqQKQv/CsErLMkKNW05eoaN4XQAyd+uxJ6Qkb8z5XVWvUNaU9EU9w2xr2jOimI02gJNiXR
T8V5Kifbq/XlWvZydi/lYBWgUehQUcqg/s//j5kIVPKxBm/YrLVQHdBUuF4ARFVLDhqI0pR1xmXX
kcPNmzzOWr0A1fSdlmglFU0DhISwgdGO48sO9exrdyJPEw5vUInVUK8gWufOBa93KjwZ9yrqZO9b
37NFeic5gqZu/Wddp5PEYb8pkPDvOiC43UGA430zCLyMxs1h1gw5jNB2nSZdy177ILQUp25ymBGX
mSa/hRhZyfPlv0+u7627DIJSodh8nZ9i1YehCcBMjRQKqCF13HvxGWOfJg9NgRu8I3WzuOfmPQcQ
B7/seucq43m1oWvtNFBivhec4htnlKXXw+SzeySnvbdoZGKsYgTj8D+RfOmrq0qak/KMapj4JOGI
iAQVb+zcRlFM3QbMBVh6koeL0IUNh2jn+rQ07GesNKhZZQBE+Xh5i3t5GHyz9/p3ARweuHeUZ5x/
ZsVDgGaJs9bbG2x00cZz73jXl3c9NORS/9VJBgjR700lTCi/U5aGcYof3e5QjEip/wTqC1rLl/+/
493e8NZygrK+jlyt4l3Wp/v1JcP6Nyrljmm++ObwOPpA+k+frwJvzhe8pCyG7u9fz3Qq7hmWrC+u
S3sKs4oRby/HTyom82c/cZ+eUckkt4unQ0mWdyE44Vc5F0cRp+OYBZ+sO8w4ibmlYMfzAjT1h9Lt
ZqVvmglV4JfoMI7SVOF3uWqSnCMJpKqd5Xlmoi+rrggDugkuRDbIvvKI4zHJSqFcmCohpMTM7SOB
ud7uAU+uFW6lEwg4hcZ3SYzP9xTAz0iBGo7WuAxR84lq+doRA5Wb2dVSmdtDpvL5qGdhYTQvDyO+
6cdvPSTRBFvEcHK2xAAm020YL2fJj2dCQ+d2gz01v5EXVjl/dR7XB77Sg8MZfDcRpC4mOdGt4EZp
2oYoXRdpd+eMEQW3P0RyGJEU/fp5hucexWewqKChll0DQ+FY19TMXgRPrvrYKtDBPr0kYhZ8oQ4K
FfWo0lN43ocMPs5SwBczYVz0S1sVFoviK1hQ43/gh5FOq+RwPo26dV5ewc41DFod+JlftyJrC3lW
4QngwNKOJnQ0uBA3/p7UDzhHNhInnftFGaoemw3VPBMXt1VPsVoLkxoJNfDzoQnoAbUnjvUYDUEO
h28heMdw7RkXjPsWA7/kmZKrUBRuux3vTpRzqjWRxEbF+QpMqzFRpLQyJlXqGkejb92dDjmT/NLZ
ynvwn891ecQT1sYSKttklwk9fdUix6VXIZU62kbf1/gGRFYjyj79jmWuCJP4LB6tIB6F1+rvcLo0
O5klGQ/pe+1SoOABXR839Ew/eWVeY7mb1UIR8+L6INvgW0TmbchGmAM+R4CR4jyUXRqxZzw+5QZX
Qu3q3YUx/HTt4JgcJCcsc6CjX/+XdSBKoAT5C5++xbhh9LlGfahiTFvhIWqed2WJgGkk3TzOrgqe
vsRmknPT4YZkgbXVGh5Fz6Bh8vMAv3U0OLVQuAmuf0zR5D58Z7Af/I7wS6+vW8J+I60upjvs7yHV
nYQTp6u8LBr/VK2soewMQbCvOEvJ5n/+l05L0x4Jjg5944djhfDbICl3lNIdG04OCVIoBn1ZCxoZ
vNvM1wZktkOCjgQekxU+jd+ezvBYMbalYiXlykOYQegHMD6tSmqYVegty01A+2lJby5E46oDzFEB
hwIrKfCDYQv+AutVuU0i34p1VxTa2utyjFEJ1fggE0v2/bUzv1u3D+Zf/9cGoXHPMzOA2PYlA6GU
LwL1ETMBnbJ/lfUuT9MR5/v0WAYtsuzHZS88sXmcrWTzzBY7bRvS9C6eLJ/ltlR4O/u4C8vPFOPB
AGDiOO8dDpFznp0Gky/9tdV5aj9sYIrw+9+h3TDQVf8opAOUlOrzK2ok34T9d7RdsAl/Q+ofMFIV
VNrqLjT7wsS31SkuEycA8e4wDMGhJTB8kOCyEABg9guAeuSmgW//YofDb8iCYFcGk7TUdDAs/Lk2
9RyqC/14gXOp2JXVZ6tNLB+rFxheFwU+waj3wZgt7+zqLc9E1BSzUp8SpqE0us4PWV1NjLYu/ljW
AbrhNxuJIXHsaCCHRvVLZSzzNJ54JpI+5/L+G/PnAKgHEtGqOy/IuaJXdMAz3WEdzO44nDiphxtf
sFJtfPxBucu+R1A+IQcXQ7KBit21PtL2DPrLUbh8o6u8OjoggVG27LKdOS7IcT62MbOcP5vxvuLI
Oh1CHMu8THU6o8S9X5ofLzUsIYubAkIU5jwz8tCePNJYZCocC631g1vW/mqhUtxjCZei8ObFbFdW
f0hnDReMdtlQWrLz/2aNy1Gip3IWIM5WLNE9az5dZR4cY+J3+G3+ypAXphtCfsgw7D8rbr6AjoVt
gq7jcHIFcIaBIC2fQ6m+VRpBwGXC615wiGLwbVung9Pz+8nruPgjhgf8zKCkCg477hK3sDZRGAGS
eK9+7BAAS0JzAGiRI8cmhBoQ5SivaqjgwK7qqkN33HtZWtSRiHglmY/UYdL1M+jf2kAmjyn7fN9w
489xt+Wzc4OWABFZ9YKiv9ChX9eYHgmN+OXvylw5A4Taxz8VZ6wOzoQI/L3AHqAKMrpUsHQaiGkM
uCTxCfDJ5yb8uoG2VjAAI89o/N3lvt47hQDdb7RkFu+qnUG5flkc1srT2oVu6czrctFMsvfXpedT
WugertEue8DVeQT97Cg2pL08pwJuyWJWodS+2OyZQhBYhZ6KpOzAVnCjG1b1YsbsLLEhUXtcbXFG
Gbpns4k+WXnbj8K9G9ooVpCpcpPrsGedEi1NJtFLJgko4xW48raiihAZa7DyxxA444r6jynLf1mb
6P/5rqIoCQuqTp6K3RJTSoq54Oy8ASAqTiOtwu56P+Wz9uQCvTPrmM/55zL3OWbNaUYwi33aks/S
ap/7gbmZ10FaAptioISzw03wVte0yw7Dbco07U9006vPSHYom3Uj8Rl5iVGhSGkkvHE79WTNuJVt
twvYnLl66D1hQBvOg1iWykDpYbWjR6fYBw+F++a4YuDVYCvE1oUJil9KZYqeWyt0UqbXf5fg41kI
DxhQZzXm1uNcjndI1U9bUm7+aOKeIw4OGZXeKB5I/ZbQ/CE04UeOhtgs0+7KL5isVDPLKHIoNN7B
Tuo33IqiJRUQQw0ztqv+yLRTYp9wvS1uGwk9gGiTirmaIcVmm9WqaQc3nx3YdQVG1VubJzUvO2Yh
ppfaAFqaIPgUjlPcwupSX9Z2pgb2My0MMEzVKKx3ARG8UbUB1pjM0iuAfvTiJXhNSzK11WuLYdV/
ycO3lV0bOR2EQwDU8NhZJ08HzuUcT3bBhL06hIsfm64SS8AKCz2lRKRgqLgc/wgaJtCOlpnAg86f
Vog5MmiSYzpo5/uRy/fIv1mW2b7Lf39RJcz/CppC8UNYqKVwjAX/qlELqm4DhtAKQKRZe6nG332G
xqvypdVBQy0UDYCiQCvmML+zXIuRsebzmxVZd/Ca0oUh9rwGTbv3MEpXmOMZV5ct//p6mWiKGAuv
vDwKt45mIFLut8qrabMQKrkcFoMVx8umZDyLUGpRhdhb9WXWIUmjBbgj0rio+LEj1BW/nTNkQ/MN
sGoX4gT5PCcd+FTWqNgGpqx3QxcAq53JRU0PtM7FG+04X7P8/9j5Y7TWzSjCSri4hUReLlPwxAqd
RdTEPcAW0A7S7KfMWpXQ8gPj45PiwWwAtx6yDaxQfE3DTH6r2fIVyqthrKR0iTSRxySEbX+WlpAM
yrWrvFgE+J6RnywJB+8A+WSRL+s9ZXIQsQUVrwHf5CdXqwBvqfp2Ib/CMnoc0Qyd/PGOL0iiJh/u
Ll74qTjh0bloTxB+VHblALkWEP3TP9ZIhYd1VMTJoyUDxF91meW1G0DEWUpGiO2tGuVZjuxTi7OM
SebLcZT4BZwRDyGVdKimOWrwRe6UD9B/MrXdncbBoNR6OgIjSoYWqhDNjZE6Ouzxt/CPxWZZhOoc
BLucCZp2BGjjBwyZNHk+5cMGEAA1jc7i63msEogZFbEA53ShRMJin28Hb5bWuxW1LuTRJDHmzh3d
XCrSXb5HoIdNorE1/BWJpv5oDhmsMYO+ecIxk5RSvd+N72Jdb0dl9AKWAygeT4afckZMkeu5HTsQ
JuMfRw3c/qI7JvljNMmEYvsTW3fTi2wuP/zzbmNi6Mzsl/vPwZagMz2rvRIcPvZixunxPV/Rg0Lk
CBk7YPW6JyxFyGsLF++y/nkpQbl+IdJ4KT2yWmac3nCR9iDHhgXHSWDFNIsFkPMsdDZ3DRrm7fYi
FettRhLW6yZB3HfQdirAgniJdgGIuGyP4cKTp4C5yoaWyAQ8aGG2tdEn2WSF/3qy9oprXEPTcf9m
shL9d+dxF3ImWzChyMlcKhKH1nVyRNP/TDs64iXkrieUP8CinQK28YbghGTvXbZV7lsMILRY+ETJ
F+x79dxbEFM0KNT+zvX/CFRg0i5vjgz4YiZxWAnlA8rqMI8WGu7pI19a4g5ndi/gUdfPA+LjN51c
2C057JZ9834zXAem7yD3B+ffJilmklSB/DlHbil13uzgboQVVaCpS0vhOt1g41EWLIP7+CA+eBjV
pUVRVQ2WJsWmhUk4+gIQTebyG+IfS72kFNilejfXKp+kauCfCVQCvDQIt1Vcg80kRA871hxb/qfb
6aUsx8XgCCbBjbMRUsn8083/h5+CqoVUK4ICH3mwXkAN6FwI08Prkt04W6f+vyduX1M/ZDgdodEo
ijagM4tqfxJE7BEKQjassEUYOqqncAmQZKMsAkwYI00GcRQ+M3qFFsnVUW4MV3g8E5vpD6E0sdW2
vgKaYhcRAseU79FRDo3psdjIaZ4IoLz8eQgrjSWOz2aueoI0jhq193DD/3CERV//J208QjaGFXFj
Uj8i1HHa+arS3UzffAsMGY0FBqb7fU0Z0x9zCeEsYmfSC2mIrukuredTQNYwOSy8AFNta9dp70wD
bTW1eueEOyjkauHg+AwfUX08LW/qBJ7X7rAwDcEZcB0hUIM86uryRsOTKR6C+o5qDVL/yd0W+LL8
DAT0tnLTdMHGZLeSeNtI7rZWXnt9/zJiFCz+CuLpZtVaJ5lRkd7VMgAAKsgMe24yCejmfduucnJu
fI1aewdSFM4ufvk+5QcMCX8md704YvCVYIp8hIjAJPA1WvElpb9J+nA9HPkquU8oNiazjAZued91
RbkCFDiiBvB7CFh6X8eoAJpLEKZImPGn9/LxN4R7wAzSq/5Mz+GCParRHCmu3TFjzb+psG9RvGZp
WwSRW2lnX1YbsHEEmm7Ih7rMN7weMlVnNETJFCUEnpYXPuhMCgjkrjoJ/1xw+uaw7ZOEfkDDnK1/
6XPuAxuNKsdsy3yEDpzk2zK2PkUN9yW8C5BAI1oD/G49TBkr2eV4Rfkv40OTnS3FdzXLbkn4q3sK
7xjswHpZ6Xu9KTFbJ47PIRq+DiLXVdLtK2ofdOzj8PJVqJibnR25TN9i0ityQyBjYPiIV14H9mdK
RolwvY++oTvwvpH0Ej2XNVakIvn91s8stgvpSoaTQzLaVlK/AVZm1t14VhFH7IJ8T4fdYtndJ3fZ
BnnKWLCFofi89aCAIW0rNF0K8pcVMXNk8/UMcMVu4gGI+VhiybBauQ0VUND5AVb5R1sT89ZId0RM
ZYUkyLTOpY0sGjnCtMsYfjXunejC1HjCazFd+LQgKw5z328wehj+Yp3knKHwvry1754ZZjJfEQbF
p0VYrgCP2cPHtcT4/cTUstAIxWCgsH2FdeOwsf7ibMlIVTW8Iw9/Vc7Vo+4t3OYxoOxkieNzSvU5
RqswFu9f3lOEvzCe9WGCHt9BwsdySD/ebWX825jqNYGzdCe8sYTgVND/T1rka8tX2PavdoZTfNIp
xhhmve0j4b3M+xWf6gawgFbTcypyfa+wWeKK/Ps7ZBfGpDS7oQjfm95ue5rbHKjn/VK25+nyLaEX
vUV3+Uvpxbxoy850Tvo9wme4Y39C5xhVCfOciCKI8gXN6AVzNoy+HwDRSQqGNW10VjxZYjrmjUCA
MI8ntwU/FpVFl+LbRnQzo5rDZVFARJXlDeTH1tjpwSTgD6t2SPC56cOLDvqNWEHzD10R+QEUrF/l
5xXmp+/M1Iw1wVax2DvO5+RBpckFVMkrRCSDlNqFsK6Y8MIDkihPs9/j6B1KYc76sZ0WRALQGk2A
3Le5qY8JiXt3sN+zaBcI8C0sPPFZW8r7eq7Px4ooLs2GWYACHPNy67VSfrwh50I7PyM/yFZyV4HM
6Q6ATQihgjgEC7rXQvvY2c5ziXeLsa3ueDCx/lUjgfAZBA/WZ4Hx+jw3riZzFtEnltDZEJX/ye+s
N1Wq1rfnlm1jrwgT5BqZsuG/d8ubtK5oLLZG5mh4TQUVUQyL3mR/SRbTEr9WWucrClpHXvl056L1
9CoR030mBvaY/c1/pipTygWzOWTWYlnJJUUQOzC0mp2PlAUdai1Q65Bq30CkEakm5kCfJdXKbM5b
RHpAIWMxZ04N2xry9llT9RqKwsGId8spS02XE4BrB3l8dd3kKpqkc2N8EIGNsuNAZfClOroT8o+w
jAvEOVlz08LNydGX0xHCpBQ04bnGbknA9xijwpzI/IJC69BMnVsAzTQoeHaRZpt3+8+vWahvgdT8
zskjkJrkWf1ISbsv9mZf5d1K12XMgaOt+CbYBaQixjJZ2ktCTsFZtosTt6hiFHxSqFBsEmwq0jtM
EEVfdus2mwp8XHuhkOfPT8vjTUhT/CfrQDEFWAk15WZwRWz5OH/qOGKwlho4ZF/AHjXWpTysHNCF
MJpc/xC7o3611NtKSXsTQGv8Jq/HO9a3YeWbYHXJ8vipKQaeC8xaFKKrqA77vE25xhd8TIiv8YJa
Jk3jSxXl8Ie031ptgqMIQXue1XhQrAvQG/xaZ4rzPJSyutpkckHeyUCZzTyBK2OUPJ+IU1nc44tr
SIhX8fsYiWHLW3/Xctdlj3gwSSVqjbEUo4JcDWO76X+7idb037AJ9O8bFTffLwzWAR0xUeDrKQ4+
vxCuj1TVgwPzLa591h24j0+KOVppqEGqfgkhJUAgHogpPTejkiahUsjiIzDn/zLJsVH2UkPFv9Vn
f5tQaI66dL5VRLVs/G+9TM/n9nbYZNM4iAoHE6AM67Tp1wQCjDDjeV4jd84vQ4Gu4UNVEwCphCVS
msRB7uVVBCv0VBH485USssEidpE+iX1Pz3IzSZJ/CKQXuhYEpb9pD/hQ9k/fGL2Gzsn3Ozzd8pdh
wxWkZmRbcjvl8fEAFgIRGJdEfazaXL3LyVHUodyCbHrDzXfm7VU4sMXa7xJk8BLfMT5a88rUCG1P
V+pocC+xKWbl5+nOCWuw5GkDhGE/OB9v6VJE0/XBsvPG/yROi2dz55SepCHsiP0xXygd4Nu1XXlZ
Lh7ZIp3wKZAfuOXxLOG1XciOfGruUAUO/q+yGNsDPBJtZ0HkGq1tMor52ODA2E8BjnbKoYXiMZmY
yOcS+XJgkLtnU9wkfve8AhFoEi0cSjPfpR0oPccbsjLFT6BZJzWjNdTnA6ZUC6sNsz4mqAM+6EER
lJaHrVxdgRrXNV9mGB9YalUoLTd3Q4/M5jaLN67/K2HQJwxMr4elE+rMf62Rx1l83SctB6u68ZMr
Bn5etZ8p8Bh83c8GrwxtfyN68d01lZ49htUKjDsg3lMnZhk3W6KRv5MMYTkMi3uGHUGUgl2VhPsy
hxkp1o/CZw4OxjfvAiHSHOwKUgN2tLsVleE/4sAtY/5/ABRpqFFajdmbdrQeHKCwXlDeA32eawZ3
vAjzlGITWYvTj8WLeaP+H3+4F4k/awhWpABstvOO3Nr/s4/h94wkNXqwA1zxI5pMwejATWHkN80S
1BZ25HOG9A5sA58boncmoC8oZqNqpsFIq9CTEA9sTW9JGDxvr2+7f4u0Oc+5cnBOq1U+wf4nEIsV
ZqjTCIwQYZXvrPniCm06oYxGfItR377fcye7fiLH1pBKWbkouMcBEqDmjaa3hPjXBQDjAiNCqoZW
hJHZMW32fqr0ixZ8xBaJyKkPpsLnKqNj2GbzJ2nY1A9OamSx5LVMtz4pxgIj2+5tpaM5WuyMksR8
VyplbWO0y6MY6Ua7Zyt+D9miSUrFz8TfZ69sHWWIpbrHq4aupLJU3iKlr8KJ5by3gqWUaeMR8iLT
ZOdhIM3iF81y815ZfqbpRqt8uDbBeR3rVTD8x38O7oX1C1Xw7YN//N0ObiviKkB0NvG2V9ftt0CW
PfS9nBkbmLkhMOhm6URLpbWcROrz8X1313v3dVKszXbxTC4hGClmTFaVHq1xkoXozwR33Df8vCF7
eWW/lgkIhKsuGuAOKGuMOp4gxzSzlZfQH3cYEJRZlmyuYXpHssu9rKXuVPKwwf/gNzBwKxA9gs8K
54Friv6qKhkdTj0ohWlujXIDFgnOVQDIoIFkLJ1wMH/Ub64ZA7aeiS8KBtzCMhCWcPuP60Ud1u+y
hv6gLiQg3xEiJxtTc+0GqXVUoCfmmbMKiDW7hvCGZ6qw5kHHHQHU4Xwa2kIauNlnfPUDuIUpEgFq
vNKfYLSSVJYZboRjafGgSJcoZi9gKLNO/x2yFjKJMFscVqlG5vUy70I29WhcucGoasr1k+9aiQ/l
Xx/xcnQY9TZy/ATohbEBmiuSXk9sd8SMvf1koVFQbu6UAHKLx3axIhRJ0jyQG01pPRct26XQzw1X
4UrD0nZDJBUQqFFBAkoGc80gcMuWBDv8o2sPnFDoIhb6NhPjuEw9mPnUW0J97DYmtWzl4MzCfHg4
6WACc4pbFO9Gfx6B7Qap1kwAkjzg9kHc8qAO3duT4DOFLutOz13aOu0jnF29UdD0+d8hCVlEC+w9
/oke361tS6xD10NawdlMc7khB3kwU0T1ERbY27dj6VCoYS2lIR4OvnrjZsAqn/WO1T14Cjvy+uMd
N8w7AmiYuAP5fxzkpoNkz8AKgWDGI/O3Df/l8UEe0HPgkwvB7qdgefUBnPxT2B8GJmzwoxvlC/X2
6Z9SW5RqeniS+AaNAHfPFr3w/Em2remC8TLKP7t7K9ooHPtkWi82WvpJOezUKXyrDMjoqRI6NqK2
todwIx8rJ+3Rtl4a/LBKIaQ4mrHPV7lsyos7W2uoOGPWUOV4VyB6wtG40hll2kNbZqhs+ugmN6pR
7F9kxUYzpI28thg9kjm9CYi1pSTA9Bz1SmpCzGZqwUe95oj3uEx6iECLQFP+6+zyJ5e77AEvmhEv
fCJ7HJmpPuV8IO5/P+6SDm8eM0ygCEsePOB2E6mmTwuZe+FBAOkv222xkzrljVaedUn/TkoNhBue
+flSGo1z/6g3Lof7F0Sv62rugx9dslhuQkksZjRtzFLfFcj6/sykdYjuW38v31yj23l1P0o99Q4i
vNF4u+yGFuoV7bg6tevouk6HeJxPit3256Xtiq6O4mCpl8lpQb6xqL9aecNdhBeUdvN+6HwgPGBc
WNsV0i87NK2TDfQpFGl/SWa2PJZNSwE2NuHoNEWKP2XW6gza/KHq/n9LcZYPG/B2PIG/tdIqc9Fd
/muayyl/BGHN8382pRPajQcKMoEMc0K+ERxs0LpsfnxGnYpotZw+PMFKe6Agqv0B/0he/HWGi3bh
FmaRhbo1Q9kVfYRsZgcSdnti1lJXQhmgNbQV9aXb3ZyAVu0+0ZJ2yo0Bg8WWahZrafOXQ1CWUizY
zwa+rih7ewUrDrH0TGwZiilhFRJ9MgpaBlb1EqvM9iP/bXW4Stadu7Rl0I4jXYeg8/wf6omFcanM
0rlzYx2R6HvcoCPU2QAgYZsrKnmej+iyRQzLk0L1qbJjVpvvuqv29ddAP2IspCEh1npnNUse893y
62C63WkF1oZjdmAzwWm9mPaKYp5DQb5cVonBtkxbGtaJ3iwhx5SJAljjNPjhp9zM7uV1v35a5UN+
hAEeKzNRtiN6TPsuqEikX0e04YgwWL2MR/fBLrL5QHPI6MrAHMzVA2wGHKnXJpu+fIAnHhHynYHj
jwTXPqJBgqKKnKaJ02kehq6zAJj8GWO3aNB8OLlAtNMPbyZznqXciWf1YtMPRrymmIKaPbKg4peA
bOXNRbv7fV2aFW6/KHnsY3boEfnl519cudViHfVuK3oEOWpOaJPOlHldJ8uXZ2lQzC74rP+qKFea
x/d66aQaLbqitL42OxXzjyEGxW325Xx3PVHcu2xdDiypYhfuExsJdqQfnaFVJM16i4G/yt70JAW5
DuNAG8EyIQPvnd7v5ho5rYTGUmn4ZCgUooDvVi5YN3AwLY0+f5+PMjX+Wn3tGr/Za6IYJ3z7SnIv
YODWT5jc8jxUkYyN2r/7NOe3e9RqR3DxMvFJejedMgrp4Gn03aOwL+NN5w2d/W+tjrpsg6PhomU4
qmLInAk8RiBLPbc34xs8ipZK0/NSd6tP9ybFWTJmSj5F9kZdFd1qqp2bE7ukXusWBqb7AuXFCkvM
W4p+K1Pu73NOo8FUumYwYssHGylLKs2or4sv1+Zqk7bgLMHZeBmVwT+kNN63oLbBdY6b2hNvJF1n
Zk8OfUiVVakXH4lmtVITH6tKBZ6gRPofJSDoY1WZRjUiiQ+uKEnaXbWfbIzZOdvTPSUVG95jQmx4
8G3llRT0+dnAMD1YEx4Z7bLuPlqOy/8y0FWDAlyp3FkcG2ntyVuB1L7m9QktiAyMF8Y6YFAOzlGO
EYMDg6Nabh61zEbM+UENUKASUPHkcdf/rXCHRpvMIEbTUNzBt+nYmD4TDxpSPcnwfeUsvg154Lnb
jGk6FLr9C9O/nzIOXPWHkLs13M9/sPXfZDn4hDzJvZjtiy+feRlacpos2qN2z2yo8v+raOGb6QPt
qhQi5wMQGBmUVyfG7kTZwxEBi/EnvRlDmYcferVAkRNcjQGNA9UUFEq8Fkap8QO0TNaT+rQqeXGB
LVmgs3y2l8Eh9Iqs1vDXsDo119FdlNop8/22yHHWOF5nFH4ZW+1jdPh+Jx7wpmgb+/YpL85Nz3WC
GHNSbrO6Cp0faB64eZPEBg0CfYwBpRViA7n+uQimDC3dNc+shD4kgK9LuCJmALNkncawSAKybFyS
Wh6+kRLafmoP07xjqedBYUOxHgxQVKyANObOZH65/2Yu/TNSkJNkQv1wa4qei28XHVLW0RTzzdtt
vzmPKkua73Ak1fLoM2bhihOkzT7U0hKR1YbO1m/ckEuu3naUEXlYnjhCLE2NkqbEHD4Kdb0b1Y7H
ZIUUnvxAt44WvVSVsYDTU9XVFwmp5e6CmdznsBjN8LZ1THXZ7MWP6xR4UnQh+XCkWpLIHfvqDhT/
YFDhlj9+/1E+eP2vfWrpXV3a78MM5PpeVanz9fHBaG0WDcVS1Lbw6t93GI40qjl/WTrZNzLkmFgR
/2BSXyyE1CgGIjrkFrsCDoizK4x2rz30fLVYi9NdTjobzlvIU/OmFanhl3ZU/6UkUpmSst9b0QTk
9FPB//YbxAdzJjSO06XoCo26vs3CjGZ7RpwOll7IUYAOt/dWfEvPOig6wrZTFIlkSGej4tXg+mnY
hDqfcMBFHvW+3JsdSNfVUjMPZHqvzoC5687M3BE0z3ROwiUD8fF+w2DxRRKp3ZJ6/Llk84hLLEnd
FAdlpmGeEBqIquB9KBbbIQCfcc/rTlR9EVpw95PZ3IiYfBLuJu39hNhIlNBXfHM2ArnwPfpzKoIg
2x6AmCg1EkJ2MIgV5Hqy8BhwcNLkufgXRMvFPPVII77lTnKFxrPgJ6vOQ4Gp3ne3z8obpFzZOVM6
VZIcuZnk5WBY6EQQpyLDMi0QboYU8WJzdEZjO28IdFJwbByp66izy5YT9xgVxeTqwjp9i5KrdRBR
CxIAkzHdRb5dwkQwd+tCBukiBWhOQDM8eGqRLHeOObclGURiGPJdvFGIu3c3WbqR88O1GAAi+9Ga
5mAGnq7uXeviYC+ylscNzweJAyjS30l3wN6yXW+8s7mdJvfwujVVZ2Q16d5XKBK+JHRHvUowmkj9
nMe7GfnBtnwBJBhqSQYZdqCo54w3L6QMQukl+RA76LluUhVOuubnEdZOViOFE9jkdkG6G0eNtj2a
UQzFFOFGJPWwSFZnzMIm68gkzOGurg2SDJbqs9IlpdvAqmchWHhySTh0zhXSYAPeqx6iSMrRUVw9
/ClNtyXQJvtZoNXaDzC/gKGnzEE/tObq0XDYdqYR6DQ12rQNPhF8jIpi5vhyHFXKYSf53QNg1xov
zObyjG4JKZjWAVgS+AxO42tOMyx5rsGquEU4LfE7Tq7ojqzHBO5Vq/oMQW7MAxfQSZ4r17ujvG85
bLE0hKv9XlZs0yzSykaKmIRYTpKphLpH4Lke/NnFH0ScqMU+jnfbkIaP00yyHOoaDQwhIgw/EbG9
pv/xjZlSvupCkrmtwDVcKEK97PoX0DVLOLwaOqODaS1RQjgTqkLXq7qFtAkRm+4zJZHvwRD/lAVW
BbOB/GN5qG8v50OILwq4rjTlgjh5etDsvaY1IMZk4UKXQB2HFUvBsYwDLGdw6fvXAmwQb7F968f1
SxjWse9gt2R1nrBMvWS/jGZaSbrC4HnVrRupWq5jCjWV35zwgm13jm4e1bFpfriUuWUxoS0rSR5E
oHKdv3/VQKewV/z3nDDDEfrbp/0qzDMGp7ihB8RJZRGeIblJAEH6/Fup4xJ3+8O5GZMAJ3S//tFZ
Uf2Qlo33eFOP6vo7axTXKfCp30aUuhpa17obigc93d9pwDxPKcw9CjIht3BdrFBIWshI7mPZ4DwN
37TSyqqXeTElfNoaw15LlQzVW1hi7TQEASHGWO5qmWnLGiamw1Vm07zeE+PWbZP4m3DWSTCy0vS5
XSKyeFqkcYj26NOfLUc4O34cx2qLic+6XTKlMRZKSaLMpT1RG8Nv8OgsVwc5PpVV8LabzdXtfYMx
4IOSWtmhLOkezwn80twguDp8eO0Uv0qi4q6mQjue6k37SRHbhtuVACxCW8kxo9H28PwVsWwh4fAe
+Y3lXf2SS1catBfkrJuhNvRxaMVS36AW9PZvVwxMuHWc8wJ2ttEdbJPCCS4jtfSLd9MnqUcGQeJX
0mmZsqsMblCyQO5Vfjs5/Nbmwkg9Z9a6FNLTdNlvheJrSaKMnTWVcflke28pUVCxheCW4KoHMFlW
mU00EQ8v6JH/YswcWSCEG7zNWvpHV7nTb8K8SWn5NJ1I+Hs5BJup3ry53z/o2fs8uMFsAMI9flXk
RINXLc4q4Yk40R0vxEErlNpt4m8bco6ZmoetTzymfFqkysDNxK3yi1HkfEcaOkLt/2kgK91Ysn9c
gGrOAAJhdsStkva1OQtUYJfjlabrqNm6k6QdC7k0y7Id8D0lY7IzPVDprLnOsfx694Y7eZjEfmVD
gVYEi65QqBRGGHO//ts1xr9dqjDzAeF0oD14yx60mSTMhJRGe/Z/sQtk1rYoXIkyjq2FY3E4Yh8v
nAI79y6F7PNCTXTogeX/BEBMxS3aaqiE1SCQ6zCAy9Xfe7UZoeaDf5iIFAhVQw6QYdJi4cl+4qNz
8gNrgi1THFg8UhfTrts5Y6cn86C95c/pnSSjlmbmi5hSvZsxFf+/KucjHy8NWPxf95LKMee0Roq5
x54rt0cCTBj2Kl3CII4xIQxGvrWiudODvqoccvSLoiu8EuNOufxmnjYCagyO8xtjnFD3b11x9/Eu
j2fB1Jj4JEWU8O2brIBuW5D71s+Lm5ihMvRG3sRlmlwLXf3/SOZVxTdliHdKK4y9V0vXz2XX6L9x
oegaI5r4RBO/LzatQBuaXKA8+bMqENDs1xTUYB7Q9mipkwviRF0847ag16Vvm13TBQGpnfpWYOH4
2G2q+j25EmzAbZ1t7GwkMM6+yztVnNM5RmuUlXcqme2c8FW+hAdKhNbubyL5mxQlW4A5XDQKHQgi
EuMD26P5Dr1+XH0YjyNYW/D+wdRA+yndM1jezuqqdIiRjZbVbwwkfWTy/+s0NmBsACAn5H7buvka
LU37/NgZ2vbMTtxIeIz+duXSZG0X4sozqT+ubg1gPKuV6+FgyYrIdVzGuH6slqePr9jjCe7vFXya
3GiyhV6x3Lg9fOoLwTTNUpTHDnJ+mUtdfSUeGw+E33pXA07dRaSbkTcHYjT2jzwZBLpRbdt9IsIh
7dh97FJAec7m0MusyxB5R2ORvAoVEuW+ISq9GM6+DabQpRGJRj8v7VS5bDfIh8JRiuiXUTTiOHfl
oZ4M7ID1GSWVcusEHPW1NSOL6oRANM+AxG75RW0oTgytbFzNIxYNtlEVFyXFi25QuQTVffPZudiv
j9jXjZCxYk2cuSWAbQrrBiS1OjelWFb3uDRb76/FTaaMPiFqmaapjaanCUFOw3ovdyz41jFdmtmU
6k0NxBCqF5X2BGhp96i6kkJMcnG9ELdOA/0E6KYXPVERN4zmXOTdlZ1ozCRuDhi4NADe4JFIDi87
I0zQpl76Y/nTehVCKbGBNXbkDpTNzzaqh7IydaJZ7XAOHfUv+7ug7Rh9efpnP4seJ/5lEj1Bq3QT
yVg3w0JMasPCBCzHdw5hyraxY1No7zBPh00g1+ep+XVV+YZuSQ3ww3b0QAwIyva26bblY6P8ClUs
3J0Bt/k0qJ+/Nb5gebl2PtJarA6yIwp85K3nLrBRedtDO9OLHZpg1DRdJDa2wPEYNigL+9/Rxdh6
ts0m0uzYSCChdf33gMU1tChnT7yZH1BmUBHRtrpsVUpK65fwbFfvU6F2Pb0FpGjCqE7n3Lxc44V7
l//rJmzwbJyJhZLjuxLEYo6Bze3dWa8U9mESiBi7LgIWgRfeHdjOc1t1CPNlosfHLHXU/Fv67sN9
DFDQ55KXRdP/mHWURy8VmWuZCS9rIHzLGrXUUuiWEDlL9RB+NfHsztbZMcVqn/TRP1h9gOj6aFj/
Z4Nor4wH7QqUGb6gfqBV8/zLCMCvkr4Bzg/m0Vhi5sQv7GzxQAhrt/PwAX/ZeO4oDBv3BSOxr1P2
53oNNw+7CO7nXt7tnon7lcv026XLhNhjiYL7hAAjRFWDWOJ96ZV0rGz2FCWbOBS4FtDHrPQO9R4n
/PS1gZ951PtnlMF9jOjC+dZxqefZ2EBb0aoNLaODCMTet2I5D0w6Za5fYrzVmlpi+G1DQKunamoB
Yxmbi/I8Z7Cc8R9mtywsamNfhwa25ZHib5YztvPZM7xbo/N+GuNF8tvBVDN7xvtrxltZNzIHxLmo
fddtBC50z581Nsc1TLWwd42awAsu+74WhBTgytlAF1wdIBr97eIczQPot95iRneG1h3hKE+s1f/Q
NWpdWZbaUy4NBMu/UBRYhM6ivgrXgtYKX1vS6fi1r36+JwQ5GBgsGIpcZSUUApqPzFWbnVSZZqu2
UB0WBEKtugIpDCwZLDR7N9ld/XBVYUJagRbl2EhQwwEohNuIOfg9+OpfZYRFo6/v1PG+zRQoChV0
zX0LShJOyVEz0YlVwGQs3kLrUDlm1Vj3h7JXa8ywVaZuAmYY69y4df5Z7jSxVBBi6+emT+G54EH7
A5Qd27H1RSk0dOqCD0PtlHqjRopHcOesUcb7hJVgsu4yp3VpwxM+6jRPu9LsusOszJWGm+CmQqXA
ofXdo9RRGl+Rabsv4NtMVdf0VaTCCKUHKhlnaSTLb0DPDRo4cq7wEtiiqh3B2HfUOqzDH+dociX8
cfRnKXS7tpQcWlxL704fEHKIshbvYhI7CneafV+tkJZcUy5v+qc5hG9AKnGwfDUunr+T8e+c8yJk
8wvdHGzpAXldHnvhfX1Q6zD13Tsl32Gs2PY3oHbQ/o3UHHNUWSFQpWZ8q0Igt/wZgrvdz+iYeGDx
m9dpV6nvQlm8LtPraHN6UA/wGdxBpj+Q3HxtZqEsvtNSPiVlJVyZs/KWwid90ro0RPfxItp1ujoV
cCYT8joKOfCmRVggjt8GrmhC+YS7OGxSN4VSIjalaQpgfHM1x/0JLocQdEG5YzCX9AnSp4Ulk//N
SPqRoPsewDQXc1tb+QvSgexOgJ/isROViXaTEaJzBmWvWjvupA4u7XNRg/F3tT9WKVHQI+qjcy3J
Nz6rrCUgndo0fs5HC7L2dJxYF4bM2Ylxx9QQFhvYck1eU/dlQV4SRQlOTw03yk8j+Q+HAFNRcjnY
hn5OTlsEsyuhFplkz4fl/odrLArn7VP+YQeLIJ82w4kDjTZYDaQcpFvW0wsa2hdkjE3HjTHcmFrJ
WECsLKYcgXrqC8/WwokzAmZwTy2k3lcoYwzw/W8ELx5zpM7WR680YgP0trr11+xjW9vtB5koS0HD
kZdp75Hnxigb9JTLk5U5tIMNIPSMMuh46pW63c7BaDX9BcIw7eLPWx1LG/uWGo8O71DCYz4aBrER
egC6nfCLaKGd1/KHbtsPGV7FMD81CLG4Strm+th+fAzH0oCU5HNxI/RKTEwz36SEmbCTLnuUVQd9
ROuTTSkZFSdV1dXHlmtffEAMbd91NK6ZUWTx/if06P/C7Su2ExFnS4DsmZW2CrJtrXjDxOAUphPg
Q+fm9Mp/9n0iwcXQFEMTRdgNILzGIQBQ+D1JhBDhyXbdW8xj9oQTB699pPjLy/IcHA8RscpY8ckq
vZGJnZcpt1OFEueGGK/TDCoEk2vf3AirVfuoFMtyfV2Nld5YNDLyQa33/nZokZq59xwHZuwQAvjl
2BDi42TfchtsC9vPdzODqh6YU4kYqz+jvx0rNNwvmOBdSgOTEfO6xkMAbmC22Kgp5DHiWZoxt/DH
pWBzqmxXyrqmonVGC5k4uVPGTlXuXzwEjSOrHbW0aOzuTsNnsmrEO+aGoZBzIh03dPnDIlZ2vC6B
lPtcFw9vi0yE24k4kJwN97ZnyOrh9Q1NV36P50aXtIggUA53hGZEXPTgnaxOOyV0DCk+wYJDZIVC
Y+whM8aBdAYExjyy+XQ4BC6dTP+YIRSIWsoV0CJwJjOg6q4ZuLAkW1K1YKjc7x9T0/tXiUSPs3JK
psDJWp1BOfhk4c1zlkYzyNe5a6cLCS3T0cy8ZHjp2p1a269USDdfkddwmEPl/IijhuMUK78ncEve
xeHjkil08KOzSkvJEDcX9Ya3QPxu5Cs6Itu1+RVWTOwmLBvDRbEUvywmr6HT699pmQ5rmIB1nprn
2+kDWa8sp4VAuAMigdQofCz0RGuDAttH0AAvMjOC0/lI1iP2IrwGSX8pze/tvZ4dMGlyP0elraeI
xm3XTabock5OZkJ+i5qi1GoI6q77nMHb7ma3mVSHKpfshOFPqOAdd4RszN0vJ7syqqFJqyWseVyK
v6sLP94qRmGULc0boEsI2YlOlHGGB6wThNW95b3LAmt9EaCzWdRI3fTLKgvbMrZ+uK6NheME6/PV
vwHACu7Eyt1wJVH1wJRkohVb4+HiEhUDRJiqZV51AC9b+kIN5PLiK01jiQl3fPdFQ8U3SS2kKqEQ
Ze1DVrjyTX5sdSgOtyLVdB9f5Bgf9D0g/RiP21Fit3RbYiCmzKsC3VachXOQTJUMaxPKtMuRXJ72
D/rTcUOWkC/N76JFI+j3PG25+kxt+H9wCROCg6AoaeD+gaqub7Z+oIKXFmqrt2qoZpxXhfa2EuiQ
nHj0SetbGHUqda6X1W1APzoYnlSW+dbZ5UAU0Wb991UxjlseeaiTbZitb8N7kOv6+r9cbhSbRLQO
j8TUkioDFoLH3rTDf5aDu8I/cg8fwQAUnDX0hgFBnqeukOTerBybwAlQDvRaPL9f7be8z92glEyl
wUijonZezKM+HrA2uivNuKF4WBuVOfYz8MVpo22gC9e5JR3vsizkV2Eu3hQ5NNPAxsb+C6WXPn0+
AwPCRBP5M60so7g5RaDeC6mvWsTzUMu7Z17D29JUISqnqxiZrgqRmXMqX9U/etS0bTQ1POVqw23f
WEs7AS1UL1W1PmOwMNrf4MJSx4kIfhG2fJxoqpXqWMiyzYGlVUEj/6m4xGD+ESSkIZK6JwOQ2c5n
fOjAISuqK1q2hZkMV6oNx3lq+C98CZLURwnq+zyvFJK5An1UOblPAiUyLFq1RnPfN9g3NE5TNxeX
C+VOfSzayVl5OFVFpzQsq37m+WRgPtNqz/HplqoY0elHUoJsE/qC8xLfyiUdVDMvYA2hVhP2IohU
VSZ1CL3aaNElGFCoi3d3JCrUjYK1kb/v+ZJ8rFwPD6qCmnelRz7cQVFlyBa6EsetPFLLM6GrBI/+
S8buGryMLIV6WONbXDxbXdH10JUP4lp2EbGeI2jcIavuIrSqdj1jNYXHXKOt3ypXYRPd2IeMgg0B
sW32rO58M4OZ//iLLADMUvg8imSsmuEQEhmAaaw5qfFKPXamd+m+fIEz3gQZNjSFzitxc0/UYFhj
36pwyF47NR3KEt9qz0sDa7vyWcOXfUQxs6yQ1QMciyK5pSIpXsNE6X05KciYapPWdeyvehMr14lC
fuTvEXiOPjOQLo9APvYnBYVG9MjAAAV43+N/9l0WGbprHNmsd5xASIPtydOAVODypieZu2gy0JyC
3HfH5NqFCrGT9c+o0T18WvxrJWcCoqxUXt5Z3gQ5fCts9Ae2hR2XEwLzsG9qQfokPd7oYxVR8KCb
sVM04v+ak/zMSwVTjXpM+7FqhjVbNR5k6JjqDOAoGi94uNqEBgbfLFahLxRqMId39ZL9L0TYMJiE
mRhxi4OPdFWZy3zslS/EezX8H/rAJIIpNU2qr8KkXcqS4vcAXvHqNjBoB3cEMKLOSzJY4xXe9dQx
Mzv1TcDA7XD/3sUVBrdJS+3LbsH/gb9zVwTkpk1SvQ1OTC/RyFr8hMI1UAK2Y9Y8PqMSdyScflao
uI43vf1MA8rQ99uMHEgdC5vE9FpU1LNwaT5muMYOk4HvX22nIYB53wEY3KkKEb/F6yhYh+S1lwly
DdT5AsIdnEd8uUlPWIQc4b4st2qWaG6aNEMcd4ctBunDNcvoCid+ykpyAlxTMAlFLP80HHU4LDYH
Ldh80d7XzBqKLGqRKeScwtRqHpRCA3y2FHRhdd3k8Y2AAQwwKRsvZZq/oTrHy+kFQNqAUXoyuX1n
J5zy+vJhpXQLW9iC7C8eDOpiQ67lrGNNTky3vCSvOUF5b8sw5ywdnGSUlz8OMWyIZepwr4XEY0Cd
pUbrXG9YLbm2wIUUduxRhRV1lWUQkyHGAe5Z9rU/ZqWfG9+Rx4kzB2QpKQcc0BYWK6TXVWhYowrX
8UAJKE/Hm4cGH5Xg7oMUmZL+0Og/gnVtuC1pVA36xqfKgxbxBrMiHZxON2hoC1/DY+U5sERd9taa
Unstee2wtI24M9kW/kng0uyeBWYGFKTBoSFZEiqwGnqKRN+d4Bkl7p+M75sxqH7bh31CTg4yEdpb
GNhCfYubw1pMoJNHxIuYP7yanhLn5RNjWN07yvz6hsWkJP7RkHWadd1nNwiY16D6auIXYJw65dGc
62out62dr804/SSsEmyXL+lW466jDxQxmlV7LNKKgwHjP9r/Y/UI9M+PRTdRt6CjG3vW2SFWJqFA
tbAX/XkzC2qSaoxLd3TuQ5mnyX3gv6N5FanvD/9nGA6eTtlFhfSnPRJ6dkFh03c+Lhx4SQGk8vL9
EDOvA9ZE2dAl19l0UzpmAI6zEtcyDcIxGoOq5WMF+JxPjJrfSFolt1IsJHJ2M2NJrJzgdS8TAEM4
tfvsmK+U2fedapSSx4V/HXEiWPwRZfyZ4pb4NW58fPaOZ8R9ITrHc3V5ZgXGD1HSrCqO34xY36Y2
BnUg9EwtO0bYx/o3dgI7p04KkKsnz+u2I0sfFA6EX0eEnOj52HoDTI4GVDVO/6aNPqtqRKSf6oPv
wwpv16SQTtzXsXs+WG8mdtQUuoelUvgRFoFTSaoKcwnAY8Uw/cvHV2zteB9RlKZH1HIxO6tJmZln
rKLH9wU+8COa1dguzePoR0RkDvSzT/qoYWoQyHapTgAOsegNQ8nh6SWZzkAGX1oM9A5gffTXNJuQ
psOS5yukakHNRndL9g7DLHh/PYGp5vmVcjCfeen1xlOd1R7puAa5HLi2A3/1BipYVGZoGDTPswOm
DgYQM776affzADEsKq3DvfHDEyf3Ad7QAKL1mbPq+QgoB5BLdJe1c2K2bVdgkzKOoV3+EKMH6PyJ
cTcXzLSwgTgQvTnrIktg/vYAFt8Bkk4PRgGow4M2kir5KFD65TKFODs2qW9YNnfFm+CcmcIiUSmD
dzNFcK2n718FFDAzIPpaxW0k14MbsFiUgFwid6RvVOBQWxzgi5RCN4Gh0ogSoBm8qNStoyR6gmIN
O7Xaz0Bp6sfxdRokQAW0mBJpFq972Hqf6edWT0Mwf8fBbzCZYsezb5R76n1rlMfVK2thn0jr0G9k
GyOD6y+wsXWOOP1OvTR3vukDtCy/755iBPBtJ67bufJpbM+gxF/iNpAahnFmuoff1rj/NFTTPtP8
PwunmSn2n+GellwaH2gINvYnSxDg55dpaCLXrJVnHf8Cx/SxOwfYI04shds1PNE843GN/7Ym0oGQ
xE8JXLhM85lAcFxplC5FAw7shfshPPkB1b4ekgE4coYO1IBhc2lX9VA4+3DbFdNKdnbxKWBz++1h
VqQNkkSTjqoCTjiaeN45d8rfp9oVrOQWrUJmhSyusPaQdtcKeCZXSTSXeX8QEdbOqdeuSKjSxYFc
ESbHwo33vT+XT2cMFaskbg+jSo/kCjzCBCLxuuK4XwCnhie4WtDXEeVaTP8CcmqK5KwDNU2jQ5cF
IHES2YI1PUOUqPa5qbwWb7v7MDrXkukBqM/15Qjuc6wU2pwqrPqslKHpHCwInOa8XwNzXlTvpkf5
Gy4tg4A8PBsZ9sFn8OklbA9fKq6ix97qY7LdGBwbkHioiTmcqT0Ac+k14dJbOzykg4q2U6mXG02O
/mC5RUr9+67JAbTCQPmplLiQ1E9UqImDiX0dlCVUsZt/jRK6n5MLooMkjQyod2n6zoqnN8U6fT4s
oR0vIF7VJceLnlLOXUGZALgXUASSANNcq/2XO4tVhV0fn0F1ih4X2tX890s2LVLA7bkm5P7gvgR1
dcZkJyPQepbAPKrkJfYO7KDoUlC1/b1epdWfE4Uop1LH2qlXPgXesXpRXcAC1fD773o4oF94HmmW
Ke9dIiJR05UibhefL/zD3H8UcbEHXXevwVMi4JIlAgL07OBk29rKyUrokiDYtoNSQI9Mwrak5P5z
tHnR3ZGDMK7GnO2Ug67pLP/IVrujcJePquVAJHyIwctbO0HqGHi0/eCm578/WwVQJkkXZ7TldOTh
J02xQ/2LJEpFo1nj90a7nJr8CgHUebXzZskaOd68x6+9OrpmSrjdq0L6l2EjSDMao4osGj89EzhV
O1ym5MTn0ZL+gRaHzrxPRYoHg8J9EsXq5dUMIccwbZZRToYGdwpURZ4fb2b+H5NEoKdOwKDpS+Fl
Q/wL36r6I5b6kJffUISlNmr7nopTK1SZbeJ+kJsLqGC1FR6eps1K0atP1MogTirJ4hGbTmi6lRvy
SqBVnxHvtK4CctLeSHiWkVwurUlvLwErxKSMu2jq7gctavEYoQ4PuiHVHg+4fTpcedq9yMtLe6mV
9Jrh5zc37j9LQw/oGQn/HTBd66m4TH1LF0RGotn/dht0MvApal2+PCCoLRn5qCEDta2bZnFNpnuv
8PEppttSMVGQocDzrWTzvRIB/WZzf7UCaURLirnRAex1f69EYDKYUor/8VWzvqwNYLqj6QhnSe2t
i/A0SC+jG+pSHKlmUegbbjRuR5nUrvx+PDU4QouY591ylQ0eIk3StwUfiQW2AykQysViff9+9b/X
0SpK0gG0b9DTAyeCv2/a4x3s+3arSk2w/aBR26GhTX8YLD9lpGYDxi7b7KJ6eDrq70b4mWwKpC3S
4uyzez2MhduotZ95D6PzJd37GJK00B3tSMT3dM3TuYWwyqc/41kQ113UOcEJp4kOIm0pKI0WNb1F
ywxjDBuuR5SpSqsAFupWlZxeaAqoS8Sr8X8TqvrF5JeLnWu1MtKiLDtE88ji7x+n3eXK48eqhnHV
bwJ/AyVhsB6TUe4DQshaqBXLs/Ow/R1nLI8EI/2jzbJRlimTPFFaebx+uJtda5muT2jQpRFZczjT
lGJkKbSRSr0i05/+feGQhiK5RNYIpR5W27S++Pj9HEYkKoDjsNWsN1kFuMcNXtZW4BZucJRrnMvj
reqOW7m417wYdU88vdbXVTnMQvvYxhFkqe/xObJGsha7oh6JJvgS2wE9+sYtyjNBe8JBMjwfD2+F
V4jOW108TjRcysD8ghtU3n1fqiBawQxR4Fs1X/neVkRMMz5isPiyPL59VCtXtkY+h+6riKiMSgyF
dA201qkO5FrqTWKK9mgjUWzPs0C5hg0UoqUdBl3Egk/oYpCTf04FRkwGzcuIj7T5TEC+xtV6+VP3
J78UOEc8Ui4L4Kp8yp2jQyWWf3kRPVN9hR6RGRUA5kGIiVnuDnn4MdQiCuHatqYJwRkvTpQ8XNtM
SgTqpRPT2J8iW+qOMqji+PunU4U8I/grDESSZgS2yqeg69CxSAaAdQR5opW1Nl4+X4+P9i8Lj7T5
7s6M8KuCkQCJFYoZH2ZIcNEqH11Uvlwbz8bKazjKlrX1oiTLMZWaaylIfnNAh0S4s7MvbujCNG/B
Meg2igNyT3qpZcRtT1NpzW44y8N0Ev5VoLpF7iHhYs8wjs2nehpnXdc5zUFUA40MPKx/mZnBsjV1
LKVVaCR/07VoMmXIbhcOno6hYdXiF24sIBTUORLtnmSg348JjrbHFdD9vTeizJhhuwe3JBQ4sUrJ
OjVAaq6eqh7OAFPiN8JXLs1yhwmi1Tl0JX4DsKeUGKFkdEBQLKCcQrfUpX4QVvzpbicOL/dVf9qo
oD9nmAcAT83Yd2MNzUVTeudhP4sa+qpuPo3OoaPGbNWXG6zTevLKPXpQTiM5r/ZWluQYFySia38A
XOYNfhAvz5epaNnnJyvIaTHT4Qom9emiXSUYxCcqrlavOjSpntozoSMuhPrCBz/qM4f8jeLD9XUH
Kp5/s2oV3LTQXpmdEVfpBMBz/FjciUjRt9IeJ6bW8CEdLxTzymog1ZQG3PMwRetWPZk7QYxXonNb
FMdb9MB27679ebxGFcSpnMKINFKh6V1BBxnKcDopFGbImFKXz6XrQPxOdl/zt/yl3/ISEjA1s0j9
YqL5fUFJhACELS7oUuJO0mos+06LG6Ojssco+h2le1o+TmwT3pjV+Q9NlEnEqRQQLcn17Jbdmirj
D9jssMbt98wHInxm3nOJeujwFRgeiTD4/gOmoUQ/+/ukgRDR8XwPLM54e3++Za6qUm2fNOdsskZC
lptKuNNjUutvbJ3bTggaZRRaMzJYq0cbCbapl0z1cG065iUn5F2xH3g6wB702AFu9iPdBLN/yQ82
7Qx8JndUBNZ/SBO99pUpkZHyCw1n8UGIPGT9BLke91HjVv/89N57NYamqY/sdSfBIoYno10EDCHB
OJjt2SHeS+kTrwa+nsHwUk9+b6MKVqYFzlI+/s4ogGqOS+QnsXaxe4QWjHD8kJhefYsmsrPval+o
+G3LoFdnc6Zdatea8SoqrikuAbKcXcVpqhmqVWhOWmpCwkNfW3w/DEya7LFKJigzVeFH5h0KE7kD
NuYyzNSJ9TwK0gBPCBUt8WE74Ql2Q9yL6Qx1XponBCu6WbkGbMmOf4QwP5GzNO+FwZ1TM+PIw3hH
SOJHyLfIcBfB68JIwV0KpQjQvnc7mHWHybHrzZfGyAPYwH134eQpTRzZb4eq7EHkElwo23cOgTN7
dbeCcy+dB/begUwimhnWyc2Nr2eLC9Ff5WJz92e5OxsLiBTbIbYEqo2i0st3qvYUAVzJ9qqXr1vP
pC/kEEH5tvydr6QR2ej+NZ7IxMQNTHnYCV7lWCvvIeCM2VHFMcGOzs0B5ZthFsoRjUUMGyCJWycC
zjNrHUNp0FArboQ5tS0d/NAvtjyOIwczx5qqTORu/OT7gIgUhqAkeeiCuzvdrgrt486RsJBldiIS
r31SrCW+nWr+YUZAcvmw/2LYih/jo3mAccTqqPQhwl+8tVe9C6a04/dNcUWyO2es14R17mih1HQU
9UGeEpsvV+c89HeahTe7xzeyohBc+7C1OdlFucIkxi7ka+mMsqNUkJ9wnYu7e1hSQe8et1WOQEjP
mRjJNQISLrYsHxH6PtE7H3TB6tFX/6SjNlh6brTLNtDnKta0oida6G/sVMBxApnny0+IonXcnrhA
RyAz6we8dH8xjnoxt0nyPiij48yzwJrnmh45r473QOjD9/qSzGrBRcQHU6RE1TFO0ClzDBNbEjD/
CTjYmnlH7ZfmqyFIC0unckmJfZg7aB2o9X6w8hOQBSSGH+aqYtOtwoHivGN1Bs33FSqioC+ecp+Y
2gWlXqTx1HWNaXNcOX4Co6ReK9mxTGic/bSmCM+PJLuzVKdCW23ODfMfj/CL3zpME5zDOGr+XUe8
3X0SMD42sto1eWDNriukkrO/JgnMiYRvGOAZIW8JME+l5shr+vdaJasKsdxpfPP7lX7Yo8KECyFB
Knm9tL+QvYUU5E7/mvHSH9LNkP08mgCwTHxfd4e63hJpJLUjTPh9+k270sTwiIv9kSHXwkom5oKC
XHRtFPsTsgxGaDFHLLx5iBeJRHaSsJjt8ipSR8OMAQzGKdJd3nefieaKCF9D8vpDS79u0NpANfz2
SXgcd3WaBqNTeeLr63AhlNolb3YbCCUflQTeVzJP/CQsU2IO65sbyQryEvqyddO4SL0mCW1dI4ZZ
9i3pJ1pckm3TNOHaChP02/s8vXN+7LK7cdXSQ7FdwUCk/iNxMzWIPlpjzGyY2mDOvoGOWAEGbR81
sJpoKLz57Dx9k3yjTc8bZAKY09ttLfNYNaxqqsrVe/tgKJjNp/i56yC9kVXtnOAIGvzXNDnLOv5F
3Eefrm9hV4LVqTl7idXn2bh6PlZ0v2v9N3PPxR44ZCqIhA230ZZLU0NL9TjT5j3UCRqYycIKpJuE
mb1GR8WymhN2k7BuQncHje1EDafrNcjtmGMplXOXVuFHhtxIVSuEzeRYWsjwuf/I/BMtXaBY5n/o
MWVOQEzWVgxx2XfOCgE5yBk+3okKa5tKISFeCF5pzC5QdTqNJgqvKqjI8zG2fN257HESY/x98x0l
8+6plCOl6RtGiZ+MWSgrKxX5EiZLEKadou8gnr26aIqcoI0DBc4RMFlF/zGrrhLk3iVSlWpI3/rq
Jr5YirG/9D9xm8xLWSkd5CDDsyjLZQ+05AU1ogx1zAUaB45ux3of3Who/f1p1HQVGT6lWoQatydP
zfvZYWCN/gz/qydW68Gzfe+syP28EZaWv8WXYEGCixe+T72MwaU05/QY33fnEMOyuBkU4P92pPF5
Uir5Ahtl5vO6HlThKZUd/nCMcWdIR9j0WHeqjdu7+jSSg3rg1E1I3GXhZK4mPAQvbsM6r2Ufse9R
0QpyQrc4Ux13PdEoztPAQe8Z1D0qcBcC5TLtGSX2Jfu/egxpBb7h9OpWzYNYQEr0RzeJQPK4z9ad
B+I8ISd9kyBrA0mxTdeHkytzKVaOZgFJwsFwMIkQl+UmGvh2s+7guthqX+6IstRWU88ekAwAr6dE
mnr9sJw7bnGtmobfQLnpJO0ytBGXoXXy5vMF6bd8HN2esEtdvE2+nk/8xXQHdBEZEhzB/d89hzd3
zqBWTxEzHVSUrr1G+whhaUs322KRo/rkM3E5bf4VNU+hFXVqg7dv0wDRQpN7V/uz1JVKI/+rdxWn
5nsiKd9StyZvkNq9ZvtuWkp9DOzvUcW8KkN3jUCFKts0nl2jU9CNNR05uHYTCZZHOJJ5p25XoerQ
Jh26ORzavAo6As58RwNgbr38UeqOtQxo2oAUV7YD046xvcIkWqyZ4SbwDfuFG4nV83ION8WLxjW1
NCuvxogTD7qUEkXGk0nIjnIrHDef+lpNb//pDDp2+KQRQvh1uhysVT+Du0+lHuSgsxvExGYm2jmh
tFbxJoAgI0JRVz2zBxInREmoxdq1B/J4n25C3P5pTfJQEr3Oekr5V6e5RkrQ/eE92kWLIrfZ6FEP
j8kSP+X5J6ludDgGCKVpfMWjdBOZJRvlsAIUpA+H7i2P0vZbc8fh6+17GCmPlEMo8fPgdYIonJMv
6RGY/bWm59Tw/dWZLDYC67QP4MYpI9BYQlZ0xmtAQJa5bjcA9Ir+EV8nZ3VCmPfg1HgTrLW6d8C0
fFwUophAMXbAUdyOkoBbc8deSBLLcKrmQvARuXmfF+uEP7a6MJQaivFfAODAv34yTp0sxMnYbVCm
SGgGGWoGwRchh+oDhHf1YV/bJr06SfNaDgAY8wkt/G+pAH0dWB01egT+QXyfTc3JivvT8CQYF16E
92IUosVEilI4CP1ODr4SqgK5QS3UCaLIdBLMxygxzzKKw3PqSxAreVEHV1Z5ispaLxw8dxaSmP8o
A0wXnZxm2zBu+CMfYj4Lp1fgQa/K7/ZiLONLVwizJNLYLrevzZrU3AomC8tEcpxtKU/YxvUWfxdi
XEF6fOZrDuOd/zo2MEb5BOMERDiqI2R+dtz2S1aBoWwnKjK/P75eMvlJKmsqGqKTjjVSHo5wVzYc
+98IyjuB/NraKZZ1J7Yt2BdqlzINldXlgUvG2cEauvyeUCXIK+O7kYz+rWBZwf0PwyuA2aeCxy2z
GqnOgtIB5o1iWBBZwjxj9FC09nQFcW7pffkVNBqOezulQanJZMJtYRUBdyClc0p4ZscMzhCBULJu
faYKpNfmA0qPWsxN9lV9SmYpPzUQYItveVTYZeOIcGZjREuFkzpjo/fDw7c9LpFxdcANtqcjER5i
w9hn62Gov1pD/e4cah8/JpvjkpQwLtieMtWe9dDxypxtXMlFqpfUnMdVa9/RulnfJvqSUfAY8km7
FXhSoid8bLfKVBJLf7RdzLKGaDRbxDWulD/zrHUqw4MNo0Z0/SPEqB33qno/rriSUYVP0vLdN9AL
cIentbKKYiNFf71XQsGjw9bi/Ca7fU32hHQXQO59kMsn3txrvMufSAW1/sx7l5hsnD7j12EqEJfi
LHF+ag2OppY766pTM7M+a8UBf/K6xb1yHDsk0XlRMb93g228RIP/u2xIXm63e9u3OcygB5qiOfTX
icUYh2jUEw5XwSxRf4p26VL76lFr9qSnhSxFYabZTnzbfFYYzzlz8U2JVxolfeQh4QG9XEan9I4N
LlSIYH9LG9kAkoSVLEpALIhFzuOs//cJLqED7KBHIO/0cDHKylL8Xrl2JHo0gacp4rXRZt4duPkN
mK8fqSeRpSZIoCZIiWmVtNbbtFr8/g429wnAitusR0QVWh9jmHpWvC+gTjyCOycswN+ZuEG5U/s0
zr+hdIOgfuPhUXsnM/SQbRUAj5Sqgfc/5OhSAaM1WJ5Cbl+XAp9OKvW/V+uj3Ouj3GPLInXJm9AK
0lshUZLxKHCnpXDsFvAr7RI7M/8/o/8SV+qziznCVkA1PMyqt3aBxvbJ7UQuVH1fP6zLA9pIj6vV
Aq83wQJOMbYUkDT6epMmsuUAGNnA2Voh5nYdYEqV16+WS1gxqjr5raHdSvsVqVypxDE2QT/z+a0F
O5RTcXU18wEu+QqAAqIYOzGCYei3adZfA52XnhlBn4c4w4WMKKpbkFghyT+GdCnkvzA7SkZtu2Ms
CDJXaqnd1P7gLWYIAk5ZDfeBbVAIw2+3YoIXNIiUZrxr+ObjRUXGuxhUQg+Mv/xNAiHfOSxtYZhn
ZOPsxRklf92mWFjGalh27LbRbbqOR5fI7on++MPnS6Pr6MHuEiqAkDh93k1Snlf8q8Ild5ZUzwjt
IWBlOaR70SL8420p3wRc9dnWCTKEGD0W2YMBKKDM42F1LAG79kCliYX8uG3xMC0d0hEv+g1WvG2E
e+AulWNYEN43kLFEyMmGuoGhdVGX7z6lSns2jv49I5ee3DEn1h5vl5aNN5O1oeaxWk7NCmU/SdOt
DRrb6HwiGtw2zJcCX/RIkoS6Pshw9M7//gGKAUKy3j/VV+6IDlVWiI1hiVznaRaHuIip4+c2BHZF
ExGZjepfpKPtGbt70PFhfcdD4VAxQeAciDNSQdIQQDnYZmVUVIaGeDYiTPH4b/JIZTb+0QaaWqRF
nKk40X+NVftq2VVJV55VmIqK3HeVkj3sHZqrH9b5lGBqOe4rzfg0ADR+8Aj0cggvLHm0C8Wn3DKl
k1DPMorgZciik4538VgrAqxNrjACgBzYHa1DN1RP5jlqsZi6U+Sq2M+hniLTOlJ5f666LQXqcGVu
6RyMGZJim/1R/LhFrmpCOHbWTrV1LOipwFmyjAxrvGunPXzXvwIiQRarf4Mg4yrcCNGiaMmBYOnz
NYcXKQ9SnAsEa7IY5quYxyJAfzqyrDbHy29aQAkobiHSJQggs8B1MbUrG5b1c1mz0/Mz1gmfk8Xq
0SrzZzlIYk6GIjR6FfN9wdvPM1gkrTvl4ztt8zzLCFrxq/C3P6bmfZaIgpW4Xp8qdCQErKqLGA8L
QjuJfhTcp/6Sp8AD1YkC2bnLQngMaWBKBOpNyOkTpS6Ysk6MTzmZ0AHCRe2aixlTDDJAmOWEkoSQ
7VWRXTu9Fovle/gp8o5+wH2yCOWrnmVvkeCCTrUDyEJk/gIwKL/T+T1WiSdJULV4wv8c2otKpfn0
PSsYuMIVmtnv+wnHE2pthRaHT3MAIjeiyWB/xSvrgVIKkZHP6RP3Z2PjbDkYgzrifvJTo9MLfWXf
M2llstjc26aRzNunACUFfkra6s2+1oLHhLoWZGeiNoXDl/s25mG5TBTVEuXiS8+bE31z63v/qPvg
x/uwRv962712iCLw9vmpPHWCeAgBxMzBnZfnxN3+oXMRjVJrY9vvB4gB/HqxZCVhf11Op/dkUrWW
pH9ISwTABJC4ZyfA5WGmd7o9xrJJnZKvxEfEt3ZHkWgXPmLvUJfsNcYGUhT3TfUGIiOBOCHh9Y11
rDxFy+Wn+VcZd3Jkr3ySPMalmDAc5NeNsOGXk4FLYo7irijLeUZ8m5uRe0o3Zo1IXr+DhW/BirP4
Vwo+7FOlac6PhAef7jWYiw5x9s+HvaH5mtH6vJGGWq/ztxcyfNH2T1Ps1KfSBPN7X+zcn2mE0Wja
dM8MRz7IC4bnMnsLqdQj2lP2tHNq0ZIuDZWzcz1+Dai6z6P3n1Yx9F7xVV+5ceZwos7WUk8CGRjz
RGLAiufMBViiZNxRTTfrIlQ3zQ/DRYY4IMCmPxOOllW96TZo0jx3XKQxW+OAhC6H9LrNS/SaPiEt
aajmgu6OWXGtpLkB78X4woGFM9VcIdtAgfpQDrTYTOflgcG4RqmnKHoHyE6kZ/THqaOn6wHnxXI5
bsCPCDu30sRt0ER2XG6/6/K5NRORf1BzOyBzx5K+VGzhrQfE6VkqB36pWJcSWFW9F3DH8gs/f260
dIeijE6wNiIRKP7gbPAV4OYif3S4nxVWegFGT7+lBPMFbWp1+XZ0KJ2tu5joiUFDjyvsZ6S5Kutg
8evoXJb2540x7+/TTvO6qqt5V3SrRGv31pcMMIuAZd97bXdcxvOBFTaAEgeiiGquI6qwdFZWb3Zr
I7OTBXKxRa8Ue8qwrnBjt/3RNMXabByn68DtET8ERxtphQkqcyUW+dTaFpqc/fHlTbhNQqEh/IKT
QZSI0rMzMpUU0F4Ra/haQELZs4sBXvpz8GYSFEYLtUYL8jLzmwKYNLzY1B7F7M4LpekSrfJUVfvW
NLT2wiQrK0VpjQYjTS145S8GdKlVExu9ovMvQG/3v0fAJKQIyglGTHOQgwq9SAYpKQTORdmapCm1
TIjjfi3fi4xJjnudZ/35JW0j31KvJUhzXahguVNrJFUBI6r/bS3lgI8zKlFB447c7kyOcUTShSnJ
i6HFP7BTBJBK4ww4ldhxSqjyAk1e3S62GBAmHSdM/aVQXFKggTy7SVHiroUahae8/LylHerrMoq0
iE+m6sYLQ5Hcgdl3cRgGCmJ4Gi/YsJJUHKjBJcsIxpMZVVXM/mV281vGbAPPq/G7gdXQ4/E5/2M2
heAY2wxg9/X0TRoxK7/uqYc6fD59LXPpqKGO0Kb9DTYRq5EZHoGSv7GShX/scvY3cL+splQGPYcP
2k6ZTwGkCxATdWUXqZkLn7o4p47YhH2U1NZ/XtLnU6H4WuNZaFuacoiIF7VR+H2dqEdqnubEp1BU
/6ZI1rnTff8DbrXdDHwNDfMNpEgglDCxPDZroD6jQHIFCpWC1+ZcinnTBAUfWUQ5aqezTer0bo+s
/bOlhS7rZzRF4Bn4ukY1Fid3n0cD/GSFoy9n00QqnKg4MToniM8VTl+LsRUHdfiPGac39KK342w3
oAFKuRRUvgHjO6DDHq0qYpzyuXmRHiLHQlPR/kbf3FaFUL0f1fFZjVr/BHEgI8PjVyVReQbhJgSl
YaesBNjA7brsMQkqFO9usYZTCoHlRjvZs9cwpbhKrHN+kZBVTsgu7Mko6PV72/OBkiJ1A+Np/RV6
2AIXkBWE5c78q5oBjsFUkyCXs+c35z1IPPKbuy8E0kAgzYFY3HwV37BlNB+Eydm1qKwlHti98Lb8
JQMeUc2tt3+imKNrYk8RDAEYhGn4H5/U5eZGCSv1eheli5NHjUtZPOjU9HY8PxRxpOGy4Rme8DsS
mZkFMnPuZY0hq5SIvrMG6Mwee2WNROQM7kCIS1mNUQ+qSES08T6D5ep6eb83W0kl+eZ9wlD5wzLZ
AiBLh+QfmOFv4tBxldhSnrVDyLhHiLvWEvabPsGdDZWnzHBoYc0ez+0u7aQ4K8Uido//noM2P4G/
eJGLszuv7XiQgn/XXxM0RLzYBeGXW2Z9fCazsh1jPTrv4lpcvYzqQg/IkIMOQclDgyzc5+gxShsK
XuTGErVoKTYlwsU8dWMoSarioGXFUqW4+kFOESPpMzpgFZGZHtXI4002XfEs6vU0NcYvxTpsyV2x
acqHGf5XMjhf0uQaCtzOFor7X57HiNagzgSpEBJFzZt1+FetNIUPv8JlDUPtk0NqgD7WDF+UukWf
URVlqEvr6QZbTnaY/Vh5hszLo5b/Zv03Tijy2/1HZJBtHlofvnt422rPI6oDX0Y+Rege4EYyDTK5
e4foW7Pku0zKiMjHc80veJZER4XLD5olFQhftiOtULNg3nSle0ZzaOo/uqiv/f/F4UewIcaJs4B/
F7USE/+Z17io4tjHdAiyv+R+3LX6RgmK5/Da7uy6aArVCUq8JmpoElASH3liVagckW8SSgUEpmoP
p2UBwAFuYWo0E+tY5b8RdcmtGTlYVTJpbpi2iTVg1G2JWL2kk0s6qk3hWoRge2evTKNZULM1ghFy
Ry2tVxtCHc9Ra1AP12fWKaDu54AWiymxx5TgD5Dl3yv2Avzg7DQAkoq50crOS/xnepzQkJmV66IU
BtkdNsy94J+VCDokH1HUanJEJIkRLQ2Dhyt29fOoQL+UDqmDRxjOKpopq+PgOxFpsqi5k90QIqDD
Fep6lW8ifADUtgayWYoqakwM7GE6QxbI3WQTeaWgfOAnvx9nIaqIBbRWMPBCHUpmSuwzgsWlJQBS
XX19v4IUhD7MROjv+/JRnvkPPXV4QW9P+zs+LSt4Rz7Jk9N7yXsikRd2oPYAl9puqhamABAI+c+4
V9on0LfxfwalByEHr5IRBURDM5G0Fr4+1Vjh145rMeihnTyQqxnq/6O3uy0K6qErCgmi7VIbS90+
Ggu8ztzrbxt83ITYg7r1eFYvPr4iu3I/QMjaoyX1ZM10pQbkXp/wqKPaphDEFHyiUj/gV4KyjyjP
LeqIOKePw/pNmDjDt8YKmNjlXpxs2dQ85LDcZqmXs8eL82mtnodWPlToTTOvGwFlWUg7NstLeobw
ebWYnU1VMVlElUf2wUrECKyhHSWPriVuK+6sSeHns+E9otEO1nu4fJozR99R6TwRYRl7+g1E1lHy
tSHWuxDtfy44BRZo+QmC2BHotRpCMpefw98S0Fo6JpAnkBBRJ75ML/TufkvpPiuq8vX9FjVpB9yp
PaVSBUNMa4CDOBbQsIE/ZsbtJi/Ic5omrLnA7bnk6Ap/OC/5X2kQYrdKlmEik1G5V0o4t2A3LBDV
jTd0MCqNwwu+BL7m7c0Nq8+sFugRNVNPpWOwEtmmcE/swms9LrHQFgojShgY8Jc4VfdH7SU3xG5d
dSC7VuMve6avooVZzfzOAHzSktHQ7ZrzEzmC1cMkVMjqXxlIObIsbRfqRpx3cdy9rOoLCBSBcspb
QyFWUiq8/zsQ76ugk/ZmdHYYKNSVRjs8NIBlERz0Gb/DG15V1Gz8i4vBKHwgxyfJxYWFMeGsZ53f
w9j16QHN5ZlN/rQS8ARXQR114wLpyp51rrIqsouynL9+DXjkwYPnL1bAzCcLvrQt1wedpBjTRYV6
mq7lJA98jkzEb6xKyWHU8fHZcXu0QRBWIzsG3EAlIDzBLZhKNpbuBaiRHBl/L/f69kaAko7hCfeN
3uBOuscKLeTRo7lpd7XNbCb5hfzgh06XZX4PUdYnl7/tVpoP8GY/s6Y5joPZ8V35nmTytuOEo+7F
QxxErZ+4dNvHGLdIQPgrG1REZt2ZH9iaYVaGkWKuS76IazLYMR17jY+wxyFNOWm+eMGG2dqSCX5A
KdqAQ2Q2/UXGgjvjfjs1oe/G/ROAN/QTzPPn2p1c63VdB/CXnNkcQ8Mfa5nNG/zZeVhB4DZZzi8D
NYLJZDWo+BbuHPlG9zdTCnmjYhe1c4KDKbTdqw/xOUKQp5uGvldmzyA5BMVwghQmLmopBAXlqBuZ
70EmncxxJ4mdYJbDC/TuwQdSC+PVfC7BdtTpDCue2y2ixJwZJ4x2NJr5cnRtFN7OCBDrMbwlqCKO
vfqb9N5qjQ+V4pSmz1b05WhvYJEG6TeZU6yG/V0Mf+RdJ7RF+Z1BEhOcMEfrkR+TRC6/L4XyZxsH
wyoJKThiBN44uTJ+m83rxWRM2rl1Cv4sTZRjbNUgWXGyVq3z4adou9upWGbgFIngEBDDNGtKu3c7
0GL3ya6fBBhAZdjdEMcTLvCRknXtNyK2LvfxulgG0RcNkbgXpe7c522fyEV5ir/o76kunreR8OeL
QobFFIo4WE5lFcJW3u2OeLB+Fzbdbj/StVPWBcUUtnPfSUqRSgqGmBecJP0+Xn74OVxNmhFdwqBf
/RwBaqDEheyHiAVY27zt81wQge3BQBEJyvGxER5rYOMFbrfoa/+QsHYqmPerBZenEO/4QporbbWk
X0I5uqawgwLJxj8f7FQZw3auk3XzigsJjYbrjsD2VrOJa3cj74qWDB7yZbA3kWtwIJqDnRbLT/+F
2pfSFUFC0BGPKubprAop7wKhN0cceE13UBteHZFCGy95gH+IdhAefCtw5j6YkvuH4jWe0pX4u6vq
HGhmpS2P3uPzgq+g1Lig0n5G2GfkktvSz9oYaqz67U0ylFvRw3wIJABLeb6BDM3vLGxxR1HsYODp
l81m+4buZruWPMkvPpsW4h4Z0nV3hPKNms3Qemq/nc0bhyRKpjqUqkrFowiQ8MC2RpaUdKl3Dqf0
xlCR3d2p0tV9klFkp92CmASe9SNAix+NkjbBHndiLjz5MA5hkBXzf/1LzQXvAibti9iQtuSLZcpu
3u+0FfOf5Rf6rsyPlTpf1nDx+T+eQSL2w0jKzjzE0SMfBw6f4IUE/eKUt5p8+8NMBN7fk6CkbVR2
HvCJFt5Y2pQQrO1jfG6z5Le2kJGvrNjvGxZL8002eH9TnJ9psgCvwyX8lXAVcFA5GkqFt9LfIw77
/oi6Zf1eSOWwFgJZ6Fvq6SFPTpoyaYJZETAVpK3w7HwIT6iBwBOdWaxgfpkBZS70hWTlVLtV2kpD
eRgeVlDn/Z//NBS1be9ItIhgVy02cl4WOlSmFFHzaGYBR3jWksvZUjhzNSenld3KCPOz9xSZwr9V
RWdliu5aOJKE6WTDah3HSXK/C3h4crKn31ygFp0UX8aVtfQ5yeDu0XN/TxRPUGi6TJ4DfORfK/wj
djlgaBLRP9AnwEZ3AHATwg+ComuiVe0cy7Mo5mDtLxjOn9Kk36zvRdT7JzMc+NyvlNZVqEI/uVi1
pqYEbP39H+tH21x1hmaUOtUNU6zGEfYBMNYhJ/D1EebbTIF38tujXNjY6dKW1ECN329+JfoSdGeo
VzBi7mT7VKGOz/G+QT+qwRbHNLj/lfUR8pv8Iy73QC92C7qZ51Gr4pqIVk1a5dTtYZD5XOWQ29md
tCTFU1xN275hvsKNLchsg6MsGAkwHgzTjSMjZRq/oB7B/Imdc62NKFWC8WHLTBjqNzRNOA075ng9
hOyyhtjmn031rTkcDp52dfwPJBo0kkMJo49lduj7n1RmStyz2LQAxzfCM5DY/QKE2K6Oi2X7TSoO
eCGv/rY2yahdzx7J0C95gU/LGmLLSv9EFd2wNkea86gYE9HwRuD3SztEujEF05/k/LpSMs1VXwTQ
MRb+W7zKdttL2pdkPjsl+99TPVnUJFPzkRaaRxhBC3GZy4yH6SbdYkBT6R65tkLqk/3Onn/gZ+Ol
njVkgDoIYQxBOcUOI0c1nWnh7ZpThHVdWYS1d8AYEtUZwBlZ/79nVlTq1WIFdOYU+MOoBzPKHpOZ
igJeYgo0M1wlzLYCu/3brala3VN4hxb9S8B01qPQbVqJcwX6kG9KfMKDBeno8JieefsxSTl/XoGU
pf5L3WU/DU4m1tYHTW7srp/rYO8RQho3qb8qe6vEt2Ohq9XjJndgT6RzYEi2fSySz8hyr54K7EKl
q8eUW06Sd8/KtyBirXEj4YRpu2/j+7WuwqgkrGLSxoShyv3kQxcX31ZmXF8RhTwhBa0duZ0XDfWZ
tYxijj56jmn1jRr+q9OJLDNaXd4hz9hys4ZvCODNn/8RWE0Z7aybgM+6D5ZxMrp4tfHkbD0gdVRb
FgWeaODvM6MbqQLwEh6m92VbvsmtRnLsoae89mj//lHFs32S/5bt6HX+KCbTjEmVlDRlizIb/15Q
a1CfNSD02In5Ilbst0sAO+JAyNzxbfy73zYkmFlnBZFcbyqZ3J8/ZY/yzxsZau8yYaqHZhCdVHFF
cctjc583XJB4g3AcUCp/pvX/gO4D4veNGh0P2TgLp7xhKDxXGE1AAtpWw+lH3ae9eE+2KJMZ0Omp
B+wNYtU+ptgsnJetJUN9NBltXPU6UBTR3RJ7kqmUlq/q6wFH9P/3lorhFpcLJDSomsCOgo+S3+0X
RNjCWTg4C9bjpFMKXNz9gx7kN8RTQ8bex4+wi19lNym4vpcfqTkABPEJc6su5APv2GtYSK0weh89
raTuUSV6lzQ/bEAQU/vWilSwWUGBFfzwpnAfYFSRmPzwpEAxX5R8jplXKTpCmVcw0R7KSWUiXYGx
GCzhL2YLH0i4me4L+5XBVU1oNXpjB/9Wb9zWoXchEXxGA7JszOmkWBhIHU23Ks2ejhm96gB0ASkp
8+Xqd9b0woSDyVuSJcHqLfPUr1b63r1I4kQg0fxA0fQ9G3HmPAQxLuMwoy0w+W5+yUMiy4cH2u0N
ZDFk2d+voVU/lo98bPVew8r8BZayJLTzzJsXxDsmwCLnezvGufjq235usInAp0Gi1jc0aMtulfKD
rdHUTwA2ZZeYbEjGn3ZZ4oNaxIGtk6in7O/G+273Ink7QSeIrwAAY+Ix2zrTxO6o+L7RHZL51pHt
X7cYBr1xHE58BIjj9+bGz5z44dnQ/a49013anxYoKfb9sCGqHKHqRPqJYh7VoTrXoe7xjLa/wu8M
0D7Fq8GlyJepnHQ1F2rrnZet4f4MPOGYGHXOBuuozn7xU2ALRb1URu+O1Kq0Z+EsBWrl8ZMoeKno
2eJA9z02oC/o2+7H+IwYMbh+vadrF2ik7wooLckEiUc3gWrs6BUO0wWG2wEy8yX8rvc9qJyhxkKD
z+FBbzp6HLHaxm03XXDC0tZxSdEgR0jC0zx6aS+75vFaaZ8AqlSuqxkCrjE4m2qgGi5KKoZ3nVMx
oFpg24DsE0YhtNQAtfnLT4LX0QRLfYvM108fuXjpHxLer4zUPtHHsmc+E/oCO5YtiQ9svf6W4b2S
OEVNL/7/zgxO4ibLWeizbtlENP2ybuMQPK3jey4bn97mDPDYLqiMjChfcaBpK5Hw+p/2tuvmcUpY
M4l0YnHVUrL03mvKQTmgZcKbAPN46eWBh+73Miuz9ZAJc2i+9a2xs1bkPOnYw5kLU3/bzVxl25Ol
Y+fFlhc17Y5sL7VbWPx1OkPG+HSzSa2ON9GWUa/ZZBhdOuG2hWob92qhfvN6h48VdFwfJf1KzM6x
bur9CiY8sQY1v1nEdqPCdkcSr7sWRNdWT7qq8W/AZmOFohtMvs7sGCV7LPbEkYkGEaKKyjoh+Xmm
7j31leTCd3zLp749VgbLqsEmZohXoCjGIdmRoXHLqO1vfW6jYanCI3WaM6ZHg/LONMU6qLzamDSq
7amxoKQ9l1iFxiAzg6LUeyzfjNOPsakPVAK9VSXhbJXxnLWiLClgDP2+YrQ9msARSsmU1OIbYADJ
mtHgNa/PFuszqv+egog/Jz4kcHeJ0qQyNQYQ0xccKs4hXuknZVedYr6WUzoKmbgf6MVZGrTsrjyK
H/abNV1a9ueUFNn500SGx2WZVyAsJsLe/EthS0sk9nZj6RCrRrzEOJEKpZ80/SyqURT85RoU14Og
3MpuKTbpK3E2U6EoCAJO44oZufebcPPvjwQUG7tk6reOTVncIdDoMgDxc7oaZuTM9pEh5qhgfGjz
SmZLV2uMyPcUkineF0/nsTgf67dqQqTmqZ15zd9G1dFyHuetWMh94SAoO3Lx1WEj8asSwm8bGVyw
OpCimhg9dxy8Ox+ZDWmP+pBs0sz2FqQd5qHOziG3ENiDSff4FWKPIRaBH1REhJxiuYoydZKSM9q4
16FbH8aGvUyLhacnLx4OhRkuyzlsKqCksIeCzh+3AEYG39Yv+gfdFs61e4ig6RK6znBZTD9Kjw+Q
rofChY3ph5jc8w31AePKqc504Ja/ChChYHnFl4S6DtH4rgfGtfILAiKkGyqcQJkO9Zt8RE50Zyi5
15deBKS4DfZbBkkMMuIdIzyjlB2zirpX8rViIiVInHPJd4aMdG2Y+nCZRGab0iZbjPP3DRAS/VYw
1lKlgKr8w0OmKu2esQQqW+LqFfYKg8B6PUS8GBgayPD2YFxptDdcLrkyFLqx8pZYJAHmWEY5AC9/
hshmBntP6GfHDUZRp/iOYCynzNaLfiYulDKM7EfB7umF0uOqApzCVtNE6utLXNDR/hHM+4Bb4+Rv
CCdSJ14b4xheQe0P2SV9caB5fHniH7eQwda9y2iJIS4RmjYeicKeG+M7G75rCGKKnV9WssTWZ0Wa
JkKlWcOZP8KHefN/59Yht7AjVO17jWHg97+H3Hqc2F+E1TFrtpEAexy5AQMvVl/rY+xchMVOZLGD
ksWPqJwtUaYiSHjbiKzDxgtwbs00fybuzthFi3j3JT+seYnivb9Sdz8OJVn6ko+9BHvwGZ/FrpJf
nMNZoVdRb9OIe+av7EqrnINPUgcZFlR5XR0/EAt5/Ba0X8lRtt6HNkNYsZfgVPiXHt9qfCBgdyx7
oT+4C0C8DdBwSooix8fo1XdyFSTFtGd9gjwRzPB2DPK95wPU/0ofsZ5LtlERXhr2bk0Kqhx5FEDO
m1NAZSnQwrFItKrnL4XuRGkelUSKB0VtAfR46Qf89OlYqZLpxzQy3Y1WwyeZ/2fH02JksdE4WYyz
tBjdLenX7H5lnlWcKNjnNIHB+ByzA8HglLSljC2+S6GfmcdMv43O0npkM1AoJFJcl4Wq0isG/WBl
I/mhYCL7E36AvEIc/N1SgNx4yMTbytBt1pGG4nplXe6y2iQRupYvO7B4OidCIElGHz+X87xIQ78S
KH2ho3T9zuQrpQzVUA56Mn7aPhhuU4XterE369YQUtfiKkZdZfEduj/TS5rLPwXIuh2+iTrstBzH
hvgCfzxT9cSHYgq/6saUH90Yn3JN0dxEVo6FsE0bRQ6FLKld32tjPvaayZcqJl1z2/ZNUVWMBj04
s5ZKgpJffZL+f0SsNcjJddKC2w5b5qTKL6CqKy8C5BkWBg5JElh5B4nKpjNlPpJyTUp5cWezYGYf
5MIniF13lX1pXo4t7j7fBsj/gFgKhvtNTD9RIdbpRyBxihRzCs8cT3YToLMbIn8RQaISdrUXoyC+
h0yI3CDkWqX2oSK+i8/wfiwlk5beDUQafi2NxCc5sW45ryXJrIWBirSfRu0GdI05lFx8keOWegpa
45afJSKUYf1U0ryR0yxqnH/b3uhXDRQ9ejYEb2D7NXW6/7EhnkarAmdnN0v1WtqUApesMy9xHvIV
N5Gkune+jc3yGf5Eh5jyjsN7I5eaI9fp06FLZ90WeSFqQcSji2kciyJWaQs2u3SKsGMdc9FEZgfN
0jW8hvIybDgxujyDkMd/snYSYs7tZBQTRj3Df+hmYv7KGK3aqZEMDkBbOAoTxfHCQXNjFRFqbPTD
GKZsFOnpJluqEAH95CeF4Ll+hAFsQMXW/Rku8SHfmkptoKRQewgPWdijuggQ6pJ0sbrAUY6SwxLE
TENcj+mL6C/pbjrCvlMGZVHB+t5hWKLNUi34XXypyrhNnFtUKeCbvmTSqd94nczHzK7NHUjcpPVi
HQyNRlZQzMfK03nr5VGY+ziZFHiTYKqvTClVfzgBerXnrSNKWMslEvtF9I+JUaRrx8szQhboyLk4
RhvofW40h0um6PUNznxOIJtGfJk8yH/7vN3xBJR/qThiAkHVh0X6fjF/HDSLFMHij3ZtfEMyMaQd
Ir4G3OlIylB19kDVm/XykgzUo6tURCZW4pjCiv9eN8QnX4/3nC4lUQwc3S6F+JS8+EMaimkBYkh2
ikNBsnmJZT731KhgH4WVr8gxTxM7BwgNKdnjnc33quWUcZzwBAldAN5VRKzSv5uMNynKhlerCQfF
c9/A1k+EYN5X7sKTDexa1HZypDIBzgW/pz1sjaggo+U11dja8WXXlGIWuzlwuxMO/iPTjGEcU4ib
ZujMoT4vHAbCwimGJznenNBzGHvOIWJqU9cSUN9inD628KPiXIHcyTXbN0FCrnOlZbJglpeGYOT3
TBhA3bm6m3X/uDjAJMgFnZVrZS102Kg4XjjywAAuW/rRMkQrL6N5bJqarv3nnNmA8aSy62koUM8J
JTnN5PTcotLTEWx0zw+uwQ8LX8Cm6gjMWiI3tgimCNd09rMGdfyjpjdJCP9A+YXjqzjxCsIX2s+E
GHAMASLZohI8F8LEtgEM1RR/XORVT39iSiwbY/woutsDmGrFm6OwWT5rpUUZiV0NH8SSBD9047mV
3XFTJNLTeo8k1/LNzREuzguX89xc1kHQRobOiDiOUuqiDgQxNv2TM/2cBxtt/nHShthyoWCvpt7j
SPtjfuMUUiOqjeMEFvrcp6L/mvARpTzTOY9m20nCsBdNHDw+55BvJJxkVor42qoJRvrU+TmoTx63
KxeDf5n7LNwZLbzBjuC4kVvxOfKpvRbobJ8PJlUhV182vX5FowbJf2Mc2vUjZnmAtZpW2v5z8JfK
N36DkEtM7owoq9cAb6DjgvO8D6/B4NNUZCHOQm9OE0EEl5FQl3loK5Bbi1cPws86nDNcLLM5uAt9
rO+f0ROESlR5sJhhu1EjLJyz+ITAWKm5Vfodjd0bDEswvrG2OFIOCbT+jPhybyo2a2pmmQphfwf+
pYpXMdU5DWK9Sy4dq/RBk/RrSXO/Rx2XcOpkOuFncdKYkgnmjC3cLYBzLNiho1F+y0Dk9lLUe5jQ
1lJtiRSklqtFS6U+esqBVqyhPC1xjML1UyVxLCadGFkKPUyvEcXQYCxbrbyDygVezYk0gNJ2dPIY
hc9GLcTMBs4o6sXxPqedZ9vGLJxPFe0KIJqK0YkJ/c8Z367X06URIJkGo/f5dJO8GBAXoKnrraB0
FvXUZx5boe20fdDNe+qIkJKjD2ajRKwSm2Y8JVBw/E6RJR4T7stbIfsZdMH/JaJune2pCMRS4Wh1
QuAUkawCWfbYOwZCIlSCsJKaekFs9GIDYM/uXywCDQTpKqcNVTJg/V2NlkoTT35iTQ7T3PMx08w0
GVD1+Ao/Sfx+1bePjPRahpvk20RlDTnB5OSG9/jxN38qd6m+sZomZDUoDhXyD5kzWTxSB5sIw6MG
upqBB8GkRyuqMPbv1valdmbVR9HNP/klW8vv8Ie2+w/1PdSKReGeNFIImY1EmTC2flSiG24pFU/v
/dvvIpWSxmlb7ueN50bkARyjS1znuAlqcGcDxJzeT7Xjjlb1VIhmQyu2apsd7XXvPMYRdZcKDc9l
0kLLJr4VvZr7x04ZIPFzmURGJ24viSCl0LEvg8wcd1+9wkYeMLzYe88CmTPcHMeI9yr3Ikzdp+9h
SoNoKXpZhrfzaIP1f6qgYgkpVziIfifAr6GT2YYjueAmvL1ehonNwgsyXX0UTENn22IlOx6nixVJ
Rlbe8lUJmqqXKQEIRnWAd6MAOoF2aM8DTEvq6AEuw0zbN0eYYb27Kfd5DiHIWHubNQjEWgoQsVZw
yq2opUFEOx+xGDTSjb/NxIuz+Ah1LdfdoE87a/EKgKVIoB001fOBZl21/VIb50+cNHweyjy144Kj
U9z113PHyKSYGaDMzyVvu2V0PdXJkpXTMTm50RDLfoo4wo/SXaG79nghlN9EuVP1uyr64w3ARwVS
hrFcGZ+iW/8stLNGze3dauIcPqx5vW8ChzmViUv9Ua8Q28Wtj89gksrHy7Ke281TCGFmrUH3j0mF
xyvuYh2uhGVO9Mcr2oAC7oaUkHyF6X38o1QYSoXKniwCpiuutkJLY2+ivjnE2xiIgtDx27Sof2Qr
4Ig3YNBT5ocS8JV/8e4+UEOlaVnojkNAzXLQFRmjOO+r6RE7VcdU6eqdxtbHDoOFox8aLRYNuCnr
kuivjujuwHmxqf2OQR0PEcuTNY66q2bkyf8WxB3OXq77OYOgBzB0oTAEwze9rb8Y3T2wBEqne2AD
j8v6bB4zsBHRKxclHJ9JeQEJ0R+M6eJoqyRuq4PGSK+R1zlrJbVYzMqUWbxzgN5p0geacoVOVr0E
UYRfYsTE0dUKFMDH9PGgo7VLW7KCAIdMupSLWPt3i6EjicTeIUJH7UTxGDgYdOjKImk+Eaa6l/Z/
6GlvxHwOZY0X0GQrvkY2G/VNy3iVj3VmW0NntDOr65lTdoKRBEdWJ2qp6x6lTEkitP55BJhVBggt
D7p/VRHQ9IVgkju96JscoNeo7TiZfHu3CcBix+CL4eU2gVefTz/SbC/8Vj2dakGOcn7X2YN6730b
rwciqY6uklCsl/uFRAU1YnJ7bJPGGNiiOELZCaAh1IrvlY36hAj7AiJrUNLtPJzHaNQ+14AjimAx
6ErZw71K6tH9i2f7kEZ88lkQkIXYjW85NNA51IzmhzabvTPutRvM6Lo6PBLyTVB09MrhmCfW7Fp+
BJbs4hskU96IpqfvESTsg9YWeavP5oE8BaBFI13fuDc/lJOTyykFEgAMvGYVP/4zT/9SAZ9IHyb3
Y61LRlBRGF/p5GasoC8/uXMjka1905gCHavR89wFMV0Fq7p4jOTLYnCqlytm/qs5vQto51WG7f42
qU02t5ZBR9xst+vxpspP1VKR7whwwfJmoL3XsBrJmCPXeOdMZLJ3IiS1wlJGklmtE6ZrXZ014ZEN
e+CGDqMtK2HP2dhMZ94it4n+SIHLyA2nmzdt/Un9o73Sku1x3kgHNw3fpVboYloupZz5dP11zrQi
HWYoz68oiKU053QKYIPwxD2i1vbTKpDXKVwdb9UTMZYCTIonmWAPMVvBkU4wrHvDt+/uw8awNfAA
1OIZzAD04W37m9AZadqNo58cp4qJjg4kEjHdy02/zK/8XUutwJ5BIz+7Be4BXgrZYqhiMdKnuHN2
s+qX6wT8J8sg6CP/EbSKSsrb8AKZJ0ho/2T0aBklDjAU4mMZgFcZc31DjW6oFQROEI2bBsToWf5Q
LUj4aQUjuCCl60Q5aCejcT4q4SzHwK8k+lOVnIcherkhP8KD4o9MYROx642M/bfiCgqBQ5u58buV
eL9pl4kkpZ0bBIlgd0uglcIwgJcuJ6N4Ok4y0TeaA853gAd1dokRXPjgRRBW2pGMjRI7BzH070SZ
1NxYjVYvh0WU7XCyMWP5Sf/vHott/FLKCF1w8sN+67BSnzKkkitEjMhhBI1k6/D4hHLDrtCyP92y
JDwBB8mH5gXZtuht3qduituCQuDzW3VocBHdcQBGpKXeu+etHrPSmMf8qyjR8DSKwkbsdqUtYmGl
PG74K10eBLzZA3AHrxcKHJLGTW+l5BY6YVJjo5GwpKCNjt07HrO6SKH1qLTfdqnLqnpYUBVmTRhh
HTFUTyskEvvaxWl/XGVR9eOrBTaDVe0aY6eb3ZQslVWNAIEcb5x3qK7aEXrJsCfJn43FO/5kul8u
ElIT3dd7LrArN+ME3MzmdV+Bpskifqg/QJ4tOx9rGD0BQxVpPoryoSDALQCzGp1/5foSP4VkF+Um
UwLMRSU8NJE7O7ODpX20ynLk33FDoVZ0EV1giXQSYjOKEI4GiS2iTlW/qfgCi8O1qkXzVD+oXnSh
BX0qnmGJiblP+FJrsGKvwL2YcSzVO42XWDkdvRSdSn3qCRLs8U2tFhU8xXTor4LbxRvNL/bWI+ma
3CtE1qyzlXSncz/iJTIWRbCUEmo0jSe7QEu5dPcROG+8Ukw5Lcz1jeYyJPfwAKKjAZEvG8Y+ym3K
GT6NykfUJCD4tr1wTdm0egwI/5q3xC0vTzE8ID60aDEn/2R4E4ffhmK+DHJbMXSCkFSP9xHmWnxo
CzztCjILxRzaHlTxgNXnLExswDU4cCsvvR0fjrXR5TL0LHYgBp5+TTYf4/WRvSNfkWnJ7ACgFlAa
bDb8/ff1a4yIQvY49FDx4gMc2k5HGZtUG6fM+IZRUUgL4oyndPsB/fE6iI/LyHW2dbQSgFlYp5WA
+POvSEZcaTQCJmycijnXRbMKbD0BOQ82rD380zrzKcjj6T0s3AUn0eVdmgZNaRktldhC9XSY7d08
DrtKDLUQVZ8zjH6q6+RdXESMTNztYCkOVCixDq9IZElRbTPXvYc0aGPN7HADx3oNBJwzltSIBYFu
xs5dBtGadQkYggp457E9ghgaEmdD1mSgdSXUWuEp9+pPYjh+OIAl21y+78Z+umvg3Bfyfz9nVM+a
odgl2XMYPyGobPMxZbOcGXM1lEqPGkS6onRBx9kRP8E1EAznL45zxBiQ1a04ucyl/Iz0mfU99SEP
7bB8WrKiSerd3e7QGNxoeNvFu0JJEGMzHsMvYabwXnintCfTxjiOXqlgdUrgYXJhXgt5AFjZBKxI
WzZP941OCEap6se335hsr1VG6yvzoJM8aAGumKh0UF4rQxt+aiY1gR2PBgpiCCq+Ii6SUJRBdBE/
PO48yNfAuDqmgNm94BXRnPmi6ZiAdi5dODUxJL7Zu0x8+1gSpaxCfqphpPmT0qtQz06XbOGgGQiB
fVOsIxsYA8sHR57o3CJ2uMpztjDJD6WR+sqXT4XcxEvl1KwtUKD3QzXGQBekfs5V2GHNqk/YYU46
Dwf6iBdgaPQ5lCaJNzRECTNZdifXtXPNewPhyBdS+aodzzG3TbstzsfPdbtH+WNFebP0dtCrlZt7
ANK12TjB9zwV648U5x5hXCubdbHhQpnxGjMYLCmkMWj+d5r4/8ro3KM0hn5uBxH6zNgPjK+IduEt
NFH1sWPGEaNVOytsQEBPCM8KEjfinb+xMLK4LMwZi8OKF6xDCpdC6cnfGDmEW8lU2yr/FwdpQjCr
dsc2QuokW8SNuHxQp3euAfLTWzAnrrjy5R0Avg3hjigwWlcqg4JVaQ+yIZqqrPaCjo/rpCCzRiCg
PbYTsD/GXG0bI8q1qcVAgeXHDcWETlT2iNWeMis7G1a/UetOl4fN5NlI6FAWk3Ar7sj8F5CjcqAa
+WfmYtJyyCda7+j8xGE3wrfIjBk5+EPKVsdrWc+erydMOPmXF23MPBdhllpZoD7wGiv1AEvds1M1
JxUGUE/PJjn9v5BMJkvSAQGdtiHTPQD1jgN22TVH9g15DV/vj7Nf+LTKWye1DXDJ6J6n3HHz6Da5
btUw+k86lgg6pSsAqCkStZxG01urkdiAEEthDS0WUDUUfeqNysHrstHzpCTICJHHBUn4u9KvjHVe
iuhLhJd2QVsy/8E7Mmbrsu+fzfrASUoj3DwO877TfJ723mJHBnPOhH0TEvBaFj9WzftP75ottPSv
nCTA/3ZD0NFaxCWekKVH5g3zItCdmTzySkKEebbaCZnB4Hn3m58NHdRrbgqQzvjgplum0+IEhu/u
MPgmcrz69BkLiIwmtfjlM8qnusGhB2rECTFqtU+LAlYOJlhNNPZBFsf4Rofa4kvW4wGyV2lE/kpX
ahHYK1yhYFNsoEY2qPTi8bI1aMXDfQSY/0U12TOJmqZ8jN4Ui5rgrzAnT9Zm1N+yFdMlrV5+dDMr
67uIRlUDVSyDWi2FSOPXveCBehCArT6oPOeyx3hLCvyDJcTIFBqEBR/h7hfTgeaODmhSqHVms7k8
AYMHE7aRg5xyKgLd4lvDEPjLjs4gkmlcs16E6dqEKq3NYNWNPcTMHL5qaa2Ed2/JVXc/DKexKluy
YjgoxkC97PSKu9mPXUo+PXUzPVYDoBPRpcHxM+OSHddBunHWgYS5aJrXCAdsN/AVjecl6QykknHi
PHQ7ldl2wkR3bfNbYsV3AiHIRWuf26TjTlASjEpXLvHxwgNGuVcvhCRXGOXEvYazW/SvhvzeQa3o
WUiVPAs+ciuu7A7XucDcC/1e+Y4ol0TvP5chMt8MYpanmJ4HfKqudlP46oYjR2rHve1c1MdHmbDY
PGgqF7MZd/lEPwtTL99BRxvMJeoDSiJWtJhww6A0yfyIczHCAt1eZLnhsZnHNriuQimM6IXmIXmQ
HlQk2EJX2ihoqqsYI5s5iPk3QBX+9RnfDzw+sZGsfixqIIZn1HYmOIMeV9q2cbMrNDEZ+wQmPVlH
n8sYRdwLUIW4Avl7vYfZApe3SUGC5em1ZMEwt2jQSUQDNatMzKWDkzEzXOaIjMYjxFKxE3W2d8qG
HYVgLLCQAbcBbcLb/p+yEqY4l5dFaXiu1VnGvCYgXSeV2Osmwuhv2m434B7/OoDOTi858vvI+mQB
xSHd2OKOFjhOkBJaCl65Rf+irsfCHkkrJavzNtRB++MhD9UcWCkp3g3rX3uIHv6gK8RmWvdDOLSu
v4Bngsld0OmHMZX12mXNy0I7cNVL2T01WRFKiCMOKBI5I4sZyYqwi5fvt997cXe4AldJrRJ3p+hk
h9t7mz1yRXiKdczG9QbI2bGCHLa/b1A+RC8BGsLm/rzq5PuAi+q17v8tlei5Fvhu24AXlfrqO1fL
AxGDNJe08stnuoe+SQSk9gZzCtXVSkjoVXlcrny7ryKSBNdjjSXp3JO2RjbVv81RqqPzecmifUQV
l8Gswo42fKTICnQ4UL/E12OwcmDPoqeSuWWJUQhfPSgsUdcqCjr01unwkT/N9cV3saqsRzuMRhjN
CB+crYvbMwwfXQ7wgQxexf9tn5S1hrHs4lfAQuIMULB9ROevqgPYxUfQ7uhYhVO2MvAPFde6QPAx
cF94iuStgM6XgVg3ou+n3NZu9MdO9cF+oEvRPpUTONcg+hrpg6PJECjAelYODAEI4xNgYcXtJP36
1yOA0DBbinzY4Yh7ccbCqbFI63FXxoiR2UQO+9Nasbqn4z1ifxXCxXxn052sE4kiBEd5XvI2DRJW
7Wm5V0bjWXWUCYf2UATKGL6uSPqS0GErUHLzdBTXZm9KmY9ZZMPdOHVC4lVcSA6POL1VBT0/byyk
WV6xkSw2+0QXtUWAhi4OmSzDYqd0eymWECHkJgm72fDuUillAb2HN8PrZupClb5dDEL1Tq2g3Iwq
Zc4bAlX8xvUXSSggjmOr6CcmOoQAyGYUEcWB4KCcNEb7usEfekoK3DbJ82RbnMz8nTr2KNI71Hjb
yj0L43b3km/l2bi1okag3kxRlMPLUg+vk29jQmlIfxyMBU/baRYPUJlxxr5dOT+LrmkORaOEQmqu
tSIjrEYaoAZM921Fg5vRt77B/67TyMpNpIjKi5VDjxueX+WEfgcR5V1V+NM1ilwoFmfIry0uJUGC
P+ziFy/y1Y1JSzMxK5ojs+mrmGJlv+yTN7OF8vKDa2nUEQblMkiMyE3KYKgauHoqe0UkW4H9YODL
kO70WDduREF3gvK0lJPjopys3tFrJ49krkWUUwNyOzo0daNOPMm5jGh8kTKNzxLV+m7Pf1Z0W0OL
KYRzE6cgoTxSgIctIlqPhWK6ASmRnIfy7yBFad0bNlbPS7nylxymdJ8ekp4zfclQIfEZ+NYnZZee
RJMs2Yo2h8G1CUhbiYkI6h7KcwVgSwkVyMswiI+Ztq5Jc46lKV6RzbaIN7mmdmw0J7gIFY9c4n+l
tQyFlSvdrJUUHLCVlwdSriXflsYmJgxgC07mOxLhoJEYQSQzvEyMQvgm1tpupzTPgOmOSUtHm1/f
bvWL6tjzeNpAfPMUcp7yU7iNugCRW2mu250t98wqL2JK4Sk56FK0ESJ/AUERiA6RzgkG3JsuYXSP
/zBz1+fD2rtyO+MqTR+JXSuahRJT04LTn/0DcmkykMFlEXKh5Inq5OwwhWXhB8n27yptJ3u7UWsZ
qKZ9Z5iisBko5kPbAsQuNtkobjpcsp+mllXfIwKH2ubXvw3p7/7TU/y4urUYDdbMrMUlbj23EJcS
GtwxHvAdL09Lgk5E27z0TNHsTJM7sgdPvI5K62sllUX66VT3S9ZW3nhi+6iec4fuLVNpP4nJg3EQ
H87O+3h0XzkUeMSqv4BQ3U/XBHckwfmx15Hjg9AoImeGKmFVqku0y+QD+m585irl3OxKUVwseAYX
b+lOOBQgcI6PjXsICOgN7lrNAaOA97eXkvoxXdKqux8OcMrTdpOc+V1oIbe+VRlL4GqZrbpUYA9p
2wpxO2gYLMxumOGvvBIYI2AaZAf6bV27l2gkOFbRUQ4bRKce8MNqcgm4FqlEWoH1RtWHh8Ul2ufE
+gqk31MjebVCjfL7dRZobq4gMt+TWIebh8xWIFncH1t8mejmYhBLW+Y3yCs7C8wEnJyrhXLHIa5l
YwiEPvfBkS7u6Ht9D/fMqEqAHNd50gH5pdjCFeshqt+rH83IGP/Jc8dOHN3C1uvQatp8xrpwQVNp
XbLij4UrU2K+aKB+L/kKBdoXyDvJ9fY0yEi4lB7lZheQRQ6kC5O1C0pAMBy35uhQeHzJ/7qT/ufS
zqkqvtMueVqz73Q/pJV7DCXNUZJ+8PZwF0x6yju8lqkfmClC1VNZhkSzcYVuNjf1UoPrUdOC3h6F
CKN65tbCsD1zlIwAf5W+li0WYv6+859nLMisMI9RhdeUkrE552KsmiuDA9Cpo1Tzajs6QWYAO3o8
pxD6SNqpDRBfKgbuk5Z8tpYXNPsOEfbSX1Ho1vh441NRAhoaiff0xZH2xgRbdj878zcyXzVxTfz8
0XDP/yNYuhcTj/qKAaYL8Y/aC93vPba/mE2KQkrtIA8gP04NSuIXtNJB15CqvxdIVDdWhzhyWL6O
4KLCkevc7JeN1dzQg3y1OjhO8BbpG9q2dTGA/qFgCCJK+Ad/W4JjtaunLJaVTpAgbjGmhHGq/Xku
lwoWH/yHsVPjG9fvuBuVwwG3iMt/v70j83ybDhWjcSXSzTCVz2Y2JpHPubq2nZLxtXoAwZOzDijA
GaalD69pFq8Uk2FyBXUTMbjUhHj2jrEcP/Wk7Bwe5VmhCf2kteZKUsHD7N6Rs3BwWZU144YhRSlT
8sggttnKpJ1o1+1XGRANWPclHrVTblZTbNSbYVaN3EFX9Awqsvrt9hEPEekZYRz1TSs0n+xZNkUV
XaEXy0s3dQKmtHDnfzwEcMr7zt4IakI0PXeSVAiUgztFHCxXOZkF5gGEzFsNRLBS3lIuVEOVJZnz
p/jksXmHzh5o7PRBR38JdYDHIFFsP4NcRieknZRshY1IhXWFvg5P0swivpn54KBB0Oe2u3llXUhK
nqil3kBS8t2bxQnBNBlcJb8enW5kCkeHXLzkmYmoX8rOdBMOX+x2KW4fU+w7jcrwSS4l9prI54IN
XhJwfHiZbg60vbM7P32sXgMSlTFZ6uOsiva2f4SDFuzLsDVe6bG2CPgy7V0XFhB+jCKd03998AEG
MqDRp6JERe6PxdurmNOoOQO1E+dbzx67X8MK97mb+7crfLNvFT9gVOsnAfBQ+xBqA78og0XGHA50
MhSU3jgCemsmOC1DKyIqrpoexh67ehpxoB1XKZrru9H5rEO3EmKi7or/aAzytOgG3MfL7tFQ4mp/
KBsQOp8rbruS38iTA4zvaiL3HUAhoNbMUhKEVnVFOMSG2qy7cYoadnYivkZoQXGitxKrrdadvcLD
CZh3kYvIrEJ6FV9ip29lN9XKS5riYCTFo/BZxtEc8dI7uAVxP2E+w1WJDE70Yvb7be2uG7RPvja8
np5X1dtyS4eL6XLrNfNGLGNvkSloiXFLND9ShIt77OP34xey4pyrQPZI6DXsRxnRl0ICwmJDEo8N
/vwmy6SkkyQgeB4hgquna7BhQSiMrw+9OH6MZNJOCcX+AcFI7js/4l3Dp/Qr1t3D7loh79dlSJlr
Wt1zkoLOKYBQ0PlVu498kKlCHbyFN3jk1qYJvYPZzaj/IXFjhHPsu36r1OSvIG5HtFaXDsKPRLMa
KflGzWVjgZDzSMU6+D3LfbfUjTZ3aL3lDtRSeymHx3tqr0hecyV/KNq/yOttpDuifnyWVRpHYKEy
zsB1XB7H0sUmcNP9grJztISX+k4S2eK6fsVi2MXwykb5p1ncLdm3KKCIJDWBQHED8NerHVc0YaAu
Ixbeqgq+2TWavaApGjNOj8iMROFX9oYECfqZOKX10oAFO6DaDfbvkTZOfhvx6jm2SYko04VT0QRv
n/xQTEyI5b5VhzaNoCGRIjIKsyPbP7xUB8DvTxOUMHEa0pAe52zNAHq3VyfkF6IWUhj8QUMYoHed
zC0VfkrQzKqPSoEuC1wFgQ7WXBicovq6zEEEATq3qDZVsJGfovtpT6gFmWmfnGdrCKhi21AYpMhs
BErDFd96ugeyUNgipHiEPMaYwjepKCbg3HzgwJ51lRPjhb6EgLwEyqhe44bOI+Gq85jHbVnwad32
rBVisFuMPNFgkvAXuVHdXrk3hzclPaNtN1ykhBl7x65ODoO1yZkD1iXDca6QXjZBv5pVvGLoAfvu
tXdhebYUqNY4UpQZoZojhBTPfyJSfGXJcqBCX6MEVFx5jKZ1EXYN21pgTRRWENOo0RP1ssCIyz+C
sCEv5VYA/aU/+GcEzoWGFLpI0ixXfbfL1XGU/FGpSBw1S/a536Wav7yIQa54GVu2MIgRf//qLVX1
bMZOmch7d6Kfhy0mT8ODLS+hOCA47OQ4WGBa7pSwHm6ZggVGM4vE0AJVrQzcEHe0rnKi9aYDuvDV
c+WD0Is3J+8L/fzVjUMqPaulwiKRZXlHPapcPhI4vJmJPnuohc8E5Vp5fhB5AGEpfL5+eacOJEED
CH6aX+SXXZhvtf2TNuEr8frwmE5mdMHngoKzY6aEWqUGaN9jdq5mtEOqr0y5UCUh8DlVwak2Ep/K
Yff/zuf2mT2igf7xiZNfF5MCMzbxgr9FMcevvmmrvIGnP/MmGBkFPXrBoMNoeER5gV8u5WE/3H3N
4hHIk05LhbhGx2flYr68r670MRB02wi/a+qJ4EO7YwEYGkKm5CcAlPq9I2oxJWz7Mtv4UP1AKuMw
PkZKH0KGLvFlhq32UmHWa2agh/eg1I+s99DYdDtq79hi/77kby8HO+F0otC5Vf7aI/kNOzTKgD60
ZxFchjee7UjkZiFH5IzvgdI1ScSFTbEuQ60OBqo2KK6U7O79pfGN1BnVTuoCJOQjsssuKhKeVpde
vQPWB1v1kSOyzx1joxeja5iCEEB8i+LIO89IczpdfC9C2VYlNSMEIbGUxJZx702ZRZZ4YwaTzYe1
Ps+vmit3s60ADgaCYUTujS3UNbRRjzSj2dsqstp5Y1CwkMUGoUyu91cU9plIX+r0eyTmdd4Ui9CV
+tRW4rXkzptQJo4pPi6gIcd0iLY84CE4hjiYTJkD3dznf4QreW6zAoS9+8fQ0IndmFldGQp5Kejr
7fv1X6eNR+Nw7pVfxUH5nU3D9e00A6FUUZExvK1SjXcJhjrhIf/A9D46dfqLKRt2v7sPE1F9SEVY
83ObU1yiId1af100oFpir8PZocN2xXwL49u80NzRpqVsYJAqoDX0b1UlWh+F27s0IIR5qcdTnH77
q08x0Jso/jYi7j5u+Bq3yXRqoHR1GgHWcIzS3vq5/x/JX+712t1RXJebFvGqKaKfKd8N5BhHRAEf
DeFwFwNKHk6uwxfBaB3thauBf1TBaUVju2YpTjJsKeY747HiX6lvFOr4fQJaTAspbR44jELTQFgn
/oWQrLUJmLHsiFGe4FUL4S/LSdvmfF8rrqfSLDMfCE1isatPdLdZfMTotK3dXVEEkwrUN2eL4Ijf
NllSueufHb2zaN7mOGNDehywatnYPwweYC3AsSKkwAXRgaTaGnU8vdTNNGSKryzqDzQOP6+5vgOc
ct1a+XeHRadYkx7f48JlZSHuB0k7NTrZDfS8gbhyInassqecWIV2ZQrhXv3ZDT0Yv9gDhXRSusDK
iY7Yk9NwB+wr6gJvItjTxsiYBqUJ8+D4E77bs5zzKnDZEVIT/rG3EEgB3qtASeIawR/tH8g6TrhS
A7k2cY2tAoUWlCb36nQGDdBOdLW1SfkIVYwoHCg9oKTghYiLXhYJWWRY2v0Xq4/a8J5pnsgsoqxF
YHgcUkSmaIa75h8eo4UNdXevV2rnsHNAEI0AP7+UmJP4l6hTLvbrDe0vs9PDoRWny+t4YaF+ENv4
6dXlgL1tC9S7PKGY9IjLcKkHA3pUFoL+C8q3mb0umXlKJN3XxPwlTYBMRRtdWouHLscfdhexhwLr
jtUcPYUN8wrM7ixWU8G3s9GeGmhoDb+Uq6ba91fCya1SqvtXO8lG28vsddGLvfB3WLe2GRLTFvyU
Agjp846AmLqX7YYS1vi/sXfN4ufKtZgD0ezNYnr2nbpF0JbCOB1TCbM0FS1Kcz2oZPp1onS+OUCf
y6ZIvDOyY7csnfOMUvmAyTuvJ6uaT3owIh2n0fUbxedc60EVS4wSxOilqL8MODSvpE6QjkQbq8IC
mlKCd5zlZmI9/P4dMs+mWm/w1DlYmTp9l5pLs6oyFuz8QOCJEFkdZ/ve41NE91nkryvcqdf8QIz/
NSHPkZzpSDl74y9FzQurRenBq7TTeQWzCpiZOjDMIzxEzSj1XIJU6zEn04QYOWQbLbSyQimoVXay
sDtpCdyQifHTCII7W27JD0L8rQugoHjVgPzdetpcdf+LhVXcz4d1thNuIgll+7qNEi38JEmxV12U
LORxVOsiILnwQTD7mVqQZofrwgXjK2De/vCaVRpqUq0Th0VTLR/ygLItqQtwjj/dwwVsNScS+4IT
lhnE+vHR8u1GutdZLRjDrgXWy3sOANHOnsVxL7SjPH86wo6ZEvR+oL3V1C5v3RyPJkZM15tKNSJp
HUIJ458Nhf3a3U2Uj/hn+qEHEehzDJ/OOXA/GnMuQunLiS59e6qfNOhyNmRahObCb88thSVdubWt
/av3ngURBj1aJo4B46no3l+jzzuqnnIH38LQ5yZMSOIDuVCXxWDeDUM84efh/HHu5YUFGXkFIb+3
oLyzS5E25J6dieNwBmzUK4ypZPDVBq39plEwJ6EwyZCblNNFLjmeitjylWWuPFXCQntGhc4NHVfE
7NzExA8f5K1SFhGIc2GkD7UpoOGs4qrSym+RdStNyRwM9vWrqYKotlNV0iHZby3heJIPgXWU/HoB
f7zjzHirfDj0k/xaFqlaEQJl0msD/RXJhlH3LPnN5iKdwOIOnNgv/idcYwF8Biud0Z2GM/1tK8RQ
LG41BD7vzHqQw9YTyQjkekXarVK8QP6KXyGk05Ro5PcFy+xRnESwpL2olQOG2OyazYrQoqBOwqxX
ZET70+BJicimoOSA6WLuvBkW3ymmNQuGxX9XWH6w0E4NoAv18ZJrcKgMAHrsNu0acauaZozKKavY
r79bIB69EdPCjiJfQlyIBcf78NgvRHN4VD2U0/vqQ3ajmERIP/SpCUOkz9XgB7tHTId6ze4HcEqr
t78xUA2jhaelumGqZ0wqyz+30py/ORJPCdOfz11g1lKWb67NA0Su4t4Ag4E8jhkkxnlnh5SL9SkQ
2KNKtOnUTD5PKg/c5u2Sv0Ft48o48Fo24QLj73/flPqwtcaQgoYwlKm4vfFpBmXRVrii3sWY/KNX
1wlvpbPZQfTl0M5omW22AZJlc1TzMVkGtgqQrl6EXs4Mt2dJj2ZYIhj3JHK1PnVvfj/n89rwJpvh
CJRleBAo2WfQwgbYlOC3yND58VXX2XEqOI+MBs8wNCKirAp/Aqg0zwyRKX4Nll8bnYhbZy/xrxjp
7EH7f+issUTGSwJvhF+3RIN+Il6qyrKzRffgQpeivQny42oWKm6qzVfdjqVHKbv/gE9GTKQwddh4
LQ/n/bfGZWFYf3R7+muRiqEp/kQGuycTh0czUf9K9OkUNZw8kOZONU3u8zSUxpPbd7tx1wGp4Mw2
QHrgXjiIf7oXPCqY8uAFdDIxOeDLwXaEToaOxvgE0Kz8nY/wFcmHrhfPEWLDl68WsIMjy5FGfFSX
sgRTKCuDijCE9TEX90FSRBsTkZ2vAEBCi1QVgOdU1NFNHONUXGG28gcUzbo4s4aScftgurx2/joM
nMRVj8HDsrdcf/n9/jrCjfAu5tll9q24HuzHwbpCIIX5dbzUT+pN8vNn8l4XTYNikLLALNmsC2Q4
mMX9X55wUb0o/H379MrbOmeaJKPdeSd3oI7yYJgToHgNbFqzsrGyZYMQxNqBN8r3+qvYhp1ADKzH
2IBQmo57NmzE/kMP9p0NR1lUoZGQruTa/SibikdNcVjKylcfCFWeAa85bPN/M0VP/BbilbqsS7lJ
h5xBz5QBzc//HG/Eu6C+d+xXQKiSSiz38f0xJKmd+2dfh/Q/TuR1dOk0jgb62NRNpcD+ivrCoLJu
TbYqNbGa4xDrx0/SOK7TYEbYIVs71Xt1jSJ1WQAYuL00DDs+iZ743t0SfU/tnTdOqe9KxZgeBlI2
NBTf+wFUOFS2SFdeR9wxcnEnyut4wVQuju8ws8xSU5LyOkUOS1oK0cPBoP4skEOFArytycf1IUOk
CQuKc+J1q43ntkfJU++9ipZS4NHYHw2fm4TWpJ74z4XQ5YyyohLcbfUuTh6cCWamkvlnDAlX3QQu
s7jU3NAmM1AeUxSfZdWkXh17JVnAxMp0hfWJ3WTf7NqGHi4WxgF0rqfOSBKKmOEzhkaFML8veVPF
M1n4WEs4FfsaPZBixH7xyToePhnCx32sX2Q55aM6tynoXVNZEuChAXj/0Bx4M/WxKoYWXAG0ZKFM
aSc67KnRFmCW+oPePdFWMogSFthILu+8O85ftvfvqlqdyO6F1Er0hYq9jPiFrZ9dI+6V4ADhOjlI
OLXhzAHhOiINH1Xdlkbb3gecmFXBsj7uWGIrjBX50qws3aUCLqE/ObTBZOZwIwjTFF72Z4082RK9
WIMXVrOnEqxPzHOWqdxgf3kcFijh4H421Gi+3vd5SUe9BJBlDrKANIPkFdG97pY6OQbt+F/VXMoZ
0ulAvl7bQWK6X5qLJUQdDbg2Vz6WS4fyMSZFiqjZqllkqK7mXx2BLN56ELm5VPV84tdVn3hl7mGI
CsqcUiPoiNbToL4mP1SW5GSkL/on9YutTD31irvgDl0zchxW17PRjoIdqd76W3cJO7aemc5nJ2ZY
AsJYMqoOCqnneG1TCPZz+4Amwz69a6TRfdhOwcx9Q5A9UY6HPwaN7DFpcldjmXZ+gFJpiEaQen3d
jNi+2i9OqxPFK27F61bR8R/vlG4tuhfWOjrDq1QiVQ0GKVg1ztg6S+lq/L7tpTgJzwPjtIPssCmF
zh4eFwyaZZNvWxtuWyXiyeCfIxNmGYa2DHgYu5fu21/CNfUeihiwCs5Bsz2ND0gqRQROYkcAUtUp
GKeVWr8JkbwQ21uxvGzuhlni9KW5e8Kmz8eN/Vz6NJ4S9GohuKhRtv2nwXcZmOAMWWUemmM5xl5L
TdzlTTLdkvOkIObKzNFs0gZ2syOH1ohnPe3Q+PgU8FN+kMckmONSzEpRcksBEIw0x/LuvVq+7zcK
VhbGJuspV0cJdMmC40KDCOxhAwc/DWpHI8mMEH8kQAgktvT28C97DOUSvzH6zurG62vnasBPiKOa
KUSUO27RDnzWbjkncan7XtKbTqfeGyfvXbV9LOxFCOfZdk7XtpoFrqjQ30jXfY62v+HGGUEc84QF
AW/gxE6IWYue4rWZxdzgMgVdDaFstq0hFLHtGf4CkH8rq1fSjrB4dC/RGconUIem3yXJZQlnWVMT
z0qJ39lgxw46/h18qnIpbTviaRrHdY4Sm+rky8CvNMi3EsD8SECi2bGqHINsEi2Fyhc4nNTBuN9o
KY+Dk+TrnEcwbgoxU0naten8rTUeaNYom2vgLZP+FshKfP9r5kCX8Ga2Qq4IBFUA5aMSiPqQCz5m
ZH7sCvNlno+AJOg53qQVrWsrJ2By8XuYfixq7F/tUyyOuvtKIEl6RXnFaEBFMzpco5r5tK64bcme
UYs71z9FOZaxN/l6fTandjHAPLbxMDeiqk/4HoFPoNaw92EHISsKSKv6xaUqHcUW4yRUYbkgLJ65
D9bFKA73mfX3KGCCsdrxwdwUkYkirVerJSD7YTbJgXheg2pFypPCgYl10/4w2wc2zXOJc6370RvG
049bfxaGhv/yx32Ax0F1wgioz4z0R+4PHxobV857MXWXS5S8Mdsvij77B1yOkj+moJNujA8HUHcX
tReIJ9cEe0BkdFmdveP6xUzEKxxtu5KwYayLbv/e44C4nP2OamURm07vJicHKYDYI+uWm7XwYORF
/kpqpdcis+IvwWmAY1/rZ3B1bx9DSDtO43IuSfnV4fWjJTKQ6a8VhntVYxyv5TNOCtVwskm0fqZe
eGUitKMUf8jl7T7/bjYfNbPlO34Ji6rG7KlAWaxcEV+4NZrohOSWqsOC01G+aCQeBWmo80AU6ZP6
64aOdUqlCeuLchLAee/PbWSpg2ACiIIiFH+liJ/7Jt7DbQY89YrYR4yKCzsOoZzHPmWycsrs/QDJ
mZftaBBfWHRf5zLyTVfl6UUouJQ/zlb2tIEIdwEauzN84NDLxnUVaWAS5Wlizs8TJHb5Vb6p5IXY
uksUN2X1PJKb5ijC144XsyFZZsKnKNq0m0DhcsQCzynI1GfWhdvI5TN8eas8+IDYNWzR+T6ehG38
7UP91l2paHm84Ru1FhNTiWmgNs3Ako/qnQ7P3BHGL3R/nr0z870FfqxOT9kzoKq4zQVnaO8MDXIk
cyTRyMYlMwYseCsQMboCLTyoepcWA+4mMAWcqubygnBh7oAHSTogEG2j7VHEx+Ooj9hnzf/i/Lz6
XryH6sWTOar1NVJW8V3thhW9y6IDiKIfc1wK4wWuboKB6PLzI5qmpgBBeIATtIcprivd6J0B5hPb
oZl5tEcdQ0RjjdirEaGuVB7M5sG6yy82gpLDdEbLeoP1hz/wi645VzXgezfyq8jErl80jhxOyGFj
Nodov1P5o1+9upZeoRtwlqN2vywUDHzfuTq6gsdhINC1siG2WT1+mDwHE3WJehXrIlCEyrcvTX0i
IRUWYi2tapH4cSWgrMd2hIFvfUlhtAT5cDDq081hLPlBhI/ky61+vGmjsVY1T2HStPZroC/cjTGD
QGgDt9HxTnKE0PMgJ9kL1sDpHPKcNWXgiqQrwsxgTyC9nOjgUWBVwTjYozNKzHFupN2XEou8JKeN
JM99F8DRRH1xpKPhmY+KpZ8/9f6DP9UB4oE5o5bIu+ywLwv4uc90cMNTaW2FFKTufEVpYjdSsPeq
ju9uOIMiSTHvFbe5Hdrg1GdStoo9vrYZWBfepkMQOi6vGcxW8PCMQ94gCMniIG7QB/eRQclfOKvA
z5rahSNLKKZmGnEVVMvedL6GpFd9MvRcwzNm+1P8smvbJpu2/3TPSYeVegGcGFpAguvcfzWnypkq
uK/rJu8OEy4gjRGOGrOJMopB98Y4TOcjTqTwrBReco0zYmH0tDgaG423UxJ7gL2n78C5tYS74SoJ
Jc6Qn1+9zIrjIKoFluUfUDmsvlyvqXsmKc0TuJZtNFI4egTjo5jx+2YZLNisF+9pFdUuy2b0nSoC
qnTDpKCvKaFERwJQzH2Bx/RC+MdWPDsliDUSwub1iL6XdRL5Dl/xokzXJF6KygvDdhdqao3e1/VW
/g4d22qIKwEztgmJAAUIR1BJ/ZCuprtcy9qsu4lB2RjnN9oy/QLpgAo59N5imlhyytBbUfbwR6zx
K0iAT6OL4K73KUOFnbNt/nheMltdTskfL3jhTjIV6u3UpRz2dJOrAP0EYcQMQqxaIPmXJUWslxeQ
POb/HVjeR3m8ByR4gomYHETih6SwF0Qc9DnN3C1veqRYHKY/DSfTtjkOa13a6SXKIWna3hHdI+Ou
/Fpfdfjp9JY5dSQw4DqmOr3aLsEfiGzfKLQfnnCixut0/XXHzjsdYikpPovPZyOaJXYOzA1TYxSK
57DAVgWIhHmbK0xP8XI4+rO2QxX0af1gvJ3Uf/9dFcn9fx7eykVd/7NMOfXbvM5RP2hf7LV9jEVl
miv3t79r20fDr90wWIypy04akL3ZNriex5C/8oGW0jnqdAML2RYAUJgFj4pf6YoGjrg3vQgRt6qL
hW0xE9fEIifQlL1oaLpfP+OZFFSPP2QLCBm/uFCLwkcsDzZdLkwuEcy5RNp7psvLvkjP3xGtGJui
SwnjruDlk1NLk5XbZ45E06upz51ufcjZ7fZYVAOZIXiACB/+BYG7bCSa72xKKeGf0n+VhjDE3Pn3
PYJ9RQopWCGjkVBggNUkIHtDMkvBICKSqIkuOwCSXo3RxZtdiNF5jZVt9SjP0GMLBpODGNv/wFO5
K1K6LP/Wn2s/oo6FDIUj9QB+xezS3R0ZNcfwZstmDDiTx9ep81H2ylLzuVcvdKyFKAT9qhS8fq7B
f80Ts1mbflmbT0NbPRAurPWje/e/AmhneLTczscxSY6tXt7pu+zCeIg+1VM7TydfoQ7m0zPxn1oz
91VgcGGgW5qMAQkwuYP3COJcAWfCP/n05x+49gdkRS3Q2uUIiGVqtc7XH/Ubs6z3Iapw+W5ENg3T
OlQunTQsM0RgSP6jjMCF8oDGfjub/9JXVs+SGztWsRuKsSOL0v6trjN4M24IXIiUMGnJfWHffm3f
ncQuDUTYoI1Bi3j1fuydvI2Rhr/StSJbTj171H6HFDb0Tforc7gvSSyscFDyR/Yuieqra8ohfwT8
KpwqN/WR124HyoaGnbTX70Rr+Vt2NhEPHcYbeDF1jU6G7U/urwdMXgeMi+IIMqgW0+xGbvcljdSl
cEBG8GZKEIBu9smu1fD/EvsCwIJyI+Bo8RDiNjVB8TcuN+wyP8of+HBEd4bAzjAy3vpktIEJWLsR
xFZQ0Vl67LBFYsyYxCPmyWUECLzoq5phpDcp8+rxdCDYgF2zWPxpGM0ZUE3s1IOLXWGhHKtlU2K+
Jen/U7O/dDPNCjPATyH1FW0Q8eqjyhctgAK+OBEQ4J729dVy6JXXeqRVIpGpoilXo2ejbzJip8ya
nbsLuOFnwnbZxPeoflNnYZJBRAmlJTE/+UQs5E7GFc4EW1J+ukEf5ogfq/EaUI8QFvNkKWJkShe4
MY3l/qzjwHTqeLNek45zIVpClupMeDG/HFu4bfFER4cHWH00/cFUXrK8l3UzCCW3zchvBVLt8tXR
yzmnBimsnNXKCVVj2moJUwyFpCuU8DfWMny17x3/0ycd3dxyhyNzFwDi8y5TDwhfiBIaD/9Z9I5K
mkyQEWcIg7f4uAcc7OtZK5Z5e958UYr036GuO4Qhfa57qSZZhi7pbfSfdDolTrsT+3uF7xRWJxQ4
iV55/NXlCta+MzPa0R1LrQKrgTKI/KJOg+ItPOqtehCN3/tOJ6B0Ijhnkt9MEtuANYTfLQye9rhN
911ZLRVgWiP5KPxAyUcRi5yxDilF29syM7cbPFySzIZI8SkVdJW+E5AVqEBJdnJjO54PjymcZQhp
dMkH+zw60iXN+haL/pZHctJJA2qblt5U6pgq4Jqo5q2KF9Aj+Ld6rEdMX7Gt2vW8E3WxWVh+Lq/c
Fu2Wij8AU8sdEHYvdyqWB6csEgE15gZPJf92n572OKaNZ7fxmuDxZMpB47lT87M01zIr18ex71M3
Z+Z85XJ6kEng1GLjBNiXXbWXF3V2INDbq6NoR24cTLTzDd/23GbaDij8hAh5Xxcjhev91YuRkHxq
CUwIR3pEyxggYIV1HGHVicPfV9BfK5NrbVfxAIETySlOCxRRGEr9gviKxm2r6M7N41htUfOKbxT2
uooymQwEt4gv6SEDXbIVzzy3mIuC9WIVfmFkHXsx3C0fP2e1wSzZLDGAtozp/MHMFQBPKbQsssIj
CygX2EeiM8vzya/CwksaTfbUpm3rz+XGhrBZpGxTbk7aIRByn9s2zN+zGw2TJUsNKoJyslYC+z3f
BuRsaxCjYzvIP+kbWLHCN9OQJnUNsQByUHPsJZ5pG6ZzaUUgvxOx0UaKlYRuzW2SedA6jW736ei5
jL8wKtIUyZ/KrpsqvsKsGXtBtLSEDQXYL7OhyCTJ6TgUlHh15f4TAfmFRfMgBgLkcrbZcNp0Iteh
NDlfXZsy34jW6hCZ4Ndni5qEa9KQp2nRHrCA0wAN3RY53XN/02NnVxWBszV/Zx7BNq07878PWufK
LaC1xwV/S0bdORDHbCASaV6Q4Oh/OYIDaNWQ8+52gpA4zng2xfyHO81x3ryVA9PnPvYfWeh7bOKy
gZ5/6RSpfWlrI7Hn+2ec2u6c8Jtb82djALt5x6bI235O2Pim85E3qdae0MtMNnH9ifIHn3WfN8G+
b80WvgfbwEVMJxR4QcUOZ3LaSTalcxq/OEbaaQg06CHrCTQVbrOBwy9YTP0FuLOctOwjuchxgDaD
yz9xb7/q4PvKX/IWEvkDZo9SiRG1VSaK4AcYRVjKQ4Ksxp04J7V+S3WI0ftc8VH/VMXLNxMZGJpP
5dsLJwrjpxXHlMZ2ffVLCA2vtb4HA6xCVPzXawtOzlOh4zzJDDZYLXsB2WzydKH8k9ktd70QunMF
meaVRrETf8NVG7r50GRwAP4wMWDNuTqZzpshqq4dznZMURSdaEZJDEW4razz5rXHy2vGclcR8SIS
ymbG/R2CP79axrR2ViPmkIWm4O4K3v8mVj9YAFO0KJLRemHjo8Zolq5ebIpGFZ8wql2iwxL4UWTL
fXhZ98JhFC6f/6KzoT9kc2rIsC5yUshtSWMhhtA7NrUGLki5pXlSKf8pD16+BBxoNS8QfrjVopLA
gP3YpBHLD6jhPGFSRGdTy0/ubuINGj0bAsCUIIxmWFI6e5oUFjibhN+VJE7F83I66GCxDep60Hbr
uPGfqbmyenH1/JGN6ivsRygEZk2vyRVEwzJ4rVXdEms5NYROteXuWnjrXEpKzEmV9UY6u/jALiii
AgaB3GZtb6LYQ+Mhz2tvinO3JUEThwjXn6/Z9M6hKxSurrCX8fEpa3E19ehPZEC/Jjtv4B6HWykd
lMG3SoMlpwd0AqGEgfHt4u7vm8demOAExxLzuuBATk1CQu/LzEkE2lbAu1na3STDA9TJV+YV/yQR
0xb9zDTEMkzAvZSPr1boASqjYWd8UToh5xmAMIillF1RGcvKf1eiar4LzUwbOvBXAIhR2FyLEW3D
+tCOEEvuvrLfwVjoQwcFhNKoPIZliiZXWqx+Xfs7VDMENmIVPYgGGSwoSrHN1q4rSk0QE88jGriT
0LkJA6EFVLLc0CVj+jGc/kPozoe591nDrk+RNZwspl7jWAw4d4+RSqtXx9/jl2+ny8S97kBzWb99
T39skpZrOwJYzRCMdCt+nzhVCsQDP9KzIvy3TYPkOy/WY6mK4/fmvaLHcC3ScW/r00Bhu+FmQAxy
3QMI0WKBxsXh5ebSmnhqesHmuXXSt1tV87dmYmWk04tncHwCuEeJcKwwjpn5mvDwdafZ9JzxCzQs
HsuQKD/5ju7WCIEcz+W1ivkI5oD51NUbg7RS7OijWhiFCcxSfz9Q+UJfZ6qlJxFjpeEE+pqLM7lN
QTuedkHbTIWjK6fFZ7MEFrhZMeqBUnyHLI/RzEsDhMXN2SP1EdFWuQkM7XN1aSh+iccbTi4E5NmH
ep1J8o/0JKo0Y5CtrJw90vj7/iBOSSjy8Go5Jr+6HO0Z/mwcRee+cxibpbwxoKGvE2YNgJ0vK7A1
ivJA1qUpNWkVtiv//fsu1A/fAtdGez90eYt4ijDoQrxOZG/CO5JwdAsLal7wgQcjujYreM0FE9R5
qsI7lcHDVB3+6oIIUSlfWMZJdVj2e4S3rMeUHfDcBHp4L9x/0409GO6vScmTJn15scYudI7Dm0pO
yjiXpdrSWj6So1DWb+S7uwPh9KMbVE0JP9wmrOqArb4RgSguIngxlMXpxzaZCamqGO/umz0nOoNX
LVdK9v6mwsISCJy4l02t24ZFeI1bBN035WXDYrLTvWkIvpPX9SLnwf7kWv0qAvqyNkZhY+qvPOB4
37yMqEUNYM8Dx7/BmhdhoIYBrhmqAqMIIdsZqbRkiW19tCAS/pTE0jCxjO/vy7vhH0JSKLCua9Mv
4xHDmwRYZS88wYnFOah2lrEV0TBuswdrmut223Dpl9MoVtrmLUtf/Bka0K1CLNCra60GOebhS4H1
EK1J71gdsH8OthGVChMG+zFCD01L0XMAMdnE82DexsmlWAmqKPTP/L1kIMk/A+gVGHkqjZLu1Go9
tEJf7+2EZ0kw1VlI7xNIWbx1AvRmGA9xDG2cKRA+2jtBeaBl9d7kMpj7+Tctf8r7wbA8AaHXoy3G
+eudeDzgD05VHqhyeyqKkStqErsm0SznF6Dv7so6PFUF9327V01yoSRE1d0pnmuG8lsj74X0tQgl
//+GfQ55jme5FY7NxFJIgJdgMO6NLOBa/N9EMA+dHNlIc3FbvBTkzGgk2YPvD4Ivj1VmbyCnZ7rB
wM5MdLJ3lLKyFxCaVnQs+EYnS+Z71B9xtH651VP5/2ZUNRfWb3ifotJg33tVBxugIqeFWpWbq6j3
DJb7B3fBeFiMPKggJRiO2LBzMbO74WB3gNp3a2Qibiq+fw0N6vljNYVI8qb3YcYcN6ECQkxHbgU/
BVHpqGEy1rBcuA+boqdMiHARoTjkzlELznHAx82Pplo6YPxrPfCmarJZkystIQ2mVyM+pjnjyyva
EKI7VXDEzZ0Acc0IEipVN0y6YpMw8rtpazJMCdeOwmlkZqJfj0dZUnFyVyyqqyPOGmk4DOCnu/YV
KSbOYXd7+kx7LRmdi+1CiW2X5YUUkGSOh0QvIskBmUA9QrlOFXPet96UKZ8fQZYs780FO9J7ZPjA
XCRi79ucUxreIO+nKa6YpfDkxxVjckkqU0MRUzZXq2OcMDUeB/ZPyBRuxB+i2zjRAsD9UrRvVBi/
DOX/GzImUn7zzI2kuCo5BLeLXp5y9CTAlJYa3bYRTndkzaygUmV+5XmPpvhmjAgfQaCvJWf2bJFP
uXwvEpUAhGubSEKPl+2upVglIAF8tDcAoWWF0o0ci6XTYlL8fknuz5nn8I4jc3SX9jvITp51MVGI
Lkyb9xFYAQzSm/WPtx0fjD8vRsfnq3FcoIY4UXrxym6ZU6ICXPkjMwXFg40XMvTs8kUXwlkZzNxC
FMbb+fSABIizzYgyMU8zJ/eJ4X8DdmD0ZkUdDeaTuxsLIR8Yc0+Cn6yM94PpQ5cOSNxK4ws8fgpK
8dkkHS8K9wap2qxfaqHesiOMS9wYJeaOX8m6B1oaZ9YsfWuQkgjh2iUyr7tc/D7PdP10K2yScnBG
q2uEL8Xw0RfUg/5NWWHCBs8gm20hfHwGBKPaDG5joEPF0+PnaLYrDJ0zCKBH4us/NFPZAjmEHnWK
wKijuR8UZb5cSypgqePyJLozR0bUaJnbSnRiakOtAbhA0q8QXG2vfhba0xDpWWwBbIRcm30tCGH/
UHr06WN0/cAeZyQbjrLuJ9Xs4cylG4V1hlj3m5HsFxrVJCviuVtiZOXyjEHNCsIdhFuA2L6AEM1u
+617cYhgYsraQ1DOSZ3w5se7pN7ZqUa0FCVctHM/zZ1OOZDNhQ+woCtpW2V4Y2UEw6lkLhUHGYjA
1uTgCLKGY0/1PnRs1VyKhULtHWZa3coC2da8yOlYcXNTJzg/a2z5/LrFw4PrFZGshQND0Tpi77rH
vERtcS4W9BuNlXwLhjcNWAfob5IqcBaYe8sbZLPlC6jdt+k0CTcnL0QNoT+WzEy6a6vjhQX/6Uu7
Sqp6nRg6Ep32SNgZ+koxdnADtf4IH1r6rBEQAeWgBHTGd6FmwXa/uIqQ+OIT9/U7uMyXBUclC06X
QLUBB1vs2huZMOuOf1k69js3ilhd+p4RQAF8L/4IsyPbLf3+IBzPtwzETK+e12A9B4sG+4DykfVC
uumOU9/nbRWuFBCO9HFaxhDo+TJ/jdXlI3wf5OE6u7/IBPsugteaUNTq1p3C0a0Ex8Vc3BQ58Kg2
bWANHaF5C4OrHF2Vzu8GJKufqRfcJSIp2gvbf9AjOfpNOOsGusLDv0JuXqOI4wupn4cSgbQhFyXh
8m4Y/OFGXlRz6vdGcJg5DkxVo4Zruy1p2K7jMflw/Vc4v2WWZECK7FY5uxWDx0prbQIQLJjfQO/9
UWsZUHScFJa9xPVaiYeXWlYCPrS3XEF43yH+HR/o2RVO3qzNQQTF8nI+Iu308JhM3Fl4//tDrknO
6Kusk3Fe8bnkM9tB6yf1x5RUUL7u/PZObY7oFlWVaOCA/qunXEy/JWblNkTBWIxzuWdymG1ok3Hc
RkLeMNGiz3gA4yqQHf/zxvlHA229vcG9PK8HGucHJSj94LZG4E+YEBVTjTvhCtWQ1gAUa6MTskr1
nn8PmZxQ3lvjbqfXI7zzC/LHV5zm1hM0y9DCY7CwHR2ij5m3yfbQeX+toaXYnHNFN4GpqGRSTNid
rigdYrx5hjDcEVY4Ub4T/fGxgWvGCnfatXn/7F/gJWFyiloQqxHyHwNVM5DZqxcL7ZovZ5OYY5Rm
PHYr6CkrNcCVje78L9HbJnsblQxoOrvUJL4RUY5dAHlPDe3N26yiz3UokT4MtsZpo1TElAU4Rl5G
83rQKhxPA0PfnVVO7AqtncBp4HMz4HvpaLj7QMgGRyskLQYxgSKCW15z+cvcpRBoT+8ymWD8R+HT
vjiMPsPwAg6fykKwUZ3AP+i17Q1sTa3NQLZ7XH14Cf+tHIotten/FJ4y/zkfwvtr+MslDNYBqYd3
RLYVdY71mczMY3D07qShxHbgKsZLCuafeQoqS6Xly4m1gc/vKtGOpNf5SP/onrHtSN6NAbK6Jpos
qwBA54wwadqIjlEeOm4Y6OwWOy9irsgCv21ldn7GFmk6xshZ81mEogwNCw4XbMo4U13+PkEM7D5k
Ia7qJ/1fkmbUACQn4OavWOJsp05qFhb3MZrWnVxhx4q8G4wMBrdgH5G1wUkOd+SN47fNSoL4FP0T
r1viPWR9cRDkpeZ8JeoB0Zwuev37bEn4c1optY3pwSD0K2gKpsa2k+xpkSxglZ7ZKM391NV6n/tY
q9krYBjOGsg18fuMPDbx+XdlO5pK9s8AU0dZyLt0WwFzOcu98Zm9LK9h2rwuxXQL0/FotYOP6fh8
c78dyk4TsTM4YeP779wZSjrxxXoieO79b1OJ7vJX3CNW6eOKD6rx2htHstFUz5Pa0XkVWRPvd3aQ
d9hwk3i07q8BiJowg6wP+KJ34IkjUjnrDlXec8zq+KWq6bJRERWQXWvhgx6ZQraQHAX0Hva/pNWU
LVZ6IlZoobNOJdnXZAW7BFes1YHthHdLIufjZHZ5tTn+h2j6kRbuBis/uiQPHk5GTCH2Ch8ib8Di
0GHU7twKRHuY54zRdFDosUK+nLeRZ4l6XdXrm4YSDCyBREeatAs+8pH39sy22XVK8hl28G3e2QV+
459UFC9Gp3g7FSywp2hSxgMJRD0mFYXCGWKpp/bpw+TgwVCf2FZXJU7tP9VZxzGnPU7qlrilfbW6
cH1KtClKHLZ8RnsDZs4mHfpkc9UVuoMvcOKy8fy1/pUFX31nXSlRG5Jdw7QkmMHm2cD1SrIcSKOM
J0c/qRP9j2R8qlvX2SvH62dA4X54r8aie4MHU/ED3p9fayp2nMUQUjD04QQsuf+G64/ArKBPqTG2
6uMNMmoY1DbzcrFwuyHUSuyjfHJsMBzAfq7JvR16UZe+Tdqu+gKWIkBwEE/arZKkYJJZ93z4+FBi
gu7ugabzYkdwfWz9uRum/7cmirW7uzRSUQ/ahSNl9XVo07me/4sylLYXPuoGyDDydo19BB+Bl1Rl
Q0vEzH7d/TUgBr4D8YOPhA1rhJuJ3Nx1fgAAC37fhoIclsV2FTIC5PMO4PUdFEdQ84kqZEHNKIHG
SHLnclpb64oCd/u2NlrZBeJ/UpwIRA/ggALd1nAJd9MHwMwV2ojYbQTPAXSRSs1K7/ofpswdV2NY
oxhdrVlKmQem+pipY+H94M+s9FiCCFW+n2N98hMG+6rU9wn3yNs64Q/vsBQFaZcAfCBanozFyp4Y
yohe6J0x+PR/tsoVB6qwYXxyVDtNFe+28dFgysZLw3W3Ez0DWFY1/2/2sOpnjMTuJR23iPUWeoQy
z0axLnjNZwP8GFAxXlXwmD9rnp9Xxyap2XnfZMXjJhpfiXNFyHfkn5CmAAcownGUcFRE+mp/soTE
ehUHnNxPD4pTPXGjN9VZVSXeqssFJX3Ief975YGwXdbXe8IRVMLGVt/9Y1t+Hh3u7iDgREPDMCI4
y+5NgRF4G6Jhaq0p5idshOlFAGGeO0xbVeeiC5EmBIAx4DZdwxyoPApHUSva1WCcBp69JZCWrFhV
J3iqSeUdnK87Me+fejreoBk4QkBWBq6bJP7MJCSKYsi2sf/W1pRzG+uKzFNcgwmcMou7AYJe5+vo
rz0OJPzMe4LJGsjh/HUI+uYAQeXx9xjjDLc1MrkLS1ZAiwonheTVigHRVztcYsduunA5KzeJ+2xx
0mhOsEYhBGzkLZ8onEGbguIGtK04ftZcIoCBFvpwJeGpCGb//h0G7x9YHQQ3ojx41T2vS+f2iZNr
kWsfBlWb1Lbx9+LZIIY4UF1TDkt+evqNEs/3Kg4fCbxOSC5Y7AdjqbzrRVpqXNTQOLnIM8BHdLW1
odVHl0oD98qI8xnBVnpKfp5rL13NkoMlwoW9QFxvL12CjCU7BG5kjCihylOT+bJtc8VAnsOgdhTW
l7gdH23z85fv83gfKcso1DXsCEHma4RZENvbZVqHbqEaBiS4Sa34LTrAELzfrspOSugDSGJ5KXHl
LSIf0DJ7qgvl0KuNRrjXNCwTJQG4VerKvRBq02HcWRzgn8R+YREQrL9rms+JWHC7wXJ9LWcqWGg7
gzURXA5aKb9OrWcL4+ChQwyeZaMLIAUozzK8wKD90j2avDP3X1q516YITdtg3s73Fiwq0krl5qO9
/eIkGYS1ikFcvrDKNtbelAs5qCgh6YUsRDAbqgyxn8EvalTRz5XXg/VFxLxifazBYVqXVw2UnRlF
Gfn6CiHB4cK+FjICbchb836oqYzwC665sYMquTuArFji3sS96jwRsq2Qtx/5jB/Vs6tAf3IZhgR9
EoGUaUh6hoA15HEa/WGuKaQAfpq6b5GKDVwHbMPiCGvAqCAEY9G6noCy0JgXRDrF63R5jh3g9A4g
x0d2DqCayARF5edSOBGrTEcCJJ9l43Mx9ICN6722XHzQ2CpECz19JMZn4Hx0vfObhrWQAtbTeEGM
7hivgIAlrcGqyOCD4KC74NWl7tuYWECTRBxaJB/TNGeCC54Y9Y6/4bhWQoKEbvDNsFlUPRfcY6t/
HMaMYduUSd91Hp86PKTv3WgQuVOBbiHNjJnRVfXen8RUzkFCFntt9q7Kb7ynXTdv2+hjPx/hc4MQ
3TI24T2vIC4EA9TIEjKA0z+Fzf366eC5tR13zmgnIjXzc7PfWR3moSOuY6GMVLs+AxFs39eyKBWF
xN/jBzfrDewhZSB6OJ3C1S1e9k4vVGI8mAzYcpfNPfujWffldkThgMYNJOJwiGjG2wEXVgDCeyxC
3FZIXpNRd3a3JuJFqZflcThGpJRCaCbna1AShT0KZtuKAuRBzpBm6dcdSmDeVMeMlqg3kadXMTC8
j3lM79OEpXQdXCSBv1dBw3YxZOJCNpGGTstW5+5V278E9ILlCuH4gKfbGTOeX9SyOWCM6SzeqM8/
BbAw44QHDumCGeRQlUmb/b5dtw86plbDvi3LiLV/EOSWgjxWn1CPU3p7mARiWpdLYhnUJsi21+aF
2NO50+PrEhSy538jdBnC5cvTWMDRdGDyUowgAiVr4cGD1hau8veDUseJnTBbjX86h3ZohimbBb+z
fEC/o+knHm6n1xMF+8d2Q7YVg1nu5b8w/hZmAdoXMjfwyZLre44nj7KVMrAE3OnJp0sOJDje3Tta
VhC00Ckae0vro3k79WaYUhWnzvwMGzfHzyrtt9cu6oUY+MUF28JF4n4HLKIcheHFGL5+xqmzveod
M2o2jiB8gAJwnZHcXjkB1TZHgixW5n4gKpWeC1oJmnn3v44vsXE+jFUBeXwbyB8ZvrDq8NNZvnGL
Je4492FlW4oYrUY01weV6odLLaTOChYNX04PyMKTfa2n+aTe3cds8JPD/vAm5PwXoC6zCloBT3y+
XaDIrQ7KmhiAZToJebRBW3NZi2eCnBqjSIfT6VLyLwa8vcx1j0u5YsmlchGAmCry0YKKwbFJnE70
1WcItSf1+ZCpaU0swyeweo5LBAdoM5ndnxvO9g91cz49q5ISS2ky8MOX+QtqnjR/bwCddLBSn0Zi
aGpApGfF3Q0TB9OmdFaVzTa4UBrcGUQYr+MmKyZUmWReksST1o/v9rgisdRXFdJ/W2/L9DfW0rJm
8EqERzTZtIgV4s4fRlz8aArgsZw62p0ORgHOKuCg3twXVw1KLbVAsKXPzHn/ndUvckzHj8xrEd+j
M/rTCv578ri2MCrQFB/x2I5TBGUnq9iNiZPRbqoDi5QC84ixUfQZzTr14xWuGDPQxcJ97VqYoOcD
PNDxzDZD9FlMnmoe6pD/81SZAHZOsUIoh19NwzCvmy1hVnwYPXspwSLVtiiihaM7UVCvGTFrlDQ5
drN2n9WvsbHD5NfP56ig6cjpwcTSifyvbGX7Ah7XIPw19gs678Ai8rd7PHXAXEd4sZr+6aPfNSfp
RUAonOwaM9ETDr16qXR0vZYCn8f4u5cNJ3u6PWWu1pQn6GG8YvwsoHb2N8J+c6RYpZo8SaKKGDTO
jaMIqvNlwk0Kk8iw06+5eA6y901idAqxt65xObnSIkjaZIIvFyG01qGagxGXz1CaOgvgtpQ112e9
HZaROzopyeMfympBDXfOSinGu5bRpBEoZsAJia/ZJi+rStysCzbY6T+Mq8FKXZojNAuMyxUUnJqW
eziuP2tACcVTWLV+Uircg+5i/sdFKIM2YqRg2ZINZBimkUAJyUwj0oA/D9gmOahdH3nywOggaZCA
SBkA8aPmu+zkKHuDpbmhN2aqfcNxIAQhCCk5Uz3YfXJT+g9TFFL2sEAho2GWONYPiHP9cAhecufn
lKr7gHUopfTxXLRresvh1K0OVoUGY1Dz6X+FrJDgWuD9y5N/rZLqPQC6Q2eajF132Wrv3Q1AmyCH
rccqPwl9fKR6hAaL7wxj82R5UOQYKPDUz35FXfGngsue6wo50a/uDJrAa3yyVexLOWhKHgoR9kFw
nhSw1myZKHdgLWngmoggp3wqeHnoH78Ewta5IkTfyD8MTWJnR0w3pIZPbSQZnCPP2l/jeVebL+eD
oeJriFtOr+H842A8UXUhJlPe2gLrG8M/aTtnO++IWfaJVmzu+EncO0rB38SYvMclyXjyeFgDPc+W
zx6P4tVveUYaJ+ce810grLMg+T4PGXoXudavXQwLztJQ1nYuNp+oAHoCiP2rocV3soAxq5tvfA2+
uuzehbO884ptsgqRQfa+dOZfbqjPQMEaO0/cRJdTJ4Yz4UvvhTa2bGE8+w+kagJBcbJvWMSpzisH
OskqS19uIXurvZKOzYVvxOCMPq3Q9aaW8Z7uvVV8i4ALwm49kQlsVzvcX+5vVhoWWhEwk3NY1fTQ
nMkEq/xYOMuAmTUYHDlLFjuLhk+CODQyjxk1dPiJiF9LvWGkkA8hGKheBF5tf72TPcJaH61jyg3l
S0hpStuuoydbI07K1VAQPtWBvXTNLHVFbnMfY4H4BhQp4lYo/W42+nvgCRkZJh67yNeJho9EZGik
nVLfoCX+Y7amFGZ6RXVs8aMTeq7l+ybSDnbmrsy6ExzUneSoYHJSdro03quq3fnpw6EEpmKTE7K8
tFI7lr3l3a5ZEI+qVkAbnCtauGbA+gNlkx/eKUx76z1X0soI6dm0AG4qlPvXAPYfABCDX63x1omu
44im5mo6IZmutYEMyuA3lI/ncE5APEg+AHVfgzW1WQuU/y16JfbtMDeahcuidz/hdCid7BaXndjX
MJnSK9/9BllOdy1BpPLuiIsFL1l0ZZuq9+knocRd4r2M95eTzfxtLkbXgq8GMvWJ8m2pb3aTlJKj
l7ubzQVpla3LY/Lllfr8pVQk8RGRFRbjBd9/fcLHAHchnoel4cAABTOBNmY/lcszS/VtRJMkxYJj
MrmCHJ1YKK8Aqng2whYgMsBaKzI8U0Fu4xq9dXs+aLte86bXfLFEpD3nkGbRCa8zVe/CCgC0gPEN
qVGbIxIc/lSd0e9EUo6qg/ISYKe+IbJtCLGGZmzC+OQulUYYgtWkTUnFs6dlL9ZQUFfjzwq+d2Ql
U8IIkTADgRh9u9Rr6Pz43IuDgTxNYgb6JKD/wmcXmtUMgrOFvPMX4pn48gNYb4i0tfTyFHhgFcHS
lzjtOn1Ty+ogxBAJw9yARnF1S+/fw4FXHBNNf0wsGIoFJ5kC2dpLpVRucu6KrsrccTtNjDgkcHIO
uK4Xq3RYGZjLNSUB/4KO3fvX/qN3Ncj17eiRCia3RAqn7P2WWyUbO3e0g1wcHdILrGDlqrbLGT2v
7e6ndWiTKATkx3YYO9LxCQktNxqmJMv9YQLNO/zZiZqwPB/FTqNfJ4HT3X5sKk+X2meeQ+aFbI+T
l/3p7jVVx4k4Ur66zmCACFG8XCL0/Cv03OyltQKPSJ3UmMTpnwRmPIRNQVfPM/cWgXlxEof2g8RR
Ey+CCNT8VSi2R0ZiAl8bvEpHC5cAUjvedI8uS55w9uFQLugwZ3DIGUeDnmYIr67hhQM3BucVI9EH
+wapPaptAlHUeXBr3qEyU+Pj4YN9RbNwS5JfioWGi7oXZkvK0ebqOpWRwcK6qk3yIq/LZGJ3J60Z
O6ySDIZfMzXh2HWqYyUmXjbXb896r+uHlGWpeaMofuzGZubJIrHa84eVL82zrY/U7itLkru2Sq+y
8HVIeWmKHGdMYgj+dcU0FA3/2mJFhtJeGi1dgWA799s2UkF4woWd4uxgEuxFCIe6uPqVzxbgEqrl
ZvELt3OiDrMNOL6z6UfRIAZOJ8DrwnwAO3yYtWSZzbstIw0i+ex/Iv4gdqeRsFdKPjtfef7KGn2w
kmGZjf90y2gH0hjS5ISdlTwRs+pPjhDlbmnN/ovvgnTiWLHJ1PXla0o4b0rcq5+7uQQBuQzFYfMR
GEBRU4LDPHO0fyxCvoUhX1IyOWJvK6NGQyM8lzqSlA5b4/4QRV5PZ2azK7aBjhNYLnckmQgiAmvK
9kLW62i9vfyjbCfxd8AvGnMAhy8BjkgD6oZUHcBUeEi3yrvRaPtTMRpqUq45Jgg1uP1p/abyjfgy
WmLiasRY/AZR0Ogr26vmKv0svSflQ6iym84tZZrmv8TRvIO4BBKwp9fWw4T+bt16/XVzUDGhi0id
+6OihbHQ6vm3zj1Szxu2l9YrU17icRmdlQPsdOP8/wCC/fXKhUwXN7W9XTcFCBhNDRwv6SAdrovD
HKatrUOO4mcO+K5kmwx9Pqv4J0QV8IkSMglFCKuGhD0bLuk3KCLPCwZPm63w2yuXj3b1bCVhLtlm
yfW9SViyxHyvzhFufCdJiZxsRrFHUoMNdXbZnZfv/7RJhr+Uf9UVWpbTkym4cOX27Lr4mnkOaKPQ
dl2KyslSWmfoIrxAm2PoOi6nAtOBb6j1ZhyoOhT/10s/hCVA3Y5lqI3M0Y6lCyaNouQFHQKVTtXq
Cbx5uL6K74jGXBJcj6ojNt95YMqiCppHboezfmY2pnfXOc408GxnllNTAkYSQAS+l4lnE8rDY1jI
OxtUT2b7VhJvAYajM4YTKslQ+YlEvEueKain+LHtBzF51ae4ajGRQRtrnDKCy0527YAvnUylFPNX
mDCAnSXtCQ+Z4sSgziFu6wKgVDGMHLvE8ZlmdwYC5PGBgTKrYD6LgfjbryiLs8crVqoqKWcYVd3c
hCPrmxbzN7M249hKBdkZAaUTNX74EI9v+9u/GjwW42MXbCVxZiZa9/ROMbE/ByzKuRGpIpmeJR+8
DOmpC5M6U/9grDDcqdLnKtCTQxkRXyVwssC16eXVO/IEv2ej0Uz+NquNf+/WcbFthPL62J5+6vbp
orr3sYI0WUSV73VMDVXUxfAzr8CUO8wF06oAfQYhv+uvMnJ0KbNB9k/HmyWfTVTaW6/tLN6HnIxn
IJIQC4Qyfb0INSgSTyvIsqG9plMS6YP2oK4vjZ3rxl1aruzluMikBi4N2HTSA5aB3rVzGzAcwP7l
Pz27SSZLxWstpG6KFXVkWFOk0Mg8Nh/RoVQ7gh2x+iixXtrXJOCGg6H1mM/TvngYBZwLyv3WjG6B
64OW59/DHIrFwez/ShpXVDJW58SvodSkXOeo5VBJQdM5zAawlv2S4Kam2NUkzIEs+TU0NhNGKOA0
FfbP8qQt1N3IfDYjwm2BHYco/Xq38tw9pu2bwn1r+xbt2yGk5BuYKYtUAn2J2ugeJasr7SOLr7zy
76QASgjtr5+eSQb8yTkijQrk6eU4EZ9+DxIjqtspdhr6E5iQEyutcDW6xXuKkO3mb1kes/Tc1r7R
csjCXS8zAM7kQ0uEgyYOSNMdQCXTzQu+UEyI55DrYNA2smAwl7gzNnPX4mZ0VsRQ6UogqZ+viA9T
Ru2dkhvRiZhNERF2eTxo7JUZuN+sskFcPLaBUgl3f9jHR19zseF+fLo/1zdqB3pW5j8XSISUXWwH
2ysmoNbwagJXowYcb1O2pHizdI+2qiC5VtCeG+C9Gpr6/TaaiQ7Onqz8QTnF/YXUKn+/ZQfKzMGs
gRhAOyvjyd3QwO3+CTFgm+OxnrimvsanI3yPvGo+KtQaypR2Lld4dvxC/AsAZUXjqj4N0OAiaViQ
/cCqwIHgPB4O1+paI2UmZbgY9rCytNdo/IBLVHxuPsFihfMdZ11hB5oxKbzifFBaeMJtmYlqxCSx
k1bYpt0KBih0qgJgut0RQY2jAOfChqwCE87fBdqN3l9UwHcDF23rxD/GP1ygeZzw+nt50OR5wiKA
L6SvlluJezedcISy7YIBfszgVoblaI/Kg+3Ih9sJeClOg+wpMSQKChZC9oNk2b5o/gW91oBbDSWf
IDTY5duPH6duM4g3WVmgFJIRlGIQuDz+I+Ig0mYspfIAQWi76/LfoJETWuCNtTNv82Giu/1TCcta
pOm0TUhM83oSyNbxM8DefZYCZoEIq7y3c3AzukPGkhd5DGaZp+s0Z7IVMSefIh4uxaOyG66SivYT
EN3/G+8B/kBRMUZmpol5NglI6kZtqknttuxp3NcY5ksoinlOLP5OUcCCOHYJov6wb+IUyltHg2BS
QEFHg38/AXyKUhHCGHoU1dAIf5Ef3uK/9vhgB0sRsgfCy2qM7Rv38pgKBlbJAIjFI/esiXABgfAT
ubi0WemRUKD0vmNWrcNRZ6H21ebRZ/A5dgJ2ofUO2zHtDkvGV2n01L2SbR2IgpTa/bHfWgmYswLI
YZIA/R3egCTffr8ypgAd4hBSKonJPDUCy/0hc9Qed5ZUc6DfizXVPLDlA62dY/Le60SXLnraqoGe
iU1uueo6k5HRUu5jG2H7g8bQRkIUV54GaUXHbxEQNKeCtLOFuqqCaoPSBF4N3qXOatXr0LbiTY/u
vutYiY8qEkXbWP5k4ICRH50SsJtCudw4sNEdN+w2OJAx0flGSswgnj5bnDu4ng1kiIJqyULUWJpY
LVJ11pcC3fYvAL39oggQMESWk2e4GlqTwAzG3O7snyk9WgtH3w5rqxtdK9nqf3BdXSXZgngWUcXc
Sn8ewEUT1/Dr8FNJBH1lpgLfwKUKAvVPbDeVfbr10Q02Nls8bc/RjDY2JiZdiJ5BbgLbSDhhGc7g
DLYbfKYhmsY/wyOlzQuyxYuHAQ7paTaTNXq6SzBPtt1xqHTGYBfEbDSV2lGiAI7E26Ws+xT/nLTQ
uYM/MxXCmTUtRDlE022h4bA/X9N3oE8O+baI82DF8gOGrnX9wmfsO1dXa5khz9gScwKsHQSZquzu
ua+DcU2VjNu/ltHGJ6egKDL253tCuAEYAKeYhHl7mXGgCYRV2Kl1kTE0Znhkj/6FvThfzcyAEXpz
GEnI+PJzUkmsUiYBDk5Uocyfw/ME19NtR12vBFPcUWtcS6gAsGv1Yums3ZIwGjP6eamc52WcDOeG
rR1cl0N+5Wb5EC7IavieeU/KfeWcUUfPRy/5t/NUgw7Rb4Xz+C3IikwopBDb8i2fQpnpnSW7xG5r
KXcnhaZNTaF5c28tWowyTVrftUhlvmAqaj5hJffwBvbMxNiynkSjWqeQ/MW5s469Y6IQKMI447Dt
ZCG/3x/Df8buIJNBby5laX3YE7RNGLC/AMmajRTcvvgqSo2ttrFPfA+mPftgDwodGiLESMOcD9SI
6qzTQBuGxBGT2APppXNTVjsPbnd8RXhxHwxCRQHKfiXfOnX08wJ8XrUTz9Tcq0KgYjEF5skBiyDt
sEWOL1fDhUc20peR4DSJ/r7xo21QVxY6G/yi7CJqaAjq6lfuS2E3yWP8aoh25Y/LwIT/1nKnot1C
vkfsRyeBTm5Rya1bLAp2NtYXAMhtQCv0vVhao77NRtt/z0+Qp9/BAjnXtf0U/xDArDpQfhXvEmty
qNI+sgb9fBHsdvENIew2hYu4hJPPafupG9Z4badYCs5ELDjjN/BbByvxVHONeDPQyisCf3b2BGz+
43rFAd77a7kuYblAoFKE81OlOQSlbe+XEMozsaZWYgV0XgTezwfmaNxH4r3jmhXsJ9doGPSc1r85
wY63NDAuk0woem10kdxkAMt4pEkfrSgnt0XhCMHjFjFVnxx0bfCB/OKpX4i8GhC+qAmcqkFa0mR2
xOnU1YU7/5SlqjRjstpmlqFyCzuIKlbpVu+YPk6MLV1YaCydwX6nTFxBVNQrIxSynCvHK4uSo8uI
l8MPXfC8m+/tTCyBt4802QumXp3a17HadHp/RUp5OrcFBxRG8BhKAa9+g86vFDrwsCLoKv2zsA21
xhgSUkhs+FZzwjktQyb70vAefGZRqXyVJEvKNY/R1bfxDye6qeiS0nR8UD6hqvFGjaE96C9aIMPr
bwVNqRWzWisGJlz6QPRDdhjO9K92Siy0kA4Um/6QibdRfx2T2A758OnAFMweZw7kkAoD6RTCERfF
T5fCitHXJxDErZEqwmgH9qzsNGdm4sfHKviWg6qv792LgQeNB8kXn9wwEVkzqY2dllFm/DTrziuj
TToxMLOItOD6VfgappSfLED6aDLLQ824qM5h5/5SVdBBu2qvavas6X56/BlK/at5rAokGpq+BCGR
6k9PH1vm5qRG33FxtlaYxUPdl5/682WSWInetBYedI6YxzEvizzcrw1lvcCH3bMmVCM74fEARyyW
XoSa8EECO2j7aZIVrQnriXKJ/9B1JG8Z25bw8zqjigmgOC8ZGLRS0WAUkFmHO+znqWY7XxmQEmtw
eVkxDLgMPPDH/pYQowxZjP0mFoicF323JVBEvWiuC0/qBcZH02/jXOexRuUk3ijYB2HsPr8XZnQs
EwdU395tvmwIMBD3SxuAKAppuWbSvV7XNda1HvAXwFBKBTF/01CWRPkzMtrf70YrMEgOf2O+VOq4
E5sDl+pfZ3S9G+a80jJ/dqP+1+l5tFXICScVs+ZlVuGmwWXd9QrJ6S9uBcDViN4fP3BccGuP/Sow
oh5iOZ15bYvNNbdIyPika1xSXhL7xAkEev4zWM+MFY2wZWLtANrizjejkmcduRRiK7wTOBEnDoMX
TE/QqNM6HgwnwaV1UCxgGtWlvYKdgYtAiG5uvvC5FEENSXNl5nP+Be1dS25cdXZa3Q8xplL1bBPW
UJtDR23gjcMfI+eEtv31sb7qiQbrfFeY8wCoR0zzJTGwLSkOWEKCP71bpGBEsybkW8L6/Ba8y/UW
IokaAfm1nkk6nbbL8nxHP/mBEFNZupIIs3aASGr+3olZrltIT62tOhVjzKl5PGMSRo+9p9LfU74/
SALbm5WP95leGZCkWQ8VzZWQVpKr5q4dVVZ8neVkW+7rMd5mUiuTPR2+JtY3/OpD/TDcdQO6z/FA
xGbvSTJY5nbsGXUZaI3vf/m01V86QpojHfYrWFR2y+AQBqmY5KLy0hqc/tnz2wwU3Mz9F7EMbVVk
M2BRdNtjkBWzCltulc5LlcVC405n2TbRHQ+k9jIVxpqLziblKIM5t5hrjAb8/MwZZHMBO8kHkmJ9
KhZEiwQk2ZTsMaKxDd5YYyB+ma+f0M23NYe63H76jo4lt3fcw1UjdUiMRB1ZP3hwikhe4RfUzTad
UNBZib1j0NxrVZiImSwqLnFtIkikvpbDQWnVW3sWoVuPhcYQTsG3LDEH6MfcZhp7I7QZHDXeibHh
w4+wwsdZOWjoI6jcCnqT+bCEwhZm/TrVPomXWdh0WBZPu2kX8s6hJBkxmRnM5aF0Yb9s9YKZrJGi
nZY5WuBZphg31cXqgtxxNA7aa4LXwmrrxDkvaay4wCaUQ75jY/wxqLPeKlk6CiwhasfuZ8zGtY+9
8Zsx5VW/3edXrerHbyV0UaLE+KgeG1yoqn0rGK1x69hlUzaO8rSH0pAdGFfNS9wBV7Qnn/O2L3S2
yj3F0hD8+s0ax7M0LlGAD8E1HIcjYJE4Ed4Of5wmvxNQhDOOCf961ug/kULJdMLYqw3Z+Qw3fWkX
6aDwcnYqtVTBrA03lI8XqT2udDfJjF/IfG1RADzXhen8wkXsclMF1UUcQ4oX6wcSTfywu5FISwAq
ikO4CojoI7yNlAFE8GqJPwY4oZunq0Gum+1aclyAeISBfev/iBW0j7a5PR7A1rc8U6EJ4loG4l0Y
wf+hAcod6TNNFh38brgzCuEIKqc6MoBDy8vJaMAD42MWYo4ONloIFa0XO4DwWmwNXMTzmUCFmWIF
YV2DCcci0LoMtsvgg3d68EJdPZtU/XirwFJa6qlBxHOb9DPio0iyVjAV8LJ328qlogt9E5Q5lJsS
cemtYmW1M59/QXB3Lv9h7EfELtEUly88I4xSZ1404fl9ortB4KrVbAbLDfwInqDaW327r2htFApH
RFxrcQuno2atG2iE2UzcW4dULoDKp/kSwWN/clzUKSYqXhEs8UtgDx73OucjfY6shw0+YNXJRZhP
0kkxmYClYBA6PZXZ4Ha68CrSGM7ulYsLRL/eV7rIlahn5jq6ZXRAqjkjvS5fuG06ytk9VIxGacfg
S81Qj5yN117o+8Y7ZMJ+QIyVecoGLT0ERQoj+B/seyoeGYIx0G8RUjUMuOLEWmA14mWEr43XhjZc
4IW++rP2/NHXf4YXrc3LpoUEkdTWc8gLBRwF7i7yGX9/Ez91SJfgl3J45C50XArq78ryC8tkOD8Z
//Ft3kuw8nPhjgHojGdXI0Qnm96Cj1lEJ8SnowvFaOt5FKpE/OFNK9CKczTe+szU2C9e+w+XI5K9
/KPcr44W7+nufC2PREPJbLhlIwuNpn1NDRHPWOczg+v8xtmZ7fPH8PSVFg6W/oMuOEqqR4xFVDwE
+RczZ/q/rEPl6sQg/mkxoBEs51HoCv82w21N5B5rA46AEaUAo7/BLxMoLMqwcL8Re6f0cUJPHVeY
JszlHWrehUy/ecwaiuazXbDOYrRBh2yov3sUiNoNweascsv9eIRF0QVyR4Cq3tBZl6onMjPhAGRq
JPnI10AYTq7Crdo3k/GDorROBh3jB86kQRfn/mV7DHjAOCSdom8I1OBP10QyCfZgrw4d9EoM81X5
abjwEtzvIW6QWKSo3nodKlPZsenS/p+uKY9JIoeYK71vaBoATqUhZVpscXe03Egz2DmlH0pRNzhp
kkvZdXzwfZIw7IxqgOOpVpa0Lkb/Mgbq9amlnOk6L1WvFQJSBwRKFNBDp7Fwm1VlP2fijOTVWgJw
cYzu5pCsOLqKIdUhKmn59nkN7C0a93LOywnR+bwqJObsuIzsI0WflJhiIzxPwFQSQLlYcLVcTsrh
m+yTwusSpalD0FBYrli7IgCwmkgs6TfP5IgHsSew+WQkiizkV+FbSQeb5zAKQV0Ew+J5X13aW3Xd
XI5O7w2zl+5gOOEFuSF4CgEAC5Jvw/v4FgUvp6yyUhY7kq/WhL89vn4bo8iaB9J31T+Fd5y4RpVV
DflXuCC8Ju9EIjI2nkuZk3b7xbkXygnVlqFiorIJ/G3sXxbDHdNbjIfjgniMwuXy6OGliWMINidt
LjyEZzcfvPxlCBMxeO1JJUfW0YBq+9LM+YnPyYtJwuSHajvgQV+Xo97VjgFo58KfQePqQPKdB4F5
AfHtB3If1a4ZU/9HUng7wIB6bWJ1DC1BHHJKmiPycrLFOvqkjFPdg8gcN+kJCN/ewY1DUrtIKixu
h3LSXTZXAPBo1+iFdPzF2dRi3H+jOaDub13fbgkUae1WnjgKl/lIcIztYlNB2G1BQS8Kcb0aAxtC
m7ZN9N5lHelLKz1ijsuUmsIeAWInkPLX6i8/8V2N170BkUhpcVv7lSQjDNIGKGJV4m9WG21i1pxd
QsfElaNtaccUpGHmNfLqMcXhDktfW4b5En1NTyKOSdUAi0pmAyCS60diZCSBsQG/jj4zQeKdESCZ
TeMOxn0ht9sejURlWndwDQmhI0L800uyCV+eTRjR9paUhBth4pkD5Fy9lMcMFD4pBRjerBVRvq0l
ThBApthw53aGBuQpkAoxCZFPgMedPM64sN0i7rRDb2ujf7uNsSUS3sVF/sI0eSczxI3VeOJcYkFj
M0XlvpNHPIaV8pOGmfmGYV7NLyiDh2OyAHspqRBQ7tT6jEDwg7+c1Ik5taTdmfUcUjjHZ3e6WGId
E6RRvrFmsqWjPuh/y2m1Z8820YlDv0ei/V2gyzHLb1efR2eCyKzokLVq2J2xzPAsBZWySkWhDCKM
Noa0yAxkIWf3zPskdObKC1Tl9AcaEJgezBJ3iOdRHQdvBFRhdo3CMngZMXuCNT0wLD3jgGgq7jE0
+SQy17d6mLzkbY6gH6PsODr1SheTrM9g2SwHvLcOh5bTGOeT3mxz6HTSv7xkpX8YwVaB8Ykl35zf
qLKdqTV0PPTpW9YinKnWkly/6qamrycsgSus/NrwAtwGPVibAy2CmAr5v/Q4yZnh486wi3INl7ho
z0TejdkNJ5Aa3iEnmvU0UBbEw1Bn09cW5Bce8BA7Ilhka1PlfIpqGH3UkUkKU2BBY+S+AzmLfKAP
1rOAT4sHgiItUFfH2ktxw7t24EhwgPL2/lXHNicmBT6ycaBb84gviMrX1HjwggL/0gqsuCFtEup4
k/DSqkT+6CRq1WuGsOm2ELFQegZuOSbkyRZceUNMctyo/sO7YOQqLptF7BqDJ8rE7tclzZHi4K9X
vLroS6e5lPFuSU972slb97dugSlb43GXYf4fkvLjSKb8OkDUfQDe9gjEfj+74U+k9SA1mtuZDszw
PyZr04Q/DbU5T3lIMbE832/IQplI7naD/dooHQIrfF7tJzLKobSY31Tn7ERBl26QvQy2Bq61eMi/
eOi6fVfMAhj8oYpki77ENZN29ENeQOtwG++2hjj95fortlDcHMta8Yb6bcvfHBe4438+5RQqLpG2
b4XtTIs5yGMPpWFC7POFFnGQPmp6jTfPYv61bMONDwU+mfOJ6D2QLU36ErN91ttq5j60m7nVWnCO
obCADlucs0CujWP3Anp1z3JXGWeekHlde2f3Q53F3fBB5iBBbekfzB/TxFQI3g8rp6gi0CtgtFG9
4UM0YGQhdsATakQMgj3rFD8tYXYvh6pur0tKhtnXADnh/yS+QZCcmdFv2z6ar+UwWL+59LTr75rU
XPkEZkqtgoSoJw4qDb0cSysj8izOpg4unJirGpZAslAYv9O1Jg6cToBQ7dmbeLc6zksPUxEzcFez
Vxnb07RKd2CFBqr256de2zjpuj5Buv9elVXRuNKiPwcCh4Dr3hH8I3kVDAtEH1tvHCfwUHK96wVD
fn7hAKx+EyN/NrezX9OfwZYsXeqHdes6TiBYwvp0C14RG0NIMkXel6FG9msrl0baAJ//NbuOGW47
jEusKsPFS6MIxBCkddnKnLi+6JscUdrs8QJ+R5LRyz9m3a6a2EBpcqrIS3JwHqUWNOHNm4cfbDYp
QSL7XqIiEq0oLNr34Bl0gyznQOQQ8Ydsr0EDM5l2VURbnluAScdTmYMRu/I9kC1wKqGfRQQFvFX+
7VTBLU3/kdvreucTLTUcfxj3q5jSxC4QaD0wuLOVt0CyedoXg7oYxgGVlYx5N+cFkJBXjzYeU2tU
xRofNKZgfU7vVhg8uOIyowLyK0VU9UHRPrUtW8FarwVKyMkuT/dGBPfUjb28yXwSAj++H9OCxEAj
3OkS04qZYjNNyh565dPB+tfFGOlPyLbBaEpODMpgv5nzlZLzuJFI17yl6e7j8T+yAgIR0cDcQx3D
EqhTViEqeB+N/VMcrO74s4u5LDCK81EP/4H1bBZmkytKBBcyBHH9Q/IwYS1KojCuPdTXB+SE4CXx
uui2OwCcL2PRRUI667CptyiY4f22bSOzFh18C9FZdbJ+MEGGmLeCtfhHnHNrJNUNJYn+CMgiqR/P
l5vLCJ6HmBweuj0ImA3uNKMjd37emPG9Zne0UkJBXuuabCJSA1iEpuUilCLc9bMwSUmEJMKuNiGO
nhMvrnXgMjZgCDWL/7dA8HL2+4lj4Evvwg0SKV+K1gMahLlkdMmTFLE5txbaBeQ4FKTRkZG+eVmS
xFRuc1hkgTIAgXyxf5lRALhFosEKL5zE3gWHhmojbvIyIYQ3NBEhy8dNn+vJlA5CiLUlZYZiAY7V
JU0e99CCkA+CvlX6WwUqdyVlKYZ7EXL/YdfztBJZA4JphNz6zgSH3h3CLzIikISw+1tcr8bQLjX8
CZ5QNpoq6/sDHDrqhRUTRz/v18lUodAgZWpCMAHfqHBUx9NNDSiVfzTHxlu1rIwOtdpvUVvWvNxU
KPqJOWQZvbXvPGhLoe35lQ+s5TPl4kf6OOL/3NAzvutaVdUnDfn1VKxffQItkbMyiaxdeLJ0cqW7
WUBoSMuP55trbRJplOksPWjO/M15Y+x1qvkeP4T8FoRGaBn9EnTJUf1XrFWCVa59XjymDRpw3OsA
+I/dRVSxp/9mvAGNPSzLGyIiOE68F1oF+MefcakE9nFx3deXvPZo5RlZEiC9Z86SKvi8iM8AoVLK
riUCjWSMBlwFrplxz5dGSFsNW743jY5N9s648cFdW2Nx7LNiITWeKQFvn+Pdefn7e3xUDkkx8QvK
XIfyD3JgR87qu13INQCW2kyEvDJMaOmsRsPE5YoHGM8wNOeW1GlQ12m/CssFOUBR9G9XiLNKiRHQ
TUydgja1f84em3Haer7KPB6oe4qZ/G+1OXOh9Em42ImqZu+CH8uwPFeqqtYxNM4Icc49GoU3zvee
WeQUHsTb19klqj/T7m1QbupgRBCfKUzRbs6Z7KLigO2Q8GI6JcXfsxR0/PpjBpnTmSeIcx1fDI3g
qh/ihPiyjQQNS2W8It8T49yGjymArTCcKwxcIZSjMjNIatwyoGv3QjE2/tREnftuf882b+Rl07Cq
yQX7Anrp9oafzD9aFtLY717gbcfVBigedjI/7GXfQrxVJpoiwKdTP2M6dmwjnfD7tVf8jXXiT8lG
5Ggns69b2zR6ajK9YvuJp/BSMMco4XAoIx2Cxg6Wdsh5YSAndh1RSHsHNjb8I1eWOIu0RPmmSNUa
qQNneX9OkHOg3E0yzvOgnimm4uK8V3YdkAQjoocRq3D+708wEN6Md0oX0a6oXb74WDe+yOJkNLL1
LNE6gvTQxORAjJLqZqURNAAidTZPScZcKhXj7eWXcD2FcgmjP75xhX+Y/Ko+i8ghKpGxOluTsl5w
eaLc4L9dIYbUWsJS67ONueVw4xeQT7qvsVV6ZUzPkxW0bVoiABS7GlicBNzK098KLMUCGsdEivOI
W4b5KJqzPzOO4EwNcvr58wsT4B1p4MR+fBkVDVOV6OEYmg+QKplytMSLyxAEFbUbR7KsWk2gHayv
uQ+Yh5EFs21uueiWNIiT8vdDe83rCOQrRkkA2FJWhyO6NPJGIN2zEPzH7AuPiwz7JAUKpp7UEyx/
O5r0r+ko6aQnD3h904qsU/sG1Atug4wzVdUk6gmhfNnlYCo50dteKNga7Bc7HigiE8H8zVSrz7gc
fR7eY40H2AI/pXjKi8B9KJViVtXHsan8gXmGDcHcauaxe7/KpO2iXy1l3C8aokv4scbgTa6lrPYp
TaDYEH7wAx/mI9jBWANmMERSU22o2O5ZMDm4DuKid5jYLp7A537sKFCztOwqhYxyvCda5uUMGdgq
TkqwGwQYXv23oehi6vMm5fP6aCEAnjiXoQpw2wqnG8nVI6+BSQKDk1JgsI6hiav1UFobRjx1ZBce
F87+nSSlyeY8kLbc9hmwOFk4b56aCxP1ofIiQzRoe4p1i61+IR1aUPblEUqjh2xeaY+SaazxrMJr
BZx5yatDsxJSxOiq2wofKXr0XEr2LibY00TkmeAEbIJVW2h73KNXT4xFmD8jpMpAFlvummJnnB7v
64deYoqXMNOfSkOvEd6zOTafCnjFD6UFyc21AmQQS9doFJOfGxdb4seZ8dfes+dTKNZ0aXQU0s0K
jGp3WXpF26WtOyQPmGzExgmrwD6hmQ9rWZ486D0xxntHPwiIxL0VwV34NOk+kZfBpEwedUGzTVt1
xHW2gVlffGLIiFI8ZuNP1+EjAfWS6F6aF76cVOSa1gSaIcfaIKUgk3k+kXKUnzCnVFCXgUKpPVck
VwqulWXvx+6zpXIimre6OcE1JADDt8TTEIGf2ubQR5KwG8H34ERS6iiAqgY5txMeyY97LxpRKcPM
MlZw0p2qkRHiLpFtoFR+R5vYCQ3j5AMLYC/eFlaiEu7uVo3I3Lj5aFGz5KhDsehWskBWFfT5c9ii
h5wCxrMMVZ3kLle/+j+0h2/jqk8/KJ75h5jTRxA/vlvApEYqbqk/P/hrtAgxxhb9qWHC6nANjj3M
OUFg5Eo4/bQJS69NXACKWy2vrpJm4/2C3yKqwwY99btsbO/VSwLcKNIrDrEu1nzd/9+h6lny1VYO
0KoqDaqmdE+Bi1lbkDXpnEjW/w0oP55zYu7Jdz5VcFCa43IgewPUa1t7goWYy61w9vHivpD6CW18
osOS6ASgbGcdAswXQ+UuGt9bBJHEX7v0yq+u4p00TX4iyN4AEM3QbhQVhsCGCpQcQDAk4BLy6aaq
GA5odVMfSejspViwm2MMHv2HDrAyyVmlSNPbYYDlOqawnK76PLvMqRmIuUZOcxXOy7bUsNnlTa2H
E+SLLPQPXzlV+UEBL0eOmqNIUIXCcLhNKELhzTTc4btMBj3As/vtNUOeEgiXThvvlGNXmqAZafn4
0kKDF0VJwYT28DwQ4LmxqX6LV4xG1vHzC7qwtJYD6a23z5URMs9qrf9Fq1cRf6Q+oH3bxClfCz0P
Hiyde/FZofubgpBWXlak4gKkO0leG0am85SgUum/Bjs56lMuC5C6Gt1PEVKlN+Cl5Kq+IzMIqmR2
IIJ/UbvL4hapR+SgIJaTVutOiNbkeFkLP4JP+8zibYtqnMoxv5ACoCNT0DUk+pT7A0C4OIKNuZLi
6Gqvd9lEG8wbLarxmEtsVHN6Ixl+Uy4w403MnuYyYzOHXcgzrN91ZCaoHeZHuYlK+MRw4htIb9US
fX1atdUlwrHBByrnSbx0pJfg3mZXv6fEbiQghFYwA9odCt3E6aK1yofT8/RuZFb3YCtQzvKlTGN0
RORLciLuJ0uguwQfHtkhN/M7Fm5jd7wjAvc6MF8OX0yrKJgwyOf/5yxo0LO4TMoGRaqCe1MQ5JYG
cxLCBuODFCpzf2XoW5XgsdUCIga5w+KNVQT3fwg+9GkfI00tThmEiLT236rHVvp1YFCWSKptQPfE
UPPpFJ4t3qDS2ZaOMwSodTxa1CBULpCMZyDOFWmnS1RblP8flquUaOcMfwbqzVYnp3u3lUMMHBcF
sXSEknk2AczOCWO1If4WNoGaMsG6IbanNt7uTv4OOvEYWmparkNXJyamlEHJwhIYq7H3lv0RHppk
A34bOwtUrbbsQ1yO8SAyab3kJdzw6jUQn4NFx486QRNGOwgCqyD9lUG/yhnebLk/hTMtvzjsCDJv
KmeGmX2XefzPJSDqKOWIvYq7orSXcLpC4hiHanNy2g64rO06naZxOtitQROrWogHWRxKB4e8N1hO
bx/Ysf9n/6X2jesZ4m7AKgwgFieFud3fZwmktuU09+/QqvMwwIexJIvXAim6UhY/D1wZvcP3/NlD
m4H4YhXNnEiCmM6v8EnTcaNg2InJjBtVVifEv37UxRJr8uNXpD4v/Iwek7vF303A7BhZ1zpY5OZD
q6lWikdwG9DagMMRbrJ6z8LFOVozef4zafX7Wll739nM+6TcVTc9L7UVdaWvJtIxdKMzgxQFGyzL
XZhHnKI8vWFf6hIXIXfZBaoTJ5Eg6RiTYIpElC9K07hSMSSAJUN4a5vBgV+6PCHAGwj1BF0SWr+O
IbTKU4IMVE++Rl7exf8MOtODHhHlI0nVeKi3t8wcK9pY/oRUbWqzqEFREWUFHwGpM+PICG52JkXb
PrUSZnHfCc4cxU8VO/7i949r5y4NXOV+DIuTDbhXORN8FhBSX5+6rnDJ4NN+3W5xAFjs1W6fu6qO
tnUBa8wbhQh0Fxgc8sGrg2w4C9wo1MJmgdrBV/u2pQHsYCA0nDgyQV2BWcITg1EHR4P+S9cnkm7q
xaAM/jsxH1Df9Dksk/SkPlJjBl/YoKCVtBnVYZiBP2/5bOnwrRNLDU+/rUezeb7WRULi3+tyyz5O
GYmkLSRS5QlwyKp4i1fvR1OUKIDhe6W19lWd+M4tjsgeU5zu1vLvVoEeOCoYn9L7rDgTHss3iG1v
wdVWOC2DkL3rcaTfpSnr5tKMxI0B31J3MBrtQMLmzbLz/t9gpIpek1IM/LrPOC4q3uIa5YNm0rKM
7HGnG4NjmDowo7BFPomp9fClx1SupXxfd66PiBWGm2v/p4NS6vu/WLG3wHtp8Hc707PJFuXlwgrH
rQbWvbhydjuWavFtDchuZwVu1k0qF7ayc4iFoEaWQqu2y8YLyoKBvuu/iZGlNbUZJAIZGzzq9ixw
HkYuVLwvOMS2dPBzESZMo0kNy4y8n2P5v7Rx9QQkMHIHs1JhNrpOn/jwNBO11iRoqVl6craV7Dc4
TKTxUqMntcwgZY+OrWSkkNNJJPjFu6eNDMRyS0gmaxQQQxLnz8RUoVwhGZZaGzYt6SscbBnvURZa
YadGrAOCmOjhlf7VYRMtOjSLv0GBabdwmnBYn2M4OI9aPFxvntaeT3LFoZqBKqqVP4WipyMJYFHr
iA2lSZtH4Ey0j9oqEwB6YmdmOo6iiRqzlemVDTGsAHnm7k7uMjGhuvQEXumsaJIGqRTJy8pEJopg
Xn0KsVE0FzE6gyticV3oajKymwnoGTXKEGBduXBK2V2oVfI/N/tHJfHUCJnnJ7gv+21rITm8lgDi
evgCpisokFL0EP88jLN4RqJrdyi1oRjEMX4AJLx1ODs8qQTkeADOzRetz+J1hwa0v/v01GwN3Fmt
91M5P/lMPzJ4+dcTBiU/7oyFgOJqAoV2HP9XDLdL8/VxAofNkMYf8pfJ0JEbfca02ZdGhFfqkBUl
9w7Nu2/ARKNDcwzMkYcK7SU0bFYXtpDE3P4q3gxwll8zltJOxrOZR1fQz+LTwnbiNmS87kQdR+BA
t7mC4UGmUQvm56GQ6J30XuZFYoWvpQNB0c/swPr4HbJVt4IUUSja0d2WgufPrNx1BpfpcDCGE80B
BQEhRytW9Jras/dndDyQaOkDONRN0zrR+GO72S0iMLbuvSkxzm4AYp+kqgbK0n4RrL9oO88AUyYC
KZQlj7Tpo3jmZuZn3UguRbVoz1YKJVBBOphdxR7Foi+dCMul6RViiIzRXKgekgZX6lutNWKJ++Gm
GXlssM9SOamKlN+uMRwQCkw4xcYSWnyLjOZc+hFkpMUEc00+Dg6VcZuOyjCapDWQpGBGqU5EEwfw
dfivX7raJN1Da43a26GN1abg9TkY4SKe8fmQUKUp3WFUKop9OYk0gdkYLJAd4ujIoe23dnaUzSnL
Nc3T4zGGBWdMIQWKf0ekhHqIX5lMYxyzYrsUmJ+2YVnX+l0r7/yAV9u4ooFWxJRGlF1Fhq3cU0bD
2yRdqRaMkoZfAZ43USlUjWp10RNpnboRJ3G+4fOL1zdmQw7HN5wM+ElF3xfwJj5+HjOs9v18WO+n
iZI74XtWTa0U9ZqC+bU0L5Zlil/6Sdf2m/QtnJrlWLzDGoeYF/a8gdgSquv8r2zri20RG6nezkhd
Tk2N2R9lImhxdJFJ/SEoYVnMfU1l9wlQjt4InMdnYK0gtbyKF3WWErQKiAGQ6Wmq99UYpVFAtURb
PPQPNlHE0Ir/BntCJJy3rZNMhAHhsQqrHlSfBglyN+76cOKzYEXjlpdaGbfNx36uKdmIhchabw2I
/6Fh6oy5wXQqrhrMxY4vQiNq7t4pKEdsgUOmL8UuSTRCGu05Y+Z5k+SfHICQzdVw7FSLTXFbaj0s
VjQmnEA94j9ea0ZqJAT2KMug/mlX15iGA7s9EduYp9m3ypgU5bujAAUR81USbiNUDz9u9AvZelQf
78lB+ZizndniKX5SeUWpRX4F2jSsHm9aRM+For72y0iq8v0U2dngx4flDorg0R8d70jWKcZxARxZ
TzlK5dKGzdU5jMqNhSN6D5ck979Px8wiexJ976WI28Sh4I7HYKdfhueyCCSEVPaqgaFTWIzgjHqs
HUhsJ99NP9ySiYqmu6lEH0XyFBvXMRG0zZ+cL0B+GWHR5qtG4sMhjKY2XfZChcuy6lNQ8OIrKDPb
IiuXr11eK5nxh6qMKBu2i/I/hMyvD7x0tRkDVZudJVuYBx7tYpuLZXki9/DcuKQUJu0msAkioLeE
bPvxZXE2bR8Txag5CEsl/qWIw7gqpGgbHZkCbZbWHpOd+M6qqhh5B9U/susr4wZjN9IThfilEqS/
D5e7GK5R3KabATFCR95Aha3S1tGJ5FHl4lZwmVI7i4P/7VwU7QSn/G9glqapAedINHMUsA3lijDG
/3Q9TeR+km4PfcQbAoop4BruBLiAgO2VXaVktz1mxhcraBu2lMFcCafCnHVHEVibZjSnqgwo5W6L
QbLtUoHF6OHZ/qRKAZZvZjCaWuKj2gFhMMBSwPtnww/ZYZ5EA85AVgPzTp8NdH914mN0ATIUo6Ks
Sn2IerOrpf/fcDWMU60SuiC545PyMS+FwMGE1r5UvIYwYAf8rfaL8wVMc0DpFwOMwcQf4i4sdX2T
HA9Nd99OgS2zt3bFu/dFDE8UUnbSPH9wNTpp1CsHFGvAO0Ff16NLmEOyMen6f6dVNSshzIwz6tf3
apwKP4HrN7AfluYyezWonfZ8iRkOBEDlmvMntFMWe26c/5oNwLt5T74EzmBpAeDdN7NzIs+Hs6n8
RdOk85tp9/+AQavn5/4qWtc2rtu84yYbEdxYAmPRtYbAh5CQkl9I1yOq7xVY8eM5SjGrQw4pM9Ib
2/xTQg4StddxraujPKj0mVX360JpuroA/iBB062PRcbXgGEz0TBKGRPawOzQXBKqayequDAFh32U
KYQFiOaeTthjnf7R/m8/5F+W1drYOg+imxJo6EjXraemUo+PEcbC16MEHYex8bETyUl42GKT4Avv
6DwfJURKksDEdOd+IfWqrlt5NUO4oTMu9NUWn0DO5q2DVxYqUPVP6t3s4oo2fG2gfjMPfqFrv8Ho
9d5GHs2fA9gh81RID2lXIR8pxOA2UJx7Xjr0HW+frEIgmux+WDV19RF9Ki4ewRuqSI2yBFRWUz7S
49ktcZPwYl+FqTRTaT4ylyXglrCE+VLJQMCGnxtBeYffnC+ylMLJSf9H5ftE58iXkKPlfod8cEby
vO6UgQ2+0Hz95AecR4GKQOR7wUHwmBiUQcWJhKz6qofQ6jmwuFxoKXdWB8CcQMWgWjplht5MX2dT
Jo0Vckuz1KIivakQCLzYGnmmMrJOmDKDGKjSWBxsHO2ZhSO57251M/wCXFUn0uivqZpZBE6ANxzJ
Z0qQk82obJgfh1fiWvkko0QHVuYm3qvu04AwUSq9MgZ0D6Oc/W+HMPdIGh7HNtQssGVRDvKvRGxn
VnSRIbLMc2C9FHI5uLKELMd+B9Zy2uzDqvFnb1+2S3zSaSTsklNv0hgu9/NsT+onxaDMm3Zh5B2w
xIFFMHDJMyYnjgw/2tiv4NLBGCWzwKOJKXWA/BiT0bDUWZEWxeBy0V//zsWkRzK3DG08J0A9tW6h
79gupqYtRVuUmEGhYO4gqNc//Lr5rKy5b/svybSvURy0u5cpeHBkWxQ9olCY1LXbmJCtNLSlyk+4
q6DF1RYpWw6MBCokLtYwWqZIDuQIdN49YQjRNDbaqJNJUQRltUhoQfSJ7vzBLFx7HwaME/WNJNpe
v3ATVULljzEwG0Pfhd+NRhHzPDlYhJBns7gcobMI2HpYh1yClK/7E4a1asCaZH20JIQz3XmgkLrl
PPIwSMbpCTm8sc/fdMiWRVoavE5VAjTkR+d0hcJ0oNBZEFfHmg71u1fDlkgvKBEv3x01mVvsj4B5
VXXuY4bYBBsgGXkhw9xaSLTwU1ertINsZs3xw5HZMQSoVJWVP13pqwU0J9L5RsNV0GxRNGiaPD9K
clGNTaQjyPEvcO6Tmn71OWv2tVFz0P1Ai7c67m1Nq4q6ZQzF6RrlujuKSuzaNQQqiy5Mnaui3XKB
1BVnCB3L3bM8wwOV0G+u+lyYcRsSGRpU0ValnH262rjPWcsIaFughZZzgemzcLSFl1ayQJZrhPrn
Vun/pDyQeC3JoKYv18hHIbulNapdsHVyvJf/uMVfaNNuE/NxlQ+Fq4av3qfLcehdQKE2IudFXtVB
BfxbHOhMd0tPDlqT4OjBz93OiJeWYa80LTE3weQqZpZSNy5Yypq1NfkHUG7DM7QgTTn25UEo+aus
oQmFdWHpadpUvIjwsudZ2aruVYvY3n+LewvCGvz7r17kV7vycvwHFzFB8zzlaK91flJP70vxMIvF
jpdAi2e08LlET7fAGWPvRtQO/EQ1t+lzrPbOTK9mdzgu8BBF8f7bK/1freiEp3cBfuTdJ5KEddNQ
Tubumwd/sJKUulUTTNajb1XV/0VlqgiefD+RHs5n1ruy1/rebSuLBgmFC0iMJdBwOxeAZjYeXljH
YauFVYQx95cG5ZmN/lE8MhOgQ6pE1mi4K+9m23qgIHHlfi08h1b7nyrP16rZcWiV/yTMQlz6zZV0
8SPQ69iyzMdW035hHUsAy8x6/FljYoEm8/fvFnGyFY4Dk/zIZ27Nc1/I+C09d6hjC4+1pJBOUGEq
6p3ztf4np9QPiOKRuNn2uBPckSewFqX8PVwgoc3tdZoCPoZiUufaavJ8oMNg15/4yFoVGnsYCklj
qyjJtfnycEmSQAgKXkilN3m1N22j4HFEOoDsKjhj52bULX7yrCvWJFbbr7+kZ9oS8dS8q5lMN48U
2bOv80m8t/03FHrJD3g5kGZMAQ5eijbRsSnX+0xoKxYCNMxd9ngI536pdpeHn9Rh8gLAiqoJT2pV
VxqOUvowEsYv2ueiqBnqsZf3rJXh3UlEIZ8g3oXzOy9A0WGgpTI1g3Cj5wFpG8UoeBfcoCBj9Aww
ahPz6ge6LLK3+d98x5ZkZ65bgtpINexVNC0f+ib/AixK7Mp5I2kOpcxAdu53TM8ps7RlhoTzecJL
13qqPliPbWYIoBmdDhR29qu0aT/EJACSaIeDfer0uwUHD86vIBubRbYOwUVx9C6fjRdO/8Kj16DY
PzrjmgtG17tGlXbrGdyIMUscnW8UcpfsNbisodm0rYMmUc5EB+KvrRVDdiiimjdck2De11dMrtgf
QO49x2sT/lQ88xsYaBIDviLR8qZWzZzvU3i7MRD8ucJZCOmmixM8U2YMd9UNc0If9uhY5aSLC80M
n9Ru37sI40lEO/kgVCBkkDXH3KxjYk3Uy7+/yinibFLLfdCyFeL5pa3BnYvHuGhddjzJK9lT52A0
fCxAQeAMC7St98pgd5QUY9cHa3Xh+69DexU1XKxFhoFQyMjf0idk5hs3OitzTbuEIPaPRq/oasR6
FdOKayYLdrB1wzyKX7nMMdvMYnfzobYgwuCsLwMo2+/+2Uc9RPp8JGTIuv+A+asgr03HMghMO8zs
vth8N4PnyvCxRO/1ecmeG0b44FgF6/YaTdtRttWOXgMVq6zBWc8JCYdY+pfYM6USOjZNIYpq63fv
H4FNcfvZsVpozRHWdbpehzHLjpGuZXwNu/wb+G28OE+zJT2Ub7KvlExiF9Cj00pmSfzVNo6WHhYN
PbP/STNQAgwTUr+OMlF/yGoKUp3oDQUshN3Nuxt8lJeLHcP9pW2zkFqO0+vXRJB52BboBhiUWqfq
JTmUrpDQYv7d8IUUuHB3HCe5AAwz4+QhP7/psTVUvsOcv2xYcgyPInLMVujd51UbmccGTm/a3DdZ
rMKflZa2K/EPB4PpeULd8DavJXXIwSm+xay1FtFmUp8gKexBJdeNkZWkhCEJwXFDxRVuPyXnXplD
kXEtBVCv2URSwBBjxQoY/2Qmim5SDq568C+Rfuqkk2v8cIB0eqqriliOd/kDyvONeZd4WJLaTLuz
248UNGsKuzRf4rsEKZx2V6HTg0eYfoyNcTDYTvdzPDySorv3FZisCmxOko1vcVPE5CBVogaJZ1Zl
7z0e+TzNeAr1c94MJS5iE4ls0vXJHo6HQbIrkG1L1ZOS2xW15qkUQGxcfz+i8GvTl1NnYYQURq/N
RVe4424vQd1mLfgv2Y2BtVZQ1twAbqMP5AUGkKG5EppFXZFzJhoKAwJPck/7IZlwOSUc7RKJlOco
TnIjZrcXaEQSkJKL5has2QC31aTYwhAQzgzzMB8yvKu14d8M4Q8yZX8ojg5YNNmGwuR3y7YGTg0n
Q//76pWFt1DfBUNvy8nXsBIU/vkAKfHx97IfHvNda4WF5K00OCd0roo5EExQHmImUhEzZECNjjeB
MP30H5oI9UM/brHnuEGAqxC9RHvwGT9YQVtQNURjPjROA5GZTarjlt0/tJK+ot0P+kDFK/Wqe2Hb
l0rnReaGzR7UOQgK6CjomrfLxvV+wwwcWVmKUTWVwrgNrt9b6S/gsSPK6di8J6bu0HdJxK+9WQ+L
RBaPPc8guA/l4d+Ety9X/fl3fWKosPEG5hH8k1SYgMZjDelDHZuexzkDzB0LMnMqGKqQPy97giLN
vPg9MzcDX2Z+YzwdUh/341tS68SbeMCrpFCgqh8oKdWswr6Riqb9j4ptA1Sf86ZaFq1n7FjW9dqQ
X/mJBk4yOCwDOZ0rFoBI9FiZxMdvgRSiSApdeFb765hXfLNuK4hAPJaj7meAWYa/O/+e8uonqPiq
tOp7Sf7MHZs3Ik/AeRKsLtOu4erS5DhaFM9UclJHK3O7xafuIWY4HHsoMFMmV+Pso0C+q64mTjvh
jvivIMC0SyQBYqD50MB39MSMorGQUzsBoemS8tj0cZxpwig1W0Y1DFwq4hflBK9EMTwyZFlWYJI6
OT5sJPAtu+vCxTfCuXAuF7EFj8UR3tOJu5hXTagyB2XfZlapH4bH/6Bk8MKrhjsOc5drA6JJfgjg
XHNIsVvawcySt5ILq5i7OFLy68f2Or0E4z8gDwFTcV/mgIcMbrJYXDg4QLHWyZ0/RRGM/l/nqhgc
efWEyczk+XRrUOb6KLMVxk4xoKdHECXja06Pc9RYsDhB3Lw5jGeZ6SN/guBJtyGwkHo6LCja1438
5SPTR6qS3YPDRQik6RifbsYao7k1UVaGqu3r9/t/4gq9aFkse/8Fora0Xcz6+mtzfCdrdjMfF72h
QWeAX9UUSDIdad12YKanQx2tG8e659TU8/E+Qm+5tWH4KF8ltCYPBKXRSxZ/pog2qmsdxk2lpwC7
tOb5F5XodZUxyVEYCGbnInSW9Nl5wDRzLEaypISaymmTr9Ek5w0UX15QSccK5IyIhAxx2qdoi6Qk
cEC2QGSegSHoj1536TDuFyBJALORGrD4lRq97nAXNyxSBNC8NH+mfMi2NQfbc8wRA3yg4JKQXR8H
Vcmhw+bmVTbgGjS41s7Rw0PAy9WBW/HiOKdL0hypc4X/EdXXKaT0qJpUFFMrP9K7mgWUwEn9tmU6
M63xhVfNtMu/JHe2P+Gn7SxggbhHJpcr1pbh3eKMwSrmBJVm9cHgRM31aCn5vOf9dxYTAhUCphAB
kZfERZVZWDdywaB7onmU9ug3uK4d79q0k/RT+zW4WytgVzYApgnzSc5trpHhoHiyplHHpVfPs0Vl
PUbUOEs5OgGR7s8QF8ZcPcAaailw3+AiQP8bpWCMLZ3vSpeJVwcorMPKvWeEJccdhdMDGetkkg8l
pshfj9zURcHeEorwpndGxwB/izW/aOgBvEe33erjKRbdNhMulakMEOvahizoZ8KOoYeBm1gaju2N
2uU6bh31at+7eqVf9fka5qdyXZRzbcQQbgC9mjT4aQH9v5kt4T2LmVN83O0JTX9JIyw5r0F9Ztuk
aEQqCHJIawPAfjE45jwuAlRiFh9tXMlanFv8LDAxQ1j2WiVCy8Vcu/jvVIYEODLCxsgWNeuAn31N
m/ybvfoKNBEV/qh2pGaX1mnHr05Z4Y8dTcH6jUdrtVoPvyMrq/I50vJYFkm0x66x8CyljmIbJHZA
rQhDv/DjTk2pdm4fjxnghUcQ+gGU9R9nAmZmmNYosq7QkuwVCCVYofLwTMydcoxhlzJCtaa/ryQg
nYZCq/JTRcdihe5ghhvgbc0RFPMrywtsdjz8zF4p7dzWcSogWGsUQqlprZAPK52/mGQKzlA8tqPI
AJ7TLzB5V1Rvdvji4T1fEpugn0Wgn0AGOGsGbsog9/PMRLlDp8fiP0/ulVeRfiP1sOcEFWM+nHPt
SQT8orPkZSXe+tk7in/nnDcYGk7oJXPXJ/xZqaA8l/y5LAI1wYaSGU8dKL5BIT/e7NyyBLNZul6z
DlWaTPHT0LKVz5fB0jGg43GkCDJN92S6rPhIG2vnY0buKHiIuH8pq0EDE3ufQHYqz5N43EEGwtdE
wQZ/iBjn8/9Nbj86TkzntIjqdzv2jp3X5+FjlvWpt7X8oRb7R0kqAuyle+6bxvPBuH0W3ZYPbeVn
lp606IfM5DTRC8g1SfMk1RWiLy2Tuv5lc65BN0AOE4VEZ+kWzEBHSaeabxBNkhcNI/NKEBMlZYPl
XjqcLiRzIZyP8bT6QWdr64duCfgyMzMyFaADmamJ/SefJ8RG3J6giA+1gsZknqNmJQcxbfpzk8aW
n5a61UqDny69VNvXtlvVsASP1Irfu/XSJ62W91+EAFvTdxNWRsX4W/56B8aKZjd9aSrUh+ctOXSx
yWp61TqUGTsovGfO2sw2XOb+01Gg+IGsvvQN3ER9oFciZ4grfvCJB1AtPQANJYzOsamb+0rt4TwL
vERFSO8XtHpSp2swqxM6G52pUY997nBkfK3M5S4cWsWNxlA1LArvPj3+/2O8o6Fisde6H63UOnNF
IiQW3jGlY+AA78FTA6K2f0aJ1C9BETiurjfUVVtz1L1Xq22ewcgcbGHjRCPlCCNZg0RxtQ6hIvrw
jJXOs7DuwhrRTAqX7290huOZNX4MotIpbsSs7rA3zEqr+3k48YJmoz4/pLlo4kiNhsHcrZUCn9ua
mOBGyRrieXfyzxeRqT5pdWDGJjgM0KXKLyXvIPSa4g5W7VTRkYMa6gzmQvYq8qwfZOApZTEDfZLQ
/zGRUnvmtJ6Q8kIjwk03gffU9GGqKAHPUsXmC0yvu+bH4rIrzDVqYH7BHvdGwtbrrxoLF25756TD
4nmL519YvyKKlpEzPJwAcPFTNh/7Mo7ThwwfIFOP5WiP5dyOyb2yhnPQFj/h30VH+UMB772cEvO/
75jwa592mtJz5TvDl0YUPSbKpsHeQsn2LK1fIgjA+AxSvzO5Sx3Bvhr4XNnt4wXBYShvfk8D3dKb
L5UGg1f9vJDYpS2QLQulCwxzZGYEI0tzWkvJp5c+VetnhHHd/fTwUfkckQWQBm6OrAfUab9175ww
h7k7m9y9YsmlWpIdb0IJfh/tIiRd/GAUd2m7n5mtH0dX9t/vwFnuWf9uw8ZNJLDbZEB+yDP7CIAX
Qx4YJvy0JvUYrEuc7vEtQiTajmQDd+/JppdMDcK3LcWBxk7qF10V+4PVfj866gSELV/YQLGm12iD
V5aeOdW7D+5Gmr44UP8fpT0+Njk6dGOOg4h5piGvs6d5raz8WfJ1jj19yA3QdCNS99u/DBDb8am8
yXiXo2AfffaK5Wq6xCM1BFOsXsdCVD80/XQOkHMyYXzJDLQPHTmucTcORgrxrxfe1nmy1t/I5Oyn
qHKv5VBx4eUkOeqZHfXrJVEsW5h++5RZZ4gV+oJdQ5ENdyFSvqPzS7i65qRxm0Mw3Z0lFgYqAiV/
gnOx/VO6ugag6lIZKSvxiw66FigNV6+gRJ0O8VoEzUyyRWG3s/BcneZT6IM9DYHRZZ+sMe/VbdDT
yKk6cKhoSDleP6/NTho/qc5gsyJAxp/wwS/9KJueB/04+aPh3VeO4jzsXiMNeLlYYIVZIzQegtrw
dPDlj8stDmOhH2iaxJN+SJmImd9HFByCT85LNWd85Zwcg1svYTMAw/bpfzLrMHnM2VDPmAhzRMHU
DVikulTkvll9xnEToGTDWXuyLGYCEQO8O45nM/1HGBVPi+LuimhOCWstO+fJGyTlB/H6delC8ViH
aV5ceeMwrX61BOwfwKx74YwGSSxBfqjQgRQcQEnN7yPaZ/tY92eT96bVAHneB7KXFgRQYUezVMrB
U6N/u4MD67/SnzHWn68h1vzdvuDVbVNmQtNwlrbDUsgaz/kSG1U2wM2PnPKXzBG8OZFqKJXe9rYt
PZF45bfC567N1AtC93u8twqvD/ke1r6MGyx664be0CLQEAw6n6YuDaBoGoNGyeiPFBrojB/ZZP8+
so4yH8+bO9sMJax9Dq3TbwtoTjebMyBU/wjhdFX5dozcFoCGCZJKg7lVJNQzGZ8D9/mij45a/ZEW
bLvXi58NRkO39QZpGxUW3eKmcXrdN3Nd0PuUeQgS9dJle2KWUfukPtMRbCRQvSxfD7wuoH/s4To/
ZefXowhV0rVMRVEEsXq7p8TZWSnbx18KW7UOPkvCBrj7ol7OCQ+WmwaTdWezoKicr/FyDGphVM54
rWJKe6dyAZ1pZ1Posy2ngC5nIOe1HMRN85WDplI+HQo3QxPjmh5JywP1X5CGVhWoa8H7E6Sd7GxZ
Z/jRHY4weJpqEJo0uzcPhwgbIOQuExin1mQRKXlEGQeIeGHBHfxwedo7PevKxqMiXf24j2Hqa4rR
q8qrTgVc2pqihe+dcjPA4g9yV8OwQVPKazOHBsb46oIBwf3CEWsKa7qHRzYt4pkuVIYklylwAkKL
OBscpolqxReXA982UBziUx/RmqqWoCbxB/LwAK36/GlcIX+1DgPPtBOhRFfpIdYPddzQsUdd2q1R
lswh5KbtsC8P9g5dDe0aEFuvxcX/FArJ5Ik654He9eV7NkMi3vCzPJfiy71LOc3AbGLdstKWH5Kp
ccXkmIiUDwTmH2t2ILNLM0VTVNupYjN46LiJyKmOpkLuFJTpFTKCAes+QdvpXQJB/1ptx8y6Bdbk
2K1vdv83hMmu85N/4679tBoCzTcAAVMgj3IlrKWZAgsUTZkQH/4VI/wrmo0Xp3L3FvdPbFfJgA/R
VHu5oYVz17IJiP5zfjmpDkWjuG7O+SXX0lZJrTwe+1hZvCCj0UatS/dqnTcfii2b3KzEwi8DO2Sy
zH/gvHCtPTesW5JZdv/59XwlluR7SzvUqa2JrB8edmrH4VtOB9SZ2999sV2Zm3sTla2IxtZPgisK
dW3wSXPT0Z2kVQqPxG4wrl7vygJWhioPwbSiTACDWJ9sA4RmsFrgIDn/tRI29INalsbRv+PRQGZe
8E0Ajou8c2CUH8ckqG5D5FVE/MunzrlCCcn33Oi29Ex04B7ouCjHW32BmUUUqfsUK2PGskeE5MGg
IMihahj9LTUmkodx91aXDICyO9yZcxqHRhJ+HWDWeZ2BSU5rB58nwl1rLJQCJWvNePjJ10bxQOPx
a3Is4MWNrBWqkxqpjSmXy3EBJ7EWJI7BHy/qKLDyr+Il7xtO+Md/7f+lliEOTU1cFfv692lvSyA/
8sUxuDftMee6cRHuC4vaIe6H8J8PSlIjGe5kpHe+iY21pX4mTip+29fEApOsjnbbhgp9AroiiguG
Aw9kspQbkWBLLIgFTNbczghiFA0fH5MgXnvCTdrF4rECC9qhBHOCkEkMa4Exthy5d+HvH33H29I4
aAaKBH606a2w0SB2jv7eEbuPpm64+7QewnDuXpPInwEjbvBPAYTX+aynijTkRrAG8NRBp0dKzPJh
mOYKlxwzeFhb3m/SgCfcx8nfN2cIOJYuS30adcag8ZxDFaWlXrL8RToAyAxY2Gb4Q8bubcpz0+Xu
xmeE8QfxDg6Te50zVOjDqM6zoX9eskCZnCGCsyjQ8+qYCqQDwJ/kjAJgOX44c64lx4iSPKLlYlHB
UeaQNvNedzRYDvXth0y4iiZViZoi8NPkszS5o6nCVrK4B23Gud061nDChEhMZxwVWg++52D+xB0u
6nN667Tvzx7mc6B23RcwrF66NyyBVh7OafxbEKP806FLVLARLk2qXI8J4oRvPGOs2Z28Xi4TuChq
xvA0mDQQISyp/t+/abDl20NZnR29Kr82aLiH8IO6/yiWjZj6a+asHta7XAkING7y9z/hpTnYX3x4
u6KIcaVNVlGQs/hxyg2bqQRjUx1FByp1Yn/DFlIm/HPukCD8LJx4lKGt3vCzvYwsGfPk3Z4UHDDl
iRxD//YWCNnGk3jEnjTrTWSOVS0jV0ffw1nAtM4f0NJnJ20pVtu7CcXlNRo0nttORSpJUScEF91k
GOlqrXdv3pWsG10WPKlSjc27rbNnYl/zmwCekEAgv5GfzkV0yIfLKlzJBW/b3uWMVaT/X1zoPJfA
vjf8bCWKqAFsY4Wikmj+t4xdQScC0IMKL5tdKrHTqU0UnlNkX9PQb0DjMSwSQ0twL8JOLMjlxDs0
XWdd2b9Yot5Npg4LMuwlsQZ7Ce7NKujO9gFMgne3KTRB3nJVS3p1CZrARmwB1EicZ/Bb46LdIwpj
737+K1Ed2wmL+8ducsozE1GRT6fVxvntbqvptfwKf8MDWMDi7cyyCdHEUBmWj0X6lRTOkJLw4uNR
e2SrHYJpzA+QhVf+sj85i7pXOMTkas5rLX67hJNOTnajRHx8ItGjPp3EY4bC3oND5fTniiHq+VnS
ub8gNM5uQttUitalyC+MXK/4vW97+2LLEp8K5wkY5Uzv+3MUe0NGK62BL9D2aBqnflIOEMn40FTY
VPd2rYcIdmp0Szr2TQn0bMcUb7dcazpOWRQD50tyq+zvqyd3VQbgcoE+tlBZ8PLc434cGa4Ws2dt
kvOSUq+EnMfFpZ3KRzDPatjYIOn8nHEXBuKw9Sg5aUelWFd8HKEAheD83+JxcIVXPHWRfV+23K4i
5RgwFTSyYAAGlFG4lTY8cBlDCipUoqRkU0i7dVSoJSDCUSqIszalLCUVuclChfZrxR61W2VstoY8
uHEFcjHrQSqo8AdasCw3NvsTBV4Bze7kxkHTWe6r6lU950nIj7IJl8ApnpRQRuVFA/9R2hFw646c
zpmFJnus0IE3xtnOcDno8rjsqcgg2hcCDb2c024lFjSxvxCqVcTawDf0Ko/zk10vgoxv5Z/ybrS3
RXUVghaiKjvF7gesclaPjtBAiBXidQxAwkfxggtJY9fQCsaYA0D0ock9cO6hxneg2OF/uencZbrC
8XXR2ONjuaOaDwXobTozAJHC635slwjCrRA9K8kAPKziRJO6H9KYX6Gz4pm+3KIzKL1CVO7/pNGS
3roBl/55SS52voiyqDjXy397MdbWh2dGi5X7QEgMfrETNlIoNjDtg3Wgo2s8sx2Eo4gTA2MTENkw
W463UUiFSXMPDAtEr0yOEJ3AOu5z1Df2Zk2CdhxiRD4nTRwodGpWviB3imCnKnLYPT6k4vXcc0QB
m7bX8A647thW+5b7/XchOMOYXyPgINaiIY1fASbW9kavG4a2rC9qbWkAgTZQlwbLDsnCKqmJpfkO
Ef4GG5McCU1yvSFAqknyyBvTdItHTWZFPF3dPXLu9Oisvyd/OU9AC+7TH8vYddFV8Ovb8voH3t14
EbgzxlhVxLa4wrHdQw1oYg7fju18WlpjGy5QzMXjszIiFR4qOSB9PfCglt0xpMXYOEEd0Rwota78
8hKGfnk57BdTxrak9ciDlC2NN3A98V29/mcyeR9dAkJbOpJIBuhnbur81DbkY47qjXwkFL7bCTs1
MCjMtUJmOCLigXBUInEABZARN1bKNrcCJsprkTKBjv/3/BVSBolrnDovjodHaLRXtd1490+uM07A
bTSqJpmJALWNoRkQKUCfiJGFgyNI0/rjAK9Nawt20uQ9kHPrwvrJj4aryvq3fZ3jOV+PoiBwllG/
UJPuu5MDSX1QYfmQOVGBrVu0ng07XqWcx/kvDeKGjt31r995f/tqvltphfqIPHqsFPUk7mY7cx+d
7xTg8mNp5FlQyVgW7xOMnD5Cf5N5OPFhttmR7PbN//K2BqAlpMTI1xsVJfN530r2KyfP/VihP9r3
qYhfzeYIOY1x7pB/L1p7an2rgA9qkRHHXQkCe48sYANdJwbtOxrAPj1goULP/tSXOduzDgQ1fKf9
v/RCwfRHsWRzBP7jR2/OE5LhnjmWkz5R1UmVvt84nZ2VVDNMMYU0w2a4AfMl7I14mw1Atl/rMqi3
AJF6GG2gtQ+ZhME3D0ew2UFlC0gCJD7qE1712BhDhWwweB3w4BCyJ9k/jy64CK/Im+PjNQayOJKR
s5HAPHwg0a7ykaneHWAvfdDC2Oijy96trS1NrIaOP3p674y8iOx3W1L4i/KFjSadhhkzQEvka2fB
k0qtmYfPbcLcTqwHwWP1f12j/EVJCqDUrHi17/RCMXl9a2wCir0TpWTAeYlKoAsgtLLiooH2IYhO
ElfYB/tnt/KY4QJzioPBLKc6UY0b3lszMMIMdJFGzQBWuNUOe7kknC3Nbd3GS8W9ayCrZoXEngrz
a57aMTyRY1VqZ0qwd6j4tEhspn+AI+Tu1Ai9OqOJdekSvFYAAcZho4A9+qlNFSs8d/WhgTgTuvzf
1viaZfqC8RU6YY8Bl//UxOod5gLj8bJxQrCTDwCECw/meecX+Y4yI2Sq89nfLxtWX+rhAmLbg0Wb
Dm982Xev79JGKkI7WEbSdHbwzdSoOmHgzNO6I8h9cIBuWCaamhouiwOBY1YMDT2XnL/0l6nL4/W9
3tUyUeX9xXsHUE66P33ofPzQWQN/KwpXpmHtofnLg9loV0/ChoGDJcQLyXMckYChNUUVjPD1WBZD
5z6VFeHs7JE/CnJP6jQe4JFmiGedCwOO9lkY64HMlkkmLaoc+zOUuPkcZSUw60qBeN2h4IBdovUL
EH3a8c2oMq4N5I8NsYkMequs/esakBANlIvRziCWugVboXGRzXcgLYDT/hJrVtmvI0app3d2Z3on
v0GWVr3Mg1O8g1Hmc6gfuej0a7vw+76AjeLC2iHvjPhqAZeZWHpnUW+FBI4KKGGxsZW0L3CkX+vo
sp4XBQKQg6SsVDYSoi6T20uVhlxdfIn2kW68y4Gig027JQgVxsquuFsHe2Sw0s+tgCP64yATXfd4
SY8f2a4AJwG3A9fLiVsiM3oMFmmotiIldne0s5Pqo3Dh/cBm6IpxNWdABLNxN/Az8VDWcJXim9vU
1f3re3quJ58EyvTpboRco+xhPB2Pjh1zSdTsBu2GHqsibjkkIRJY+QYr8LrFOpcncW9AkbrpwDCr
ClvJTFyH3BlOD07OaAKlw3MV2QrqM147S7ZC5SgBD6Ahe4ut0hQI2l48cV4RB4MVhdbuboxCeJB/
oXueg2e0Z1fmXSjr6VIi8Yhn5NKDOIHxZQJxP86l3eT2sitJbxdf+/uv2bk9ev0kdA4vv09oddEk
m6W4iXqA21nV0E19PU4WVbVrcMzffUZEZp+8fzMznRew1hoWdfPVFP05Ouy3mSY8XUdO8Bg4qN2n
P74cnzXWnlevZZ2lyoRNNSGc1O5dB6kxxB8led26tj05rRJiQXANe7ESCyBmB7oBSFn4MO0A/qoU
g6anuJiOgAVfGJgrBooc0qEigIeGGpE/lRDWc1dLklpF6fvJbvontC7JNt38N+5dcHMN/NYxUr1D
WAnZQ09pzcyQhVLEHtNo9QTnE5fdIw+8PeUJ6/lOZWi0jJBE2lYkQzG2zEUKlw7EPBx5A5VCrRBP
FX8IDe6NT4AuyVPY0f9ZALBvgpKqEpUtAJy5NnYAXblfG2RkLiaqY1tkfoa5iLGL8IEm4WEZ+tgP
LikgluFzZ0eNPIlFW+WnKQa2NrnsweFHwwDbGjX+yKTe1rZ+xusoMab02Oiuo1lR+D1gBm1Lij2r
17aaqssKSR5hLRn9IS/vSv22Jzd1i6MqzgGmTYVmTU88Kg1ejj4YVKOzEATtbPDVEVFa+inivuC+
6UynXsVFTUqPDm1jlw+sUN0sP1b3CxQHPaWHZKKgETLp30+1baEf2E47MS7Y3IJWQkCQgb4FTUkz
8X7y6wwCixVPYLI5H9+HmCfeGOyXCHbwhAzUlykEiWl3sSMOKDOegDa+rqIZbmk2ZbUNPYryemdN
PPgoV/bq0R6pwJ9WcdqHtMfpKrj8cxgEW6FtXjfI5zqCztLDB0CzdTV/4s6o3S3dJ6/Z7mceMmn/
Q/p+Gak6sFll2pMgO21TethTAhN3WBrCoONHki1ENFiWfmOqdjHVrwD+l2rcGWuxPX+h4+N2C3m3
+SzEqCvmeGW4hbvDX39fbwvyq0ayqmWo7VFe3SSLQ6Zp/kSuh7+kTOG8O5ctNMQfxoFoyHWWJHtQ
Vr7Vbik4lDGZW6oWm66ZNPJh9yLTSnCgyINC50wDOBwLSyrE6K8oknht/XFR6dowpWh91p7Fsqk3
MPwMYZ21UzYA2Jtcf7hfsvwJQW35mT5JrNSiY8xwQwTWxifJrH1mVi7N9wAYiZSLp/AsXt+LT9j/
OD7VnbX4TRnpqLDHbrwjmXiybNbUFb4SoPp6Xeori7+0YXD5+dFY1kHhhomD5pwYcOimu2WrjEcc
eXYfS2jCPnd0o+fIZHGE/0qAzBWvAL1qil4l0kMI3WZawdRsFROz+R0abt7yUiF8e1cu6u4eXb13
tnVpj0I3NmwueH6b1Fmddf1giYFaKeUeGE7Aowamfwvac+uQo71VH4OOJ0zJtXQhAuumS3viLYz6
vJb+4isCeBxHhbnUFueqGOVxhi9xV9YRcJ5Bjn5kAOyUmOrFX+iWmaFwKb/t3411OiT2FaFL+IrV
XqX6fIKD9+yG6Gf5aqDPoi+aFOdjKzFitH/rIwAHhleE19PBvblBRJSpo3a2kOyPjXZun8rBjVGW
jHRWigaMt232g5JkUyEv5hcGGNuB+lGLSJLEGa5aHX9gq/Sy+6A/t8vGQ7VdOb0b0fUQf6fpen8b
YJ2FpbnLeVRA5BOtXYQMLSCnwLZkuJFsLLPaplNzVnm/UShgQQNius792d4Sb+wmbnDpPsSyutID
4CVK+WIst/nufgGUiFVKo3IypFBAr9YR0XmgIpKvwl0oNY6Mk1q6gaYT9Tqg+LCYSZYJWLQpuUWm
J8ZCLZHRmO7F2TaYBb28jRJraVG0/xihzERc9gbDB2e8DJKh0rPkIZDQklf3hOFn9mi0i90ghr9a
KGFLhaHKO/XLV91tMLXBOfJLAWMt7Aft0gNwxLQG7+Ax/hevnxJHu6f06vhL5owytrVWe8SLrNVk
vPXqlTsnBbDqydhQIfItI6iRm92HUJry80N7/+Zq/y1JGVyJYJXzTwMr0J4pnOg2NSCT32wtPxpK
VkUqbidieT7GOy64tzpp89Gfo9E5axVtP3mFkdFRqXJSOg7jroUOjkl8LlOx1M40dtMwcYdLvriv
LKz8fCIc0LlnkMq7BoEJp2izEciJWogVjXooEGf+DeVbb0UYgfJR8bmR9KsoikJCAWA+kspqOqv7
1D2fqZ/8U9aQMed7KV+0y/ZjD+NAe0IajwHpPOHEr4+S5cPrRIa/hryD5FezOCKiAOE/TsVEx3AU
ULHQybiJVZpuYieeIlGDlOyPl5LNwWSNbUvdeLdHjPv0wdb3H9fOnuEorfyQqS4HUHg4uyDPpu2q
EBUoiWrbSWQWqwvykit3UNuU1zSrbN/JD/r7USlMuh6xkgJkUbwmI1xAsdZfo3idKBCJJt6Ivqar
8/0mjYlor0KfEc4AQN37SNqUuEenb6knO9KRdprL6NTAecd0P7c7OsesX+YKbuwItT0DEOkwbbwB
75zkpuY3SxGgKlHSjaMc5RQFIhhMB3V5uKVDYrbVvZEl9fDN5HsIr3YS6XJdNAV30bt66zMRZGi9
3scXZ82tbhoLDofxgwzB7kNovxVycrh/lCL2Z5RFTYWIOC5xadl82swTbNSfSrxVyu5rZEKe4E7j
Lw5DQNrG3ASg4ginLCXPbGXPH7D7NMYABUVbddX1307OrPh/JM+z8FZo4ALbFvr8rQqV+mHFMFTr
0nIKg/Qm3zhdFdrhPntZHOOq0jvOGFHFmuYWLauTI8b73uFK484cfj4TXeq23MSoqkmtWgj2fR1Q
OVA0ZL2p+/S0ia3tsLg5kl8cV8drIp+mrYG6Q4ePWKL7roNyhO68K87sH/zgFw+IkkczfTQSuyJL
mHvjU5DGlmnQNn1g2yLAGiKNLAvM9Ca8e3OWeLjl5v3DeLH2IWWsNk+5/OORzZEERDBqHI30w/MO
Y+RyYKZAiOKTJ/zmfOfNEzzuTLAscunNh8RQOS0F6SHp79yw6gdciFWcHs2AhNtR+/3ygSqi7+S/
ZnIJrqgPcGNq2IbV7zL9duVUhmE3ivDdumGIwWF0/wKBO6te7WAVGOXuuQeXoMCvWjKIOyh1D4Zw
R311QBn2I9Y5+xMp2y9hmNavNBUjW1S8bYG0QP0ZFxAbsHf5lIu868eZ0T1WiC3y6GdwEwD//s12
piJn9quE4MXHny/1BCK1QR0WFabqF4iw5YBj9uMXhc2MVMLA4tFVSBwx/ewgtnp7IuZdT1ACNMaD
stTeABH/CkTL1eJ8DS8ohMMrStWD36ycl/fXc0Pfq0Zx3Q37RnbzoB0NwP84xh7R9YCj84738LZY
irc2d90V3irkaI761rRRZcT3NfB2ylhv5k466u7OVKQWoKv+JKpIEuZ3pQMAw8ahNMxON5WoyIhe
vtCXFx9j4gfrIeM5eIJ1IP62fPgiH1yux61XAFvaFoiLiYYhsXEPECEhp1ncyqZXJYfsFDEEA45f
iZ+1o/i04go03rBO2J2s/pgKXNlNs5pOgClGTcArMsgGWpelK+UL7fFtVNL1z7Drus228PLZkvd2
D9w46XNsF2W8oxNxpYEH1qoIA/POfp6bsSByZ+P6Bqq1AD272j7RNyDmN1Gsxy7tuyvPymZuGPOc
FYzyaQ4TASj3gumwc7YugXVTo6n2woSIEBxG5ZXOEgsjmZXUEnAl4lh6BFejiP+G/kOp3JYUfGbp
fITauxv3QIYAIMzjvxgjMBLGyifs4KzpZ/VirCSmk2JKAfaD+T5uRpWwG7IVifpZxyJJ1xRCcNZ3
i4RFvUynU6R8g50EK030PU5Bzp1VeY2Oq3z/HX7ilLFZsk5xDPYKQ+da5qkShNLqWdI4yYh+tNtQ
/G1fKu0Qb0VnpH3AsJwmazUUusWvW8enlROiRdpyD7Clsl8+6uB3iiZZSfOvEaaFGhV072AgQshV
9tw8qqKqsZSCCAFjVNnodaMrkRWReV/X7iApwB0k7A6LmZFaj/Vhp2tTG6+EUXQqwjMoZGkXqiXD
EjYUHHw3rLxfLRUNO7qwrEorZepN/HlB2o+lDG5T3CnlFi4sg7+uyYk2qax5tJ045cERv8RBGbdv
5EkfUsTUpBpZOvBcfKt7zWRndFEVc9YPrpty4s6tcBHbYvL8KquxkG8nq0KOucM8YUA835KDS/ES
9CtoFra/RNEIDvTccnUIcs2YigMq+hqldN3/tPOSkmJcDAD6NEv7z1GFwSd7FdX5g5r7uutDR7Mv
bLyxSzjIvICiwvJDykABH1m8rT2JNetkIGK9zyvEU0Tnxj9+0usCKVL8Fmlx/7ABrNLsHFlb2MNJ
J749ai+dhJ3q30e1J4UZ+G2lJDCa5xmoRNoTUqH2efTF+zlPdtuBnZ6QW2yZoVCzMHc2C1dmseUO
MEzIlQhf0I3HEzrW5HGjbSHuRgXKqoGKo05YhvWnvwylaGet0mnRkt1fSYaHt3L8Af/xN1yiz6U9
Ww/nYC6lPFhUMhkT/OjNPXd43GDU6NODeKpbxDRGdqFGmF3T4MGMZ5quKuorh3YxTcGRcJP37wsd
ZF5aZY4qVpy1hL/xusIxwRH+OQIrpEagq8RAJp+yrzg4Hij+gjaVhvMwvCM6LAv3iSFmWIrPI2/q
xLst1onqgTt6KOAskXPEMBzO/DD79EYj15NtSKkK97ABJuixyJkRcMxhPv7QWAxYK89NI3Cgq/tS
a5L1MyO7i4ZFiso5O6OaaxaMU7+GwaVQHX8pMbe84IbZstQKc8BKDJP4sur0/lUIvAaKgK/wccId
U5fAxuXOA543h0XbrrmdZCGTra68d+oYPooPYCOkYha+s6urd37QVEkE+XR8VtcOW6c7jZ1hUL/H
jIOGglpXtF0s6VPk4UpCuBhX+33I5NM9DYDtRarsTNH8OrmmBRxzoTfjJoY17WSHrU1bVVdJK2lh
v+saVh+1DAdeijp1GcYWuDLG/g2RD5WyPUp1O6bL0+gY7dGj92aZY6wAx2NOEkoaW9Ic8OrRfivt
E0N7sfwEKBIMHY8FUMAl/LXp17/OCgB0byR2tsBDFbw46717V0yZrc3JeR3z7BzftfD6nByYhxWU
4dedXYbWJA9iBm7DGnNTeZVZu8vQnatdFAsgSWwz1kx8P2qIcetPVe7tZV1FbWPZFoTh6nkyJLYe
5E1r8Z2LKf5DbaDzfvbZNkZEkehTUC8vvoKF5PTgk/kuqOzK8feLI6RFUarfsJ0A9PAl19xNwsjk
/qN+tbDtn4rwREQihD1yUmoTXO9gMJDvNFHB+906MpbxHYCDOXYtnL7Kk9eSLJsMEPZRhwaYpIQU
8aDW+x3gwFW/jV4Ls8l4ViUq7HnS8QgjrF51iLrcjnsrrBk0q1AUqeeatWsPiGS1ugGbSNnuBjkZ
O09RBEof+pF2g0QJr30ob7kW5gtOHA8Eqx1kkPyJxNzPefw5zbJkUTKjwqxRFyp5v2/j4AcCxIOm
a8xUo3O3BIs+SoULK4Mq7W5205Ej22LLaTkF/5uazOdBU/cuhJDyHFNsUf7D2NSKw/07LF2PxP4X
1QjMSA+ehcgzD66EodTixTu26GlehjnUsXnO4a6q6Enxwc1EFKFNjEsQZbBT6sPzCbhXw+Pw/oUe
e7ny3+fDmjGHPGvi+uHS9/0XACbV7RFw7S8UPI8WdVx7nTIEt6MgghlXabUzqil2SSRQJyH6ZJ61
/hrEAaWMBmnVnoWulmn3ZfFHzIWiZ5iKIbcV4pK82WilEVjjr60QmGXQne3YAvtxkp2LUlJzFa9q
MvbfH39VGNeexykG1eoveOiEIOWRb44/mM4KaFGAVbAEUTwFD5VBXqjERfMWAyDJXyMwCBOR9ZJp
m7RMPWwhzALQY0J8Aw0a2GYfpUDl16Pq7lQFwbltysQDg+4ZHl3lgQfnEC5b3aHuZ+vYN/kBcL2A
EIlN3/kncT+r1J9S1B8Y7mD4hdusBcq7mteR9o/s1S8k//Fc5xBh4Qcy8dMgNDa588jOPGceUY3W
Bo5JgkFRTDczljWHmbze+AuaSOM74bTBTdazzqGbkcNwxwTp26MrKvqMwVCKKqUbjW6do4wDAnK4
dSEgCguUl3XezfHoYrwxS6FARiwVNckrpCvUKOHAPMZdLv9xZaq/kTTMUD76yl4iDDrC5zDYxjxc
yapaXNggKzqxrxwG9yT775cGKkX+CSvg1cD00J0UYb6ca/0mshXxOHYPuPtBeec2twq6GhimweRA
hCamrt33vUQixjU9ZSjobzeELsIqiGCJVCjOSUJgcHeywKXbDzlWbzctpOzPvsKFoxzQl+NuoLJt
woZUHJtMDuKlWvjrZ3znhxAePtoAP+/4GT5KphGKm45J07UTHy+5v/myEyrbNgtD7+NG+lLjjwRW
xu/sAcw8yCE2nl+BXfB1IQtOKHosc+ONU5qXRjvlZrv8mblEzOrlQyigx4pde1HDZW5GOR3VCalI
Quearupo8QbxM+Pv76by0DQc6PQwHE8/G72a9LODSxWSc7KD+w4SEm52ihYTilZ9rEZlOf4Mc2N6
eD+d7Xdwg8YEA26gJyDwZ3lBCrT+pOgZ10wSToCdzLZPzxu+5UtXIjYwRqDZxYYpu6iNyDBv6Ub3
FBslIeE2tc1k5jFxCNWDkQ+rNUJ5ts13RXxKwhfZCUSO7whV00Q4tUXud7iMBvtlcCBNdToB++m1
LbO3ArnDmGPKJZk311+b9A+yP3iX7NQ8q4Or3Y4+RztJCC1mia1mOd27z4kOx1aLZusA+it70uJq
Ur0/BPcy+vI2L7Jpt8dhDpxCw4j2W6SbuRNGnpgB7wEOTKPmLFN31sz1MQe6HWJ2PNe6t0Yrm7Wd
MiFZlO5WA11iacWURPO9XK7Fy/grb0UCViMvzHQbEU8J1/f2K35jkEIzN6DCdwGzlwFsA3z13nqm
b0HmV1d4LumF9+DqCJ0MyTAJRtnCW8XRt7UG3PF2YuM+3/05zN+86yN5yUTdl84wRA1NvH4M1QyO
NVxDSl91cGPeidVPV/yfur/V9wImyBd9XI69j0hG37LX1za4aFXuZ97dKw2pTG+vFFi/wGlmCnfS
TkkZTV924q6QpgnYAnDpP1ghyTExMa0rG2EMbHf2YgGfxZYEMr+O6RV94ED6Q+cxqdkd3xEXjli2
UiU2U7Te1fp7UpiqjuLGQbfRO/WdWWaflRC0DBhukB/HUjaLS5F/ziTO/EQxHzIL+WkzKWYVXgfu
Jzhf5rmn3O2JIdqP2u+jMYOhvBaO5j8l/HejgniR4S9tt5L8rySatVYfKQeSYHk0rCbCHhowj+2l
68UBRDyCzsIZXHtJaQiu3HBNbBjl9J6VEpvr0BWCFqevFpA7sdJGJkHnmDEi3Htd+2FJawMsh/75
KAlGgrtDYORRlnaJBmwiZ4p/nzmeXLkW2JjIBtutVUiGD2TpcgazHmTRlPSpDJrgHFvUjH9Kxk3Z
uHL6c+k8FFKiYC13reED4KX458Mt0EEeHz9G9atTsdmv2Dh6beLofnJxkwVSsuM8J29UYVui6T9d
wIF3eN2MoUgvMPVK4ZKUc1MlB9LWrwwXxLU5mGkwxh5mCOwKj3Lz/7QBe0H1gXboPF0Q98/7P087
QfAXtJWi4f2JNEfMS2G6qfEJB6Lp5+eqC0gBjt0NMvn8kQmqU3KSIpDN3eAlkW/EdEr8D8xoBNv+
knrQK5sr5jzpfo7TGQaB8wpkb0kPwEfOTrIwSjNl2ZzvdumaZknQBuT9Bk+ZHf+MhJ/XNVKDRIoN
mqRVrN+3baVsqjczCSuCwYaDdlsN+RauRNR106WrC3nBBG4vFhHxQ+/+6MDYwfzArPdu5oQsDusG
YUiB67BxS4Yqg0Rxem7Nl4BuIAZA/R3vwUQqnqDu7Z7a6iLemUAweKOECfU4jfLwr4MvCcYwMeOy
taQKZICvv8kbsb0MKcRmNezPJK7UchkmEewRj1Qh8F1VXXwqyB3Rmm3NB5uBvIJoNJRF/4lA3U2O
pM8UGdZLmrMOI4eU/dzdOr+BK+KkUYGm4b78NT7nclApizVRpKRK0TPXs3qKxGyAsUoTUgFA0vvZ
AdYu/U0vXdqoCpfgDGJektWmmgOn6xEnXxf2HEgPQOnUrPiUc/ZpKBKdWnj9w+Km6BjmtnXVbFMe
Apg5484CT2NHhDMF+NaaXzA+YmvMZ5qb8/vhHJFfjYjuN1d5ibVF2fnum01lAwSk6QtQ0tGc4gke
W67FwfL76hXcptQhz+HIukMgchzs4GUJPKZo42tZ1TDJJd9SbDyUg/J0j3RS4ymOp5GLVMPt4LSL
14n8vATSJe5HYiuycTCClaETlBd6B40BuMwFjunswbCXtT0+v8nqWVdFnWZQS1kp+2KaqfwrG0KD
0bwEX5VaC43gqR4dlDuHZ8plRerHeEo2NFrDv7wXKhrbWxYFelL6xSu9WLLcY4+BeEm7bs/DA2Rw
wBhu1cn4KUab1yBEyEe5yP9tdxwH6FElPvBuifE7UQT0GeXUkS8480kL8TjN8FQZFhvA+7orybDz
DYNyNTw0gn6HMyxCw+tUnFXMq6CMMTSgBn+hPh5Y66fn9xW2faemHAHNZIIfwPEEEhJF49+rkiqD
o0d2k93dcwb47VF7ynrBWWLI+uBJ4HaMsLfT9jIlzCrTeA3mGMCWjKNkzlwa3aOO3UYYJmExM9A4
gHS58BrOV6/x6nfRjqYEkh9N5wJ6KFmEjwhHeXyFeNtIFpYx6wg7OF9i/lRiT8XPkpYnSca2i80X
a5qgZ7qzTbZZKgBaGRMWQitLiBEvF40cVtrxauFWVUpjb6M1IEqUlu8bpxdDdqlNW80t9XhaNGkj
7uIVYIxeNADyf44GkPbTOm+0Qmh6Hhwjm/+l6PlkSTVQ/i96snIfgpe00aZonwbZltBxIWgPjsOO
GMzgaG0HZCEmuQi9/YCW7I6jr8uvidRzPqO2uUwQpPZjJh151sts70m00Zj8DASCpLdreQIgPC3t
n0rcvOX76MxVn0wsudWrYVqe0BmiGufyEEuCp41aQInfDDBtLnG9t5LUz8TtzMA2svTNIDed2lvT
5Ayq9ctCGUOEjNnDdKBATwj5W5JAP+u9XBKmGSe/lqUiIHIZ588eWpHNm179UjwHv77QSikc6F7B
LmTFVhsTjPI5YpgsqE/ce5+FOUg5e/8w4NWtZEvv38Y6CkyXH4Xox6+ubJgZfURlTTrDt0q/qgHj
BhGLThmfaKieiOj7fdTbwf36JmvU+7RDmjxQP9ez+lRFOJwJ4dtLdHyfaVN9HyifiApSst9QxYch
vPOckdRVcF0HsY8fpaXvZR9wY8K4e8LBW565pjvBeFPVQliF8Mc1own/XTtSEDzmOt0lztEAQHkF
y1nD8p+dcpRrEWr/XnaUggmv68rqLGDonphRgkOf6oAuc1CMXleWphSs6fmFMtUY5jctO8McspAQ
azsknB4o3e3mqRVpzq9irfIwjTnXFmJNr8IM/RgQ8yhAsYDyE37H8JmyyGMC9evnCAeH+Bx161YB
qLZu2PD7AzwkmdrW02ZjI9HRwl4Fk8w/BWAVVmOO7Ye468uIxKXTRuNFv2bLiAS1JhCi49/K3HbJ
F+QCvTm8ZcSXlmsjqJxggkVRABetBaOIZD+/B09TKnYBsoUfoVIJjIiJUf+D7ZhkF06K0zFkUfYs
nb5xdW5GLk43fSHIRxWTMUAPoOrQrr4m3+hS+8YnIY+vKW608SWbJaXyvOfVRdmo+T0XVwhHwOrr
7S1JzoUNRTmMGFM5zGfQsj6pKsk2nOgdgQ7Jdpf28Zso81mKA9Wan2yDVrEgRshd7/9ydOwBw6g+
nVEiUxVuDRw1Joj6FCGmXc1k2EPvSxvt4ITXt/eqU69l4yM1fsYz54uWTO0UckDZjhxg42r85OIP
81ELMarRY70xT6T85HnmRTzuEaUrBwltPA0o7I/u+3u5mMK/WJ6PgrAUonyIpLCi/nBCqi++3/uR
tGOdq5wI2+mXpRUJd6VeSG8IW/X/8Rey6s5QAU+q272Xi6xus9KgKt1qp8K6xMenuXbJNs96CngG
iHV+FNd+OtJ43CCQzvIGaK/L/qVzV+77RaZ/kaw6UKdhVLvV4PbBwn4TcmxjWDJVimpsJIM04yOr
DQVfOAaTADSnCd87vgr8zbn2Yr3SSB+hgzLpfX2ZYkv2u1FVx4G1E5DgEJYOk/qhNEjgf+8J/OJT
IHl9LmeLDi1X8niWqzTgzf6P5Ff9L3OTdUNTS5FmoHD80irJp1fMouy3bhbM1OMFrXhYcC9aKQuX
uPfb7vusSiPyVXS5u4LWg4Gg0ZN6WKeHBl0Zg7iWtn5l3KGcR/OMtxvnJ0L2f/mIIZM4sX7kxvp7
vngK29BFSHXnT6D5jRhXUlqF1ZHu7mtt9blz4ucM2QdsqYquzOEC4THQT4jYirkeAhPLJ/yDZ1rM
hb37B082hdC/WZkY6KX9qOR2dD0O5LPozVSb7G63p6rmdAPp8C0C8VYfAUX4VaAeVjoqaqL/Gjbm
rpP2fO/MeeHfxWDJo+56Htfz25qQPBGtK2gfPZZj2UgH+oRLH1Tg5ZcWwGZcEOrGk9uIrXMK6ufg
BOn0wq/idSTws8BZ+sBR5WU2CY5OAPJX2bhiT7sgMlMwX9O/t1iRm+TN05HhN/p5Ei0HXD4h6gwS
QtUm8UUYdvLSJSL3jkJw/vqKF9SyITru0Hquz5BiC9HXLHIBkIA/VFDNyKJ72DbAECKvoBWyneIB
qc96CygNBPEY9vP3mXbve+wNMzJO74eYjcmEBPDXg9MS63Oj3yas8tHFVJXOMGjp1rKIChUMqycI
aN908EoofKIOYDLZbdNyXYOTzUYloSuIR+JqlyVBkjl14lzCCXF1jtcFtMci+79tJjGqFzt3iAbO
7bfBOq3K/8Rw4Dy5oh5109JozkZarXvdVIpceCGU2bLRY+ncMFmatOlBiohg4CIScFzyIUQH/iAx
I7k7TbtX/TH/TSEozB/mryQwrd5FArq/0NisvEM94jKQMcxODgSnVckMaSJl7QDATY4xhcOHL99t
U7iVzomUJLukk1v6Z9xqBaC3XV2+7/oeVCq1uUVCC8YJp/brD4XgZOPllvfYFZeHzHZht77muWUJ
4T23FQRp+lbgQl5rxkCE77lXRmiMcCrk7r9oPWCEMWutdEic75noPZSTPdGszm2/FMX+0VfyxdC3
gn2i+0XihLZfouFz9UQkvCV2v+Fuoz8J4Ri0yhYGmdDuNT00R2+82eywi1YTlM/WOIFdoHn1zgGo
shWckF9kvT2POc8p4JgYmQ79BWm4aDj7L1NpkF+G+nYnwPQv++eb1XVkKyKSq1osEXNaPRNYo0eL
BdAlXMqlkjEKtakM7DD+v3Dl4g4zVpeXeyob+p/m94gBAjRNwcF4J/KvYLU8HwOS1O5YzSWamsg3
0TsAo339K3kRGqPUEudgqcfMyevDEQatW97QPBRLTyN6/CSmj6mTHqmMO0FbVHcnUJgPRuk2ZJW6
kf6E6Tgn4AhSeSIstwOdS9H3X0ysWaj6brL8WSTSb1Api441oDnlUSFQtfUcLBt1+rE2K9ju1uKh
uW/0HSVSZ1r8pbsi6/1XfYJmuItzdhKyCnHey0o4tphjxI9K0XHC6SJaXmz1qLQ5ohvOd2gK4c2U
xHV7e5U4njHy1e1S52Vh83vaOufqIdlK8yc6fMlpYbfE74rm8JuQ0/BadLEE+Af8v5Z3QG2q9X60
3OcMxvb6Rqd8wZAwT4khpGWBiYv2kUUjgvpxja+X9UNYx+1UsJjTKLB7iAyEHVCyTDhrSajnKCTo
vsEHGeIWzdc7PoIjllNOFoPEUdYCfSqJ/pzT0CJBfiFLWPpm//IrAisoBt48lBRi69XOeQSvbtY5
5lcvA84HZPPboCpLgq1gdHqVUb+UejLwGvju2xqUJngRaLyJw75GW/RAD0dsnY0CA2nYDx9n58iH
VRY1D6talbw4M/Eq5evSpkON/Gm47PqDcL/EV8Sor0hzc0b6Srd4cQTHZYGIkOsk+JHulFtB6ZMh
d5PnmQZI3790wab7qXnjIgxnfRuSxSbfk8HRD8NfgquEfQJ97os+srfw7vZIUc9idjcbakcjOMmd
iXtcNTNpzBI6mhDrvotGeN6t5jI0Kf4Y+haEdysK6ctD4YMQE9pI7TYRYyqA6qly7uVMfEMcwfX1
SPgiDqTQ/5rdM4GDuJJkEST5hmPcYg2jYeikwhLHR+murGZOW0cCNxz3NRGQ76s6T+tmHIQw0tdd
P/kNRGE6crWl3DmlKM0GtwCKq9Xejnezaa1Dqf3AyLCIr58JmBpx5hjMPWrw6vvreta2eVRGQgYP
1R/KbjHDBHPrlHBim0rimXAAXFQOoWN84Hv/EyQh6IcAQcHtMbrcQvcHd2KrP6w4tkC5o7J5n3+F
F1UChKrGIrSgQqUZ7g/RY1gzrkyv5HIRCpTlHBlAeE3TvryxMqlZMOK19CLvLs9d3Cu4kOBPhVv+
A1ri4tUP9ARpSMOzMqb/SNtXnNPiKnvDPKMRi5VLmJaG5SExY7pUL7zPX8yucRdAznnjQg1sENdD
RrmdHaLY7hjJh6aDA1b6zyLgYTQE0anOA4arfaGmj4R/N1Rxj8Ymsydoc2+/7cK/6VNmwDDGR3Rt
5kB2DAX2WLf6ddqU0IFsnqoaszYXBO1FzbNrF+TEVYXYlVdb5x6zTKcnucnY3Upd8Iz+c4KDN6Y/
cZIIqFDvi91+g4t/w9o860HaJ0+Yv/x9O5yctZABHPSbuwdXrryo3mmneoX6ZoXpRP9bX04dmo/z
MzOf2SF2Kv5mnntC4QmjvUfmkLnkRpOr8kFp1bomJErGjANti88LmIAWFRS1kPuAI9Zzn5ykRoCz
8ReIIYh2TC1PfRWOPlm5vgjWV48qdUer8YhzcHaIsvbBvojdHVlENWFGENV2CHFXFS6MlkZaItgx
1SlUT+hqvgX0TZCAVcmpb7nnSjz3k7shQBpqhpvln2cmFedjYMPN+z1uXsJi+mzfyH/6oxIFnTd4
doSXPLHvaqBW7Yor4KlBq0YJW+6BeRJj8sZs05U6lyiO/0biRQTphlk0bZKlqMYL68SP+8NvFGcV
6fSiw3Yg3AXwfsASDrSmrAh9Vjib6uzLip7TFxyw6DxAMOZ5dfuGWnb6NE6M1KfbRd0G01XfuI2M
iSGG2Lb+0vYIkDVuuBg3ateNAozRReBNQcZLbvptBEWiZG+KKY3aypGjETe7PSi1BEl1akW5PRos
3KyDz8rXCUN6/ujF5rdR5NcNMedwrLjxBn4rw3+iV0b7hFwwZ4NhL0vgADCEV87bCS+cmMMuX8Qk
aaZnWIonnvVkQ+SGtv9tFlWKvshWV4WxnGZNxLC0YNBiAUUHL6vVcNmGt7l3nzKHoML8H60uOhEe
cuzENzjP+ShoF00DMx9cj7v8mqKfCUaoePidLiFrFDr18BW/p2MnRPCiBvSyvHbSEE7KCXlggMQb
PoWjX3hEoE6/bD3V9ijuIHgTKodsrZz5vBHfNd+L0BMrpVqQwX8aDCuu5cvTkMWlq25B4vuUgzFX
vDVaZh7ABGbiR7C6ZNSpxCXJzWFC8pYNCqPcI4jNGc4NAb1aZSlJhgOtN/yGRtaHEviYVNuSwEHc
XRM1fa4m0KudCI26WYiM+wrk5FHKp7p61tTqytHvs8zyFlXud1v3dq0wZssYlFYhyTJ/RmOJFWou
+VKS34uXkhRs3HZ4KEQDEoQQ6LDq/8V7SW54eMk0xjzl9KJTPFt4R/9xdsAalImoiVNAsZ0/yc9B
ktsEGua/N7w8PakMG58un2WDagZwL4hXA8GvW2LBl3lCphFjiONMPUTNrmq/nxGoLwUmMZGVxkXV
1x15tv8DcDoimUllUNLn32zUjNCQk/nX2zcmo7BJ3iLSqy0HWwrwB2ZpJlyGFqsZk/SloZyaIPHc
Hd/uT2ir5gNcFBAzyQIc7e3LK8WkHrGzv1Od8LV2lVab5ocGTYPHadg336Vhg33nuJAdNO4KwU5G
ImNW439MBys5BdFYSgzTZ5nrKtPTpAsCvlygXZWPqnCR0apUX0NjiBF8ada9gca26+yKH5O928+H
SUE+1tJu6CMidsjZJPub/4BEIP4WotbOecQA7Cyqs5v2Zp78/SdtJnhegRcjlukZQMf23fncshKP
DF8DIkMLHhZCweO9nSdtQpgi2qKfU1iapPmOVb3hGT7aTf3ozojz2//UxvOjuaoVjOJkuMRXQws7
vfIKsSbks9C0GjgWOxl/jx/s6H234F5gHAq8/c84OZePIF1MUw8P7rR7HUG0q++m1UX9gUC+a+X2
TpL3VQZsVPe18Oa+Jm9IleYGWnXTOVQt2/ix/KcEK4I3PD/XEf2GoYGMXfNShiXeWBM5eIcJ8w4/
2GxyV5I3lOZx37CfghBX0s2boFBxBO5TKhcaO1G+hyxko4W2TuUQYg4772XvEJIl5nLCMZ3xL/uG
ZE4Vudft+HPKAf8l3JQuNPAeEelLjkxsUH3TshJ0mf2F1N2BkD6QTMOjZ1FRA45fPaT+9ChUkSwe
B0vbA4KX/CuPW9K/Gq2pvZXvVp9JG6eSDj0lri/AOM0RTH11j3NlP0RcoiQXVsIOuDQdN0YEIElH
8jMXWKXMz0A+UYcf7fslbIiyXSsbC4XPc8761pJ1XcH3VtLPb3lXaSWTlXgKx58ZLfoaupxRvsKJ
8qq4Wz7177BQ1C00F242RwWqb8V3gcbX9JG1O5WuqG8kCDPu/fQ/iTW1VOxf4q7WfS88H2FuwaVP
tbIYwaauWlo6+HFZuMS3JvJOu3/peOqjxCAO2/abKF3O68QTXbbbTzXHhv9R7xYf0dJsZGMb7UWL
0MQ5xexZ40nHetSHXmXLqQu46J2a7mOJEJAhN08hcJo+iPOPfP5rmWmgW3djejkDbaNLLftr5LNG
TyrIgWWfk7ceS4cymUXg0oXmKNau3p/F4iI8FHt7kqFeWZiF26Dj56NyYwcxDPHUay0Ei8XXgTmH
jbbDG7+lZ0EpAOhe+m5R93nwZsudMUbJJhlfJbunSQi6aB8+61HXyLpsrJ4itOfLMM6cuwLy765l
06h4x+SYsVnrzLn+8WkSxqLtEuiWr8h8A1VafoAinZnb6cD/MMIb2j/jLX3PsERi6V9t9qxzVr+w
wz0Kjqc6itGsvcyW6eCm5ohy7lMNWV7/N6xBQi62WAZJ0sUADmrVqnKnxlqCs8CH9ApJ+UQ+wIMo
ayXcX1e/VbmEnQe1Qyzb7lPxj5ow8e08I2mKrRUEBwOJh1+/lM3EvyRMbdEZI8Wby+53Zrh3ExzE
kgqpXK39EULQypNSp49WUZ5F1oZ4BH4xb6O2Kyy8f2rzcIjht5l5ZmLQAeGGT75JUV7XCjCwgK5N
tVuMjQEIKwBBrQ/UpRigaZBCtFHifKBGtEejthje/I1yI+9aRPgKJMVzUC40RR0Xm+9DBAQyeWhM
R0Gk9X4J1Xd7tnhvPwWjytN7rEXpAqjf1nXPHKJWmzn+sL5uhx3gJ6EgDXbZb+fIOlrg+MkfWhW5
71fcfZvBgOIw97EDAnnAUCUQQvJ2tE3C4y5GeFwGgK9Ndu1J/pe/upye8dkZYnb+O1XQugXXKEae
Em2FaRotNVrhORwDgWVwMqYh7vMw5qsOmD4kjWTIuo8zPNXXD/+lTS4H4rgbjAOl723Ip2uXa8xG
e/D9eSLtiEnkADHMn2LgWdRolrHrF6CFOWggwEQdQpy0KV436aXD+Qsdv8cC0dvNnE4tAfRatDQa
LX4aR++CotZTrVqyE9XeG7pBYmDosIqrmaGbQmIxhI7kiZHxscV84KOiApHq5kB6Op/fnWuVjorb
pMOkh0OT6dM5mlIqCNxYWSTSgacltWR48ptIB81Cu4oLIF7PAFRc8gvAPeDvJFZMJ2nB25hLbZbb
hwQ9s/T5L97ibhJfN1AGxhltYWKmjS8iq7AJtJz6SFGY9w1WYSbdKV6aIcZ0pncaGR5ocuX8OAy8
HJSd3ov4qrlZypP8AXL2Z/XAJ83ElWOulz8tnX5e5xVErcJPmKTW/6SciJ/CdSw0pXBM2RHv4ITd
YsX43CJ+lSpGySnwWAxySmQ9U6miXEXr3wTOanVyyGC4Q/G/02Jx1E11mwGmg3Fxa8D96fJxG2BA
nHRetYcdeTF/F+m4SLGGO5IF4I/mvdUu2T0wdTOn5zWdKyPL/XUGUhElZzNVNDLWvuwjjxJ++6Jc
ma0ULnDikoqknJESVVIrY1F6O+NO1awJvZ2XiBWkQBq4WU4EoYjzMieWY5Grf589X0QDWwWuAIeQ
aDWcULLIu7Fxa0GmCXQQPEgjLe1dUeAuP2hfNPpwfBJZlbN6WCWpdvo9ElwambUsAZkRTVEwR5ix
a40o8CiMQsLD03FFP8WvoVkYuz1fgG5zFMXkllkkYRsRUENCkDhoyze7nt4DVTDBnw8gifbGxqjb
JsVgHoTGbqt8MoQ4psjNfZEL4KaPx1GLKh+lgojY+NuUpdmpJd7VzXTMwP3eRjzZspIWZ3mHdR6r
iaQRwYiImkHCKEbm7iHGn2e4BDfxEFc6cBCAKSVox0g9/Vb7YQUhg1JaCTz/2fydE6GHTuwj77QE
8HuwK3osCqEfUv9yCJOlCyLBqqjwGLO5o8ULOR9BJ9INak9j0JwOOU+xv4E/pXVpycAOFaN9lr8q
CGgwiG0yBxca0QU/Z/DAXd8bpwA5guzeuUhaBI9qccVciX/WSihf56LxNH6Qq4E8K10S8liy65rK
DpX56E3N4VhQ7VqIo8ymsWF8rSEiVWyRoAFjl9bU4hotkMMjSFZo/y5KaBnvQ5tDh5Qm33+EeXVA
qBDdjpcoC8b8EdvdnEerRqX/itQYdaHid4ZsyJoVAwrebK6zzh7nKy7hbx6Uwq8I35Ptnj9moUwL
/gND4mJQ4WNxld3fdVC2f8w53lY1bWwyMd5ring57A3TNRlQPXSMIWaMYVzLyIufFR/Ki7/oAfQ+
ACOeQSCpPfuj3OCwyemR9WrtruFYh2qJaBMRbmHKcZ9sfQG9ZlrrKCJENWtaOhN1Dm/SuHNQ8fNk
6ifpEYupvXbPaL0gUy2f8QbRoi83REutuXdXC3ZYC9cf5zttLvTF8gKQiBDFuheeoZoI5iMOZenF
OHmBN2i0QpziLCqLx797ajD+NbXYfvNDHgLpBQ9myLR+Ibox1DQ6WqLFDlNyFG9xd0KExJQZZWsP
lBkqytoeLJe8yhqFUypjhJOAn34CIpKHEwotr5lV9NGtUlarkEL2t/+QKLYQGXkUHMWAZX1Orbqq
feAVGzEDbjZKtl7PyCHatOoaJtrLmcmYeEx3Sy2uppLsZbv1t2xQ4ezL+8Zl74E1SvmHPo7sovqV
slhAnwVtj04bId/qv0bq58mP6UV3R6Ptz0ihD+dnwGHPQ7nMptlrPbRkgw3rAXdhqSStYEy9Gljw
TlptUnF/r8WzWvqtUOxtIAvPdXeg4+eqPIGbGm8rc7afG5T68oPMNNvqppOlRykncrUdDMowQ+j4
y4p0w6IjuXxjOtFNOaC7aAoRF6FEY/Zia4/kt4BThQsi1GwMD+luPP1ssmwkXP6CFuckLNKxzAoy
vnQ7HEMVNtBxQO6PtzqthZreLlFVcTuUcpYuP5uow577KGkF1M4XlTE6d/uFoQG3EUZCLe0ygZRn
BuvHlyzRDXvj76N2BFzIr3+MGvyfvInXIsd1pIBl0QLFlDzkIJCzyt8Y4bEeWadnmKkFAoQLzgyy
qL0h8rSURDsX0ZQ1tyZmEpP0wunKexsCqkPRZA0TGUecYywCQD1nlPU+YwHtyuI9PF/amGZZ2uKr
tRxXQZ6b7q+Scwbrqzj5fErvh+bW9ckQk+8+kta3So5GuHmXWJ47K0X2b0XaXw7xo6mtfPoGYw+s
3VEwJmkEb3IjKTV9+WSlQ0q8gRzZLLiYNJSVuRb4SJsgUc5Cg4WAr6+O40a/zcNJih8Eg9/0HCG1
mTTfq61WZqWsN+N3f3xIiIatUsN0RgYiqEzcWthYmzLt7z1mZOjQ2vQUGfqY9pXocLKJWDFjtISG
fVqsYE8FAqObC8zS2EmQdwZTzKEcGlVWOZjMxjnRsFU5VXWq5bkAqUAVUYf3ma+qGJ5tV6Zn9zQO
m3ECKLaB9Bs//00uPo8hUJt2f46rWdlRj4OViRN8FGwVmoHGI5tvYPGYeuLNVV7ZJkB7ImHzH0c4
6q6JncofFRLbXDs7zTjYeJ3OCpQf/7FDQwK7ObBiYENR3A45txSizlfdsGeeOEsKYxsPaJelnjvr
uR9k/kl0O1kJ9ZuEJneWAwGjuliEIb14/x9fj4o+gumEo9RYo52tQYUIwhD+Y1oekRMEMTd6aV62
CMlB4h2JbTEswRYZa4AIS6n5thwJGjKcMeXsvaEKkVV4N++X2NlmdMz7cFjoqiOTj+dYTNJeaVny
11YMizJ/O3cHFAkvgL0K+f+V2vMqai+VUeyeh3m9o4wGViPtw4TLAdARPLfiwhnYy7P3W/nPLKUF
HwbzS6a2PvcYALrruGWaRwwE6VDh8hzNzUF469N3f9LQshX/H9O9gu2jbWLlPhISwNGdKADgqiCL
Rwu84CVZGxpM/4J+BCBJ2EVs3lf5UYvncyMSJ39iJNh6KTiurCrAUeYzGvqPbsjFUSb9sphugdll
Rap5150CbcDgK+Y7JREPcUNjoZbX62C70HRj/TluJzieDCeZmS2XKzzJ/jgpK9AmUsfsSkVz31Oo
fKU/aYNJDshBvCm+89uZe45Zi+riA6NE5rSzTIAZnFVKHbfmmANJNT0xOxLsIuLvjnaOsbThypwE
7mflMrFNg+ynYzJ+0S07wgEw5MQEuLuW0Xq0uckSKiDyTTy7/vSEST20CRyIbtXNRoruPqMCj5WN
6HietdehXNsQ0xfmJ9MoqQv1e2z6nVfgvBSa6jH1tVW+jF9NaF7j6JssNK5y7mEa0pjROyBIua1K
SpHI1wfWqblsB/pQhzLCtr5OkjA/ARX3tx8lTasliGjxfxbKBkyLaxNUOGuFPIxhI7niTu2Gprhu
XhAp66pIoW6YwCgXm3noBhsqBD+/7fqTqkLQNvKCwl5pOGokivVKUPOT15mQA+cUla3jVQsZ2GQw
sZhndORlgGMAVOZVtpvGsbj1Zt53AFwlheEr2MuFLKhh0h8OYfuoQKfFVpM6jBhReJCHMEA1mypW
/NfIyTt2sC4G3vkVHF2oEkZUi9NQpTVaramGrxnns+frspeMZP+xUZC5a9wZgkQx0jjdXy6ye/um
uOoeB4KqGJ431VMBxYcbImALCS2fGIsbSdswjSsp8ySSzpRoWVg7L+dkH5JhqedloCS6nrzDWb7q
GFYSsw30k+1RQqObKHIFIz84H3Y2e/FGemqxiWOnnym8gIg2UHs2d55GQJrxABkml2UlT8ZmD8sC
wpEKR5w+IcxLsSYdm9zGIluJUy5FoMn+lePZiYgnU2QTyCdk7tizVcYHODBh76smPRw4TzZzOyOs
kRgPWlmQN33Q9FlhUqLjvv17uuQrPyXbSMk7e50iCnK3EGHFQ7VfUwfOp3LIOyCXgYceEApu4e3a
To2x8/FG3E3xSiGsYMuYt1nstRNzuBhxHjzM5nd3vpEzlRt14OQMGOBtzTY4BVbLlgTH7c9E1mnF
nrQOuRLZvh4VF5bmK4yBpO9Ep0cTqrZ+VH+peCT3dkU2Py0XstYT6Xvh53fTDgdkLhDK01o0C+iU
N61UWMT5IudltO2lUxeqHL8+kSIPp0B5weqN54p0wpLxMtyV/huhdNK63veQafnhZMcHt3jKwAcG
R8pwy4Yvv6GHrOoMKBy5/37OaT0PaeFCU47+vEw5YS+Htpvh1DztY1UH+l5cDSfD1Hj9XwOrbyEQ
6s+8khO1hOULPuZSraaLLK5M9AC8hTkZzQJ78YhZZedB4i1V8LA3lp5zr5Jy28jpcusjXd3IbRvy
XHHMXiAwevCXDGd+4OrhYKKuXdY8ytAT4HB4CuTBx/C3hSARG68nYrryhnLgEBwjYvNWy/GRTIL+
/kfNSB3P8OE+3g++SpnzbzQtdkxZe1T2YYqGUPhN3Bl1/F+cefCM42hl0nMT0hZK6tCWkSECtN/4
XmrNuyBL2Wtspcb/W355Oao63RnhwOAEM8HdDjQrj/ii5vcI6GdOr67wT8OUqPJAhWVWZQ9zt8K4
11FP2AZkSnByADJagTbu8UvF/pcpy1RmN7mjFWzOO1KFkYaMrpJKq9OvV3M/KWkmBH1/X5h3Xtxe
4rZm0tm31u+vlK2Jtmfa365kpU/6AlY+dM1GHYUCdI2oSND6VkzDNJRKjDFkF0IKVCaNbG97lcEA
f2DE778abzTJGbXwflH0pjhTazj4HpW+sH+ZcReoy+cnLq5oCKJ/RtmnRQ7PVovcLNpGSvQlBYvF
jGx9gm0aco/8BcQehzf/izo0faHozCt0yLTY/uVjImZ/z+2yZ/weHzzKqvb1KT8OYqOx8piD8Uw+
lW+9S210jTSSVg2AzgH/CFx/JpUHKNipMcxpAFAOYGGHCrZsg/V5WLsMHw+L8ceb06fXkak8n4iK
NC0pUObXyozk5q0LTyB4Br0+EAP7OdD986D3y0rPbVWQXPoycMiz7g51zXNqqirkzLowKvzZ26nJ
0pITcVm//8/EmrcJGyAFOzZs2qnI/S81avP2KFdrmvFAPJhud0LLYlAqdd5NIsFk1emjbiivNksk
wz/PMLAtWImXR6s3X/0a3rm0DhYIfR6iHl4ONoRaOXmSJ1gSofjbIjdmO1vGsT191op9IBGksPwM
xd+WoFH1IK1Bl+MmjRRe09UGoyU+bGJbj8w/gwoLPMC9VxVd1DIKuhGtD2QZCY3vNhBvIA2tSZGW
6lSDcMQpuB8AZN8a2x8z+ZOs06IfiSSoOC39nmGK/3lh3dCbmA3Noclbbjyc6Y2BFdtXonGd88U0
nJ7JkDor2NeUvAybYY0JFKMSJdm8ZEapM9vlwqc+UoVSgVsPzcb9e1D12ISZe+yLbt4AT8ug+5zN
8S4IuX7CnfbS+ic2H/V+sdrJOFyuRFtJO2HGP5rEWZ7SYChY7XR2FDLdqJrY80XVAG2m2PA4Y4tm
FUZ3Dkih8AeHaX+oTZvVtjOW/hwWDKlR3/zb3gbNH8maIOFp3vVjdJ/J01DQm0FbznjlxPJ3UitH
m/yxU7vCs8h0R16E9r4toKtPOzzlx/QWlGK1+WyDRbC0+vRI1JJ30IoBi452pUrWEWPA3QtyZ5O6
Sm3z8V3USvspsoae3jz2SHl20KefMOCJeehu13pbPeKZqjzVuTBIdMYfr4XkWXE9fhNUQmgidV+A
tZsjs+l7Sm6jItnvOI6FCS8s9B/zb2vQ0sZiKYk3VIPbpJS+Zf1V1pn+HzGOqPm8VYoAGxDmucJ+
c3ckvr8huf4igiNKCZz0x3GGSjgSXr/U/9Vm3xYlfzkg2XdP4B3aazUzymtpr/ckg8PJDdrpI9r9
CJrxOMEytjRK6r/ZPMjVQG3q9/9iOMD1ylEdbqT3Y4eswEYrA/r+DZDZYZs9fhZAWC3Msies3/is
Gz9U0erY9ZXP3CCZfZwtEUjQRfDCSDwNM0eJ4qxSyV3S9UqyKPKXp5fM3wLLBgiKJzulpdVFjEkA
H6vJDVfwJ7sY+H5x63ETW8vI7x/DzbhGLh7BPJJP0U9MbZg367ZM1Bm2MrfGgU9E5cFjlVJ2lKUu
fGzc4upQ7OdvYhZRu6gAhxqDBG4IEwSiCa8zDIz8bapXBCPC27OqWdhJb5ps/HirxsDpc7yIvLpc
rS6VRZLuIexvc28ucdaiGVNDUZXiseUWLkflTjzpGY7UdmxEfFh1j08iH/izUHg9yPwMNgYInchs
59uJrRQcZwSx1yDjRfZ/OYmvrAX/yLiEJY4GOKm9UxhFjQ9pwFa5gXfFPNEUaBxkKxyHXCS2wOAH
O3vpxFNCofRCKtSDCbZ+tEJQkm+MCe0dOY1ZK1Vy8pw3LH6cayfdymV0a1+Kox+yls6aCmmWJbGV
Bv4cCnAgmzfuT05/t0V7pmDmZ5un0TwDa6URZ6yK5/eORANuSgOdGpqEOaGKhF+G1QIn5asSIykF
ZjZaf3aAsyYTFKo7RsXBYu1L8SUzUVTe/lSlJM4RtS030hDohRj3PxBQFvTciuJnB2LKw6fW1gOq
w0X5uu51qMiDvpMKnSMA3fQBTRM8vT+BSsWFjR3nZUdTHGLgwlvmpJ/qO+t0rrTStnX/weZHjwtG
6VN/FjMuZn9XYrJqb0UOrwEVGk9mgU7+ZZSk9mHEAl5p+Az9J510yJmAb1/CKA17D5AQR/O7vNCH
tSeLAzgCCkj8/ODEXjPf+zHzRLpdhlKRq5wJiXABktSyt/Q6bYK064jS1aTFoPiJwhza8BtOsfOB
bBLDW3pI+Pa3zHZ32lJyYLSjMBWFUMjmhY6c7L4S8ON29I/3LgWjEV1PD8LYEFuXbb5y/NI/IKJT
r+K9OxMJYwYOW1phBIO909jYm58v/5FUUHywLoKVizAQilD9pfcTT51QU1N2pefdoShTZUtNaNSt
VuugcHvAb78aIq4yg/PN++IhzMAUXwdK0KTAY/2j76sozO7yxB6CivOBP+dx2iEeSD4i2shCawot
+tMs/9eByb+FAoBtbpEHjKabb8Rs1GRocWqcEDk+D/gvZPGoNTdef3VGRtUzrJroi+qFUd5D/6Yk
Tv4ZacuHEYCDjClv8Wb+kDQIn/Lfm656tSQC1Na4lHfhmG2LvOeHoOCG93J02wWUi1WJXvwPNhwh
/MK8bCjRj5SX8AAi358HEDT76pT7abXfIOtNIhYkvRfIh2iR2sk1ERS0cS8fgTBI9RwfWa8hukPh
jwd57fnoUyjw+bXSY88YcZL2b+FmiBHz0zhTycr7jgOwFIOEo3bkkoSHLLxgtAgkIRdgb1ZBTvTI
JlSmvlGFJKzT3RO1SmyZBA+4X4wj/ndxSv4BOGJce3BvkyyDVeTYf9RM1989aki/VcZENfPfgkrw
DHalkHPuzMDcAW/jX00mpwUg7vHk1XTEL6Apoe6MnM3fDsJjmMYZzskUKLQzo9cZreU7y6Y1gg43
E6LtT+eYLsrVv3l6V0OTXSWZOZWq5MFLZszDLlqrbDBBeio5mgGnwUzIi266dfr4MZ3zas8ygBrI
ky0gQYHiRmmdDAVq5DcMEwUtVw+w2wHc5D1r+OYGnBTQJbUnSWuc32SIfNHlJLRiELdzc/PbgAyD
sM9p+d+SPIsFqRwi+I8gYbYDwu6/UkXbNzXMxTlb1KxWKEw2EZnYU+AYcARyKeszONIXTWJx8JRy
zJXrncA+aAdAKXL0T7PEAzDk7CQ+Cpjf0HK8fj63pocTwNt2OcGuoTvTymIG8BjZu+Wv+vmgaIDA
28nZk9RG7K3twtbxiGu6s82tBLjDIdQWzrK1N1s6CmU13X9Mw75LIPJfiAoHr64cYSedCz2t2Mcg
x9CYfGLyBWHgP50gNpUhxtHIQjQVg8qtRIy9w3/QhPlRW8/h/ibRxZHb+37epMjry5Ndt8kbV+rK
QNRtIkHSMfe1V+3NRW6iuPRCJieQtLPgZJnDlwHCGZJMoGE9PcCBhzcCXW8YQZVkRlpcAXZGyhc6
bbmHOYt1+aweTuUPwCpBl5bNsRFWxAkj4wEwKfWCvQe9kPPmkqzNPjagnsjRIJZ7bPfEN5CcikRt
6KcOk3F7Z9zTDFFkxlxpPhWWo2qwsblhWc40QWh1BtlX4ELBgabtS3TrpTgP1WA95wU3ojC1Acle
nKcPk/2P9Z6c4EXU6FD2GhkOKbwCCU+4MVKafc0oXBBPSadNBIoUwORJfdYHM5oA7YJK6gLv44xs
P4RnCq43VumQeA/pB46AChnYWMgwI6mHw6XGtbUpZ3OM6dJhuTk7Dz+dat0AUC5ytwBagO0bpjYZ
Mnt8OMwLKJTzobgg2sHNPEWlGovdOyyX0reYSRA+JTxUdLlMr+RHaeMEGeqWqgbFnhqWij1hv5yM
KxrHJxQcLg7H6GHWIFHoaDkg1BjA0BAvcHCthmapEFf/oMyVtkVHPBuf35A7rglZOJJqKYG7pqv4
N+f+DtdzfFwT9+aFc5TsBSvyPxSC0dJgD2YzPNe/GKSJhlJHrz6T38NdREC02ZIhHxnrvCTMYAmy
ebD414NyE6kExq0J8kK245Rd0+sHheRJZou3Xov20D/8ZC43RIibI6jsnQ7cPOod1rXsaISdQc98
KUMCW1ZuzN2Q45FSIGO39FgoVnWgSI4O4aA6OXBBEtjUUz4mvPTMyMeaTGZTNT1x6Gbncw/8xjrA
gbw5zDEDy9ROnvloWUuiX3cuTRCdfmpkLUud1lhRtAkQzhToiBuCCDMI8XIy6lWJ7o8/H6oj3bgf
DV37LR3wEo+ruO0pP5o/N2RoWXnCCv8IJQS32dO2MgAgvT/ZaL0s9d1EuCRfNFuJmFkWE1+jVZ3l
u/VPejzEv8WhNe14uGPOyeo/FfTrV+sYkdvmzM5uPrgT8BXeIDoOtrzMHxkRwzwDHdNfEDzyUb0B
/7qfEFiQkqXWyXnZ7K/yETENGwR+Izy6OZ+bPzfH8cDHFgMtisoAMr9JvAanT5OADmgzRBSzER69
BifGq/MFW/IKqd3PFQDBZrRG0GqffVtmGTjmhz4GoRlqS1Kij2jVMqduqlV2Su64t8ymiPMlHVZL
9cAzZnDVCkuKl3M8X7N43TCEMKpNcfh63cAmroWhG2HG0x40Wbhp10t9xEloVK+ZNQ4HcRndO+tW
ghIxHVjePzFR7Re/ABhVWtAaay8odwtlMEn4meK6XrEvzyW22MIrxMS7AaH2ur9VHpFVHMXBicvT
c8tdgyqoKja1h272rn7dk+lDI0CH2YAhhxfo0CVc0scJI4TTyu21mdWmr2tTqyxrd6Y0x7h0s0GR
qSuO8zuKA/BXzQ75HmtbL8+BtvqJ7f6/XkRnDEGtubNutXAKAKPnnIhh4NvG03UlRHYYndiUD8cR
8htWUCVfg4m6EHksU8rh/I1G+LrOlMHebKHZ7WKxcib2VkX3DBIOtgHteEx12+cGQblyKP0HZmES
iUoWpggqEzaZ7k8LfAuSvM2aNS78bRdNEigI6H5qGtacbZUw0GOH5AuZiUOQzp1qUAJ/RZ7rSkBJ
4cLYnjcNcgP/cqrJR+DtqiGTsVS7jJk6rkH+EFbpkvX7erVvQFo5q1AxO8Z380MjQQnfn5G9RDx8
v75SafKJXjhV+s8+AWILWRQb3sCoqmpF28trIrwz7r+/+yRjNR8kKQ7SlEknKqInSuAfCAwug3la
S1PyJq8LQliBwm92uuU8/Y1xQI/Rei80VKEKBVQHBfTjD93Irxrn8+FCf2yN2jo1DSV6qRKZ+rnC
veCC4Mus6HqQ25KThjLTQCSBQEYqK5CpM5cAlorNqZLPnip/jXbW4uh/LwVoJJzLQef9XVHii7mL
8vLeKthKx01YXyuisNoprn07NHl83GDe4MsKjPfFrg1EyBd3DI+7i4nhRPlS1Z3AVdKM3olQdQy0
iR0+8KLsdyL3WKbtvSZ6Zwy0nexVoBtZBkzmxLof4MwY36QyufFKMzsGB+wG5lr8Y+AIsHEfm1zQ
MRAdg2JYx1lHBRYeZ4QsO9vvg+wOfwvk9rCBO1ow0BuUb4oPgHbivWNNqa/hajc0Y7LNLbUvT/OU
19Sv527iua9eeZ8KsL+2LBEyvyg3OMwpcameEwSGzzOYwgk/rVWptRcFigXq+JIj12+Ee8QfosBg
SsTXu++pc0yPU3XjP57MSeZHAcOCGVROXzFcDok3PPFAfCS9K550b8yLFymatSdEAv3tIEYb/VLG
3fkPgvdJp37tiAEKYNyIvTDo2a3bn9iVu2DZyOXZSjbvX/AaTYVjowezGWz2cSbvepiaC/8gkmBl
iwPUZO040U6qKr0r/grVgvs6frnkVgao0kzZxXHPIQyrpHb/C0Y9dsDxvdN2ODW1Nr/B68dGMhfj
fsUfxObnLNEJNQ3QQMHr3UjJurkc07FebFhu42OJ9ssSQ7Yd5jUACaJ1gnHYeNTaL3u4OOpB4ZDS
L0uqRt6eoYdQD1nFLsQS4W9NQVrdSjZpNmLAq4BDIL1QKZwSZU6+IXjF195PzMXG7zwSyUPD9wUM
WfSWnTIkOkLCcVGiDWgMBV2MGBok77o21+j8x2fQ7o75jhNh0qNdx1VhGAxPQO0ru22Fj7caRj3A
XD4kYbXL6Ru56MXaEGspOah/1oZoSSW2iv5YUuw4buc81wn8X3B1CyWbagI5eRGPegIYNDv9aUp0
MbERMxW15w17p+HI4igbCD2d9mWoQkXH5uHBfjcbszDF4BZHIJx9HkyojNJtwiasg4oGE+IIWWHq
8AptGQ+qGlt3aNd9e44urEeP88NCzYzVyr4xAXyLJrkMd2lIjXQ7RtRqtnW4N6OXwnk90o4JIpqE
uSa5E23virRBIRRUt0OW0EXo5UgGLws5nnvFB1/b2BZ0dBuWKQKxUahYuhhN13tUPGQuusE6wP/H
+st8246CHmh0s1xXUUNMrDq+bRnjZ7FT08w3Ez8r+0wSddtX2qc1I00hOOskls9+P8O3y4C3rN8O
j11q+to0iqT+xU8AWis7+yEvciaZs0fAtUnbiUULL33M91aki2inO7dtfzihKQfxAkrouINMmeni
L0echb2NdellbDAl7D2kbq/gs4VRA3muTf8WCTFLu2bwKrzXazkFIMBeeCBj1vNTDKB9v5RidcqG
L7gn9XLAiD6qjd7IuwcQo+THb6ChKlWQQyg5jGLwvAZKIpEbABIqt1kYyIQtvRtbxMJwfDtk1zS4
8Wnoargao635Q/VJi0E73T5FCBjc1V0/dV++o62aTAspwMAjW5p/KtTBb8s3OQXG+tePKYXQjFpj
hJPvuv8D3kE28NtnPsQKu4muULVLQAvlDBbD0wzrB/sGLj9CJpqGZbRwBMxLWn6bI+XNvJyud4Xi
JNuqw0scbvt15mPy4QTBtmLS4eofPMsP47505p4nMqVXzr5uBNcWlfJEpuQbv1FlmJ7IGhwJ51aj
GgiV9MBsDiA85NK9fLenaJ6YbHxGfOWVhezHObry/itc5pWUaw5rl9pPwBAm8kuObpd6VoeZnVDP
vDX+z3O2uRotb4M/eWOGiWYzTgww1RsUh0HItS4zjSbt/syZiyOW/UqXkWh3XJJ2hBRjvZTjZRXQ
Ua+1o4VVX/+SOs9WKnAuMs5Tay30ySCyUiFbRL8m9ze2K+vjWt8O1nNLN+v/apYvkmi3eD3rBdd0
KBjFKRhjsWvE9GdvYEODDAycOhxDFGQ/9RbO5eKXyGEW9tIbpJBcJrjz9gKSWJvQx1NywcUXR6jj
VzJF9hJDHgtCg1p86akUBcbLfc3PTdf3BQSQv02vvOuSY5BsfK1kaS5qm7arpGMwp/85qMwo+D2G
kMSWDU3GxH5rXqIijozP8qNIq6NKKCz0jXgv3yz6qCVFFNiLhPz9af7ehP1KKt8J3e6KzHjj4baU
wCKnbKL4ygDB6qt5bRskB85sTmHU1ciWitVty9HZlpbbzAAO87DRbRg20OXamKIK0r2+JP/RhuUP
UOb4i82obfrhLP0kH8VGajSPk6ooLYTa1Wg1Np2cXDQ+oHEaYUi8iLVirpn0/WdE9Qc8wBlYaqL1
NVHdPYWFzr4J8NeLcxzYegWOO1C09JmCvNg2UXpTO9X+q955RJtkdPKW1RRrz+1lKgRxJTXMi0fc
r5bCMDypDNfrT3Cc9KKDp5zVRlGBJm9zLBoPwRr2YK2qdhEj57Iw8K0hg6stpSjWWmdlTB8GgHis
Oo03oK57ZdtuZs2KcPbaHL5gd/MxB5gviBtm4bU1mkuM6whk3hJRzFFcTY+/mxbagr3ZEEY+Vz3l
lj6/KNWJYVm2Wk7jUdg50WEPfCXI7hYw2XxXhFDB/TtWcIxy8Af6DBpGwTVTUT8zeFDtgDYs2dIp
AFqoB7j1p3UYr7ouFh4DHFeGCknIuSQ2ryp30dQ7KAQHRkikT0/8/VJW4CqsDuSX+V6HI6gzH53f
DwBDL8L9I2vxCLulGUq9G77xy8/u1PrddIA6bbK0A9kkRcorDr/wwCwmyxc4Re9u0G8xB9sD49P6
U5Cy0tp+I+4nW23hbu9uXHSuiKorForWJlTRjDlXC4qZnmTbF/eCxtX3ZCpHek/iurziPpVaIXYt
lVs8qk+hAyFRBaqsiKDWEz9nfK1OGUqTNX+5QcPCB0Iz2+h6L4F0P+6uVziZVpVaxltnvqATB7HR
Hk1WFUkHNJYKsKMmQwpcdlAxpVHhu7aadBXX5NxhpNqTYMnVrLKwfhscohjDDm1lXT6GRrV4/inX
dj+b+snirVQjin39U1qHaHvqLEfISmv3fudFNGh2B5yzfYz4eqGg8E6BKw0Y/Mr6Kff7q7wUs/Eo
KBiPpHSdqux7W967Gqs4lUxBSv3bKJmXlxSbOdo0sAqoR8l3I49ev6azU3vsfGvZiFON0YNjY0We
PL15Dh/PWlz0kTDReOthnqERYdf6XaliWq/JvGVJ3SL7bjEMFo1kx3nruB9n33nRSfagmK/1E5t9
eiZLDmsj9d6ah0B/e0X2rSyJDN2c80I6Q4CRULwQhynbrL4mn1Q+IT/55+TRPzwg81KFrrFg33kE
SFbQ0t8dnJIKlT2Cjv2Bhju5VC8wyOmRZVvdyVW/Y8mqPCw6eqAgA3U4Y5df3EcvdKw/ym/gko10
tgwfeIsO/t/hAsTqgL+VENpTUtApWG0drWxabcDoDyLNKmK8eh/lGh53DXD9EUjVSaQPDw2NdBlS
/T/P9y4JOQ6TvBfQgvX+Lb/DtWA3W3sjQUcuazokbHvrcjYlJorhRia7QGZUQFHSGxpJ2zkhj4y+
kFCkfmaqpv5d2305KztjH//aq6hI9Re4Qoj6RSce6okC5+zOxDGZDz5eaaHuCga/0KdAgXYZBEeM
Rmkln21dOC0in1dlFzwDPzgTrHJyXe0AFtiUT/E1LR66R4IuSxNmZRB/wP9eQO+RkatyyEE1fYf6
xRSRno2AkChvaAczLpf7+BiRSAH9BTf7GBM5Dn90q7873bXJBGm/AH1pOFoBN7J9iQmIJYhWC+1E
P3wAT3fvwWJ+NzMUauJ9dYbuyIcuJ073RTpf7ESyHnf0wsZTv8MhnSJDiBcRmk1DAOZX0mCKVsd/
sEuLBDB9QTTEhzeODQN0cuVvbkjXvJXcYcqwVlip2N5JAMLVG8xE4BAbs0r5QFOh5z5LEbpjQ6cy
V5MLWy6yEyE6XruTYgj6EF8fd2xuIX0DikDbnLxCGPT84YnRlPhkxBHYYD2UpJN1oe2JOROVBK5h
PpWN+5/2DczNTE1oULA7i79p/DwY9FCnR4W9/KDMiFZIJ/IzHJqUBnBH2Ow9ciLSa+34ESufR1Em
3ssYNi7rS8+qkdJwsMsWdB9yFjejrNK5xsEKpqgTXmsdGmxTFZ1Npd2TnMjlTPROnzCHe/cBTJz/
zzgkcyyvE38Dsa8UXOzXoLecH6GODDacoIRyP165+5TcKCSIQgpfjdQWAmT2eedu6G6wVBr2vgAw
gG9nVlO7kxptbrhQRNNiFl7tljp8mipqdyJi4b6p8i3ryAEPWGOV6ij+YWEhOdoOQn6uU1s26YrK
HnJyXbZlmrDLnsOwsYxX0eGzISme0PqVI5wnPo6WP3NfDx+bT1RB3jTaHQFfwkiLubY8SjR34QVd
VndaEuP1tUuHZLaOLINZLcZzNUr3htjY0UIZaNyC714wDaNsq6JyZNc+E8HElMcZnOMbBWp+6ecG
+penGYnFIHbT3A0+dfs2CZuBZpadKB+F1mScnF/VdYJua6KNeNHRzvrlxWk2HjrlPmBNu70mbJe1
7B301N6nYDZRri6+3tdLusX7/1NE+w4CWzkAAhe9ltojcRqeYyIjEBPNM+P2/c8oZhecKJbjPzFq
UdgqPqbGTETxCoeHTf8COYfEZj31PpCew3mm3piog0kREVJsvagP3FTk+yLYo82pATTpqh5oTDl3
aJGitlLtA7ZnucGsS5GeNpydSsFuqqiXXOhjx5QqDkpxz29OGjWM5Mf+7a/qb1tDPvyP9yfCgDX+
ymxfx5XRhW0E9IeZQd0KordJh6mxFvNHSs6HNVFL7xARvc+GcIi9PyWkNHABWRvMsUOQK2g9iv7x
YMDIGU8fjD7lzrKgkOwLRrdj6HVTKIYocQFPyL5iLcjd8W9DWQsRxtfzML0/SiLId2h+N6if3gry
wbXRDBAJaEiwtsiOj/pZUsNjVTVuLaSQQPvUUpjSmttcmzI2Kl8dU7/DADWEMnRCecfJvjxagDx/
XL1PsaRPbzzx5bDj9baFuZU9VhejPPphUlEUg1xVWg1E0zPrUtnwB5y4f2by6lk+Hi9zwB1NL0ge
MbQUCXYJ0zpVkqArwfI/G4p1eJ8ukxDPOXsaCwpOtcPnAUEJMRglJbC5RfWU1hiZXpnrpQzGdCyI
Fvd2Z4Rq5LCtMt+ES/fBsLVBUA0yC6FzZIyodZauGRqd2hSXa/SnXsgMeyppgj9DMUbRUv8Qcgck
XRvWaJIHdfLACvwuun7x+riMgRoDfTugri5yhyI37zkzomQs5x6UYWK9aWAXMZQqBNAasn0zgkKR
LkxPAT/P2FDYGTf2CM7LzvwVKH9y1Z0AZBncW6ICLJ8XVqma1TJb6KqL95i9xNsK4VxKeHfV4pKG
vYRXf9TihPY1h/UGkWpPQa6q6G+EG10iMNd8nTA5XngS7QTXyd4xH1uqteNGOKJJnuEINAsonYcm
ySFAkvUyPCYwfSyT6y1ZYAwq5aMAy6OvoHl81Ra+62j2cAZUCzIGEHszXjvYTZzGkZ6YnRF42S1Q
rtdeV8mYNTkQtFnIZgoQaRwVS6LMkg/KUfMqs6/vF0nEwvwrFDDiAbq8vdPMK/9nUTLB2zm+1w8M
Ck14XibLc+qJQj5IZ+RMpPdxep90zQ9c/xJI60jZP/RxY/GWgHFbnnrJ75kUjV/5FgjaazC1861c
pVXucqB98birnqm/xu18OEOMwIo2N7ybnJJo0XBClTEP1LZwb3j+dHJs9hvKl6uiupNP5FEPryEX
VqayOsKNApY/5LeARjBw97GhbgavrabKMIXWfrqrMj1GQverb2LJTo040phGi8+ehsub8pN/BnlH
srsfYzuwOXpKGnimVXdopnbRvk5aQZcmfVi1hhqiCv1vS+zVYZzqZe705A70Rxoll2Ja0ZmjnYpN
QIYAXn/8cYuwvZtXs1tox6nQYmUsMgVgGDeqKUWBVnydHWimP4TMvLwjD3ay9KUwdutKXnqOV9Uu
GKaZkDukFICfZFSfWp35h6ZEskFejG7AjmnE/whN/2EKapXsWaSoN52OXoYqTwexEWcfNlE+9XDF
lSgBNXmjdMHSq0bnGM7m11bDoYOxrYAVUOGYB5SSLW1bvalEkdqyuhiTwxgMI+KL7fPeqaB+Ym12
jVxaCjbazlbOh2T0AwyLdy1cL75RBRWys3eGepSjM0jBDSxzLVFesos/FP5Ac/fFqIW8cNyW7xos
GIfo6i2x13iTqrAbNQOaVu2Trxn8XxFkYr/ctt+R8MNccGCGAl36XE5yv6AbzgksUXHsWOd3mTMF
IRl1QXoiPZDV1Hri0yaym9sclHhy6CaAcQhMzgSZsdTXZOuAQ+Z4fsflBwAt0lxFOFWzz5JBLsKH
+ZgnSxN/JW+n3T31e1+MqJ0Uz+sQGqN9rX55dz+DJ7swqt8O0cdHb4AzGB89xZG3XC7M2h9FGgOm
97TzzApxqP6to1GWN5R4ZE/ivJbY4D6Rer0a9DC5ybWf4VYzA/tJeO7VDDDPkoyPR0Dz8S9ew5MK
iqjMz68KM6vksMn9UT1vDvom0sAJUPjLSDew4oLEwOFDDpMsm/6j2SdANUVgB1uL5bnbs24uGMXo
2TkGRgfBVivh2lJI1UTDD7sj1ukjTImyKEs0Nk80/y/B49QW77YffVY5ACZZB/ZsEveTtZKThrne
0o6esSY9rwzx2eliLQlwJi/0VaUU95fUlYpwkaW/PonGW3c0PAho8UNB2Hm1LjECoYJPTgXrTEFS
IRRW4Hhx7pQnTFSJgnLfSFITzy89ephBITXVSr0Bkc2P1JlGCb35OIlRWlh4+6ijzVYK6inofBIh
yFIjgaYt8khXsz8dVulhOnpiKcFHmmHX1ylsd+/sPVtrvRxMKb37ImCSj+kLx8PrZp06DAA7geSo
2xGkrr8/SfBqdCVJQ4VRcJ6pI70nBnkmQWsLvabrksRlGJjbH1J/gshmKQp/zBWH9vfCodhglsou
+qp/flmX8S0KMtmMCVkmst+DkjtfrI8nMuYC+JXK0oxpw2FUQkxgwMOPs5UdWVKGZbYw+v4FX1KB
4Ri/FzYPh7tjvVEPrLBxd+4S3FwEqR9UauLaVnLbgi4UQj2/41uB4xFmY7BucgDtUaKZzzUbanJR
9jGiuniFMw1T0sZ41huDBYr/Ea8sYm6f0l1j69ueSSo76RjDVxWia8q0Ijkdo2qOO7mmNrkrCeLN
w/bAvMZFuIFifWk7qlo/997SMvK82O4AbWVIddLJfHUTLmtuK86UiKzSaGWNKCM8rFOsFhMRemnj
/SyxLzQsfKIZCBoDt7OpY1YcsCOngWbaly7XbXQxt8KmlavATvO5kY+5jLqYbEegMJJAYyg1GeIi
sU5SrIFjh64B8Wvecb+gn0H6Qo8NaQrskQ2Zj807yFd/MtIHlfuxdyTJ4LmInTDtpYI6L5NZi2hl
GjnM73xC9Q6bx6+mf0AwFbYUwbqpYkfTS6YX5C6YVRV/6BuUvzw6tRVCk214svt1MwQmZC+L3BbS
MeccpHug2h/xS3jGG2mv++L/azg2f/I1vrmKx04sh8rY7+2CRkEyMCIYjMbszAMrDOyOXJATY2TL
6YT0O6vcfVavvJVsXlBDYp3l5owPexWJvtkzW0SYcXLHrGyA5l2o7O5mFZfs/4XTZ034oZkrI+0s
djoOY6hGpPvKoDhpHiMqKlJwRyL2ZjxlgWfGRzqCtG3xE8Yz24UWHipR2gMu97fSg560+MGNlxFS
d+NM85SZLI9Fws/PVd+flhD5z1Ltq3RHrdJH4OT9ODiUo3OEvz5uX5J5GETl8frgh7RrE2qS0uiT
72mblsnz/r5Hl0HHbWnWPfU7r6qu7ZIPMOTOHN7yR4b3Mov3ylw3KlP0VRJSsAbDLkeIgLAK/H9e
ucgE/ODDgxo2tX4UzZPh+HEE94A5J0dhFwEbCiI8U/UP5H/yzt8WuojzIcR1FYBK+gf3XDqTl1lG
amtxKP627RiXt8K3uW+HQnF/kpCi754rIi5hZ11jrAdXIXNl1HJOgIBbdofACGPQf3gRtZgNz7lr
3k1zBsD5TQDFIsln3gIncOotVoZzHVpDpkj6oRH29oluIw0SzS0std9sr4vHtHYlVIhyuxzM1Ig3
zqusw04AEk21op2JI58LvIoNYXz9g8QbpOo6qIqKRDg94u84jH02bpLwwIZW5+Mk5iizp0IjcgVy
kHRIDkd0D3wmqHSgXEnjpYsgGvKpfPwuXk2m2JM4R5JesIaEXFkV73Yh64xuPWRUd6WARdySD/ax
Qi8u6YwAQVg+jFU8C+/hrXu93vWVjama3l1eOQ4TktaDitX05VF/ms11ad5Kfp+0Aa5duYWceGYS
/oa2q2YCrImi242I0E3Kw+PNpXT1EkkqAmURsWH4cSJsrehBaP+NbuyVsoBGGfGP8/euflQ2NPIe
O772xwKfdD6av7Myx8lWNu7IIjEE7AcH1Pf1NvVS6Y7pAWI9NGVsNjmGJBnqz24Iy0ksyn3mtU0P
lGPx6DRm4COFhHHraXJaj+qowc7VmvHGQ97uKnxJBlt8b9S+kGmzUVwfbLaNZCckMVFQt3vnvyzc
NW6xdnG4uFo1/8gaJ1qgouS8vEWKmqRCldRKGHGwdQKV4poo5S56tS6jfQ63HhPnKvgt6tiOQJzv
2Q4iGuXi7iVKSCGCSfk8AUHpReNpex8QjIkbgq+J3cTLDG9gb+G0+pyViCBbzic+wLXvu0fJPfKG
zhRJZOI2KbfYYk4kvOKAsxXHN+Jy9qaVb7l9Wc9IELjVU69guby9xiizbUfSzWzn6MHIcg4vpKCx
06fOrdO3TisxtS6n2cUJSXVeHK7H6RXjE58sUnXd/YsC5wIR9xYQijIKZWCpIuo9qGkfummnI2hd
ehB/nh75TbyYQc6JIONOtGVmDieu2ivvuwFZFyOjgRDd50uo69nE3Z7hKZgL+d7l+ZKEnndsjvLd
GCp7KQ9aR5s0d5bTkKnTdl+wcLsup18wryv4caLUxftNsmFLYYNVhxa53Q3yBPJCrqX3iqJ90Q0L
UI3qENzGlQ9hRTWySC19wmrAxbDdJUeH8Cwf7drPMGmWpAFSmHGMqP5UATsm/zWcpmQ/a5uoZcWt
wVGX2BXJ+6iwBL4dVX5NYSjJVZtPob7Q4f5baDmN/7EwkTsorFxWFkelgqUKCqcIkh6tKfHLF2En
/cU5djU9LChhu3q9rpG1HMNYHbIhODEzQYOzp8G7wO05A9solRPnUUqHHXMcysReBFs90XvXq0dH
Yu6/14PbCgKkrsFsdYw3LMarZhlIKihYB3nCXGgm9h6cpUWa9AQTI+9sEL/SYMnDQGkxr2OXn5Y9
YFPJwiR1tJQ0HKzuAn0zMvqMNdWQFJ9xgex78YryFnq4RCpIB8uKDAtuSG6v10sAB9FOfhszONhG
JXs6caeZ7QQbtzFrDegX50XgQ4aMVz9tcavs+nRxzpK0IQxyozIhKUydbNhMCOsAcfhKQptxA6rb
FOwtKd3yk5fcEN8o6MTTVylP7v17yfVd4zOMrhfbPvf771ZtYp2suzHC2ibhwqg8KR0Q+POfE4YB
qjwFIj0GuP0m3ZAKvpHQTAdc35TfC9cAydSuq9zjII2bTNga3ejmsa4wqMaLO5cW03jEe4SICVIa
sWpRSY863xaeIWqb1zpbzGTh0zI+mXVlL9bhSObCkgfJO2tJg5mBEtGMgC+kCk0fpVxKu/VrYcsj
9Dq+ZJneSizHZxVNrMTf8ez/4SQpdeTpOfJtV1C6TvDW5qWykxZPeOuZF4dYxmiAd2lYzxZRl1yE
j9in6HWi2Ep4ihyn0QMmJ+CSlqlU2fiuy+OKGYby2ygYXx77Bd8WKgpk82Oyl3EuAfAxNdpfvF5v
hQyd63s5kzaPEsZBads+RsXqbLZ3nGm18lfGpzJTsmP+Xsouvf+fnS+pNTfKG3jaUDqlTYnIe01u
IXRNoYgFd2QHTpKOSl/zoxUmPIaV9j/+QTvcmysZ/RUmjiaN8uzfawo9laYGECY82JAOqzCW8Qxn
Y7b661GwZYfHDmLSCn26420aumJtv9Wh05rdtxH9lexXMRMwOtdMfrcqxpFBHxFIl2VUfeJXNJ9c
27sT4wc9Ki45/EGwtHugSNEdvMdzv/Cg1JFr2oN9WoL9OS0g2Dd/UlHOcjIuBMoggIM7LCZx0FIu
U0PkRAj9nQWLVoXWTfQ9kYOPrXLGdpgqlx4vyNNiVA445IBLGYy6S8sLxhCTd2NdlNCfT9p0g1fr
tYSQdQi7wrZ8MYOD7FHre5+G3M4diCOS0mqyimrkKFOeTyQAiGGLcOM1/9GODXHLoyu4WuQnwd8m
MCflUcrnL8w0dqQFyTJQ7V9K5F1P51skHGdHcBM9t15n/ns4ctbBZO4fmGbLk+IcjZNwUFY/UnNL
3kzupuU8PyD/ty+JGX91vNQKYuewChCDQq3tCwcypfjo821E3vASLMOVw/gpjaG7NmpioKX6fc3e
BfzV4dn4gbPVl3Ee5Xb6NfR2lytnpfGBM/f+ZdTQGB+UjuEVyq5lWnpvD3zK2TfVIkCZ5TBeBFNY
t8IDEvzIIn4ET8llj5XTwGlAYUe2zPRZzE7efTrSjxBBUho+IhNJLMOKbTD0HFN2SZrnch31/zpa
+O8RTVtyz+j5fX4Ew45KD4/Jm62vL9ppdV1eq6NQdKJ84KFrNBLMFZBuMEbxbABa51i4Yad4ydB8
qqCD96rgrOh0ZBJkuTG74BmqrexYMF5pLRltRc0sUAqX6YNP0m51exBOZpiVZ4tcguKznHVok88Z
vFM/EWyWQiRpk7/893TyVgQyUTyy8BLnFOb+kRArNzPADoEuVjYbnYV9xPOAs8NbcC2/dhfHVLgU
hqzniFizI1Sj3j3x5xPpCbykqbRdESKzWLllbUWQ3nub2FfSZGkBvYsOSANEAxw85nzSGdFHsdWt
1wxOwGqJZzaA65n2BHPtFX6grEZJc4nw3JcTRm/c4MOafDJLUOdXN7tVuS5yrW9DvZG+qfsrVPUQ
lf0Zjoicmv/2vioeADgi4bkDbFg7og6fDxiQmiliwL9fN66DrcHQpFnF5kylcTxWMuP+GjQA9+m0
N0C0n/6RtyvuNuvGKeihlpAeRB/wJMRvu//PA2n+VgKNzFxdZY1+yyuK1u0jKm7J8PBQXTEvDmIR
0EZhJWp4LP/7QJ+N6IPQfr6JLwrO3CZZ6nzMdqPghw8eADkmxLSm0G2Ve9e7rcOFXIF6d52LYgaL
V/t1/yu7uBpd36enSpMz3b5RFSaKI21/bWHCF9OVuZwEJltZI52nHBLDViugbUVad8SPSQ6CnJJx
ltLhcSxcLy4sghRWdgEi7iS+IlYTW/mxeX2vFa6liAYp7KahTqZb7TLzy7uTpyV20ZxgnQqM4vvF
MGYzhF4UrkVb9VuWA3VpJ4UaPbmWVYBi0cpAA+gn0n3ST9PBddIaT42m0Ko3p+cOP1lB5gnSSv0L
EyhlsC+PqEvfcpEkQkytm01n3Q6EjGBTj4fYhqiVVy8u0pWCdE3jCUx3Yn6VytXzJBgP+rgrAW2k
D8v2y3i1IvkpxdJ3LX98g6eYKjcodGua04s0ZcLXm8R3P0VAnBqbUj51lSk8udXkr9Hjc8MC9aO3
mH7BDa0qxvccHDQ+sCtGotK+QDQ2tA3PTBl13zqLv+N99thQ0i7ZuMpXkM9DV8t4AP/0KLj4sPbq
wIyJWLmdf1iHMC811shvx9aYTfswGLGTX4eD722qQmL/J41HbxGlCuKEbl67rMCg7FsknKrohT7M
tP2LAdO+3MY+Kk2c85CYbuaw1p4xXTKHhkLGrkRIJrBJ57+dHHaQcwa4RRY9hMs1tE5dzYJZi11b
f2YffKWeo/SfNiq9NOMum+dHP5JDXWB/kRp57LIU17Z4/mJ5VhtfAzmi/VptLQYYfaiB+J6/nBpX
xBTWGyi4t+iqnIGkGSk93SmKJ6PADlq1vRbcVxvFmHCVznJUJutFgH7zRxia+e/izaHGwghjqVgw
763j296wwd0PvEgMIygd3W6hFqXYS8wX5+J4/O5ObasFSFTdRUgYaTN47R0aICa1CkKZZ7YY+djV
dKTzGNX2mLrvPR+8v5nz2aEOs4wLlt/k2RZAdLqs0SIeykbXkC7+JtRCsyYtAFOh23N5x8CkXmpS
Jxj6oB68MBB2zey9p6c4SIfCExdGDVop1FlKmcnnYbMEZdS0GNBrcoliwzYwny6rvOjCxzO5JZXg
61KXk04SFsmLO8LyrLybvQBmKUjpr5wDRkXY7LC1s8nOI97Bb8cKP2kONsvYsY6EijTNrzM79OrT
j0mGZJ5KvwENsMNboDWvvaHaHnYB/lEFjH4EyE77nkUHa9Gu/lU5k9BZaquFx5+PHNzD/g5H8uRa
5KB0pSlUvYK/AlPeQNmAMxWFS2x1NlK/xBLIpmYE03f7jCPbgdtsE/5FFZwLZRtIldfiLxl9MkDs
4vdKi7U1eJg+sIIIw4ZWfNiBCbrniIAj7TRXbljpwpMa9te4uPFXMiq12Co0uj8p9gdkxtc2PxGT
HTQ1GWJSjz46ymNuKiutFuk19M66/jqaCMZGHH2hg6qYyNzVKI2EHgzWpYqLXN76JZ5tXbGs3alq
D9lKO6PH+AxnQGB0+QJKA0A/BKnVQF3lEf/vB8NNxyxmLqyzqLd65v8Vo4fIG9aR/0TF8xKcMPgv
Fv6H8GAkuyFzD+3wgSM7Tv0p6ieXN5YwZYZ18l9NAVXhHVJRnWeszSli5+pSXe8hI4rIFa/OIZIR
hqaWyzEQwRVHBnU3csv/IYgoedhZ9dkI3q7th2YiJyyreXhwpJPla7e/LG7CvUH1166KCcmMqmtm
LGmWhRJLWeB3ZGOG2ocrUDZIofxzFJXJ5ZppX+2BB9At2OMrX6+e3PMHz+YQe83EBbnDj3dURcns
30vnVKPIcy1wQbNqmmSSkCscky9PxIq4JG9VHdqy4YmBrgyOrz0kNu0G2mz+wc19uMBfD8DSS7t4
53BkVl/cxkFBBJckTKNsyLIn0T7A+N+BNTQlBahRrR5uHUNjffkBQFTiCSh3q7uCZIwMGwyDxJMR
jsj0Xg1DwvPPqbgzOXiAmX3uJSsT99TXgqZ8o581WqtVgw/GoQ8SvGEtpdU0EF6KDkEo7xz/85hf
PNlHibEfzzmqG6PccZ3sgoxwHGKkhlQN5dZXaAm/BGeu7mzJ9i8KGSMNTqT9kdGAPdXPmaQ9ZUko
aqTwh6C+ma7VUs3DTjEQhdYpPW4oDLWBlqaP2DYqnC5QchikYE59oDW88VaYXpZ6UKJfogjKFl0U
90emgl7Ghimgmr00M6c3Qb9YEsDP5Z2V/rs0XBm2zA/TT0/4OvrjIF5MEm10mV2sg6hFHavuVv9h
wCOoKVS6O6/1U5Gj48ACDJdokBusLmfeSFKD1Qd2/aMGeDKSf6AyXyJMqv699AoiOiueo2LRWJjY
C37GHC3+6rBsvajoNL05gtNnEt1EJerURgzfqML57GKqpkdXC5Hl65Nv6IgP9qlmct7sQoACn5M8
MgcpUChp6cmKN3fFz22JKgqBceo7C3eG+PkWpIOYMsoWRWPHXFhDD3O8ONuGxFE6wF+XsngBQkQd
/hC7KmteKS0MbfuhNyj2T6xFS5bONTznkwKaIR8fvzGlJFE83PmEZkUHmoNN9+3wZvWsqbe0Akzx
0o4CJTIKGYz+FaucczvOV3sXZ5LDGnrPnv2RFIwTjE+qh6hjIdSna9DteuVXIoOUxhdhTZfJSRu2
PPvxKzcJIB8Jl9mHeColh1wbneMf1rUtzk+hEcsw4SOXfwirUPJJRmSzy3lfFIIOmGBEICXCAgv8
kBZjcARrrQyhUeFIZKtye6AFslVeoj0ScWLfHH2xuja0xUpUjZzcFocyY3lYq+y1LLRuCjGwENPP
OK/vk8hJnLUOwK8U9rSD7rvoip16zbvTmFWXPEQK1j1RVh/190MhvVvCQDyKiLyZwqu4pG4azUAS
RmYrHGiyAMukPNHtSw/DgKkpT/7tXzhcs25Qf6A12z2EsxpJwLKZfGS1bA8u+Y4FzHjnbLU0FZyF
Ke1yVeh8zG/0K1f+OLYUofFiRotj+PNHNNdYe2DvigUuNbYmssOEkw2OhA/fkDPz8r1XMcXwoIZB
PGnnp3nhvDxynFUULE2Gpy4jCnpog2KNdGlbrBeJNt5Wul9ZvpafMY3rFrXLrG68RBn/kkPFPOhu
ZjdM41bM3UHKv2nMB7NpFXE/5+UOSPaFVP8L+B8qhL2XnzPtwbAjdmCHmAmpIvFzvl01yaYfvN4m
giM0hNSok6sMYao+KcO8j9U5X8NmwQcrfI3/X15i+Po6evF3n9hfoJ1NYJIV1fxNqb3XlxkUPZf+
2RieYGtcqnBqtGTW1iD7H5CHhMOMnE4KPHEjBA7cn4soJyi5rbscbsaZn1Z80wCfzg7REqH7IYnc
5jLcyT0rFkt6gw0ZKU3b7DL3wdmq/rnYZDzW+4PkMOkIRt5Y1N0947MKAu2NTT0fnNIiuOtJi6Gt
Bvu3kiBWYFsCSUQCsyGSKpszwVSbollhxiP4QvjiExAN2sguQ4/a9dokDMaC7DlRD+vG87kxkF+P
pKFIKXAgkOIUMYiNC646DpEX7cjxBUOQA9FTEssQktSbqTVaKWhhNK0YpfxxWpXBdBEC05zAq2WO
7/tOotht3ShfAqXtU78HAC7tNEFQlT9T50kfjqQxFl7xD+gfR9E4/9ACmYVXkm8GbcCU6IdxTR25
spnsoBhVry+FfhA2zQ7aIwAwZPuXKVuOSm4VN+FVy8kQ6IMRdjxzIncYnAoKwSkN0yVKE9kpF+eL
6ZouevvnylXeWSnRPeDuEquJmkKy2Tx+eb8S/qiyD/X/7cdGDnJURz6102XH4Vlr7iTwJCYWjvA7
wQiJv8TNf935HArHQ9B8NPamkT+JkyfoQtPSg2aCtJxYUKg1+ITY6eDaBJJwQ8ZkcQ3aThQ/O+/A
vkCZHKi9RbpojCRCEj63ocdB/iHmih8CRwqEraqed0XbgtsSgkmTwRcSm8X4/6z41TOAalucjfRG
SRTTGa+RNcDQih6wtdM/3MDxZnbt/Q4AM3HLUKliKE48UbQScl2i6rWQIMUDpZiUJSx4PL4t2xoI
t/8IGH2ZDu4qB77NezG8yer0tEPVpWPdL6JdjBFOvhQMQQC1oHs9nvaKkpKw0WU6pFcwM76uQhqq
JQI3OFVNWueH8uLsjdj38o6re24wRyPrmvkECn7zBkd+XIyYlAdX+vrykthGh96ePsC45qaWI2GP
opT3ooP8oP6PZvxyC1kr8AGVbJGJ1QNaHe8HhM4YIN2JX9baGaZRynuJpJVkcz1jbIGQlPpNur5I
2+EKfzcxUVDK4YoeGFKSWAL9XG8LNhK0nRpvoESTj7w1amq/oedjAN7rkNysMyGNNGOfkUk5S2Xh
YaqoSK+7OiPXpcwJAG8A9eeyTA2Cfl7NUT0nVoWxtGaLkZQ33PNgJVwiqYC+13Ni73L2/h9i8syc
vBNT2l8moXFeTZ7Pv3a16gJLv5AMlfbYhg+z4+ep6Gr9hClBaPqt83UwfNN7uOtSkw4Lg0CnkJw5
rRW6YDsq3rA3J2yJBLz5LV1pQj7OO6gdQpPtDOe1yAGXa3tvD1QnZ0bbmYXB2v3KhZVvdiWuvg9X
dmOctPlrbTLUx19Vx1YrdyFLQ0AnTQGZ3eEZxb3YVzdwIr15yy55en+AvDeVpzmqRqBFm2ZUk/no
0CiDMJb1GgxxpbC7K9mU6XD1BzV6j7n76awkEBSxSmLvmOhU/5MEzcD0+ZolBGy1KZrsuqAdLQnT
LmBW3wRPEc+Eu0nkn+MtTkyQD1xCcAaqIwNgjYVijMhhjgJ9b4AxoFGeFEokyxLqv/q/81nmdWjO
6Ka8YYjTq6VnhcIIXU09nazlY1uih7NF7mmJjMD3tjk9tuCvx6HuGB0bqhs+KSVKg84vV/9/cFQf
dwoOO2HMJYndT+UopuF3nm9ogDWt5afsojDLEOCptssewqqMVayDocPItvBO2g8VQrLIZhg6ew3V
a8mGS8+z9KYqqbhLs0TNcxUDMRcm132+ScbvM6JmmpRIlpAwEkyRqUeaZLM35kJqA5B6ivX1FAiZ
I06eqx28+jtJwVhfx/ytRjayHrqgqdyRlIGi5MGzbDgHbYKwRrU++j5Yl4D1EHCiE4rtHe3JHOmU
genYzgSZIcU1aJyJn2EGmW+TAOYl6qP+8qlXjNR9Q6ipmU5WXIi4aBN7rvzKVYPgWSHaGEdxRq5n
j5RHsq2JKfEDeD46Fo+T3YbFdNUKiLkWXEgIqrVxGUJOn6PEHiEFTFH+nAkuZFFw4rZ3VQ9zxp6I
IsUOSPfWnsiAxm0QcJD+t3wrbluInDgBJDDNpxtuBA7HUQb5fN1hiQ7btE1Je5Nvt+AjVglyNHKb
ncTdACmVIuXU5Sgu98r6IWBZlLfAy5s3qcAe3WexqE1/AcG+SfBMUA7bChIgyju3CVC2hyQx8Lj/
Otqfyyv5WEWmds2X4zsMIWLITxCaqEG2wA9T3SrCAiGqNqkwPqz0VsJ/jjiyfxROY5DssdsAW1aj
6kyQXYZsnNl3jnzaSPu/WbhT1CF13ezHZYYNgKBOB6XRnUajtO8ybgleaGjAjmfJCQi3NRCAiOMq
QzO+LL9ry6L7Axy0mFhQ6+VuxWg0HG5gaAhSYSNGIt80ZOqPkt+fffuuJantwEDykszi01hgr/I/
GAW+2JFgrNXupxq1sMj242wP/I30l90YJ+FN3v7sCpfjCUQClWkul7PO0j3ZkqnN9pPblSxzPVGf
5m+TSlxloTc8QOyiMAn88wNSerj6JXi1DSoWnppR7SbfVBI8Zs15ztvvB3ovY7LgTZmOmjtSs8Tv
9iRreCpkySQeDqaBJyse8N44T+ELIF/9008wBwTNxdU3rb14ou9ighpA+Cm/e7+NsYRyAlOsNmpW
FWk7E6ZWXsoAkOM0TRldckypBPhLg/13sGE5dKDf5SSbAfQT7JgeLVpb4D1TxnpWWUoBB5pfeyb3
3gnadpuFsZcTsF3oMg6cKznVBxgoKxW0SyJnrmuC6Ivm/ft2yDH5q9d04F703EHcnzcwwoXAWnuj
dlE4fYk9waYU5EzGXlLykD8267kWk0NRFK7dWs7QLeUPzdNxMvUA4g3hod1fCrAQ37chw6grB3nd
oYbT+YpuD1VYwujuuPqAvNFX4xY0r/GNXY0PfRFhwdOn5mx5ZxZPuH7LRSXzxpX7to9g3trtuiSR
XRHCB7reTw3RjJNtqyypBv3fM/+AofVs9gSWCRKoC55CNogtN6O29/uGhohqoseRpwoWYXP7CM5b
/NYV5jcqGaIflzmWGF4KQaHNaOn6Fv3lUH77UcgYa4ou+Cgx1t5eXjKFcsAN7ncw0mF1KO/DEArw
HPL1L7rHv01g7yK4lnz7ZSqiIJeYz1sVXKRPI3vnPahhML4hTmJgmTNFlwj0XG82HCnVzDfzlKLR
FJS7bMY28HGkMdf0cP2kYlQdqyIgIMl7NnRGeCN87rgA9XUiMFyPXXjJLpJLN/cSQgHP5jpECg39
deACL0Em4y2AuiaOKdgZOKtfeM2tRB1nOiG6ZEKe5RFhzYBnV8GNr6y1CusiumGcyisNnqIGmqxy
0ExGUlm94ExTyjsdR0ULtX8hY8DNFIYZaC3E//sU+LLPR61e09DoGU1S+1uZbN4o7WsrrJeY33Ub
Z7i3FcCEsO+pbDLuLeyDof/66iPBOnCa87udUX8uDGNRlGSQ3tVuYB04pLlEG6h9/Tddhh/KoIEn
qzRMxNDr5EamDcy0dSIGfMiXDhQNGvRlHNPekOg0MO2+NGvNcenGFwB4GqEdWF3+KZJS7QXl7fZq
X/WGy7JrPwZXrqJpYnjzFSE4AO2AY0Vig3oEd1IkFD9lO31HGn850ruEPch07rX0QSViOTJlcbeh
3WiwTrNTRh8OR/DbdbSnp6HG65TRMYoTLqQ9Pu4Xv++fJbHdg7P/+ySyu0reKkaJ1LHodyHW1UGD
lKOb49hNmHARoA7wlrEGKKYEjiyMmZDCyXI9vmzRis2TpOF1VBiO0Cg56ZU+Y4KyrkjagRRQa64F
Y0cJvCYVhHm/pqW1cKkNjDpdJt5rmxne7Llq4Qq9EOz8i6qUmGPDz33Mv1aSBMYPrWLRjUY/cPQo
l3Ve8ZnVk4lyOpKpEjd7XnOBbkZQa2zuEgJAqj8I3MdnsuoNzQrZs50N2Q3ps95ml0sGNVRrC8Ho
UbSw89ttWgu0zkv/d3OJMJoRdkKzM+CVRVj505F1I312SbYnOLhxyJ1jRdWphIL/YS/NEsbJqe2H
ankhlmqv+aH0PpO4Ou/RACHB6UWgMc87Ei3Oltzlwo0XqD2bhSAmEKb3dB3HJU4OKkT73bAoCdzd
CgyuS1svUPigg9PCLf5e9lSE9qY1cvW45kk+nFaq2eTx4m+QFx1zLw4UimoWMXl8wMjwZ9q8+JM1
8W+DIoUtwlhVeXdd+XeJA2PeqOwqsG2NqKMgvVFUFZhLB2MJjuU94KaXXqxNbnR/GWyXv6h2vZD8
afslWqkug/oQpvY5cFNa7ZSy4cwzD268xo663z8ynNJ4x077CWKe0ZMas+T7/QNEv9K8XgJ6zIQm
x0pOcMqTd3on0bnS5r1fKC5YWHkzPLcWO61tqick9u+j4Vbmj7GA5+ZFu09bDqBurOHfUnh+v7AU
56Zys3kenOlghGmXDFQsipG2PZqrMP6RhHHeazB4VPI/mm5FrQMLFh4Ng/uc7rHiKT0ikBHo+GGn
Lwdht/Uuyr3WyML/UEN7hIXUWTpq3xFN6x/HRplmXWsTFq78MAIUOJNc1D+hR2d4GWZNdu0rJ77c
ZQQplJEeb/t4rcGRH+CXGULtF7dLLPWBp02sQ1o0HrK7oV5I6tynAk4dIB7pds3wj8HjNM5cvKIK
dm3cTZh4Q4yzJTfRCISJdkPMbk7n/YOCxJrO+DFnzARlVBA4bgoeUnn3sYVDmQM6xRrGQwmdMJPq
EgoJxarrecHZSEGnD9crn03ZN3Jfnd80xEYP3unGjoN5mIYyIzm5W7vJhT3eFw77gzZxasH43uRp
znzxDcMNEkjDw27csbwzw2RKqSMBcQC+KgD6pe8Z9SDDHEf3d8F+zkSquj0cJd6QBqCu7SkXzgJx
Fa8QxM1kptJ2NE38EomMpx5051IdgKFG049icAuoV9EVZNpA/LBY0xbDxBbruxkblpaioXS2IhCF
MBk+aRAMoziPjx++BlH84HNr75SImdNHsEBb7vGFjINwskRViWdBwJVKy5GDHSH6DTrFsznFvvjA
h1e3Muo/fixjxlpuUa9pRNQHhcYm42aP6MKXw6k6HJBP2M0Z6cYG7HgusUHIZozIqYujiYClplFP
7MfEvTsuF27zbQhN3QyKHllyEYcmrW0c1onqy9FZD/1yCojIXco35T+Qb0iTsPhRkPHVDH7SeQ1f
t9GBzqI8CtG791btVI/YcI/bJjU4ga2q69G3rb2NznFq/76dXf56dGqZEKmMgWUOeHAQvF2wnFpM
jIr6kBTA2JOodOtJIKWHI2Am/4Wvrbh0DWXOCXZsZ44XmmipHsyEcqNHR/3mWWVzg932zDGhEbiV
HbufFdW1udBGJxlyYadWcZBf4Q4Hrd1+GJHugwdL3tzBJeKVIbhHiWAPgSh5+BtvUrQdXERzw5Cx
UP76/RSoEpDIRKkAu/vk+ZSDSiF+QNLChUA/jc1UgYtUGzOZw/4HZALodS2gFGGVMR64G1ubCAF8
xdlDmIRAsl7gbICya0reJpStzHBMxEwp5ryiqAtQzukLPHNvfuXb+7eagHxQO6WKP7/Xu6jOo2jT
AJtosx5GtjH8bcH6Ypgr7kqSgVbnqrQkuMP8H3cd1VtjfkpUZB/rXqF6WMEE00AKmzolgOqbcBB4
Ng2545GIo591GJiT7o4wuz9wgsJZQLClNpSgN+0G1V9Cpo4ws/npy8QoSFevGZym5/QxIXru+RCc
Qn2J9msKdcJoDza9tpi248tUzvlH//9YgF63gxaxFpMomHZB4r/gztXd4fnL7HkwSWWwu4xP62pS
uSVhe13qAQs3cDj2uteNKawCauUVupY0LHFetgHrruCaodKCeXSo2KQJAvYNTWNRBM1ptL3CibbR
NIlALpT4MEsTEgNabR9mxw/MHDjeZ3He8xOHtALwtWgLRxINJrbRXbCoIDkRtLc/66s2bGyUXw/+
7xKauT6GIUAEF8z2hRlMl8XyIzNMWkFnSLILp3sQxkeyX2MQKddJzJ2vXsuxFYCRYGELRq0CuF4B
cJmAqOYmjqSG9w3EaoN+nVdE4Ez11h6EFdjpOxZirJdVeNGHXIzuACKih+sZ95/IIqlXlF7b506S
tAv5dNfXbw9qS8QPjIJMdXaD2kIyCrLpebiA62YsuRYF5Z97H0sIip5izF/H2Q1jWwHA/zUW41ZL
AZPtGunozRbLFrvu5hWHFZtoXQrS5D1cA6bg0YTK5wgzZwZQnE3/wjYT+PyeRzQyULu/VNa+y2i9
Iy65hkhyhNQbLapPq18SoP/BEMAQ72sTN2GGfobirmiUqGmFgP1lo6jNrBt4A4jShAhQr1bOmPNo
LsoWn0X61U/dg0V4ulxOnTiUo4pfneUNpY/+iCWs0zbhhvhhYnVZJ+6izXMf4fvU/pyuPY+IZY0q
rw5N7InhkajZ4zIc0tux+PChD9nACDw6pOLuuAbTLQdXzAFrB1YuwxoWQVcItp3LN9q5QDktNfyZ
7WbOSXHUxHiA5IJ3YfNZwqBbRoxDMMPSL4m/SzMcMcC1lsB0L+XTZE1Bvw6NrzBnTHKrbi8+2tF0
ihVXRCcPQhEBSjGBBnLylFz1fuy6OzZBsFpUIO0rgEan4HS1UOM/P2T92XeWiUjPhJLHjcfYkIXD
pWJng3oNNuYAe80WQLuHNGGPuPTHBUW3/j6YUlF01Kus+J3gWR6tfjkvHHcXcHrXIUwGgRoS7gVs
rrPLXxGj331sgqmZYl9WmEkfzxU4ptIU5bnyxKqWzYnMNDhPddggUup7kjYbtjN80GxsyWatRCbn
+bjP2F6DAEGPipJNJCHLh+JhX3zbYufoAROGYzvLUS6Umw/cduwj8bzC9F/DMl6vfX+NegRDDaEk
6N9/GWBWGImJzpAJzd/cYEsdpAGoFDH5eXPLFPwOwgLhdTFRD8laBAUCPxkcTnHg3iCt2GnSbteG
DQQQNSkcHEGhMxfFKzSMpr7zpi+hcn8XXILk0TJy3JsMDuMGevE7rfy683xg4xSZPE/E6M6blVtp
lwq4STFjbvhAyRVBLGgeSgLDUlOV6Jjhrk20SiNxIUxhUwAX7hInVnkNXwUIj6VwnM2CR1nANd8l
yxLLK1ArDfsNWQnd4EHpKAoK4lIW83rWmgGQeseo+4IPJWAUDDFgN29nfVW6kH84mg1kUBypgSFR
rM4BXcgoKPuIkIQlOTu4Od6ZzDTuZK6Ol2qICjXeWzzKyZkckahFURpHgva6XTKgCSSXBKSrzYJc
mZyzgRL8wwumEol2ZyRZKQFY3j9C4GLjhnh3PNH0xxBno4wrhj5TnOfMuhyYNKKcLuQT4xBkIpbu
onNdLtJdFYO/KkvvwdAWK9lT0qqsl57tL0BMKndzhb0A5rfKyIAyKm1InaCUBYUe9D7CmBZdkcPJ
9Lmj+WA0zKORDePr6EtMwvFoMGGt6LzxiRs/NCnu472QW/DIqqINBmZP440HnhK/5wZkAcGF86YW
GdsSizvnM5ryb0qK0LPTcwDFULDZyBEa1oicDsO+QWMnyzJiFlLww9rqYeglP3bhdd8dgPzhfmIK
2a/b6ixeFGq3WvFOuOUh+bWnwCdtcaOOzd5CSa0QYs3eC7p0wecF6ZS67d11T/NyPoBv76TIt+ER
SUp2S3ZRpxxGRwNYxfSetK2+wlhIAphpo6oZf6H8NaXncROfrmesb8DqFNwEYgZ4jbZJa/JQCdFG
vk2/eeB4lfOeueHrSesO49zwvL7uDjyC3Hxji8XFIOqNLiBV03EZ81yr1is5B4v7Y1dyCMidykzD
fewKJw7HFFQa9UBMaBNpnourYCDbULguxjwS+5276jHLEWg5GUL4aEmjpSXDzuZwHzgKkrfFGGUo
EWAUNk/8cxddk0F0RklWoF7mHEE+/7ypfON2xG7CzFCy1w6oixscuJTS245SiZ5RkZPVp9yIy6ZL
Fg2I0SsYkRPhoNJKhPFu2aL3tb/my7EPhQah5i4TY+zBRFxyE0hUJrMFdDI4vWa7CnZO5leAvUT2
Z74zOY0Wbb3r427rsOkKbPfiRJrtbOZP/9/VH2fHsxsFUGS+YOBxiLcALSxHWm6mrxtU37zoyqQS
Lv82wngwhAL1wTSr/di/y6nB7pe0YJsxUyogMH5CJ/OciVfHevD4FLSmAP7ojDlUHpRZSeYcKg7H
XD2JeBbkMsPzi6rTI54uIRhhZL/IEuPMvW5Hyj3BlTaYmhs5EtYkUdusnieAbu4G/t1R57ekrLSX
jTsLVwSog7Dyack2TLSMHcUPfIQx8D/sGc4eXp1hguvuzGrXsLHFBv1YtfpyUUytOLWz/9k2mHrJ
zr8x5XLKEqE4ymy9AYi6DCr9WDAuuHSVXqRJYjYhmgImFtLsdRyNG8/TP0Q+Y1tFIXhh6/4YJIbf
7AzUlxuSdzldJ/Kkyr8pw6/qPl5JyMTMDxHLvU4cUZqs0SH0kAGHfFW6lAcLhjeiV3Izf735imxv
40W9Xpx+u4XXAq0+MDH+pkbZk01h95UFbRb+Xc/9sdnYSb/lkBZ+XfxU0KcL7kBAXV4CHeIg+Fyg
PBngQftT4Ic8wudpRLqv/cPwqcu+Jb2qRrvoIh7vrJD1keO67vnfi5r1pqc8EHCP1zkDgPbWl88h
0DxZk3ZiOH7W5Up/0VB6R6RZU+gPghIbfl5+MGUJn2EWvLxEJ2dGT0EL7zy6yOsmOpfN9QYmSsQ/
SG7Pg3pcLlMefxetEXGkBlAJyzIybQESgnXKZncRgO3Sjbun0qhF/Kjjb+7FexsOxA1vlu30hYYq
BgaZizcLpzLAfUiws3CPAeeVx6uK97fSq7HpGYC3yjXVvOw9J0Q5Ud3yMCsCtOIcrrIbc17GaLxu
ZT5tBXnAfuV+3KVPZronyb4/Ec9DEaeH4NlpiYWaK1PH8zuJnsUaNC+JP5+38j/3YyZv9YW0XnpF
PnHlQtMnxdC1qSmwIZ41vA2zcn3q2j7LfNHzFzVC8JBKPEDQW95AKnjU01d27sCGgL7GS5zrlWA3
M9GaEZMaqsWIBipCQkbmPrqp9B+vk6W567/ni55i+6gMAWA3JSGW8MiydsDUZyv7HAJPBZTrhcuE
MLAOZSrmt/Y6Yc8uYGs0RPHjgWs59VpOBNi7fEm8XCcG5QM4KsNghm1m+Ik6xsfpcKnKZkS9tkb5
uzO5CfS6aIXvbV+Lltug7hE2yYnHBOh2l1nz72zf/jvdRlI2qDEH8tLo1uENL+w05Ox/EIYyNa3N
nLLQO4PmuUv386+599hDpU1tOp1dPTX8OHFxgZWWYgLHjSjbZ1Ai/9lwtDXAMC6s/X60IpOtjaUO
G23jEqj4GyEkJHBAjBPV5kvlmP9lfinaXCbS8C/f0/DmkoZLFYylNjgmMkL/2tFTTx203zEHzwdz
CSQMtA95KxA9iLngu+R5SDV0Au6bntJvnajMUF/Peik3xlyxTY8SP3gov42l7cnBmlbj880aaz4E
Em9FQOG6YMZfT2qARt6EE6nO4ZRuhTkPLYK7B7mnbXpjyZ+2tbFt5mrm+y7OISepL4oBZGzDfGHk
x4Gv8B878MjWzdWwM6XMXbuasU+olEMRRPhqqyrEyhd8QYjwMqzD1i0HiZzAZHQBf9K5Olz4LFnv
oTetSDsMIekjbinO3NvfUKh2eLOCxOkM7fQmSI6j0AUELC2YfOCGMSPIzgNyzi25KzBIcNKlAx82
LE6DzJ/PMaOfdRTG3Lay/N5U4J3yuK8gKj+8YOBn6iiQjxoYDVn2R2qcl7xWrHhaR5yszVkysiRs
YNQm22wsp2+sD+fSK449DG0sWt8K1GEXCVX1HVNUDnmVyIId8WO1NYKTEgwproiY3UEQ7X4inooP
JkHDeIU7aHCbIp/wdmBr96DRkvkUBHeaZajYrcLoL4x9HSVir3rSEXYqhrH1CS4ptkdpxkQqBs+u
BC1g4a9buKM0di9+hIxtEH3/8AS+u10U35bbskZWJ66Pupvoeg3UplUFtHJ7UBMtGnYAIcCowenG
4Igi6L03hlfolerdfyYRiRlcnPm4FqQ3Ca2mEnrNf23/J0nm/HmmfB033pGVYhGe/29CksB7vtQB
oYxlpqm08knVU+pSjighcfyktp+IbSs/fPgiVmwg5j9D4MFPblmTs1EHbd9nCmtwCwxsvmc35Kda
o06f4AMuz8rDPDk+3766D4ARP194NbDY7a3jy0mvtkMVkOPLbsnFgi1FsfGKg/I5LLgAqZANYMJV
rpztkLXrCcTR+qrTBREpA3/Rnf8Q2vpS7o5JCTGmuD+Hp1xEhhi42e2VVz9faUF53XZGO62iNK3/
+mrXHUhA7XjYiPW8MucabBhQ8OEYL/cRS5daQa7a6E9+p/IckJa3koxkJaAnz44nfv5peKkJ0W5I
37idxzfAu3nuEBLBbonhl319ce0Qd5LSzuH65GPWkar6dlifMR4kgs51MyJwYsNBmAv0OFLeEdwz
Ie3Iwb9z7DHkoIoGUVoAnMmN1DKWbJxu+nsQQpeKDZeq0qrTh+zV+IhuW0Wr+Y/gMH6YVxEmLT5Q
hAHN40Jdp6v0I/mNclqPav6HnMYRNTU2PIbfdmdDva2OfzqnuAys3bkUT0o9pPSJSlWsLfaVGD3x
aTYeEw8pZXmiihurVgoBB4yknsAgbpVDr5yiMJvbuBCg3E7tFkZ4K2gRGDtaHk1FehPDMD8UD3Of
kgJZ/R/YBiebc1/8K6l3B7qT31ml7GeGtrk+CS28jrBhpwUJSj8GOR/0RrTtKV/QnWgobpK7XEXU
AYhxMVNe4y5RKKgTpiLqECNQEvbOdQduXc8z7QVEyWpNEWqSOxCr6SfOHa+ySj+2tybye5//wmQ7
/fJ0QLP936mXvnp5vfPsuIc7RlMxg7EmtpcUo/sr9jlF6lQ55PXlUSA8cKuZeIxvTjkn4dutnxDs
40mv1lNhG/obe51AGow9CAdS5LDvEb6mUiAbmlhA1D72mxfPSQtgkUKyu5NY9V2ssi1Lnpm5Y73Z
5DS0GU02Rx5h4FGx6VZLYkmjdoZnXAFQum/djprx5CkrCX9Ws38DlgkczF3jXGg+nRiYxcBh8AH5
CPwkSuDvZf5NdKxdJIWsi2GY6F7eB5vBwrdxyvnYsR0EIOa5HxkYyqnpuDYX9xoYuO6199JIR+1S
FRXqLgEcWNA+ZPo6iz3xLFXjhqkN7ajyWnycFT/FQkJBosPSfoJaxIQ7LPbp4lHG8NtVqfX1E02+
IKcIqbwjtv8hD1ckeNw9Cy7ZPxqKX1LIYt6vP1UiXwCg/L/DXPs6nEm6d8rikX7CI2slzCES/44w
E3cLExvU1gpTgDyo86sJyoRsLacw2MVYLz89d8WDLcn1wcJBVHXZQ1SaFNmtHJ57xfXQ51+2GAYn
sCM0EPDuRZShnOTjW/pDMC/euFvYa8qS/xH9lh0L/W5B4yr8RYfa/u2Iou4keTaMFRnLJbHhNuoj
obgUHZJMV1GiSXRUAOVBTglBpDQQAQGUbfBFT3E1/7ttHx/UaLz5n1Na6S5AsGz0+0Kg9foFutQh
EUF4V+46xgCaYJSjtoOZFFUG/AH2lmWSGVTTyxuTaGkBxmKBAQewfDHHkjqj5fbIvDUxHy1OXSYM
sp+ZjeM6i+KN7q/Rud+uDGZg6Xq0LTmbpTE4ssxxauFq3jJB7A7TcT+Oy/b4SIRmeYlEpPHGE3G3
CxK4cuEffLePMfPmKvm1r4M4o0SvHHyZq02CmY8OUzH83wR6mHJqUoXUXEeYPcogJLip+pKJ0vVy
7AYn9U5DW7DnssxW5Dk0RIrOeXj/Ft9dn6N0CQPGFfenUo64uIlkXnPGOLozVJSZQbE7+n3Jmza9
YvXZvGiSQGgPTdlS6m1e7rNTX3gL7V6sbq4r5I9InhHeiVJrALqI8YzE9edrJ/wbT0Kv4GVdYRDa
n6hZFvVXQpyPsB6AuPM7C7m3fID7YgzQivo9r7wAq45+Ss5EVKE1QLccs0gzUa9GbqRJ6WGp+KcP
AwsiO0Nt5VmPi9CAe6fPdQ39VRjivIXLHdHhyx7fuSNbxbX2Dm4xQ5N4y2tj0tq8DidMBMKio3so
kJd8KlNSg/3HdqGrLIl9dZQsXH+yHwPCHeITvvW3Qds7lB5IIZ+5WdXFePd3WsZY0/Wl9MiB56Rm
Nf8gjo2kzs6lDW2NL27VvwVEwu1qliIv6vPrYMYjY89mbzeWqv9jnrU3sze/fBEMvfR/bbP/A51w
4j90eyV3kGQ8xiUzU9GnPgo/xTLzLhQC5gu5hsgoZX1l1EYS5aHjAiQ1DRPzya0J8Y4j/6zgbIb1
BhWpyQyDH1Woeuret7ih1eto/tqCj8ZEGv8e95AejoBWnnZIv1bE1G+R7873by1pbCydoen01Lit
WPJYwAbIcEZHa+gLmIADX3Wo9jtcpuJm7kNkHBWiRFh0VvuOd4ZKbuGkGEaUaNwmNi4oRpyBnf+r
pqNkvekCF6RNpnBz1i33JOgyNahwcrATsRkdO7GIs4CAvMQsFUANtIjkHY9Tc3mP7FrCrbsIAT5a
bwcvlwrPwMcPUaBjJfMQN/vA0LObpD2QnPCyaiTeojhYtm0Jlxa1SdlAu5tQ8jKQA98ogn4Nbajo
T96IP+AwTp4TC47WXoBbLo86SAY1W0Ri7erCcOSWIdxVteQEQ5X+QR5FcgJ0tDLfkAsrjO+8z7Ql
3E9wo+gsYuVLdcNLODxcNLQzt94HAuXqzSTGfFPGvobrkGId+XYSfRu/ZOSNrYvTA9mXJMotCdvd
l3P8jjaLBLKMOtsPYpF3lI/uXh82fFOgUI1yjWCePk7xHyd9lyMPAVaUdTrHZ2v2RXXPOCE0LnxV
d/tJShgFlclyo7N7QKNMBCruxyEtQPTM7xhoF4KgsZUappCQnwOW4dGOUM+xfENdoJEFeAnwBcn0
MuBrCeTqQbsrbjPmTIRC6ctOr9QVWBrh1kG4IsIKrvToMDcUPpP6tNQOKdHPAxJYxTjFzaUtD+iX
eKIJ6CdPXrPdp2UiIUGIVovNFOyhzqIogz+Dz1Jpb0RGkoNw9ooQQ1ZH1YxuaUXQDvEBdCaKzt8Z
jBtLCHayqIhLZsWsPKn12akfw/qW5wDh4S9wNRX72yi4modRS1kwsFp6RG5Md0X7VbidEUXLH52e
rzOGwPcuZmV4XauCAv5SzYR/l7i4OQcz2i8AxWDtDpF30Px2q3/8B5wxlOoOvjtTEj7kcrAslPCH
NTAEwrnInC5XcEu1eMfYdIe5AXApa61NvNRtYNiMjKP/UgUr9dJYoAkkj+V8HJS3lBRviTj4df6w
n63wVJEKDug8GyZwRtkrdpDrpdb0uj1KVrGb0Hs6/4cfAWzSgK7g1MLBwsA833jCw/jPn14ODDcn
TYH7pr3NPpOlrqMviG9GHalg3cB/E6y4g/r0NZd3ZiVVcY0p6mYExB74TcSKPg8s++f9nxKkJqLF
+NnSaPUYqnpuH/BnKo7gDtdjDdRyxH1yH/Nfm0xQEESedy6GK1OAiTHMY7QkqUNIzH8XfkEHBnhz
CFu35hHdMaPpvgIZBaUvBlu3t1U6zCxjHaO0nCz/sKNI9UPeLcAD+SObtdxPelOODq4Pp9w1Rf17
Yjbj7m0Cm91TVP402BT1IOuNmsWAXdh8baYDF0lQmf/ApOjbsJz1LTg4eEaFAus5PoeMJ0HVs51d
O0RGv2PlWuu4HNGKmJ/1nylVAgHTzuzl5SkYk6YZttjyH6GyVmFr3LHwHk4i/rQkIDwZG20PC8J4
v/0A/d/4J6gAXz/UOdwUkSztYcuy6ZhNq5jO+TaFsvJ60onKabtEeB1m8irlr+bDlX3X+T5PWM/c
emQDFnULDV20gEQmQdcrUA/hIZNQARKHWvWFR8Ne1MuElsCxj1NS0zuh1hDIZsWZy+amgGTxNDVE
2waiSliw7z5JoJgZmcPILeGV2EHl9HEj4yGD5TiwPaGSp4C4pqEIXKIrt6e/nwLg/ki7EwWo/bG0
2R2S8IkTmEKoXMpIsB8aIxIZEtZCr7Yjxnxka9W602vsnXNVjhIjTIFTHMusol2WthFNUb+WN48L
3L0HXcYG9z1PUwrwdXFoirf+vOmvfOADv2TaRz/PPQINqKqLOMK4Nn4lEInMAyhAhMVg4D8b5rMi
8xjYkk6EeJXHXGHW41H01DDDw+w6CKZtcsSAzi0/qDUYHhFOJjsKvHTT/dB5AtCDDvUDDBJolXSv
5AxtMNqLWwdeI2aDb9wqzAJ5vZ3d/9zg9tueKFPwMY5XP1aB6xr34VrLFEycZNW1RcyhZCkmE884
OgeMEzCSIvppu//g1kHA1xi0LuF0y1k2HNNa7HjgKe2ynsQtfQGfomTHtVkygkBB4jeODMu8y/oi
LpB8mi2P4hC9NE47B5iJZh3S4DOgPJJoIYld+jRfZc/trp/HjErhktlX7amuu/jq6mD5DQrcuDNy
CsxzbrocBsZwm70yLWFvO1od0W6Jr2XI59m4zQVTQAUwGv+ixPSpAwY9Yad5ivw5RtYfKI5HZFJi
b90JKRQltqVyCq/px3GOBMIf4I4Q8jhxMTr4/Z9Alwo02yqLSkA6Bkz8JkwP7gk5h9eDaIh/oweX
tcOygKZ2i7bsbalCaEUlCc5rfhLylu8jf0ExBBLqyHmpUlEcE8aXVbnj3CFoxE+8HU/HhAQq/ncz
keD8hXQGEJNNi5C+1yvoOfImRTwIiYTfKaH0Bieg+13NZf/utSCGt6eZvPpGBme2WBLf+dAzB04v
4QCpN2u1AAfGkJBbxdJj1DHdlGUV+6GUMNFmU38oLcAgVvYXrzeT3XuQfie4EJCrrw+dE1K3JBCC
VwZS7mQcUzk+DYmminWF/sm0zKJenyEMvNhta8lAyAIhNuQ28dq8SPDQ16RYSb0g0VhDzlmJ9qIE
K2qWzqMRxG2+vGH33s876KNc1lX0ukzqpu1yZkI/Ngd7bLCw+gmTCv1IJDyfgZKjfibHmHZRtGn/
B8knAKiZK/PwbZ4QOpfujeNT0XB1Yu6RAYJc4IrBwCZ5eK6Ol2VCxQq3PnU+3ATMyxaklelu4IPC
5U3xS0KJJ7Bgc+fME1F2rwPcmJnMyhEQtQwANWYQ45yiC2BoxOoNghGkzt6HnJEXuykxfVhmvX8U
Pe80ODvlXZNHy84hDKmRT+yujXdqQDrsOUUMhutEjFWVFUlOlHqhhYHbZehzHmCHiYVQ+dytH3NY
b7ODZdrEkwG4rWed/qDfqbwvzgSdBzP0weOY6EY19WqN2V6m0h9Qwml5BdI8OCM/3xVmwRCBPj2h
fJbbJgTF6VF2oE7aCTfWjl+4O62ZAEvMET7PsA3pEkDBC4qwDirVCuZ9FDYTObXOWV20eBkXK7MH
kJO5vb+1xEwZb49sJ6+bASmNUJWE43Q9OKQ7GThLGjhoPlhekULxB6CmAIl6sk6a2Q3oK7VPROND
rWH65a1/g7GKE+GV+6RWy2uUmFe2EyitTXC3iVQQqp+HC9t3TmntNhEU5UQZ55KE135W4odPTwCb
nj493MVvO2o8Tbk35aR7b+aUdGfLONx76mIM3chyD0fTSEDvMyvqkFrUuLQdm/rQ9aCNOvI5aF+D
hTKmIFzrH/fA9h7iRXKZB94okciNC9QzRd+oUn/ACXbPgMmMcEY9PTlWpLhgrDJSiI/ECpJR+BVD
6Q7fqmggGDmG1K+Kum+V2RWDNYzszSVlfxeYWsAnHqPfGlimBJWOI/mPeVQDZvAsR/Ia213m5m+r
fF0mKUSiCRqefhmzkGj6v3PXQRpHASPvc5e3ITw9xiZB+Pt3BWPJaw83t5CDaZq6GMj8CnIQ1Tcd
vGHRsfbYvNZm+aleQhecRD3KVGyPKGmkbY1xocaVUPEUonRa2M9NP4RC4vx4miEeP64vqLnvbr2u
ElcThaSILifoaKfDrIS6rGBSCC0RiOvthtZU2dAYPYpJe0pBm6pFOGqhtyjmlEoPKtdcXnzWdy1s
ue4A7UcC3gE1l7B0j2twgHgHQRrbsrE/+b7RtgX8PgxTpxK6G4oTA3IH97uI9ZKX9o+GGMGUn9y4
U/fhg8qnhM7SwQ40lq8xVN/z75Kf39EhCvOGvTLkFonGLRQO0KrVzoC0Vd27qSdUl5a8vqBSPuuT
wPvk2I6h3xEbQSONuRgX9kKLWC10oTs8mgNXwoy9hRmHuwG17NVqHQSLHlwg2M/vi3yuHxny4smm
sjFy6PHG3UhCpOYdDyK6HZs1nKCavxrYTbbV5rWFmSsW1bCL51g3d3XsP8/tm+Ks3CF8Iy/xhZZP
QImEsQlpXauleij6VfZDfRuRSEyc3cxn6/iH96y3lGNAjxoNyAY7polg6ZwwQ2L1FgEwGqdltZgZ
K8xPzaX9WG0LqIXYgeLkXWU/D2csFYdv2w4MdQqGqzxggY3vUaW+v8MYT1GZZh5L+aiZHuhNUUCH
XhirvfYdkvarTVPiZSgbsYQVjBD/0Y1G+HSG0chwCw7zQP5NK+tk0ROXcApF5isgvb6lk9AEkqUT
WxICpNB5TaHKa/mwa7axenKilhpK4ANxWvLpTH47lKkLuqL9E1oZQS/tok4rxGAKjYzbG7W3cILm
B93tfbJI3Lrm8O9xbz2FjHTE4dUVAD2QYLrJK16rzdVuuNAtTm7QJVFtA1h+Tof1RW/noRYBa5iS
NBCtNGmLtv4dpvTOjuH+pyu5WQYCSnw6eqsV0NiODGSlZAvNR6fqt3qPimJPAm6YFsLSSzPvn40g
vTWO2EGBcfdt6EacHpBkAuH6T5f8IJFC8Zo5H+vwOJ6KpRrecSx2k/Li4FxhGprp16X6smklJxcN
hyE8h903KBAhyL3Cy0PuC847ZUKw/FQ3hMqQNCysyCkwsMtLuIErbmTJ7lB3RccfqulPhzbPpHyl
DusTjBUfqOdV8GoC5JZqA84alsllMjzGaB/Dt4C8vu5mkC7NgO+RX8YeME5hsy7+edofm/xjL1oL
0LXXH/NSi3YlUgB5xXNz4sqE+LESLg36NbKNehuAJIsrnfyC9sWL92g5H+gwLaaOt1s5HWAhA0tz
wGyTBuDHVsD22vLzXI92TfWwsFO0M5ZHuG5K9yjwJ7GzZRhb/km04esGOBFKRLqz6RYm5/FYxjh+
kBkWKd9wf65pBI3ZSfioBDPr/6IdjYvnbjroZO8Fuzyqmm1yA58UjgoYfKnuA1Fs/kuS/LW9OxOS
cYVXJ/U5u32ZmUc4dXvwnMwXh/xq+A8KyldHPS145Ug32sM/nxZVk1EmP7gXzI7kPztvQS63ESJq
uyDkA5cPQ8uzYXoC9sdHQEs3Ep+IG7UcxBacgYtduUMgvmwMCGODwkLjuldsxhHZyB2Kr/9oR3XM
GgvQhLN8Jkk5CgK/zbIVIRI6w1PIQqW7+T61LpUqQdZdabC4JH85bvYBbUfCvdLVAhbNwHDMIbmz
cIad5/fPOUilkRx0o+z0cvOKBkhFupogmOmzPW5dDWh58OkrT/P+WfRzHY8IWUHsapqKzJ34UhZ5
ewfOnJ8ORzcCtcmmln19j7OWktlURSKs5YIjdF8eSi9o4Vn7RKz5AvHLyQ3ZGZa4XcVJywy5yge/
WCCP2iBNnaSYlEYsxC+Mq9HsppsmSWPJffb/SmFNjt0hxPyNYT8lFbgnaefsnrM+CFZhE2eCaiVk
GxrzXtyvjHZuDYDsO08JU4x8DTIyNFm5NGlMMAVJU/ir4ICNehAp433gWI7u12of/M/z0Z5W6zde
rPlqRJJwW6qmtJtyzEa0oJfnzA5kdrxTt7Ti3OY16RohX7/SkdZ6E04aaFn675PrTDwj/L7cl6mk
3gmGUzokKM4RAoSqyTBIOaw4g3BqtxVeopGH6DarvegXqyWnk5KuuR5dDpBb0kFZRzOSLr9aFHbi
zG6HRFZzHczBlysR0xtrWjcZy+tR8PCBFS5PbFtXS1PJu06c2vzx0pFi+n7H6GYnFoqBD4gfF8Va
58x3cNASJtjVahm34vLcpPAoUigLOsjDR7uIS9B6B6LW02I8DNfysJKyZVZl90M1eLUPMyKzOvJ7
+jqrtGRUawvjvBvDb1dtKfEHKrqlzUwt/4749ZfBasr3IW1jDg/DQ8ISQFa5dygWghvLNyybXeXy
+2nAqM09B3T0iqPrU3Ruy/0XWIppzbHc87g2XHnZJJWwwScF3oagoAMARSns6yBXJp4rVlK5bUBD
rUGR9PiW0/oI9AZQIdHlgzrq3cqAb6CIx2uKlx4kQvTswuFLDdRMwrtlWxtwFTn5eUiwzZNWDm2q
deyEaP38BDoWG5pOdwTfVKeZuAKx2eq8OVLD97VQO8pTJQD6f2v67rytG0afUlCyKAhDCPNyKcbr
ojpZ6u7RZYvP73nPcABk6PyJTfl6U0jmAqmfJud52aYUKSHL+KzVqTZuzT2XXvjEQsyI/QKmVtXD
O54shHtLIgApmRgAy31JvTcx9kq7I8We4N8aujLaJ3rD5cYsLleat1z1Tg5MB4BM0n5x482a4Cs3
TI6IXKMRVnz+IVQF/J6jT0G7V4cSg9vzTjWc92KC2BlTHLD5S5blHQmC5oGxqgszB4unehKCBwun
cmhbSBgyPNQwBr5ajr6/1PfD0boCqzYvazH/V8t3HcguXpgo2qs5jbcoLU57IKi7XUDrzzJBBdAI
VwpEcHR0QI8U7l2reVKOZD2LKKrYStbH2ar9SJZzNNhY5r69kIeiHe9JJWamFAo8U7qFsHJrPQ0H
fqQG4fEHN3Lbalu4i5kA1AZD5QaFDcrhJ5LGJ1uvZKdP9bAcUQGa7+bgSjCpfVuRLeWG0h6FbaPX
YqxmgOCpW7RMByMZ8clhwKQnKibhsss7jQL08Vo4Cfr89NBks+dzt+uWBKVePEYL/0NUUZmeTNro
WWGiGn4XOUIXOFUOFckbYvMIaTa/AW3ZVBdfLG/GytMkxT3dW99yyfT/qnVRQ3u11aKja58zQITQ
mlREUkEeSWShR998M9nxTm9B5xWah3A/433t25sz/94UoDVsisi112NVij/soHmWVlNS8dfbm0v7
gde4oiOuc2yEUG7pYBDYm6fvRzFbWVif7PWrGGN1hEQv/qEUL76vZN4GciOZvCAaqEVHdvc1ySDJ
sdqqtpsHOvkeJ27aesyqNcZl7eEVTvgpxetiLxXnl9L6OwXz99Y7xovkLyJlt+CkgiMZhq45uHZZ
E4qtzjNlbTHUbkbS7iBRVGF+oQZPnSAo/mnjlyddDyVKLJl2j7vuK4F6k/9N9XtJqLptvU3wGpGO
yWbPB7v/upQ7KSgd04CmvSqarZL+O8jE4E6HZ2eovVO3HQQf9Ya2nkJe4OgBa0gbv/6hyJGlDNhM
Afa8GsWYtCB2lxndVh11aN17eblzJJRXL/aluDXR5k+prCjPrMOgOqOpZQ5t6cOOd+KSmPH4aGl+
i5G7/5/pAlG4vHHurgTS0oM+pmoqWDyiIkVYFHZ8T030eRMlICk0ESb5+LtlxDMgZs07KTqS7imA
KZsNxWgw1jH7kcIHa8z0gGQcd9HlODkFhlaTjE+FQynIjdjuyOKZdZElO+LKbQwfouSLsUsiFJkk
q3OZEbGtLRM29j5nImintRszN36G5BJrYk2VvzTywepQOekx3pbox7uUDNi5h/q+1B3SdmZliwie
MS6I2uQp3fC1Fm7e3CK4LAmp+wpTkhEx/ElmaWIsZR1LTATK2DlCDmw0z12hGbW72SILcBqBOAVO
fhkOSNFC/fHR+iLiySe4Bewgq06jnzxxs5kTKLg9avLiH0tQH5C0SDX//Wf0AwEUc8h4vsgYLU2I
xcU5Inl86DImd2F5dUXjLff/WFLo1xXzBFpMKCAtmA+vHySRViBKCkmhhrLHhr1JBHkjOF9qMKfl
QS8USGulPEhAebOIviNkjuItFPhqO31wGyemYeMaNqY40HAj72IpWvZd5zVAyW99mWuLBGnH/EYM
Y1QrYtaUOdnfI1PjzXpJ6jm4Y9cuMCqgPWqNFjuN1rKzg06TFigknOKn5laVrLHWUqnjg3nGR2sA
xBS46AbYN/NPDOjgzEHnmzEuHMruRHp9hLmK9nvixPsC8SqQD6SXpcdoGkGyp86kIPUkKDnkYw9z
BC4y+kj634Vdp0FIcGM12lMJSfsufcVA4yrsz22tkfLXsWsZpTpO2QCwXRa/PvRMOdWnrL5K44eF
RTybpF7lCEbs4auWn68u9GSbPY1iXmxe0QUZuOgVFXGw47cLzA2jyqs1dRbH7GdFTtjw3EvB2ecO
cVk2Rv/bKmLkAruEKWvR9u+76lfkmF2AJpqUkaYRyPzblQK8S3CqmDbmXBK9wJzW7PpLDjJwyE2U
/ghsI1yi+R5o62WbQkjMybzi3zYZUMGjPlS27y84vpq/daeyKaIMmgs6eB72UCxI6Y7ClXbFBhij
ofJU+vDKv8+LGitx9WJ4gr6DSFt4fxs71uLumBunZJJZccTPoyKUWqFpD7ZpSd3xSHUhTtZyc0ie
V5NEDR+FUWPSkEooAs4FyD+l5KSh5UTCZSGo4I9xXXIPLvt6d8c480gKWwO5FxSzyvIeyw5TxD08
MVO8W05BXtQjn2PfeTwlHHkF/iTxMQh4LnixikPr9J1wy9Dl3OlgvwM7XhYYK4rtbgJh2YgcggIl
ENU8gvh1uJf6w6MFDtxvtwME/ocs3idaKI2eIDq78e+V/l18lxiQMC0fLCLE+hOKkdtft44HW7JL
JpLt5GbpO0vCLekKtpVEB35xCcFNd9dJFvEAE9DKbojvgZPp6MYrZsVeh7YUP1/wxDNb7axS4yRG
hcI6X0bzQM81SFMMne8Z/nSPzi0XM38zLukFAUDlXvGWZP55MZHp8MMxlHQE28854E+5bAHkvw7u
ZYQINdJYhpfA6VU0EMax5Ml9x1xRbQF4hsj/d7jtLxF4jo7u/wGEWM+BBbHCe7D/6eFbIsKxYisK
f1WTLgXpQun6tjxwG5E8TUwQKou8DV/Afu81/gl+ERgWXkQmQkaJPsZkzWF9Ni3GlO/lLwK5w2iV
vMLCzMsZRpZE2TThkphPqgm20M1wtiWe+V0s5u0aqbp4f+VhJgXW5Vq8y9iFndsSIs/1WyI12Pek
+7vFkIWk4MY3gPgKado+MWVxcDC12qIg8A1Xtiif77e0dSCbgEuEAPj5TTyoftH9kBU+gqwvUqGO
7hcx536JLGfh1cEHI629acv/OBcQVXhU8n2FP8RVGncslCrR5Fc/dyAQWGijZbwuyQ6f0FtWEaSc
bECYHgyFUB2SpEuBg9xQPOUE5phkOnMSwO7wwO3qOhtaXDfgUh+wMLZF4q/Rm2bwFGIaz2zJT7cQ
6CXB0IPLNbm5kx9bNmcAtifJhIpbBUrpKfPM0I04GqDgZORYm/dEKOxA4J2VZb+liv5sF5L+6AH7
zrVeEBcaf8m88OTQn90gTdRsrrvyDo1s4HMlx5053pOqAlzDeHdMoz5Z+O2xWNs4ePkd1jqY+gfG
xlq4VwPpdt+1ETSfYA2RS0OqN1sAV9lXuFfus7/XIJQaaQ6BcfnRZJulz5dvHDdOC6mKAAWdNF2x
/E3hK9Q6Y8JAwq/YU026YCXaByD1bI2tLT9jtXUJgOfo0bdEcwHIIm1p2kgkj12LDY6LYunPV7PI
biVIaakQicfecM8+hgM8W8yopf9ZIYpCEyKEtMOpIvtYAiQ3JzOJgjmE2Pt2xddlku3CIvP1stHm
eS80Ic97aEhE+C+OVea6lKXuAgeTtd5F3LF2MOVOGuHpoh8d40dNxsQxGR3oJ7BtruR6Ctt5Dshc
h/IMqDM2cTkxlGrlShrfOzAYh4RoBTm2nnrIk6ib2ycncf4MNuax7vRiII0A+2Cn/VaE9evmcbar
Q5XwFXOUvosM3820koFsEoh8UzHPZLBVi0ApsRwHO581fU/V7Cej5Y8D2VENwZFNbr/pubnSSm0e
bl06N7/RwfE02eYJadCbt9QTO5zLMTqarnSbzXMknScqB3tOw/xwRllnp9AVi+uvv5D8EgvHYlaB
EueuJoHZpmu+dwSIQmoZ6xhcu29JqZCIwI11J9+bERhsqFzY/61XRnUWp+QnELNjmsogQ6kYVnzA
1l7+3JchC40T4j2Sc3OXz2U7miS1u4afLmugSuUgdVfYbHf3aJQOrZXiLIrb1591p49mYSbWQCWT
c+nDJAjSFKd9PummlfaRrIWBR0dSkhyKXwgwlMVUQEmyAxR6fNRx5BryRY95CLznBvPdSJxCbt/K
etLs4Z5QI1wLFXVj8jRVcrrqXohvNaA8xU9FZQa8JocuP9jiv30F3KWR8OiAKf3IRUJZU1y07a23
5bUWNEUhXv0xnrY/zZHEAxznYb0PoWj3DKGm00yOmcjHz3NioxP7tzg4vFulpXNj461PbFxCnkbe
gVDKG9Jf0v3XyFJpuDng56MXdZ7ZK+UxyNWvbZCVej3QZlDEgwwOrfUVY2ejO8483KNWRW/iYnES
gWFlzxsaXAPanKV+icW3ADyO5sQe2u60vPiQCGuOB5Fpig7Ig7Nsl91ylgToa4FM22Wz7fX/yeuj
N1DqJN/xvCLtRAC6Ei7N89wy0wxlDVcWXsKsFjmWKyyZgNoGaixHLRLktey7/LZy436OFkg0V8FO
nLZjMsd3TwFkE4PKuu3NfFNoJkPpigJDwXeibb50FgaNK4Ep0B38+HMxktU1kWQjTmSTb32tyZ1L
6takxKmd675uaJy6nYTHp1MXsz06nkN8BVbgseOjmKF6oss9emwKsxOATBPDYlJk9jDR1N/CsCbP
CarmS8trqIuHOdhqq/Y2ORa3VntboufhR+fBshCb9Gt4Z54yp89yBL1a3v16jhUgyOrzkRyhdHcP
wyMp7zjomjH8yEWXm1+GEYLX2ozkVDWmwBBpK6SoqolWRN90PPUqXzCJ5FPhJFiHLEra9RenUv7p
AMHVnYfPUmfsCOGbkA/hp2+PKZeYXRKwPBzWquj8Azp7Fj5OPg7FjIdZTB6HvzPjQ0PBf+5xyMLS
DuCmqs6tPTEw0jejHolNZ5eakECsFqpZVeLRJwo+IB2EI7U3fPVxxPY95cwk8iCQ6EC/CuMPOnvO
0rZLsDzZF59RV79poZfmRLHQ6otd8ajcLs6nC406rVHKafzJFr4vhGzYWBKz6QXI0Y43ft1xT8Qb
6/WURqKzImT3R38PLopPf9qxKa/zNVD3ek30GG2niE20r3StZx1d61PlnOvHoCWJgOSSoOWexztn
NNQADdeOSp/IDUazBnuyd8F/rP2UOhk8VDPjfWq3hyZYV58ouXTWaXB7e4JZNL9ppl+USct+BGxq
cbGtfT7Vdq6sHmXgRnFioTejv8ztec7nYIFEgitPMAcRNkBRtIJ2jjD39xgN1HnDyipRmanUB/jJ
btLnwqLBPJaqlWNb6E61Zr74D6u3mZzimE2EpTGJbhMG31lhiiVts4jvbVmSo7x9hRO7ctk3fn6S
Xb7hrvRsnTZ3iJ7r9rynNC3AcYtr9WGDhNdeSE0ung7NXBZF1gVQqQuYvJF4kMxjPGOM4CnGlyEF
0d/sUbYOdR+0ViMb2vaDjyOtz801EPrYLD+lYDt/JfLW+S9EtDkZ/dVQxCbnAPHy4FxACbZEDJTf
BHLGJDH1UuOIcmvOUhd2PUivXIIEBJHl8OAkcu20N5H8vr19WgPY2YkZWVU5ROe6UXaDV19HQ64n
ih+FlKHUyWBVqrBQVTSyXIviVaI782PqGZvx3Q2aJLUaEiod7v+98WL2LsRezIpjAVSpTiVlr3Ba
4UFfHHJ+VmN03umekpD8NLKQI1ZsIP6uE3+3ejQsQ1bA9TSl14LmUin4tJYMtBWvKtaDnNU2DPOe
7K3vsP79RtmDlBVc0X2DznFmdCsFfGBYd6tC5n+GX0O1k8cV2CbNnDITpVWJaUiM7q2mNwheVBAr
V0ur0A7XOOVXRWer0n7wwFa4BtqYbiT9AwxxM1UjLMyaqv9X19fPu52pGH1nSxQj+ttfAum0bAwF
ltG5ZkYyQT49Y47ZSBy9SVL+nl/ufKIhlCa0PMHH2XGLCgSzfGaaaLuAiN7qiisnG83FBrz2C228
NGqNaCEp2GoDUnkE4TgNsM3aGCKFQ7r2RfOQEuLLvI+bVwsajDHW8hcFHFhsTEfyXe4ZcldaUfsu
u2NY+7PW1hM4yXwLCFgffvwWP5kAA3oM2uz4JDiPgA4zjgoSwDDqyc41PXVwRrJQrJSje2YTmORI
E6SjtSLLfFEgIY7dr/IHEV7LyNnYN0n/H/rIV9ksQefazSBRO459oLFzu/GotUrt+Mr8NJm6TKbd
T4aLM3a2VnfxubpWuzLc368puGCTeOZ964Y8DUjnzQEUdJJHLeGKKgFhSkx/FO2gywenAavzKVav
76zYXaivw/F8CwR0I25y2YVe3dph+SAs8HO/RfZx6NNqkWc8FJ4PTrEJs9x46F+hrmD8BR9fNORg
ZXXZVkP37lpJZ95gv4YshNBGutzlf8cYWwgGytAl2bBuLM2TjGkeDep5e3mshEe43iWG3SlC1Pzs
mPueNG8m7baQ/ll/SZWHv7GQ7Ml3X8FdeabQtZl9Wn3PoredfHh55QH/BGvKhtX07Ki4fE/JeAVv
/X4OwuUp/bBAd+0TpUZeCyw4SJAuoKR8I9zeyff89rR4dM6b3f/IudtcqkNfBQrD2paUSn9q3YmR
qNFKNlGcdM3+7LcfuNZeZkOJAXDrwmJl4yRJaVdP3Ye/KlM6yAlpDkbiePAPMVoYEf9WaN66sf/R
wb3S0Qsw4ViZ8n/w8ge/J3kGj7GHFltu67Cy+CpPp74EEVuu3hDS24h1Fws917uZeQstGfor/O4p
RQX7cSemDNi/T7HEu6uP7jfhJ8T79XCSHzq0CX5uNR8Uav0dgNtWFhsnJMbr3pZiTf4httZSW2po
sTqIGQne6Vq1vqH4j3wx50BHMklPbiY217j9EWOYU7h5kHLvaD7l7cCruW/m3oGmlFN8Xk1MJSuh
2hxTcmeWHFoIJ01mn5Ai1sAWd+J3p1W5ntIVcuwKNbSrfGkP13bphyvzmyy6z6Xeoh581bIiqs/Y
QWgz6G++wah30JMegkFPLu/qVx+08I3pOSb4vRlsI998RhHajBLUTvnKssNTtuDQqtfvvZw15tut
L9NJH1V8TLQGwinley5/sOLPhBaeSC5VXaniGORoGTdT+ETFiUPNjEoKMjDIK4o41KYgXTukyXcz
s/LkfmQI2tD4h1uuVjCQkTbtdmKjUIPiXdObvAV4kA0CeuIOfdpDPNfVDl9kkjqYUgrzEhChboHQ
GjE5npnA6yW8bLZbguqGmD6cFaM9yxwmtQbJI19bIBCeNoEsAHXJfNDGaVVV7mYlUmf3m8Nk6QOk
GftqGt/F3viC19Pegfa02jJ5u8T/rTWtv1pdgX//NtDmW6RojIbF6Jgs3wEzgztvFVDRtKSQA65a
k1Dv+2Ml7HF8kT4SRo/guyU2Yt5fB3qtjuCrmtvFVYgoD32b/LI+oCePZuSz3CBGB8EMLAb6KUND
/310y5H0+3p8iBBKybOYd27Q8SA1Cch+LjgRsiSuw8mD0m5VZ51LsILo/rTwvwrv0WNzRRkTjeLS
EWQzk/QcC3apA3KSQH4Mrj+8PJ6q8MHnQM8urpUYvyR8HMxM9XMOb6ayKRhCDZ0i9uvwCXBCdTat
1GAFEL4hU8hKiuknLQuDyNIzOEDgKyzyd1OJif1aFiXBddWdKcEsigAgF8uef32er8UPW+OE1l6n
NEoTaBsVYsROoVTqnz0CgYqxMfRzcqeGyum023bzgQ/4exNmfCJZVSl9LUsbpW33K/EuNWsN7/+4
Ojk3ZEhp1gvKyg1+ZYMZwRr/vMfMczqJ6A7aQ746s3im+DKa13L/KSHJynEzGZqZJU+QFJpSUHRL
oGLP/qiKdwpEo6ifwz5ElP2ibRegDfZ9zGnN947kVZL/upEOwApRWa9JWD3mZvXJ7HIjsDCzQ2dz
9tJnBoWimMl9eRo2YfjzPGRTwjYJhd/AN4paVmtU6pNO96kvKPmKG4Qm2F//tKGYPeT3XbnWxSR5
Cw1M40ToZTPCKeG1+cImQVwhuLFb9RU6ZwjPI/VIFTra2+1HeTxXQhu3EYsq2sA09NcDdkkvucCj
LiakXtRnDLSHbh3aU4W4Sni8o7GHMskt0DENi4MChfXX4z/WG+SI88nHfhBaUiuVD6wUwX//cK6G
uzSmTrFpXbBd7x4RDH4RT97DH5auwjA+1m8UQI2n5Byj3BSWyVangN19FX8dKCGtXVoHvH5h8Ogt
ZAL7XV1R/llncT9d86U134i5q9pOFIVGRgpCAJfTjtHhUicrmnZXgbYTEqId/NCxtqMeJ2OtSE7l
q8I2clm2AguR+/dlhprhLbueeeS5Z/9sMkzfKuhsTthlPoYy4npGebmqMvgK9ojfWIjduA5tsiGW
mCIjP+pBUjlmfcdZaCN7ezAHwfuHSjO6QuGG1v8iCzglqogC3EaV627gFSwtfs1MEdtNVrEyTYCw
bIIhX0SD0Cdi74fbHUJ+UbUddiJcMIA76UivzD3W6lRvWLNVUSgVkDPFwoOalb26ZKguyVvHtQ5o
mcZiUF88AAv1FlTN70p9sUL9RpAr2GHC0StrGZaWQLAnX+y1OLk96jHNAWGj1Bvp98510pYlH5wt
qWdfmzljvp5/hnEjKKJA5FkWjCuawxClITOXNIguAIYl4hb3j78hdzZMdIqF4klWioqauzMel5zN
TAqVYBY9Vbrfy/3+oCbMz039EwbW0iD6zf55tkuBxVnQMTq6+0qbgfkaQ+XLBBDGMf/zWe0RjrtL
UOe6CYFMuk11Yg5h2klGI0TbK+84sjepuUJCfr2pt3F0TjKfuw2GF6hJf/2K0BjPObFP2IgN6DS3
+2TnIFiVeuHKaAJnyx5Heu/kuuOiM613//xvUifPM5ix35ULeuIotHdmBHVYiB4ltBIVYLW4HmGD
XveiGUnLRBy+Jr/UahElnvy4lUa8ijcRO+fa9/nhuWWomEQt03/wICT0khAHgeVSZ+ttqgfi0aJF
3P3VAvUw7Jg+e7Z2DOisFOToGZFrROyZ0M2YHw1hTgZsYglztPe57F5ddNz8tRlPvxPDI9wpqawZ
t3DHvgdMhEGOER6otGBBa6SY4dttSouKQJ1QXN7HWvwB7xtrxh/u0sRrqEc+Uy6wlaD1Xc1qxTDZ
mUtbIP01L313CV5hVjNNJjn9swxakhd/JRIYliwhyI2wASc4A2fFl7uxhUeXofmLAB8Z/FdBayHY
eNfyPhWodR/zVceR7ArApPQiHXG+WUIt+NPUdoPcARTkRvCNRfYekyr8SRfqYVUo7ndu9lQU6otI
EQ9qhG4qLGhmvY0BFHcef1GwYE+prK7iEmbx7EGDZMAVIH39h3yTn04wKpHqBWnxtCpoyiZFlxFq
zluZqvgJhnTmeYdsOXnvMSqZczM67pmQtm0NswLQ1GamvnKKaqYPVqQ5VtltQv+AVP+KW9d4A2EQ
lENvFnr7M+F93iGE2rB81YXBj4jeDGVi4Bdn5U4/r6SLF7IhHukJpI4BF/QMfNZ19HDMm4hqTOZL
ewV1o4tgW/PziJ5SFcQbUq4TKECTfoFgxfL5rlWXV2SI8T+ANGcb/xA5Dljcxqy1bflKnsV9lz6J
KvyhVU4sq0/6JGqoog1H0AKRvsfmD0dpzMlYRtq7EZjsSV9yGEk44WKpe+dZS6CEASN+5Wlwk735
3B2g+68+pqixKv1bnNIAFV8kvTylgHX+Rz8vREm81N5sQymOPpcmqo4R5nbe+k9vZXZIpU/vErgP
hkgmXszIMUuK177VCM3W5M+9uXW/i1srAXAQiyxy8lXYdSgsf6yJrum2gZzl/gQA2ZG5QmtAMslA
kT84ZUcITa/MaJYZYOFox462IV280n8CSS2q6cbcx564e64Kc7MU+uKM9c7K+0EGFP0NEJCZzQPT
T3tMXJdJvFD/PFS6nHpTvsSq2nM1e/Dd2ExCW2xOEoX3gopCq8/SJifYDrIaqM4Kc+m83Ga6xCo3
dvQnjRCnk4YY36sTWpc6Nx8WHbxf6CIZcIEQemD4r1QCeda3upiIk0r8Ss9zQfjrUxBaR6hZvDWz
WmdI3rUlJuACvf+0s/ExtaZ899wHY6iA49k1VEqX6M7CY1Rz7+EoDVA7HRhWXqOjIA0n3XkJ+53R
YeOhJ6BbVhGRn9XStNPbyY40U/J5vVmMsuFkEKL/XWQGFPFMJnE79+15juU1aIw+vzBxXDnW9VcT
eM2ff/Io3oDsPuZp4unNMk+qNJgn8sIyGvfCSd+ESk11uzdIzMUEC6Suh7G9IFGakQeZXiT+NP/8
q8ZBwfpWJ7nvxS/H3o5zXlDQ0W1hNx9cuVRTjv462/PrI5kiBkNXYAwUVY5oErkFWhcEXSYsjXHm
rbyomwFiL5wrx4d5/V13LTCF/b8+LTZsM2jCGFzfeGfSBTGXT9SB1yJSAX5GxPmwKTvlEWWaHPNe
2XYIRuwp38ZRDfCwixJa5WCeVj+hbO4Eu7pb/c+k1nKEu2lsLOdiYGJ/sg9TKdp07GzUNWJzbzm/
f+molRNKR66cB8pCjZb4wFM4IYjjA3NIjEFg3VY/4yRYEPXPT9WyhmuMrGqxunIfhZRU5zmEliEM
QCCf3KXc0T7iHx6fv1eA7tl7puVdjBdowh271qdHh1Enz97Vf5vP47AiokfM9Z/2ztr8G95tNB2l
qt0Q9a0sif1UZHpvlBer8tixr9Ny2eDXTBnXWgjiCbWIRjYemrg9A5l+7ZCTEDv2W8RSRUuPIr8v
8Ibrp0IUEqjcUnqcqu0oPtAzVXLdvSyycAjfa/3eMlt2SgSsU2Q7HVIG/zjwR00BVvTX/xdmtuRH
eh7iRoRyGg/Fh6aytrBeqpqbdyU7QPaoSeEMFeRZ7hJDaRY16+EEIWnofRn7sNOuwb+eDaPQuWVS
pJuPc5ILpjRTYjg0gv72u3ZMwUveTid5rj36LwvhBoVDbRc6FHjKvcQ/Unw1+3qq5z0d9XmgVMq5
FIObcxzj9DICfYWGjrQsJj9n+9L2BGp809nyfQ0zNi/fHVXlA2fstikLouHl1o9vBC7NSb2t/tX+
Jo4IPUysNAfjnJo72FIhFj854OGXHWIzz3OC+IwIte4vdkzUceJxXAtK6tNw6gqLsFY+675kQ5VY
kEmH/ZNdT4iHAkXOSHEDsr0XaTwpv9sYikz/uo2BV/S+xDUFMlwzbuYZXPsbz4zKEVC4sCHX2KMa
aGt06ScrN4vidUl/318Vvrs5MoUr9EllL52IP3PAn7c/qszuHY21ZGwxiZqONOM8FDqLL2M0bOEO
BJifmHT43jIgkbel0FYsE5/HcsbWprOoYI50nvnumAPMUwgFC1VcEjdMz3TIoCMX+SDsP7Gzd0+O
flfZXQiGTXgKnWinNppsP5YQebqshA/63/o/HO/62pD/Bue2dtIQaqF2BKGjvk1EiLj6M3ITOKoh
oMsi0IFrs6WR408uiPuT2N/MuMd/BMmpGe0dKGOCxl+laz1lQv8IXs8lNIAhVRYfWS3Ys6G0iPGn
ujIVNqMBS8PZl0M+qjRCnYYUbaB24vFrjPf20qTDXtz3sCxctZytOZLnbj/OIbkpsxzk+of3coNP
/4msfiqs2O3I4N/LPJzkNFBf6L9KdoDiks17myEoUJEr51bZE+UpoGEIzTn4ap4y+H+VRnwdaDP6
xoVFv/EZxcBgiHAG8NZYnZ2p76BCAqSBO0L9tA42dqBzVaISqb2oDFsBy1IDSQO5j9DUBodS1iy7
FQJXTVDDpdP2Xu8OgDn+eXgYmfAYFkL1tPE3v69qZjCJKMhzsczBkdxpXQBN3TjrWG9HxV/MjbKm
bLv6y7Oy9DZrXAlNZ7/B/xztpV+bqnhCSzdbam9Anpa62k5g8TEvwEC8itHXuypnOl8qxIyDGwPk
MPaIXZjorFkj8Th8AQTv5wHe5PsrgwPi4rcnKQLTWAMOJ27ac4FTZuJx4m+H7QmxwdZNnQMAMf4Q
qesWxyTKqg+8cSB+8n3qlts8GpgznS0LGiBZVDPyT4czhLC36M9liLNPL17h/KCWjezbwv1GXGC1
yoA5RblrQkPFm3ar9V8whrUA9jsgcxkYiZSlT9f3AAm1hBhRhwvufFpbAs7UaPvztqZLMs4/qSdo
hC+Dcb/jbitHRjPvhHvP7HbY4+ynO7v060vdhsbh9kifAOXpdAkC0jwDZuRcBtvOnkp5ezYOCDP+
ZKZ2cGQSQBnYThzmmZkb6dwHHDLQpj69tE0gIAALsNxkkJmWHrYZIr08JIcyIjLbB9IyOIWth6El
mPA88T4BPJxqC8Sr9usyiijlwIjzL/6R1jg5gnJjcnx2kk2QuNdmYgxOQCeKySPsmU5SoIs+jsLb
LTOrQk/K2gRLqUJQEGRM7Pp42ziGxbLruwdnA1Dt4Lhtj0fUDD07SdGg4EnYUHEVMZ8XghJBNcPA
TisaiuL671ZrJHTKHwRYWDyfnfqdtosNS/5QsPTxSNMAYxply5UrRqAdDGslHfAYrht7tbGhLEDB
8gmyuwc6WTkD+oE4/7wajUKf+NfHSCalB9BVuLeO2ySrU2oIYgeXPrSWYZqBDZ33mEmOaZQ/WaGn
njmienBPfJRIljo6LUuxpmP7MTjbIM7FG4dECsrrsYl0+0aBXh0C7e7KRygES8HQ1pis3JuqV6cy
OlYLu6QOYQiWDdipxuMD59YmQ/f2oAO7bTfSZFRZK32NTVb5TVRWGIQ2v341Fhl2Mh0RHaKUC9Ev
tUR0lrxxt2Zt59394+PItKolKFxq5/Fs10AooFaZJSMESt2pGN5eHDPmwshUjkLpZOLHI/8qTIzh
4B/2G9zmyvLdJ6IT3BkjV6bLCX2XUuX7Kv6+3WoQR90rsol6jlOygfVRiMo/XS4wQXsXTmtdYy9+
V2IK7puUEXfcVfcStqRET+Jb1aHmyOyMXmkmoeMZnXfgCF1YXZo84pQFeI/QkVCseI3HN/Np+qlg
XpHsByVXJUBpSa+QdcJGIMjT2Zmo1o9VW7GN0pcEUnzUqg5wcsFX3g37hXF/ekKhoIHzV3qbyPsS
1zYbMW7nlTxc5GymWxr2Lcf3ZjJMBx9YLelBMwSgH+s80tJ2HIVE/oMlojHYhRSK6lAQAJ3sqsXL
5EqbJQ5QBkvcaeRjLD8GcBWrQco2qR7I+0T7L0orc35VnppSOgYC0xsrTxrb/9ADqJaZXZBdb9m3
k6Z1JCbksxv1BtUN9HML7Ty4P0X7otx0XYb8uH6rakmZPGnMA0BzoslQbwNAFQqh8jugeKTBLMNN
PyKNXV2dW59Jb464gb+AauESZAVR9F1pkjb2zbMO/iDNjcGnwKy/NWLnrXkyfyh7LN05eGlO0EO4
Oc93NkMDNG9a143loJsL1bSAhDmQDJhOyEpUKQHOkGs28M69jwbVUKDF4Bq6HLAaZMaSdtFfOx0s
O6Eek5pDNy/VApQ/T3TDwn9pyxvNdpsX1BmXfSI+cTFU/LpTp/2xUYv6TlSN4liK4ZhUuaAhLvX4
XEY9OkNF6ElaPIKdMHsoiuPOE1QvPaM/rtVrT05elkIc0kegc5hty7sznDyftGDSpwPnVv2Ry4MI
+N4pq4LRC88p5Ty0LhRnNe0OhX2tVrkqd8IxWRaTusOJoigZKZ3ceBrrXG4KH50gamF2fEOVlpRk
viFSu5mEJjVqmMf4tLVTlIm9ua6hukfVqGA6hqcBrN5Xuaw9OsDwq+kqYdfe7OGGKW1g60IIgnnV
8ONuKv+XySUJJOVXm528ScNosvIg9udKFe9EFhj9HmL6cX8xRT3Gm8onoDT6cGk2WmWTiFLDNd3Y
La9T9Xn1aoYn2l0qwVPxrX0UqVLWolAFO40Vy3Y5mXuOKOyia/3npirR+WtBhXvqCpI9kLDK/U9Q
LaAmXuEyXgMpkHyqr4Za5q19sziaqOrDiJkVsHjSvMEKPseeNb+1C9s1QAij1DMAgxnnlvHTC2ly
HXFn/ydn+oBC+3NDwvSTsNIh47cCfhGSMd1ygLy7UqolEnP6zbfWQaV39ZKSdoL92QoDR5ZI35sO
xcufnZi+k60ApA04WLJlVlyz9jiKH1tKkVYh/RsOjQpFbmyB3e/HgVEXen70BBPC9N+XsBUdFe6J
gMNz2YoMk9nhZGbFGto82KyLrLzCoCIawEcs4kQXFwbUfTNr45hgmOxtr+rUXllQArk53NlPHjRJ
y5A8dSGPxc6UDnF6nMbovaqkqmPOyIMClAQ/ITDpVPU0cltjBGilgzR32EFXi7lxjuxMleNQe116
LJdX7iT1jCXibwcRe/pVMHjKV+3gmdaS7O+XA1uEU2tiXhgh6YqeOUik7RMEoW1UunjFncrGEIKH
nsrjcDVis/ymS34ZHmeyMDOPL/PWh50IuroDdcL9l2+jEHfVNRXJWAeJsGZt2UsErvN1UtlZvZBR
d/ya2nlybFM69Q9FE7pzJGJ1NQll3QUcUB7hJ55t3xh2GeBoVwK3aK9iLKGDsT++oJ9WaECkpjhj
Fz/1kSiYW53c0cJf/ARzp9vN6TyNhGDYbvVt6wNCAVsfIogbJTE+7w3U/Jqq0BxbReulPsfQlhA1
ZBud8TiFNknldKdEY+bibMnznq9S/4A3H+wk3mFytKWBXVYbHRxjjNbVhNkJM16g3P/m2pWiTV8U
T9uaX3FVvTMOpWSECWLj5F//nSWYRcmv+bnU/tTO4wBOMvIxNjwBy9VHTPYOGHu4NJDbNZxc6E4p
TyM64DqA+WskOPSm3/Nl7WJrcUYdFUzCaK1DyeQfkTSuz7QOs0ImtaaFOxum9gu5FoneGcSXnCzo
7JI66UFeMwvRavWeU8eXUN1snLbO4Q/4USGbIjRP7HoTNkweHZG9OMtAm/0uJIpLeCl847Qr2nVb
orDQD3WrDtdgnlZaVPeTo3h3oIasPpFDhw3kX+OJfgZBMQTRWJy0DiNB/jENrM3PObZ5XXpMvlmv
MOKoriaNooa0jt8C7XZGDsYJRAOofQBk8PzIWgIgrf3PV53udRYAxhZv9u7Md1vNsqKWGflH+dMd
4z6DHKdFbT+Ksna3D3CYn4kinofwoVSFytaNQFgTJDKAlKBQ8E6xNqRUXFk1VNxBvNdhJKeyrL8p
gPHJSChcE5RjKtsD2/ttHa9XDXAR8Mv/943BDgpJn6DCoMnnwVCrro0bIfd9rdMwfesMY4PXzpMH
rqnApuQyYjaRa/p9ID92XELW0SarNnSgc6sXY19vilSf78mj3/qpWp8M0Iv70XuremGmWkJwZ9Hb
xcueRs4H0Jaw+lDsafoev60eern5BOfcHAZv1VO/Z10iVM+Jacv6dDzxaBP6zjM2nYNWArNY/8xu
oN7YXl/sEWZOewXVVt2ZwweIyGF4wG44PnR/atr0L7Xod5SAjYdfkt/qGZn7kSSWDjeNGegd2zBE
7276gDk6dd0/pNLK45PU60iEdDU8fy4crJbFMgoKJQ8Rbh7NvNhafckaM0qnd9cAyG91A2dWL39q
ZRMagNI5U1YC/DgBhD+K5xGDhps3xZ+ffuDseRFtYb+dLZqHbGSsBStmx7wXs4rvT3mwVD9PaJi4
ukPPpdepwdyYwXqThqAGb+tvaSz7Eyz0exoTzaT7MnlT5Dt7NAuj2iXmy5gDYEbbJQ9SPztHzbsc
rvn1KhVm8nQ3EWxE9vICmk9eqpH6BusWx9M5T65uKKyIUCYeH6ah+I/4v2BTAGhUA7ZUavhciUqt
gI8VcwCC4zilEwWLvRdaUcLjXtw+4/+2rHvOFhtpeY0yBLViBmU4GgfcWImQ8V4yTkuRcCWI3gR1
/F0r3NiQeELuVqQj8pC9jSdEQAobcgXBYml2V3T+1NbmGcNSsv9JjKi/McO2suoQGiVnM2w34J8M
pNYGvPFRav8IcZStkc8neDy9ekpjmvkkbCfgq1LNsZGaZKoy5wdpZSPSoGJBDJUdacGYFH+gQXQv
9XqxbPUihqgHFBkYRQWNXuVj40qBy7K/8K+RdqMyYcdA7CV+093xprKqRBsVrI91phrNjPADv702
isHbx3FowPWUg3QmIg9F60cpnqzu3/2zKtC53IC1uurfWzabZJIrQYAJYyPOjLHMxkTQE+aJscKg
dTfYcmAlcBBv63YPSwYbWAueQoZsES3GGAJh0fLoT/bT/9xdrFZkGtRLcjh2TAU6TgkCD/PC6cL+
WdJCraN7+zK+3/dcaXLMWCd1yid2BDAreN3z8zAPtEFoBcb6oLZiE+gOWGlj9pLo2tSLEjc7koj0
fGDESa5bD+MXmPx/FZhbqjAz/dkqZjrCElpAlFRnRJGNkoEd4K1qhfDjzEw/KVmd/x3KOezo+X+0
DQAhfgTy9vXzJNfS/m+s4hocaR7UYlhsRlUwVtUzB7x9McjR4339Qv9J2kxNqJLcPtCvFEmEgdUi
L1Gav7BtXAKOMdHK/5phIEQopfn00zGeKafjqwYxm/mfkv8OAUBOb+wjLDTKAU2Kj/K1kToYel2A
ccgXU+BF0rJX+WVQ5LXtjup9/B1Zdnb+AwFVjSTW/Ex78k/TniQdJK0bI+bunwntJmaGoGTOd/7l
1WSjf7UALmInbDE4MSnOx88GC/rRPM/r3c0LhwKyJBoqcLD2q9CDtfQe3mXigD/8oiXm9koAILt9
8ph5aFEvsaudS9PVZOHsJtsuXszorB1v3jHoSKn5Wav7Q2feq483DZ0I5l0BmezAiNDZ0fFIt5le
tJFJcIeVgFDNpJSFz3dVIJ4WX03bT0b55QlNew+qjAPCDN/ysFjeulOn1Oh5nzegnWLHWYW9Un7p
upkp1Boj24GSiQ3h5cVdf40VZ2TCprhuAb+jQFFIB/DOsHmDYj3NxIkBVUCX118B5d/AvUDBo+XL
rx8IYqoeT/9dkm185NyBRNz6tiiz+hYtyrwoKPHwcuZ5RXyseT4vPYKVUHP0s55QxeKxpW/e8oFY
hVGWCk1MRdwU3TKjGtdXVJvt5jQIiNFNJNhBmaECTd+xi6o4VkBIWaoIZO7O8Ca0zYz+RghhQDMc
GSqSLLaj7FuNYwCEWhbSFIZH0F+QwZ3ET3GbqPOMvCcbasIXouRgivQu21daQMyfBrVT5pgkK9MT
J+iBGTTIbb62Y/NuAhPiEGKD0/R+GbQU2+c2fBzw2INJSOXM5YhmwwOpkBhDBneVzrwqma25xLz1
HmGJhcMZ3Xo/KLd1PiPKSUabVwKbckKeNyJlJNeoCLufnLqPE0sUwVPgU8JTg/6oaHaGGsnvcDR3
P42IJ2hmUpW9VBybavJjqTsGJIl7wBwUglJ8aA9wgkGES8Mkka5Q1uUEU6CVCZ/auqfQcqtubrP1
Vvmm3Fa1GYvqFMPY1d8qSNXBJD4BdljSpzjwv/zTInlHU36+j8Fmy+DsPC0cp9mOnfOb83q19gx8
Ekk6veAenakK/msWw6Gm1e1BLgHgeQezHMrbuxstla5YG7WpMENc/7NCS/tb9aGaigNpqhOJl2lm
OEPemS6YsVAWr7ze/iw5dRcaBkZdRgQysrn9CpRF5JEpH2uK/3XBcdMrmVh86T7kExkRo3GQLAOr
jVkVstDK6uaYmSIW4UNW0Nt+IthUEqfvn6fbHxMaNSpOFFHS87AZ9ApM7I34CsqWYN6zXApl1GNW
XhEax1Q8as/kjoFfr0IiEbesC0EX+mPQbSrqJLSnJbHWhjvEH032dauPauHk4Vh11YVUxrxyMfjL
XRdRsg2dfg9Qz6/jJmKVB7uzn2Ga/80F8LmSnheGOvjxjvwpY+7iHv8Tm5h/P2Y0jCzeRw34IXq4
PbRINv7ZOKP85iD+exTTFco7FZGoe3oehI+TRsMwQrd6zjJ+7igK9wycz5UKZHgjZgQOWaAjJUmL
tuKpZsxpPrTnaFRJ2lQyCqGsXU5Uf1YcUXaySNoQMCPSMj7Z514OJxFSzx56DbaHtm+BKUbkGnv3
L/iNwliISxf0wPYI32klMc7/OQngtcVTJra2LlKGrfbdMssUDnPUGhRcqVHzMQ/onUNJbEykjMos
zwKjdbv1E1utUtxcrR5BT1qY81wvRlrztGY9Yrb9WHwQMsQ/rOIPi8Hk0QZcHuasxOHXTbWJpbsw
iGya3uTNU599OOkX0IzPY96nFVLFzh2y0pnHL9hn/0vnyVKvLLQPEcXEaJdkkAGPbxfjX4xQ89Ye
JWADz6Y8Y9Jknn8z/CF/MH7i63M1yTxCqawkGWIBVA1g92Dsy0rFxjoGV68DEgw0kWULBQB+A1Pf
e9gWP2w8w2atv/q4qoYav+Kshjqmj6ako5JLNLigWviBnzukQdj0erXmDjuo6/obOM4QI30LWh1k
YNNvNzcSdN7KQYroAEZG3AoqracrtuiedI8QcSSSizatalTUrp5+/rQ/DAgCmNTW2QcsL10DLqOb
vzLefQd6UbjL0VrR3+JCC6PxRtGNLZVLkf4MV9UPdOAFxG0nluKG+7JMHeMXHCKltM20KTGTF9P8
UPqwJX2jGXm1NfHNNN11z/cPvhT1DBHcIs0pC9q9B7ZHz1ToEpYqrOHlOWmvPGBfv5AaDih6GliK
6z4x5BSyOHFEqvqhi88nN8A/2Up9sOhxyMFU2IZceAnCAu/8JayrKUCRb8R1Cg+5jgbNA+B8LUDw
dCB2wlSrfXJZ20akJmM5gUGd1PzlVUMLZGZPOAAAwkTb2Ez9JdCiZBpk9u+0qqp99MHly5qh/TyK
/P1L8nWA3A7S4aotZkk4kg76VehGf6VP8V6119mG7ECIynLeq5zUx60nqv6bq6k6l8NJT/wYXpGx
dgwjEFBuOYZ3LdEMsPBI5VQl+nnGmfsbZq0lWb6T5N59An+AXQoJ/9xDxUeiYUsdYUgUd0amCayg
Iv5Hhpu9N5UJ3nx7Kw8YVmhVDWPBU9gtAtPjFwPob09KAvMrnbRd1a8eaxSRtmeujcwG/5ec/21K
G6PPZlH0CSGxR5CWB3rs0vOrARd3753tOq1IHV4IuqTZHG2J4wXrvIJVGqtnc7Mtzn1bUfC3QSPD
ELtYkBmBtobTHUYJ+rwBgvFzjgTaTjgADH/V0uRk5GnKxV1OB9cAc6ChgSt0Vx+5f72kXFp/8Mnw
OjwxRKv1ygeTOCXahG8QP55f3QvKkYAxzv975HEtJOZGMaYgQIEUNTCrl/M0yG38QgYC/mYxOi5S
1FOeh3IqJozecBU1dmeAydUFkSDL1OkH2e2FhY/P49zt1sRhiURCvBUuD3b1kCdHTqNRf7wjHhrp
oLFADZgwWHvpql9E7hTyXZd5l61PKuRUaQ+i7LCYeBSSesUNXypFL2hQ5sIlfjtlST7dBlI/OjPM
ANuUsLCflC5HIbd97ipsdDO70EoX7H188ZMmpoSb3yCKz/QGLwQOKOUb+hp3pvrdAB5/uMJNP7Fv
d/rYoIK1yRNK8kM2DF4rqbY7sNLXCDD8fY7wJ2+WOAbNxlQWmNdGUhiTOy2xUV8RfQsQ5OW1v5Hl
iGh6whmLt3Wi61bO307iZHPKViguiyuaJhFySTnMNRHGMqOykHD0m6ZPqNNOX9sEVmBCNJ43kIoL
mmarVB6g04LlrjHc4p+yKVx/BP+XoUCyHiAGtpjLBEiJ1Us0+R8ceDTx+b4iWruR2Bw5iX7UeqHO
vEz3+FKzZYkYF10ejxXD3P25M5N+HwQ7ZC31axGNDdOcX/7U4sebW/2sbcnAQIVtaEO5kJTHV9RX
hJJyUmuvIpgfWf/G3sT5KBMXu5Yh3e9iPAByzCOudQgsfHVZjV1Up+aO/wwaKUoBuIk8Z0w1bQgK
Eu2/8RXUFK5ooQ849tAUiwaNmkgdexTyswqv+FLIfQkeZWUD4XElM4Ycb/0riPOrLj+98k14GgRj
MJBGgdTeCxWWH7/gfCiqtJXOIS9/+LlgRtK74r4ifYOTXbnxyxOcEXlgsJ0PLP5W6X4jiSVD9ahR
svXZFyc7v2+Ekze/OKclEnzAZcOp22XtTTwQHQwxDjgcMeznj4xcBZaXtPxaeKzJKVlAS4Hr3yfw
udKFivZRgOVcsnYThHu7su84yGdYdKLaLrFQMYd8Xr2Bd3tMCgYkzDvSgkQhe6HJ5sLOqOGGB5qF
sfCx3Vo2WTWN1HcYkIdASc07dPMP/Ge3w4CCcMMI0NGrLq9oL4pD6UoSChk24BV5pCBnkWK4yZzx
KS39l3JX4DtSeXw+Cn1/rKOCd5xD4hoU7sdWi3EqfsjudqSO7zpLsikD0/7IHSkOd3wxZn8qWgg2
60tLqADjkDtjCdqsDyMRgfjmfEdk+YOczhmkQ2zM52v9f+rzqJBooLDv8d89oIqCS/WRYwGnGhEk
6BiNwXSssCXvb4f2OTpGO1RN4KAH8+0q35aGT6kmTHbXvrspZjtOpyik1ODMicCVtPsgllqCSdee
7DecZtgAU2daMubVnKgMpjZQ78NO3a3HW+5Ij/oZjBaegliIaxUAeUl9kZbmbJWKpys2gEmG6mnm
eb4IarnfL0BRXriv/BlaK8xDFtak9spwgRUpoyTax/08SjZNma4nWbCVyLI77kmr86W0V1jOmRiI
wgkjhfHtXiYd8/RpLeyaPbTHl/ufs5G8cYTVfMykTdWrDP76s+IBT9EDMQdHTH1vwapETP5TCBkO
1lGev3xRCdEWFODr9DP6hKf1QQ6HlzA/Xo5XHkB/8m8MX6NwZigbKdULnGyp8dXzNSAGxTkM+Z0s
dY3KJXuaw4UWJwz/I0TrrVOAqQ9iDlRkRsS9OrYT+mvA8udW1acEgUg82U1xWMBBqmk/WKsESdno
sAvShivapiXkIGEVYR0sPnAbsAHtSY835JbGkUJhnmrtdKp36UqRJMkYxjRAvs8SrWI52Jv+GVbN
ZqzcJ09kEvdD1oDf+KRqPXd/RI7lyDL4UjsO8sfDKFLqJe7uGSlqOszBWBhGotAwDcM1s5Ice1lh
JP4X9tJTT0ab58AHfCHa1VdqzZqJ6+tYmBg/UHoB0PCxJ8MG8G2srgGJaDl5x3I+X0Ljs3gNbZRl
AbEuFobpDfXCsMpFEwG7hWk3qbXja73gt3+QRa9skTojCrxcapWAcAqaa3aLxnI+7zvuu55ftGx8
jOg3kHjXZLcaI6ojPva9P2vBfQyHVyEOIsPM8sWB434L5DLomImXNzuWwuYcsj7JCJ4mIcoPs5Su
ijFQqgaTUhKPWqt8FKWpFjTI9F4Tl38CFQrT9Z+o80e8PS4X13yBPgnmYC9W0y6040xHdXTjdfRe
jnUZOi0y+4KuXThWja3vZhE6qPiQla8Xd/bHNhAJ7TXVGqn5ELXWV8gkpXz8ED9HzQFFou6RRkoT
6CvEnEtqaiKhCMlcjzTcudvG3e4l/RWvPVwlyYk+WJV+ggZoFmPdRKIKR1xtB4/T6p9JMF7z2IEa
9CJ1CJYSWrnQMoKpphhVye5nyqZWxJyUIoLfqg+pLWyJ8nJepuwDncORvctxAuA9H0pPqrPNfanE
Lp7GvCFriiLoQ7oaYKOnGJhsV5FviHr0thoAuZDm5tJ3P5hO/JCcZa7vji5yGXPBvNo6HCY6qKei
7hHweOT3j5dqnCHl85fHcxpNUvDB88c6B+GUPUCjUk31BMhM1wM/z1G7a62w2BHkw9W+oqwVLXHn
NCchfsh+ZdaT6Zrc73djdQzE62TVNZYWh/reuFNZOmCbv9SsfF3+Jv/5rLxYKvQc9ptDd5Ck0jSq
UYndOmMJaMb5udUA/zg9DK8bRDBd6MRMkNgfQzzHRTb/YF0/0WrTgwm4v/sTi4yG2UntwDb9IESb
efLyVuKdYGVZnYQn03qLdvZGgFOfigr3zYk+T6qZ2N2zPmITIXIuaJ3xJNyEFuMxveWGROJOMuKG
X8lOp+vxobHOs3sxotMZ0S+KrhpjZTT052vkLtWCqNYmxa+tT/k54w6xe8sY8x+IQzEfGxdpKxte
YppbuPN3P5Kv9QDCkkcpbEFjKWNCFeqAsYSfWLDpQqDDO8GPCiWFbFs8jxLWlTf4rpUoh3fDh17m
B+T/JYzgNcwpbhGNryPN4iuKJ+QmpZ2PZN7zwkhaFGx+ogj8BFYVY7IXW/+7zeoDFpPiGGmrybMv
Kghzu9d8ZHAuwsywSAX903ZfehETT3X2lF8gCfpgJQanDa4Ak6T/8CEzLQFVGruFv0ZXOtpEW1Nv
yCaQERuV3np0g5At2p/Ln6TP1p9IsLlBKCuN95FcFWF/6UlauOP4bnThvd6s+859YBNGtuevRE9J
nT4B1z5x9mom/436EfTIkCKWREjuJTzayLnmhucNORtFspk2o6bhk7ABGLvD0r2oEuQt2fAg+NPa
AhcYsO4yMl+qOR4c6F+wzhDh1i5j3kl14zFc7wMNuM/pFLrtfPKOH4leA9Fq/C6E2/nPdqS/o/gL
e5x3zlQz/g9RWubJVRP92WF6/RLCcx37odOP+bIlRM+hlFeaBJJYOxmBfcTuLSZjHao0ax6KDoNp
YtQJgBBssgy7iccj8lggDsxTCfSX7YDliyo0kdCGGqzukgunJpbNkJ4sDx0g1ZXhvrdSd8PWro9g
B5JSLmTYvwqeAZ78rtzDid8OOYb80FdPfC0P7xz77POI6K8WSQEHXAD5Q796ffxyk097wgVoC5bF
eoioN8zISTVfI8lAwmLG8/HDDEEjGcY0tRv0EFvuGgwKene7T+WDZ2pTN8s1B3gQ6NWrtybB0Tsn
zcTZrtoeLlL10KBUHhSt+Atuk6BkXDy37UEWLDZGIchNeHTQP6r20Wup/tiR2Y7EkzVsf91fpDat
KpVukdRvXloB2Vvgt7XXgDxom2D1rOtZz5w/X4F1dkJK/pccU67TU0ZcRCv6vd2nNpdhC/lcKWb8
ggtc+CYVl7Xp7+cEtgj6E76x2d3YQu4yY8FWaS7vDxzi6JqeOr8ydGBfctOVZPGDxwErOdmg+Ref
9FfArSQe7gf1tBXpTs63CNHMBGQCBpaXI/qm15KZOEEM/JwpBGZovJG9npQRGeVa+CjqRAwp45C7
OzFmR6bCabfh+9YCOI6Bcc6e5uYOEKLr7Apv/W/q5dyrNJcrt35ptFMdZOELIZJfvBhLvzgG1JqK
cPaxOBkpppfeCtKqr2lhwCd3X4opC1Y3sfRkVkpdFOzDx+x+LUfo2mWcR+AGoDrjvb4YnJCaPlC/
12HDKt5y0Je3ezqcjdadbafMQA7KDsUdHypUZLuhXGGdyTJB5+J8DLP8SzksOC8FYS6iCtx6UKd+
IuhbVPHLlbIKqsozkcpoohRFdm+SVGuacQwDQoUbbfpz3t4BcTkc9olw6suay8Q8SUHKkX2f7iqk
mM2o9EjwgR0tfOxhhiyBIR2DugYr2B7EgD/aAHjGMiBYM/V59x1svRQZ9RKPSsTjseOH9md6fDG4
eP/iYAN6azaNbG4I40LlYRxXE4xiKzBsL5LbPfAkBEH7lYerpIX0uHTRuK7TqRBDZrTY9m6e+CCM
nev9KHlf2W0LKjzjupj0jNc5N624d5L/e4FonsVApYZR8PQnjFxRTDBv9DyHt/FPXOCaC0eSwfTg
ReygjDkWtHo6X9O488x9d77NhSQWdKawikIqy/kRoRt1D2RKUrwxTfydSYELtgW5Z8JJ+P/K9piH
K2kZDsDyjT9JH2C/xj1SnMzkVSHJTr1h0UHU4WPD/joJ4f0D+IYb17LFdBK6TYNebeRpI3hih7jx
vlawlc72dCt5yDB0XSQsGUTIPu2wEyaLEulsdy5O7TCDJAqYe5JLzHMjbjEKcrEMBRXjmcPmy24n
rKrOamGbXB8DnQePct30G6cNBY2cUaDiwCxHrnaTURP3K9Z/L5zPzrEFNhgM2dRDrcBPFC9kPsaA
nV13K5Bnm1TuD7IbrIm974sVpNPLUfEYSTg5wsh8c1ErjCd0WloEiBNmeJsyD0T0zhfPoCzWr6pW
G+CM+OOIvkna6l79jINUqIczbGZ9bRAS+bhpIlBPQZCExPM8WpwjRcwiVNRrSHJ0jbdNh8RigU22
OZ/6ElIwdGPUZPSHfj+AMgAfGEW/6XCO0f4CNfyLJieZOxWRk79lQyh8+J3ps/nrRxjpuPEHGUxA
m9YjAFWI9Hp/rzBwRdd1UC0qhVmLdjN4pr5za3yan/ROcIWBeuol1+QtagjZ5iTdMOD5w9m8+jjc
BWz/JKuQRUEwEdxL/839zlIY6Je3V9bpQPVt6dvme6/OuqaLnzrEXiANzIVpjbKSXvf06NGezOMi
aUzxk/uePS7xUqdAPbXqgYrKTeyjF0X2a+gnmCwVlNj/b7NnWT3vVSudoMPvnJFfhxtW2Z3AJuv9
opsBVxFGjQLDSdJjuTppRmaGHIwBwpPZ9pAbz2Ei1KtIFfrrxPLkk9FM8FrNhJ/Spzp0/6sq2+Dn
F6ky28LAOHHgcUAgndMmTA5XesN4S2cSXqoQjZx32SDtUv1X4+5dXTNuCgGHryJeujJoBpoVMQwc
MjaXFxYoIyVR5zLwD78n3SdDT2Vsr7OfPg0CWk5LiuR1t/VSM9uW/U+D7S2f7dpfMbWaD/OcCFPB
cIULPWki/cWlUeC/rarye2cTFAZ2bR4VRtfIGw3rBuQyvusrJXOh3QE2IceSk7OyjLCrmMfo27mS
22sZ8qsLWBxuIZzAMkOCOd2fTvDPFAuejkAyrMOq/ZqIBx+aCnTELBHKN54fdoEXo5/ukmC97L/H
tYTQwKPgkDu4RnJ8ilGf+Gr3hLYpDOyAmhfymp9Urh+HJgkA7wv5omSCtNogdpRyBodhI5IN0M/i
MpQTxTQFgA8CXRfGQegU8ECPk3XfH8eSLl53m6TgNetgrpWPdfY7/FyI8mpft2IpLHm9F5r5CjdA
ryKC+behZVCWL34ALTj/yfNTPsrD751ULf6Ok8kmNfF1lIvl0jMtEPq42x6WD4brKAba6OaDgCdg
LRG/Z+QUlc8Iw5Fw3oHPNBgCncvKRaq2lVwAedC7VUjBnmYcHXavw8ykn0OMPmL28VYEfY5oIX8q
TyscaUJmO3rpe5p/LkpLIGcMaGwLE5dnlkn6tE/2RlCQNZCQ+CWT7pPyBmuma0Kr96+gkQ2UHZR2
PsGo465mZGvWS2knUU2FJW77Kp3NmRwvU8UIUgHVLtvmrWa110nGm4y1yHAb1KlOpfM+nugi1wfC
FxP+Rvmcf/EPiKyh2mFDSdxyUynQ8nRN8APRtRFfUQWdAkscjKCtCIFnJbS4E8n70rMog7siCzaO
B46Kntd3LTourcDK6SocAmrzq8WSk+XyUMsjqqpnthYJY9YML/0BtSETd+UTWg83bKFrpzZEucuZ
1I6msOzqlQGKC8A2Z9flC58YgXu+qyyFsCIHgMmKx0oKv0l7vwH1nPWy4wnTENVvF04cFzbUxzq4
D8OGJ5XTbepiBulLetX/UGKt3pDc2lgFYUQ83iJAp0XKJwlEBkDaIGJiHFjdvoB7c91k9f9Y5j7w
nzNfXM57Cdqq3YZ66bnbkyTaySUHChm2jI2Icak3YPb1M6nOXHU/K6E7sdeAScMUtJAnNy+UtLMi
x/Yhf8Ff3V8j6BtwoXNyhPf7nuaLil03tqP9MfoavXsdOBQ3a3TS9fPG4Phi26ImRasU217xcr+i
YIKXgvu8Splo8Kmpmu2u/HE7WebY6NSED+vEDTq/17m5bdjbP9JjV/0MHvLVpMrihMe/Rmu5EyPE
d9zOekYDCoiuNCxdAhTyQdzkHUMASmE+sY/FP9EoedM6nVMpkrqoAuisqzIxq6Ocrp7MEqMmkZg6
NDheN0+xQZQlSMKMJNAdx8WbFzu0dBakPlE+33Aa1py0iNEwzLXSogf2NRBh9w91L5VSZI4nzyYT
MyiSDz97S+dSazw4TToP9/Ho4+owLVdqvPx+OKK4FdcSoPPjnlhwOT4IPRP6ML9WvuaUMjevw/Xw
A88b+7ChzaF0hxWvW9vTyzGOD+xeZhO+y1zw8Zi2Eph6KXPSP15Bepb1uOJENhT+JWDYrRE7jpG/
HRi9vQItZvJaa0hFhwVFbaJXPFooCxBEsZFYA5yQfvmR1+a/sv2uk/XW7ylIoHIjKXcN+F4bM27d
B3N5bDRHFszZT/yVJNd7hvDOEnW5hoYvuMw3I9OMqUT8/rTcxwpNR0wbdK9mdy2kNIVwtJgRXcn2
5+qOYRiaUgpOKBHQMtyZSM3utdUCSsLatm96iUFNmUlKYIVz/eFWbEsbvYW4TcsRF3I13GJ7jhhU
1jHXXNfEw8L7QJ4etNSb9ZhESCCMvigOnFqCRlbjRLoZCdMSVtSD9eRDF0/kskKnNqws/4J8fydn
NlE1jC3s94N93pliGoVBsQ3iadxpuV9RFIEmhuvROxYcABt4aPr6DkQERowyLJMJCVwexW7dHqM0
o3lwg4ykW+mLOeyxwP7EeQMTpxlVUs640QGPFNw4JmvvkiKGCw0juHzcHBWxRy6J1u41oC5dqjGw
M3B64rJtKVFPiOv60R50dho3rMYQKlncag+grxcqSClw2LOsKjz6NMuVJdQB4vQ+4NA5ysnXQX3S
fva1b+CLLBqoBmVuZkBQvKb3MGhBWfCW21JAz1/66upvVNBTzi4EKnrdVo0qBBToE9Y/i4cd5e6F
31duor+OJ15Cbo4Q5LudABqYXimKO+GBhfDcHITJRhGTvg34kOIJzJpK6/JmgYMH4A3miaGPtLfw
lG6P12eqtJw0JxmdL03JtipsGcn2SdAJT3B4dW47u+SmncWLfMs3K20wS4zWUPDeqtL47ma9qcGr
YnWMeAQUmS5VSuD8irPfB0QTyraNWEvW2RS3f/Kfo5m1M0+pHpw7DmaX9YpVDW7oWgakX41xwC2V
XxMDVPtqXc/1DkrQvEocy5UKLCGfRvKfD1ejS5v3z9i11bwBFQzmXNGoFPUhHBggeARzxNJ/8lDS
UXy8oQxSjfbmyuaOVOoceh3JVvH0o9H1lo/9lpA61pGpqWjiLXz7Vux3C/bIQPHsbDkfCEK6t7io
Fp/vtFzuoVC/0sUAmsTNbJLVSm1VrbRhEOLLnah4vnEyuIAQSToZpwVN1fXwnbe23NDpktSHlkP2
a5gebfCbeJTuQF54RHXZJRvDC20b56SiYQa3tiirfbfyQWYm6/Cet5UOFFOosv3ZfZH4x+nBcxuM
WbhaKOswrBYmY3Pfd9Uv/PIe831t1NjhLrfXQAgGXrodWnI87bDupheEH2edwxqT0B3IFwdbSzHa
0wjUjujB+K6ksIcQ80tb43KN06xCSU6Cmzop1WWIoBvB+RK45r/gFs8pCjIdmKdfTo+GZmBbSz2V
4EzZBY6/ppZ9lt6su5onnj+VJKTnsm+RiqVMS6jBracI7LfDUjs88hQzP0OVoWxjOak5hrhgd/H4
UT/X9Lq5VFGs+J3ZdKGQMlucFS5c9pQVwkdRf3lz28rlNvn6z9JzkekKYIlgjm9Bt89mSbYFfK03
TLpKnoG/polmFCQqb8nOo5S9w9NLC5Fc0CAo9RlZDJjbBIeFMaE8bSjCjyT2BVYbxsVoSA0F6i2U
iRkuDAcCo/mvIWDQ36a6o9+kTubSktED2I2LxIac1UVvhkmQc7nsW+7aZ/mi3XVZ99LUGkmzi+RK
DwD5JH7HhXBUyBzuTsSdPCeU3NS/tdFx3iZKJ7V+haOMrWfrIzhqQNgieL/hWYBMmmgcgOqu3k3N
gQNqVmsaHvBzKC3vmNS7PHuVtS4EBMyHhJSUTZu4WXpl0mNwnYZcLA0vAHkKk0p61D3+pfsJeLy6
KKbhKQu7+L0TMSl6lq31Z4pjGUrTewfdKXn9IunsfJocPj8/GhQL62TP/INrNlLrhGerhQ2/baRU
LAa4zr0tLk6FqaJWajCRqKz6ejQpDnlAmM0ZSg38SfGfGAOrhrxqvoVli1I83/wumVNMvF2pVWW+
WnU7u/OeRxm3BpZEtz7Cp1r54vOJVMaiYdCBmXicSw8HO0OKvG77C48TPhAnkUZ8VH9kQ84CAWba
3gWIHxKBrozHdVZ0pB2INcB8RGDTWNvs1+VcTBEiwNBzaF/UQY8p868dOmxULyAp8/tgQX6uCe+Q
9nbvPQZrK0SgXk5PWGuwmikZuwIe0A7QRM61hvMzQlqwC8UThPbKUcMPoePYzLQDQsPaUzzMTien
yx8WXJMyMQyskz6b30TvDu1v6R63pWF3iHJNc1ux4VKEw25jMzcx9DdNVo5gLW46vxGsbdNt7mNa
s7LGZjeLlx33OHQwaOD0EI3wcJp0sNoibxOuXtT/qPIpP8YByjNBUO+IGrkx4U2mSFDUOqJbkIfo
rEgd761qvsZ0EH8SLTHLzdfNq+nNoA9KvFAL3xxzz6qTZ7Cx6mWY7iWaFTUEUTeIzXrt7YSw/xn5
zGsPu4HA1+ClAKwz4Ijxmb0XSAK29vOnsaNlfHjqIgptlBD1Ic2S6bVYl1csDr4oF5YJ/WDUPpNz
nmlDWYoSYo9TyN3t6e/XusZAeogvGTYj6SXDnVxGMBFyPjozkd73PxgvkoqSZprequoagLACnwnv
l+kqOOZxeFhVKiJBWVirE7aOepd5u2E/lKDCpMP4RgXOX8IC7d9Y2QEkSmDpwm1Fn8NSD6+CLVfW
u9texN/lWR8IB/eD8Q7rSeoQmHnJeFvTfeX89qY5q/Au3j1zose3DL0Zf+h6SEubcwu1Xt5DFXKo
dMunw4va0EFL10+oqpUQQ5sNczRjlAYl2JjKsRmWI6dZ9cZdjbXatmdNwFI4Y9z4VF+czslc6300
1tyxzwEIxppOH4Cj07A+5GcAJrxINKvnXqpTdlu94L8guEezTTU/uHNPkL0mfQ6n0dtrzyATSMJM
fzitD8yvQbVO0qEK/55xdNvTb3ir+FtC+jmKpNSV9UZfqFgPGalA3hbXwPR+b4MuftJbOwLDeOl9
L6ZyNraWCrVPWDvLsf6l+eSSDRGQGR4ff3hik4ixuT+o6iw9LfUUoTLb7z5IYZpPEys5KyjnGKGK
EfF9mIIkFWjmxG3Y8rma0sOos493oyWj1WMVHaKDTdUKKWJCxCNHIco0G1BmXn9TgJjf44JBMxYG
c7wUKgxR2bA7G6GwM5Rpp8DIDLNi0Wj6vvIWGq2pyKvkHuBUjhs73axAyYHbsRFZXyJS9G4dGrLF
Grkb1ZQnNtVG0hrBc1Wi8J+nA4I1eGCLir8F49LFPUK6h2CvxHIX4GNmfv6/rGtO3NPdyKmXWD0e
33QQwhZh/RvWQ+X6CLsX/Lrbg7KNqIL6lHQd3/tNNWVilEhmPY+W0bTsygbup+KZoCOcZvQbaorf
Ul/592ZCPjsillRmdBYysM8eIxX2yb8eZb+zyG24VCprslO6BAZYsLBKErwwhumBFBWUsIngUTGH
I7YtU+cESHv43xkkAF8RzqA0nOKfinc6plP741exVLyhbMHT5njxqP/GfYtAKB7afxB47ZCGnqOl
b6hVEr1XW4hNn9giunYENo5+K1mGLr+BUP7EVAHhR4R0IJZw1eCVlLbGYJ63Wyqyg6QPoSIDDwaM
nwgpHHJ+8BYk1gLYYVNSzXqPH19LfNE7XJngoW2f9L++W8nKvW9qroyQN5N4WH5uFkD34wSbd6r7
T/3Ov/8uJrA349OuV5Bib3ZJhTkZbUIxPYPA1+f9GxdRUTT/s8Az6ey5BI0b1wgCT4qlA4J5OqZt
whEodWPgnakSN2GrKel+8bftDRoPnDSA9CuHOtvgGSDDYcGW2kkIGbjCisf/GS1dZD0l6i6I3P9u
Ldnx/lDuZjQVaj6baXFTomrKMEzRrAi0kiCD4HXiHOR/82RG6vk62L5+MXpDVCBGwqdfRa6EuvBV
eTSxjQqHMKYIz/OHdymJMbVO93UR332KURj8TmMfbfdFIgw36HchNBOPFuwvonklBdicX/TbjLuh
rHe+rRWrsrhwcqqhNuCwbMBtJOURSBwFTmL+7uOCde/udA6TXK14FdntzPkKNFqZRsyfOtVqS4JQ
R4/p8G7vnl+Y2aLJtsXZRsG2VGhObb6i5d+I0qH/RwzTlx/tvakzny+tPGVUgX0jQJrg2YfHp8ID
z4o+kd8mNtUPaAIJhmbF935u9F3aFYI9tDat66EJsFKx8jgh0PdBk8wos0Hm0rbnju4fUWTmAUHQ
RmPpdI7Xd4caqZSSrw6HCu051S3/yUKAo8GLzxfodVwBeNGVr1b8FAXApzSrFfbRIP4v5tIdIXcn
4mhbpCSryLDLnCrs6LyI61jr0U0fW2UhoHMdezs8OLmhgVgml12MpNEClGd/tAuqaVhGsKM/gV8a
1YrVGXvea2VY5twF2LQ4kGb8V8O1hFpGHSNw2yf9k/wV+iP8BlaZZlb+Fw4ckquFF5n9zSMtaQNj
yK7FT0DYCG4PTXpAsJydvn05m/BEXHfAuwZkrFiLVtzhAohws/YIimrB1AUHPW8ETsmx0gSLSDKr
PzCikwb/8bOkLwvdyYkmakI9Uy3yfyYSykG91Mwra3vfpOC3PBJrTKeJCIDJhE6JRggmwSWYlbuG
oAosE8bnPP8pq8Vo1jl17XCYC/APz5IoVIsiZ7Ym1w60PN6T1uqR9RraZrKC/GD7hj2vcYqRkCIK
5/hlRqm6/lgRrM1nmc77y2f+iAoDYGl905PWMylmiCp9inyB63agaJeF29rqxZYPzzJxrE0niQkW
bRppvRp1Dxl7WPBYQrZyNRhKrIV6jicmCIHx5pbYAHML6nGMrPahYD4Fla18f+Qf1xMFJ8jk1czR
A/Jr6iFpDStrTsGxgMWBwLSwr7THuBeFkIWWmpAH4wC6AplbJHtV97Ftn7Zyhyb69kJrEkcE3czf
tXUL7kQlZT8WjzOk40kyIhvHrxDRPHfLwCXr2nmmXPCuyNXe9ALYKOTmke5Mbc30KrNzHgowlin7
ElHPrHoMiYL6ry8K5EHBmNdawrSVrQXS+kcu9UKCMtl/jsWmcHCa9vUrABN1Vl5K/D7YTjvkTVoD
1dtaE6cFxmw01ndPBdagnnPiE/YrLYjMZooHJL1hBDAn2Js+9QhtNyT74BOV4wDOIQ+7bmkK1uhp
KPYMaSy5Jf+KO2UkSBtwNWcMJ1mojHmL3d6o+OJO5dp//YqGhEbPTKMLRrckqcsnZeJhI91V3NDH
AFPHtXC6r16Fzh//zB/aSmYM3/ZOk7o19PmCMSKHhJu50oIUqm+giOP1ERFwCW0q5uIKSlnvpAEY
oV60y9rNXtBjKypNcu6l98BXQTb36yes74J0wTJEfkOABmB3ExfV+CQoim9sxFQQaI6j1EuttMCk
hgsG9Cn2mReyd8ju4JKaNPoOQdHB3NfDeD/3Zr4x/VM46pIroAoRzcY9ak17IMl7R3W9pC2kN4Wj
VCpZ5902iR4+Yo3bo7QO9NlRCBUHpYoV4U3aaUpqZKvsgzXhcXSYbTsFEhU6Z5/mmSuM19iNcE+E
u3Dp8QOVJx6CYIiIn/u2jaXZ9Vq+9fm4HhVUSOoFyeyLZEUCCKZLX4Cr0RcS4Pi7X7Tx+2xVI+6W
R2wen3mpPjpPN8tNfak7SaU8e/tfXwYzzkuShqoD4C8f+RaRm4nAwLDj6StElB8hNWEzSRNcsFOD
+8pRKL4XnP1w/25pGfyfmj1m09VMeS6U6Iyn2T8p7OfeJN2nL/Hjy9PKDuz4jPV0//o2hUFmqDbM
G/wmeaJzbCt0cbaWk+1yz22Qyt4uNpE/l7WwiRhbgjpSqcFhd0Og9SPj8XitGmBItRWBzDpgj5P3
dmM8jyN1UyjeKBOSAjxVeFv/bdY+4PG3pIaGDpjgm+a/Hre9O4Lr0ZVNNxVmF8nLo0ofSaZ4qibE
aozx0/P1jba5VbfuCIAkQIDoeTf+m8BKlKZOEPkTUH7tn5wz6auK68asED6PBpqpI6OBlxztSuXH
//6KbTsTTG8iKi5dykas9XR19Y9yXnmakAEp5U1oY/VttLAPKgPv75EH3kp3wFN95SdmX5xM2h6/
U3rl7a0IRpuD0M5HBMxKh/lx+kPrNKzdoSSOEDd8Do2v3fOqTfz/qc6HNzX3XnVAIDSvqYIftbU1
KQpTmZ2ow6iDV42VeTRTJ/oyckA3/SP02Ojzev3Pab7J4dNAe1uEFzjDuWHmwpnXUgUqzNC2cNWb
Xen7+drnsyW6BGN18YPK2CWIb7i1wGEOGhPpDi6ioLCUf15JkkuatAhHueCkp6H8N/2tJc9iROdE
OjKNNChrx7PnvpVtgxoSQQi4Dzd6TAa7/XxqMYWLXleQM5M9mPS/bCWO/EajGSDDgRMCEww0RYyG
rGBcnGxPfn4CBb/iKhhWH33B3QcYAIWIWwiKoWbp16C0Pwg+BQnpBaeP9vhjSJlUvI+nkMd1u8NA
zD7vZ8I0mF43fFNoF6PuC5i+BpxGfMaiUSgNsaNLYp04w3T6NzThsWEv6pflGDLm6v+MEe6UxfnB
uTIaGt7JdpQQtmlIIof5jgM21GfVC4u51HO/jKuwog17DyH2N/qR6usmvLF3Ict3i8JrXJgoig9x
OEy3lG29EHJ9N2n+4pB7eoXVvM9mNxLSP6lod/RAaOyl0m0wJdgOMl4YXFMq/aNRS6SCgTuZ3nND
Oo18IoMGo9rQb3mklfN20jXO+TnwUF0p3sSnPER66tAx4dxiL/OC3SdPd6VkD10cEsYAxgdO0XcB
lBfs2vtxeB24vAwqxHtLuwW/6gJ7vewkrolQo+DIw/Eo9lk9lgxDqeZIu/bcYYxOcQo0wPsCaMvz
ZHoUn+so4sctS0KRngueOobwQ72uhwpFZTXDUnf9Zx9JjZvEj5te/Wqip6K7go6ocO5OZZgnC3EI
HZw+QautSvgPIoYJ7eVHbqeah3x8XRNQo0qlscecIvxHimzjSpBwsBAHeZTfXDQqSxXOiNcta2dB
67SXWrB1MV9ciJp0pEjX4UWuAkRP8usy7PBHPM5P2lpCxce+hMFks4I8oulw+ExSaShPNy6dropg
tY5yy6rUHtzrN59PV8lEDncOgwc7GdIL3eQQerq1/CLZJ/VOMbl0A/srODcXQ4aEcZOUHLdaEhSM
6l8CNVJVoCHi+MpDv3w+Gfk4qOPiw+/p2M3EKJ+UIJzgZ7jfowmhwpYEqXKpdW8QQ1fqD+OZTpKr
sY6zbqeFTaZLwfQpqijozY9EQxLq2pgYL1vnQSE9MdQFaU7h5gA/IRvxzAAiDB9Zt7Ud+oQCBCTU
0jWYc2qRuzsjUPlv4/S7Hbqrn5qM78f5qOG0HSwr2ODesAc2WkXtetAWsSGiIDoE2sjTuQItvkrd
G5ltoPKWk8r04Oh121xDPkCMIsF1Ug7w76yiZdJTYEr42orYqH6suW3ocFWc0EWLAFHfzirov11o
8v4aV7+fkv2hJBr6lRVr+5nFeZFfrj/5uhiVSA2GHcziU5Vs1A3D9Ogvm7KOJqj6sghi2xdcjvDa
T2DEdGRoEXr0GPsPPw0OzZLgDj7JJq4NGjhbJeov0DsFMzDf+k5W8Lw22XSTcNBJQdSaRlr8WHNy
Hk5i1RcWEhmVJLJm5TH1/B7Qdgdj6TcvXltOKqioTX/aVFW1tqwr1EiPvOAuiAvXufptFEaCQAGY
bgg1vyrrqn8pWWdqHQr8e9pWHo0udqcFZfhLLx12OwczeIZeMrXA0kisXqpVduajkeC/juUP6TYg
8FPyOXnTS6T5ILRN2Ox19dMIffG7pbNUXrexjsW2xFQCvv+oNwIQkQLvUEdFzGtsfS7mvb9ZIfVv
43vobc5BOBaS3KI3tWijkDrCSKbLuxIgusd1nXomjF6pPO96oEs5aJ4nEeqpXlCzEBIOmMg0H7Pb
qE+UgPzjkDCuihRRn+Gy2BsFQyzdwDaXz9T1Hbwl0Qr+QsDhXCm0u0qRLYaM0+THtz00yqFvyIks
GATy5oNql0roMbKvxFLQ5DN21dfWUbPk2VENYDg5+9sBhQEuq55R6QoU1R9IKCSC6tX7Owcboa9z
dMC4UJXgrHC+EwQoQkl8uNCb3efKrceH48mw3DCe0dDyoFidowY0zjgPdYe3jSK3vZydoqYxHiIf
Pusew3JjCMkpzeZRdgtPi/waycR9wDA5Wb/uAHFKOXn3xhyAsXBGaeTHvtFzAHxN++DzIXkmT/vy
NmcNHNAaYYCNTnkAmjxpahWPcWmymWiLPZpUj8nUUcPCbwxkPlHyYguy0RrARsseNktJmEMPOyMl
YY2gRE/kfDVCfyOWiDQAnjtXXzdHVbctC1G/aN0Sn3j0mCgcxOGIEcYHDkEJckRvC7Ol0batYGYC
8G3sQZqDp4RGn7IHw2kVCQkcMJcmNUQU5z8ZsYyL8UFJ5Gtf074frBXA2l/wFt56ooOI7HMXX9B9
8kvOuXGw8Z9Qmg7usswaRZZ1Wk9AWt96dgoEQ3gwkDV0VSCNuwizmS/2S5QGHOAeq/AFmXr/9zB1
vDoQU8sV19ZFJFLyDJ0FYsHbHNdyO3aq74I+PiqwhCE71cJYQkRTYxrHEB3DVf+b4urSgXfMfg8+
GbSGSMqaSteYeZnzY46x4qr7AtLhuL8OaKk1q+mHFncv8j6Pe1pL/sQ+7m7uZ4f8jO5ref7lYr26
ZmTDEtH+/aF40XUhRywwTnsOvD5J775CbjC+4BVzrYOp56vgQstphu5TshJB6a8r3qNEos+DNVkl
D66kwsPNjVUXMpcNFbqW5BXM8Re17tCHle8hz6FMH57H23n/1rD3eNjb7qk1mIhbMI9kz+ef3wl6
lpKRSGTSXIzh89ZXQUu+gjmDvXE+4LjMnsR3VzXe9ko35i/8KpDyKCxtIYQ/+Vjmt1R5sF3RoPYZ
APTn/NYQnbvckTBIA4z5+2RlqNynBwZTkliMdseJEA3ppyoG1fZEGVYUqzgM1WnlkuK667XwkhLh
ehlOx2xIx6uy58gw0NSIfNTpylC71Hywb91QtgthD6ASwCCD5gZ6ZMStoAM3XfwHhONnnSq6nKBD
by1R4c8SzkF4bpeoElRjZ+8SaRdkGzTm1IlXJi6qnMCSMrxHPuRKVRea2CbPnBHp2RHWNf+VorI/
a78q5i1u6nqEOVoMzatxQ6q+Z9akzRXkVbs2x4A14jvnz9Si5C0BqSWHX7PcnkZXLNh+tXU1ZLG/
Wq6WS4MQhmg7dSEIFWBD/56i7xeKoDt7251/7F72JoGUw1ZwMGXl0eodNvIwKJ1e3aEuc7xMFrDQ
0iuBhItdwAcl4LkqccqaRR0iE4RT8xZNgPhHV6CurTC0qgTTbSG22WFUtoCdGZXx2N9s78mfjdE9
Zvk6IQcYc9Js+Mna4oT8jyo2ARD/oLdaBkpOwfSjyLV2swXX2ZvXSnOVcsWHMq6DvzFzOwePxCnQ
3rvF3agFVgQWbk/dUjF40islmpsVM7D9TPR3WPZak7tm9dgGwSEEY7qHSEDUoEOERaQk/lsZj9R3
C5kpjLJ3j16YTD2L5Hbec6qPJy/kpfLRT7SW/mIF+DyAZnu3j8x0oz5x/6cFpTcwWxqInhO7rQX2
RTBc7mQkHawyUxa4bjK2jP/9vq951oGuoCOzBc9TmZBFbsMTtKTYoJMzylRURUFjMsBgn1Kwql6m
WI4qI7F9cJvNbINLb8F9tIem6+z5BzbBnh9iu9jp7e4O3kIoS0roXC+633SEk6Jpt20AFwqNrQT3
6gspttWUiF3SgtRRKEWlrppR1oZV11LK7ZEKQl9TVRBZish+ypJQTJiRz2gDJhCQ1yWBooRu8ai/
VLSIzMF7K2WJfi5d+B9JsX0TiSRnZPkEAABC83rcDSgrUTDhvvOpTSvcvsVNqCNaOyGpKFz/dCAZ
cxoBxgXMvK4fl1uCBiSZxyh2Ze09iZWm1i20WQ7kBlI2J9R3ayJQmCSx1uQ6iRNA5WGAVfDCCPBL
8TLlRsq0ZD3HxHW9m1Tb1A0IIYWK2FsfSKifLlasjas0U+K5qew7X5XqQJkQRCI347zt21/tZ7aD
yFbh/ynijL5IG7YSKJgsqQf0yBkEuNUHSDCPVcff7gdphVdH/TOP1QV8dAiTylZnuVG/lQ5zGaEH
b4qeysTLkcbu69onfkTsfx0/8W82sBLPC8yuNV7TgKZk3+csPbQP2UOQPR5/zQ+K56jld/NPwa4D
y72kySIhUsCpsGOZCTsFvFfpU6r+yQ4t4idiH8BItsz74AGOZY7S+x49GIh4DbaRyUxeqGVI3kb1
blLZkYcgVfpqDl3p6T7rXNx89/d8PBTbKeDsxxGRl1lmtliyqbD4lUZ5J3fcZqsTGUdo+JGUHtik
ouR2vqCcwL0OlmHgiomYSC3C8DZjmOGr/nWtXhBKZGKGo53zdcyyNxZPP3w8ZDG7QRsgfOW3+GTd
hSO7kMDvLTGXGfsK8je+AiGRW8C9+4yPT1Yjg2gYrNx5nP4ONYmLS1+Q1fmglFemJx2mzxi2ltd4
QbWhgfXO2rFQvoy4xJMIjG/neqO9ytVlNROML+emvUaSe5oLYiy8AAfABoxTnUZHlhPchRJ5bEax
iIyoKOpVnh8DjqywfN66IUwfdRGFAduV48SZxgnQonEBDJ/JSWjXNq8TaH/359FcJVXLWK0CaBh7
SubrujZcSfKMfiLosLicfeBhC/7rS7JL+D4YMNwfB772tbchMa+gXb34emi8LPMcCyI2Nrh6HnSH
PFDB9y4QF2GwSc7XPhvV1Y09tjTt5y7kV/NgOJWjR+L9bbncxbSsS4lKaGkkwOGuqnISxgnXHvIW
OkkvUfM+XAi5DRU07S7Rbljdfa+YKDpsy4M8dPwfmW+1iDM8b8c8aLIs1BSrTgnR3npYlNVEP/P8
quzHkKhli6b8sDYfnvmq0jBvqApEKSIk4zAsPihcoA7G0euYOsPPt5Jl2El3mnzGOgEQXks64WKU
ruS3u+Ue8gllBMcK0NflPUDGFCWQc+/HoPWlXMswVkzaLnpc8u1KpsIP8g1dvA4R4YlPO0eGaVlz
7lSUxT1AC9ZX5dWL7aJmtsCcoNZVB4KuXzgqR2i2Kf9glsGoYSNNtOkjYv/fnXwKbKByN8fPVBe0
62StIkrYVl95gFbp2FOd9UMM40VGZOCjX0FyyjoKPCI6Xt9IOve11onyGshAurcHUS4TYdENiGHR
iIzuLrzLhzNWQ6fc3xZ5Wrnp15TbA5DV0pNn7TX9JBafBbTFXvj/2RzgtBonXVpYrepuvQcBMKHO
UXVN7I/CSPpyI+6Gk+wMvnfI4M7wixCToLHqpy9Y+D7oQHQPLZ9JOW33Fw8imDY9qAP1TnO23SGe
xrraehD8O1WAITlDBnwIQg+SyOlgkqr+hlAyCB00VMVvpGEJo8qybEB/jJUvxMQ9ydAJdTGv9FgW
Rid8uk8ycgl+3aDomP8UBLExRCg1MQD9KMidK5chBtjo79rlQAdTe5ia2EDR+5sjMRHrDxAiCX8F
nRbikZW2xKj7XD2cRvuK2Hl0RpkRV+Hk1tNXbZd144sIYL9y7cb0Xz0rD8ODuqqHcycPSH/zU6A4
ZeWWJW4tehgqyTNd2Z3cogw7tBZtGndwnT5MhAoRYmEUWEcMiVe7pLIgj7meXXe+XLjLZbvRRb7A
AQMOMbbnMWVSR8QTy3q4Q77HWcme9bI8pc678LD0RjBSddO5ZrkponPHY64Xfy5aQD/NjVyxlOBk
fsb9ZvDolizjgqmeh2v272eOBWhiQCFgbB0KU35cSfKt1DoOIfJL3kTDv/FDKc0P9OAzu0+wlLqz
i+6xmrv9a56D7S5wyeO9cioa/nYryM3O5GDv/x54DewZD1r3f/Y65VsPox25gB6sWC29qtrtN55Z
SSv7C7z1jdS7Nib+bTbPJXzF0ZQ9Hlp97lgG8mydglwDtbwXPHOSPt7kUQHuUF+G25Yt4Gfjq7VF
SeCDHAPd7RjMXYQxDhcsQOusHIGdUPoo+EQPljiKce61bZrKpMhtEffc2Jy5zC9gI7pLHU62KOqJ
Wl9FKH9aBascd/F9ljutM7cZCOJwd5bL5mIwzUrux9WFRuRCr59GIcSpR/nWoaVSi4Qx2Wea9pz3
xONr7e/Oa4x4rqjHF9pGvwyEvoBeV+QThkdOwgbsTFtt8erOXxpyzWU4b7n5hNd6O0KrdtKY8HJv
63YWQoxhOZlWsxH9XvuHNVa1T3jVetnYL2TxIE4AUZZ1IsTmtWXZ0MuINa57803C8XXOx/sDnmPv
b4g6ku5Y78T1zUUIV1wrPLjPFsj5aqhPVj2iMeTRn4djlHVcL1Rm/IIDlLNG3+zVd8O04XXAyS+p
5isWZDzOFGtNOdCuVGHmfRAekMBgDUjh6WebYPJ0BaegscHRpNHruWj4pYEPma8TE8rAOvbYSVtf
kLpa6dOslRcoU+MJLaanHAlbhvHPATYd9AvqpVrQjKzbC9Ut3goJsuWilgFHtpCs7O6wdQcOL3F/
fSHFNQfd41kzxrsBTc+BwtqQ51r8PDGThrW8oMNbz5EkTBFVyc4KOMt3XmMUoGdN3G+Y5uYZxjL0
Zmq1/Y5+K8bAdRcNJFZRKYe5q2bJ/P2o5YWV8wSOiZdkDZIOBau1a6S8tvMyQl9ryKTaXoIQkkIj
jsyacACcVifuxFPV/ZUzcI2eKuCLqswBXV4uT6qXIUDMeSH39GG7XtLTZCqrmLSAyAqjdXzg8Jw2
SuoCUzuaIAi2dq4z4Dbf67ElnvEMKLDNxXGS7Yv2/UEpHllI5d4sup3Hms5jO0KOM24ojASPnj1f
3gIyF8O7YQs8TW2E3VWqAx7v/MPs1qFd4XaDxlMSJlLk/ZWZ2nw537+E75CYmQDhf9TKk2OfVsxu
Qt1s58apbsF9CAslr85l2GEDkGcdxILT+CpgLL9Ti6gBRNFocFZ+jvF1966Xi40fKvETgwBFh/FP
SHK9W4EpRa8Z21BpyAcHKDBZX39MGus4KQciJkZ/nMdZx3X7AT7YrYAbK7A+qk9ZNNVYKe6cRyPU
q4GDasArJg82X5V/q2luGw2965YccsuoGfJ8mC25zwCZIYwEPk2hp2DGhlk7ooJS8Xf/yRplXdpc
VdY+17oPRrspIeVZo66CiLPs0ZSdndZljpWRUOjFUDgcRpNkJ4PGhXQMeWzqKsObgT4pQfWsjim/
crRrZfBQpsmmhxhLSyIQAsKTEOSOMz6D+Q/qO90mYAZJWpj8jHvPM/TrrxMEa+k8S4UrQbnFrhtu
BOIvAiKPwn+Hpsi/G3USigava7idw2nKumRYeeoobB73Xl4eJNuKFnFG9jaDYftsA2Fq/zYAFq4A
aVWzrHZ0xlF7n9srywI/27Mm0sKM+JM2nBox+DfCTFqovizEoSPY1QFrcx0+ePLVwWAN6QuG+x/C
I//n7S6cd2plq905paAVmQxAUP5237H8AD3rwlEgGb9zHvFH+vQROywwdoj+W0BRAhXTXv9s84T+
Y1ZUPUUejGQDxlTatjsNCMr8WaRL8knKzdqANNIfVuykFFQnzVkD4kxSP/s7NwxReeiIOsUxH3l6
hsgnWdOHTxNW2BwpcDqyiqpDEtUQSPEs8BL3iU7kOfOKgtyU2EmnECSeClzj08Kg6rISJzDceFH0
7AFdxK6dmYb8la0S3lzFvCJ0q/HUsczCFgW/8Nd98pO2BkdlSdXle5opHJMEw6aeAKEc8OQYaK+V
JRuj/Cf65s6oQxFFw9fimh9MFkup5hGDcoudMs7Dg1R7I2atykG0x70aEyLNqhVdE1IU90uIeofP
Awq+0LOnrE6vjT6xYBu2PI+q7jlsWvKIwFofshs9iaXXGWIzCzRqy8wQYAuisk+/Y87V9pv2HUX5
iH7SVQu8UJxsPA1D2JLKUrH/qV0msivJsIE8CJkpnYHp2yUuSaQhSxBNjFrTaJhI4OH0WufzprBw
AzmVKafttW0oerk5p6jiM8vznalJSjQr+eid2PEVGUaw6XwXZsvrMQ4Q3mXKxvLlGKr3JMf8d3VB
Te8GKrtmrqg1EXgoMNNzf1fGEooGMfI/F1ErfC8y34bJOfsMeoDfrNxcPHIIkYnxgeQZrM0DPoI7
4IGqGsXtr5Nkxxlcz1jyW5HFSA7VYLqtDif+Ea2SyGP2iXDGA1fTohx7VT2hkzaQgrCuRTxfIm2A
rcyK1vEwDRycsOxLSfIEkO6LrNwwYngJhQ1b9gjBNbKK+MOEYaHIqH1mlEg+4948RkX6psZednmm
tBRv8sOj07261quPPhCQgxHq8YtO7BPUCukeN6ngW7cIlIQAjodVZqCkMRkC6095MDf+y4ox7okL
VASZoppFjPJNT/gkM3wDl6ze3vMrdJWmWnZZbIpZ4YNKLkgMDXF+OgGr2ROVJJAXKLVRMUS6V8wv
jX73ayQW4LELmvVnbQzhyZ6ffdv9sHrfi3b1eEKwiPoS8xYnwDGNpj1AHypfZGFjShziXm9BE/lY
sSkhrto0PBFylIRwvCCXvLbwaYkmgRjqQHGc0RASqEhj/qDcvvStT44Bl5N//9I+1tmNSJPEn7mu
KMdPvqKdEWtQ2/s2PN1nRHKJKLEpV/1CiIOFMEKBhSupXaDhyIUzS0mjrv3ht5+ywKJz9Ru5C7Fc
MKKUtg5kPIgRV0gFm7Xg2uuQVc4nqu0Pf7tEsJbTjQ1J30XNBmigRmflhADZdRYUIAuei0z/KZ6s
4px2vjW+KBvxkQr7VNSsZ25/5vE2Tuslki2KwOKhBYlg/BgpbZXQWxg3CUpCmXVbJnF4qTUnG2vu
ZxW1SG4TPQJkm9cj6/GSHRuCRDzOiaNYkPTLirphYJWD1erh1MutUlcZ+ZfkM5I+w0CLlIXbBwCM
1BM7g9B5IN1oDdf0BX1/0zSjMXXbe5o/Q09wbEVtsU/EyQw8b9EdxCY9eRdjmji+ksdCWKjMkYGu
Xvvgv23D/vX/FY5Ju79EyMhd2VeSUuAbPam20OkVRgbN3YgTFYr9T1cYf7caelDEq9HN4G3AbRcp
ri6C8HFPSBWKLVjjUkl7lNcjaP3h81X3GtGPnFoP8AorJIcryZgQooUKTiBvggS5yt8VGLgnCZP3
s9E4jp+UjtbZKoS4sTDlE6gW20JPu0NRdUjodWYUJtghAbMrz8X/8Rlu0ZO+TOcL/Shrpi9vW/Ym
C6ZebX9ZjyIxFnJT2Ezua7Qw4gauYTB7MforbIaFn0IafdrFv29Idm/GkrQ1vftZR3SMM20fbnsj
h8gw3cquBGzftfLWPckc7v/8r5ih3qTaSGPLxib0ZW7OgkR59o3bk4ZVXxgBwHFq1VZ/7FobV7uI
DnZ3ieQC4wtKduqqL6V+Fgk99U+0DW+GHui0sM/bqbli+AIre3QZrOfnUOhK1Zy/eJZ266ctKoGr
PO3Ix7SFa+g7T7YQdicrCJtNWBwAHkQkQ4oHrmTdfEWFNv1CTkQSGtmJcSMwMhKOtCw61wNNy34U
xb/Tbb1cjjHbdSHXv14rbbtSDIZrzODH/L2Q6gKfp8RrtegoUYJK1XgGOrVKHWSx/dVRusSk94t5
OB9dw4pKthRowHHzc/bxvNL3z+we6cf03KA2Ol2nB85qJ0nr1AXZtp6BNNVGDPcMKigigSXmEYIB
sqlJ1Accwdp4d8ij3zQS7oN4gRWch3A8IfVJULzQPheRydgrk3uCS/bM+XKx5y/bdJljWWFRJa/I
JIpwxa5GM7bKGS+lI5azjEGtW4buDB7Ov+OQDOUceqcAj2qzvf6vZiPYy3o4TgNYf1Gmoc3Sf+2f
y0I+RcP7iogb/4Zwt8IOWybSZBzFsyu3J7yt+YlM/XZk5eFddTNonfFG5lQgQ8EJIcy00O4rExEN
fnTKP4Y4N36+toIfCmC0dpre2xjrXO5vCYiy42OXS4pJa6mIYg/9zLftKWmhI3qr30f8Lu7GsPF1
7LmR9WSeuJnvycTL/c0UDbverQJbaBucvEbacuECHauLIgZbVOz3lw6U6igx6X095Ud/+s0VeSEL
o6NDNubO0IhXFU/G5n/hJkFMUkTgIvwkGk4/n1g3RO5XvprST1YLTdpk8WDiuPK/lRP6sMu2l7N3
kdPm5NnWcpijyqAYl/CySMwhkMeGw3dYa6oDy5fP8wFwvios5dgHIG0GY2mwD4jA0GLbYkn+P0wW
cIAS6kyMyqOiXoniFePqVIhYLXlvuBnwBbaWGqXHvR0Gat0j4OwdUwKJofQIe7hYF3O6gNBoxb+B
SnQLatykKbgohzvy01N3Q5qoR44llmQ21potGD1A4TLqcySd/oH1HgSw50EG8/0p4M86g5V8JTCl
2FJZcnv88O4bphY+GcR435/56LICwF/geBqo2ZES9uEtbglgUDEvkiKvzWH7g+gsn3+WCTb7KnWy
iiAWJHSAkMHCd0vypr5bkoNiiFitRm/PvbGGy3Wl3WVUHC+fQpkjOlUDMJ/lYkCbLmxCUKxF/8em
AzWYNBXv72cyt0VecWMtMcHciPOPF2HRQsi1+W9kF7yfd9PO4q+U3itkO6QMTVvThjvnjDc9+ijX
PeRrRAqxhKekd7zkucKOtyH04utlBFqlSQUgPGTWQbe0+6TtZ89FtMcQeWozT41rOZE3m6d64Qqa
xoXgEpb67uzzPgw8BN0ReLabmUsc777IrDyEhsJZ1qwS3eG4YLil9Gwv4HX+4NjW+rMpfp5+KnnZ
93QxFnqSHvG3FMJVMDjRgvFDkh5e0u67owaAYhvkUOpP6OpdPNcZ16XsW5hh9XvY8QVnbsj/eL+U
L5AVMV5yzc6n5bHFaVne1DrQxIUeugySMWiga7Q6w/YhqnglH4pKnGAzMPcjn1DixPyj4dKb8C6B
rXdoaGCDz16uEbYlQheMaIon7OO8TnZxTkBQMUMP4MNT0ZFSFno/2/xWPP/F4BxVZniDLaC6jB8R
EhaUnur6Y54r+5hepvE370ctBlX4boHZ4n3nhleo9FaCxxGnCnKSCm0nJHUaYSrBIUjlfX7Mp/2k
yFZ8TX4YQx/Lp+4tctYpgGBcO/SibmFLXjOS/fTt1YJa3E6wEtXVvRu9GVdEvLcULjZtf3t8lzm3
0BONn5rnAIHVDLhcA923F+XN+/zfLVBRO78AytP3mxMWdoFfhSmavHAQbk4wihEbkMrYwzSjlXZZ
G1RdMrWCHIArFNmzYSHobVXH5rWD6QwpjY42vxOgeN2j8FvhgOIPdvFx6gUYr+RCgtGnEQVIzYOK
Ux1d9KwVd/Zbap+F9zUn8NL3iUUlNNBs7Z1pKjXds5iOEiTqbxPUevARuMxKmFVbxi/2BipD+uGC
NQLPOnMkaxskvwIa1HoKqAs+Jv2PmTmvg7TookEI4IWybPPPZ9/MkEvyD4p+/cFCVb0paQesbMqW
h7vsRd+4MeeDfns02ZnuwJ1R9Ary/2o68VYSO1SKVAQ4zBJWqUh3VbbrPbXD1rRqYYnOQChGQkqr
r5QtfSFeGpTaioYXlmFZNU0wQBzd5x5FxJsF6KY2O8SCz+Yi3BQhRkz/LXIcNtmvRJ0n2oSrd5Om
t3Sh6qeDSrFqmFmJRzv4NLN9xQgYUap7FURX2h6/MH7oNFvfhpbw9p37r+/jSynaBq4rkvPwhNfo
fpRN5MvVUygdrnzulRnMrMadUdEKX0lHK0fueOsTmEMpX7xKoDMR4BajM6ZtpwP28h/5RVct6tJW
m69gT/ftmJONNFNA/QJMfvcT2I5iY+f/F8q4A3wAs5/t+9ETWT05vOb5oq9s15v5PBeGWv9zNOen
Z/8aruUoTl0dvYyw8JzF/T+IGASROko13P2e02HGe2ZKeEWBizQCroGtUuHyHJ/Y8pxCr0/UY2rO
aoUIcMjq32anLhLWaSPN2xCEshJDjmJ38niDy+dkL6maqfPyflYQIYPaOfyP/MMjPplN9muB8SE9
JkA5eYmr+K+rRjZuNS4YRqWJbdJmshsed6hnJ9Ir1tpT0w1s/s/HJK5FltqaaeM7LDV39Xbx/0hJ
sw8IqMMPQh38+1Ki7kq4sZ6CqkIyOmKlWEdJObI9BzEmCtzSMRa46L77yLmBdDbMwH4NHVLbkVoZ
4a0Fe4F8aIiuliLGQTMf3YPDN3fHKfCk8QS5L3xCBEmiy/oVP0MA0XWa5QquCYcXWe9wBdo1x4YT
u7zJZ48qclsOnGIByGT0AEOgWhcAjC8UXd+zgUS5vhMtBXb/QiT7OEHaMw8kze3/cZk7H8q3EnSx
vSIqwJVA94l02fqMDuj9q1xJKFhOzoD1+t3OELvyva5Rg3cVBtiW3t21Kpd0+GT0HKougv+W7Ng3
4eFiiVCzJ8zYMCD+aIMvkAjnX4TaAsfYE0XH3yQ1/u5OlrqcaRo78yeh8TWOEXcQRmGBjWGI5DNN
nuEPIBNmZ/q6Bdt3ewPuwg1u3pmCaCH749/VTL28IAczOO6p4rC7OkRJ5W8AiXby+/7Hb9QKPl+t
W6beIyoiNCcMg01KgfG9FCLasXR2c+QEHmVkTsBay+G3m4wZu7JYDLI8LFst3XuBTXwZQmaYizvu
m/nE70GtgcLFXt/ayL7ivb88S3nPpR4yuzj7EBbptEQcuvMrauTO/XKmFd6vTZdk0OPL4cJSgykP
gGnS5dH6cToX6AAqsLv5/R9+zfyC3XyKE+tbwszbMs7pwe0dK/FB/eV2ew1gBpy5BCT3EErpw5cM
ik//p4LaM7BTyRZ9g+YIY9ICNKIWntiow8A0z0xBMbIGLD/ZyvF+i94F2e/WLfm3pak58rMdQXrT
ZMpPidRRClPozQz1atSk33fXyuHy/3Q1wX9hkBHAM4iFl/ytvVou6uorfkq4hJZtDujbNG+ctUOX
0jWf9itJuc5IO4dG1Wm2CxcXPs8IZxNcT82c4fQByPOe5eyU5cfP/XbVHPdgG8Wc2GK3ssIT5FHE
gtbERTddpX0ud19Cy+ryUfIjz/H1ousUBMpKuAq5VQBGEzWNwKMPIjJtUcwZm5jZsfeUrWdy52LB
eCPgxIC5mr/4uEBZ90Fa61gIsoNga43J/304g4m6sX8eGPypDZgYZObSvcHhUAuyY/3tzSQYikQT
+rFn+sgHfTqf41HNNplRoPsFAOQ+1MpB7xDO3brVV1Rif5PNn05ZqKFrkgAbymf00Ahm0XFznf1k
KIyD89BtofyqqJ3RQndTeliB1dCwMWcnDxrV8UZJAyoAgOGsRwGTXIYvnwGri4KJbyvUwLuK6rrr
4YDJrbtKtE9O13+ggMMdakd8Ch+J/FmyMSUIKsHIwWXnqXmYoBsJkqPqvzt14PdrhUiFJppXcOK/
5zXZQSnJVEqK8eoich88mQJ4yyM18hfaPy+CRR/mL89hjkLm9GC60XXnpEq17PPQxvBM7rgR4B4v
9t9fyZnN7sIybrTdbAMlv6IARaeC8hFkJqSQrtLfDfH4j9lELwCjtSkNbyHXROELpbsZ4oPUJpt4
2Jf+JloXlLKFGM8QemCxyvjflxf9iMU0CqAYzm91H97BU/QHKfp5HsLZC3RSL0k8EjSZguk+JWRf
7herTSLj556vvC5iv+Y1k+FNJMDS0SCM1pAj2IQ8M5MoR0/kRb/MDX8JE5cYInZ2xvaIFHmxJhjg
t4K+On/wLL2PxLxnT3OY+bTTdu0p+4JGbVwEymdG/sApOKDu9M7jFM+54yhRIv91gV/G7XHpHJ/n
VV+BC0l5ZqisuAPwGE/Juqx0qmmao3ngvNWhqdaScDDRafUeOHrFXfYhCfEawa78jQ2sdJhoy9rw
fEvf3rn9PbyESIap5OEwF/hmMUlB14+WhOM/W2wvPZkRNOformQElwNw7OHtxd90hDp9Ca0QtOQG
rMUhu5N90EvzS+8QX1Qm+pl3IK8POXLgYEqOyBQqgTsO7HdmtP23V7YcmVIc1Wd6z+zBG2qP+EAU
2CHY/mWmI8VvvjcBbWup6yKX9aWxBayWCNbKHj1m1Y3qyX6aZVKPIbq+E1h5KikzDJr9FtTgLh0o
HmiOsFcoLnFbXNQ3wG9q39NWbMrC4Ae5sYCOYD3ah62s+mujr6BBQaDt1IlWLo7n5nQJtoxDbnII
fLqMM8r5qOQ6WJpzU4uklXyiRPnQfrNaEXyZshdsmLLm7YDJrwYWusRIEYPIrYKKrCm/yMojuJdd
xexLQJjZqSPyxIq12Fxog1kdnubZ1JYjYvro7At22yKDKvNVk1qipMv841K+MWu+6JPK2P7+YygH
PkQQSR3Tvhzo5FFHm2wdUVV84XXbCrNt465Y/0qgsF2RTAUOlHX6z7/WXvzAHAAVH/EmQkPq5Nwr
4fN7Xq7tgHDNZ0fV6cnPgIGMe12UWIPhJLRC13qb+JGpno7x/CKLq3aZN9Q8F9Hq/F2sq2tN6EqK
ruaADKLv0Eha7zB6srJnTGyaJeZBKsfAp3a+sZbvak4TeiQEDWGIGS9weE+AaUsIi0h1CXKXAaXI
3BHR32ToHEV+FYuPmSho9I7LLqrQBdjhOKIYJ406xrj7s26aTSBV405hR2OsJbLzD/v/LykdRrPc
Ng09lPC2Py5674K4RMwORfNiUX6Yx0zWoAt0F1Qh50XZj5q0pwnxU2CBbWvS9BOxZcmWF5K8NT0T
sRcvau6qJ/fVxAo6y9EqzNCzqM0aqfqi6McgPX1SzA+TJUJG4LPEuQMzzb+FQob3VbMsUMGqpUsC
ZebvUdPNUtpT9MzELZdTsO/DMQ+MKkLkErqmBKzQnMfU47mdG9COmtWKpmaSl4P99vLEz4NyIuAM
6MnV5Xmb7wDrlnRz4zs7V/pq1X0EsQwObzUOp6xJwAEVI2pkPW8V6tkk+h1rOsOPLCowQEuKb9Ik
hybKqpMe9KLxoeqM8pmKs2wpihlxfoCdyLZ88SDaTxtE2MQxA3+PKSe00kY2Swe0+sn2+cYhzBcC
WNk4jh4AHcGgjC6Ao36d+gwtfdnmJYGvPKzGhXgXdeNSEce2l3cV1vqhVR0+V/ozjeqBFlaGAgRh
tcl2d+4atnTaSO9j/lMnih2+WOMqg8RWPzQwUQwG1eZ3T0XTRQGhjOM7JJPYoQt3ogJ8LvtQ3eUz
W0944iyARK9XiHBw0xXe6XJ/8OXC4XHqpE6e3BZqE9AO2YnLECJQmqIuoZHcAfE3WvJ0SApr7Bnc
/J2TayOvPYcFSXFdJshN5Xz1+KvLfNBfCDAlxMNjNA4SZAJuftIEHu9qb57io6LrEoHW02RY1P67
c6kVB/aM8/pFrib+znsVZ7h5NxSSiBewqk0o6dBAw13ifMUqQlonswcDKpnVNWZ5DhkvnBsJuD/n
gJ6Nlhj+TDgil+3O46l6zKmy3N2RQBoUJt00ZcSGPIxywLI1qN2QXWUmc18KrtUDz9L+LXCPnKWg
6TDCAZmt1BUADxvaalsTnnX/ZIlK6H8EjRdsH+LKBmV5wZewTglhhtljYA4EsN1cDLqZyWveIjyr
f7KVG72cvhRuyxzWLDkp5fUIdUrYRq+uTykDZyics8hvBtm06bV2562L7kwAYDv7pZ/zbaBuFMuc
b7qAzu7rgKs7BKiIRncT8vUeouBi5wMPb3xPeRvye5Hf7vr+G8UKgrL+zbbIwqBCZGrEq0NPN4Z2
fPv763+I0sDoUL1MoWOqtKyad2BeOmszl672hgyJ+X4x/SiD5OYjedW/1KZwsdjqkNxRWDpujaNu
wXXaD4u4MKq7pb9e8yRmsdoLmfk0vU96AaVd7+n+d5hFeM6N9+r3s/+VT5kfFrxmjy0wX/jV8P11
KI7CCi4MOOsWve6I1PmA+DOqLXVA5bQsrrXOw1zxn604DKgghafEvmD1xXSCyUMKqxSCsYD2fg1i
isrfDnvjuMGwap4QoBQjuXrqZWLBso/WRHBi4bC33G6Ff9gTf2iIZZ6ieW6QR+aqwTNxK46hIEHv
wNzMcKAwl/CRWf7pIynr7ZqJ+Amn3tv+JFRDaQ5CseWmjSYpUuVmbn1/oXrfpfsXN3h70fcyfPEd
hQJ6Myar5ioxST4Qlhufvm/TRckG+W20TUVb1tpIvnBGblEoXH94WZJMto5W8txvQNy4RozzAqyw
gpVL/wzlg+MnMJZna+v68a79aiQqFcRIx9us/f1MWuM2Og2B2x2Xk77fDfBnmopUCDowJab+KKtt
bR1hVEBCNta4QTpUT3OAo3Tb3NcfdkoE9TRFoEANiw+wwMBjFCh0P1we54CKIRcczGqJGId4Vg8j
CHhqih+25x4icu9G0piZ+rvjsHIY5YPnn5W2eAmlAdBAm4ELxF5zHAuKMDlsdZmCpJjUkWodI0kF
qHX3Ql0JPXgXpWU/uOCB5jXbDE/254uoWXfOg3Cxg74BC2ZYJLfSVF1Vkms02suu0NvYdpkwrHky
RT1khXfYyaIU9+8XPWeOFUd+n4KTehDYvksJE2fAA4QRRgscWmZUpLkSIMip/INeL/FFCcwC34xk
Co6CH0mzEU0ieRBYLUkeZHUHWYpEh4CnbbS8M3ogB3rM/wi7YM5s4sy8tjF2uOs8Tc9ci5sIgQkc
hoNFbOQaE/sWlhHXS8vyDUfaWlnrOlZArROvVtbduYCCH87DoTWXEtgjG033IhFmhqy8cFj+Qky3
Av0pGF/9fI1I1CnKBs/nrU+aafMK5i9xrL1DT0bq6FZojWTmRPrda3vYqcIxPdLZBx5ZUuAnB5G7
s8lOsNwMeqs4c7GDDHdVg4rQOmI4dsKUpFV1eEveuyAsKb56MRPRaEdgga8wGKSmBO5km+3tZ3CX
rUgR0ZIfOopRxwK6zw6T1UcWu3ct7i22JWVeGeNNYGsXLACJkgkXwyzJHGX1jrnvSkAoTAJGXmTf
ZgPvohftlFnJ/Tq/VsRnRdqfolCX2YdjwN0xillpm7Kr1SV7B6TXR2iBvxaQrrVKgXPAGxCM7nLZ
5fLp0hEWuNrIr6oHDXtoSZxCUI0WMDuxK2oM+WWzR5nd627x6pNjfj8ZHFhQZo3FR5olxrbR+7WP
iV8HfniyzgPp9uFp4NKJJEBBdy8uBTvjpo8GrRhGcHatjkeFp5ONFocxg0fCiBKC5piBk88h0D36
HlG9sYAI2WoyOUypRYW9DDC1MZoqBjjuxnG3lUBk2vi0qjfQ9ag7hfKHClGIiyalf92QiTTjE4oR
EJB9xy1ufexKBz9YRL9zR58SvO3DuUJFAtY8svGvaPx3sx+2oS9e4i+SPAJyxqh4uMfuVFSTr6lK
4fEpQPfHmwTgf1jWw1J0tMNO9wW802GHpCLVu9P2rMLktEnmtfrnW4p/H688JJBhsoG75wXlzA05
C4VMlZ7WJ+xSGhhtB8jJENHynFIKT4kDal1rPES2SZnKLMnhyB1P2n54UKs1Mt6pRNrmNBWUPeOm
4VXOdyh75p2J9tVMEzLQt639w7E2tjkf0rXan+oBlrGu7FI6AQf9Oe4qASiKimLQvY5OC3FmGKQ8
+i/QgrN25zeTOARt9KAZE62aKptXUbeFR4K9Y7KD4V1s/E3lIBHAMZJePHmjCFHFteuqS/8m7jIW
NIcyeviGbZiyGuzGZa7GBbuEDoKSWESZRWKuLI0bXJtFacv+DzNdxQjLtHJXFE0uTOhcwHD1XC4a
zRW9xOP7B2/ogzzlNJqy3I+etwcW2wqQ5ix24I4JmjhjA6Ydbqo5N1yLc8qD6KlISu8kTxt52xGd
5lJluiIg4ktUN22qIGKw+zOzvPaZyYpA6BxUIfD7Lr5JLmLirc0nAVR7QhD3CDc4/NJnKY9aqAGF
d4I8Y/Lfva+rwXOVcRcHJbjQAU0IbXsINW47OffNk9z/pWExDW5aA4Uy9qNaamcLvA3MOKq37Ugk
1DrA6L0ssGWDBrPQwGJfzt18d+MFhdMyiNencjHFsoR+cojGnCbKag2gNeYG25dIyzSolIKgwlQi
gvRaXipnTQGgfYYbS1Mx/HtxhaGVuAPvws1Z9XICKJ+XUtxqB2/Z8RFOB/TH0TOsfk5h92RrulSR
sDP2vO+y1yjAx0I1d/EhEXumoAERX5fkLVBV5oOZwujS3rfuSRJUUxC9gKVHKhEGGZv8PwDOpEeZ
XYUM/+HMkYZE7FcEtwjT4sz8s4JNWOhg2pz1TehR7Whtxc3S2vbV7H2aaRIkFOtzjDCN03RKjmMx
tWrw5AAkJLcwBkqeCZSw52mei91nXroDegCyrY9QyA58JgcqGHBx6xqOX+FE0Uz68hdy/o98cj7q
yZzUDqHdIx1GE+wiIlngzgP8/VP2DLlMmK7bsfJatf1HgtjHvsbPF38RQLa9viRjqmWAVG4dQcnK
zaBUsDJzuhXqPpkDixBHHhKQU0XKDz88vMJMsp6LZSk7oIQY5y6sosLjIdr/JDImiTYr/GoF5UI5
SPKXcQtHWjQTqZHlVo5r7zEtBl6H4SaR3rP73PKw31OUSKe6zKrl3Z+UtGqnple3/sW6b7JWGnE0
n+9zoOQ39gehJmoh7kLjfg9sGIsUAGhePkFSsktAd/jp8M40kF8pwITlptIFRXojv6enWKGOMUNv
iH+aIrFw9Ks/hP7MDAlv8KVcw1e1Szkz0inltquYhUFPtJiU5PhNxAKd/eMGq3yYZbHXtATSM3HQ
7kzodI0VeF/G39ochE3ne5Nc1161tHsUFUVP1tNDaKTb2NrzSZAc7J+JWkg2DhIZ4/9UA75VzR4A
1r/JNvWndmmUzUclx2uLSpzPFdPqqJ9zPF6bNnWl89koFE6Q2j5pSfKdfs4xsLlAp0Z9fAGDHL1d
DdGMlHnpiNOchbhzGPCYQYfynG3ZldbQftIGjYB5eUNzbmT3ls1O4xM5p3GtfOMvBPgM+xWMWgze
fdHHeoAD5sNjiERTldQoA786w17gRPTqP4UoAauM3qKXOf9K0rDqpqfkgkhX7M6YNXKla/47DkMU
Rc6pgLDv3Q/UzIuGk0UO1xLCUkploUyyIcYM5+A2ud00Q/DrsAn468ChFLjYEpom546Pu/x49y+s
xE4IvnnNSbxoNYurglU4H2R8UPc7r4DUbk8ts/WVEcg/0vT68vGptb5Q6OKUgxuRVQHkJOQALDoy
UcAgwV+wCBLbf9Jiold6gLZ7/aBzTt2rp8VBQkWDjTyQE0+6AgfJPSwPPTrTfFtoQWK3x4AGRW0C
ZIxi1sDTAPnPVedK9mRxi2ejaXk/oj/Sagwwz6+4rsuID4hGoOIk+TPTtVFociXy8kNh2fW6Iger
1CdZFt3kQNm7ZpjdC0VynVLgJdgnGKVFDq8zIV2Xh/mmvyPb1q76fsnK78TLaE0u7bqmPyhenuib
K/lJOenWOpqaaTzGHXD5Z1FeKWRagxFv/u8MzDKHvZRUHvPihqsKrdFFLU/r6BkqpW+tswvria+d
ikbGA5cczn7KNWWpcrfxFaL6TASxC015NKuSVpz9u7ENhVR5mEtU/muy5V+O+Lz1/2QHfshxbIfP
aaqxFljmVAxFV11vhZII8ff8b2Tc8Cj7XC2KE9KFBgQVodCy7u2ImRn8v8sSGlwu/ZaY4uab2hkJ
2l26EkYu9JjkzBMo9jN9cCp0a7V7jez/70zvC+OiR17bUtYTxr47LfPaujvnkO4hxdKywV0xa4zW
MoJA1kpKLunn16cuzLzbtGJnvO2u9A/fO/qji94P4DKCnMILiyUlj45PHR+sOBCKK/G+mBi08cvH
x5ilMA6/6dBDj60rk+lK2Evx6h75DH0R0r3GgTr3kBvDjh6gPhjcf5GYnHAJawgmNi+lEPzUzjC9
r3QIEiCJmTyc9QznrF5a/4FiPwEHZmQkBa2Uss/X/QY2RDuHH81Xpl0o9MuvdG54geQvGerFfoKH
SM9a22553J7zmV8kd0wkbcAKKJFSE0JAAdLcX61c/PAi5ghz/Z40XwUfoQVdWNtR3Oa9aIQnje5m
DoeZouGh4fNOwUqf77gyodcnykBZr+nlIsefBAWJT3rPI4MK2R4Mee24/DPY2OuNxVlc9D6NJyQW
gm/LUIEB3v031FlUq5QqN91ci3LGhu2G8STyVkDGlVu4uANmWG2wHLu1e712Wx6hA6P9Ju4i9Atj
hHS9ugu54rhqd5IeFmHTogM0ydmVtPr1X0zES1mnwJrxw/jgI/ZqCwRZsJQ1ko5mj/iXF30jtfzA
aiyWDMDFEKtiARQndERCcf9/PB+mu8pwH9r74fdq5/UN6hwi1h0WMu6AwxtIdC7zAIqKZyl7/LiM
lbusKFAWYiuyn2imuDElN7tWAF2eA8/B4xNJdoCNPLZJhbHpAxmXvtm7J3x0UFVHmUxXAIJRBQe9
fDxEeIeLADnfcub8QuJ7ZCe/aJGLdSbXQqZjQAIi9EddCUMQGmOlA36+reCrowvF2hc4aqDk7GaR
ekyxDYB1CQNlnJu+XEy5E7T0gLNP4kTp1KQbO1An1/ucuTFaGB7jZ+UXEd+UVPNS0aaOmp+fdZk9
4sdGSjjlrSy4Zil6iowI2OupR/s3J54jYCjtOXe0FGfjYLALP9ir7Rq03vzRpZY+m0j6yj6kVAPG
tIR6LL+JsNsBawFoRtqNWQ+qQqfxCzZKgeK/vH5PpuP+R3vwS1dk/5h3itcYZuJq6XaPbMPCxHoC
1a0UxfXjJ0mchEVOS43I6wyTwpM4XzKzfIa7fa2+F70Yp/kxnRqjCQgSB98aD6ozd2FP0ujAYV41
CBYUu/Km+XXPw/rTp/6bXEkeT0D0VyuL0H4ElyXKFfB729dNXlbxbH/8osL3VNe4EdtPlTj7YxSt
eIelXNyuXs489epwtTg/rkDD0fzqq0JzfJCmvfMwTNZbhTLxpsqCSySu2yXjtATftSjc+c7mbpVR
iIlC1rrizJMMggEHUzbMFNJi7AHer26E2EVx1Ecw7WKxReICOsAUqFbyU3WS7i0EZOxsRtkNAU9L
kIW+JgwSme0SSaij0KgurXX948aLtNmPFd/GWx018PdJ8f4FEKNB9kfKmX4PyRiJSx3CaM5/r1lo
aSq3lbcioNk213f93w9aNU/LQKXVZHMqF/vNp17dtRz2b/Fm79s/6CEhJuQS//0HrBy4N4vN6Yh+
OS6hPTyXb2+2R1dnqFQg37G2JokYCrSFueqsSFIfFihaWtVV9WbTsYVJNmjkFLefOHOuZQTZpk8f
0q/+htd+/xSw1+c+YJ2iUkto7TqEqQtjnq2/qNucoG/EJ5zsFwFbMQtWcrXvh8GUWzrzAsBf2pY9
hZfSHIBky/0hDzqX+6YZwlnJIXBywN26I7mizHKkXsJ24ut3W5zZ3v05622zpOmBKJFcGTOK5aoY
f0P1q/oPmHtleWmuIf7+6zI3P6CMLiricfw5MSUEakIe0X4c2jUTOssjaDnuVExvg1ulh7ud8GIG
s1WLeA65YSiCMFtkMlGZC3rxM0wkfx/i8SIoIvm4kBjnrmXJaVjqKnlUQs0WZGPfJg9gnPtkuw8/
RMb8Jlj+FNCRKjDjfNSLpCls3RA+A6Oqdl9UTfN6dIqK8MDSVDrxcMUut0u37iWurKfR1E6+PbYo
DvZIn7OimVrERquxGr8CEP7vukQnFq3uyP2yTIpJbyyMwkgQCkTJC1QQssbXj16Lgx31tKcU37Zv
32uFB8APa9qKb2MUS8WQ+0TM+xI/DFOzl7jYZoBDnS8P2eqSJgvtUIh70PkPRKTul8+gKe8HXoVn
2GSgBh7JsOBs4Zs0c1kEVxhCpz0A2A4z+Pv8RFx1a25xidwbSuxrEThYWgnaQ6FnDRTdKfSC8t8L
b4jWc/hmxQqpqSYBxBNILvHJp34cWJxRz7QzeU/sdRrr/MR/BEjiUgdUwVw0bSo6I+mR2vE3z40h
cbRInokfu36KI7T9OZEYeU7HvyHaOWqOaYSrsFEAUqD0L6ZZrQs3+ENW25KbClGokgfveqzCwD5A
uQ6geJUGoiL9NOeXuNBT5pHF/l++JOAUZRuiatIWmcio9j1uLS5zlw5pX3AUJI6TKvHYeofYowy7
/3KG/oL5LFoupCdHGXWyn2CyWFP3ILTsetIhG72CCAPBw2aX1YuWA2sRR6kLQlxjWBLf8mVE0Xcm
TNHSFLIPw0xUuc+lDujSP3Kkt672IqACIAQZW77+ToLY5ZsEvPN2T5lzIwTpge4tibfdtO2jQdpU
/gb83u6+E7GiKFDvlJXwXgjGoEQQq1tlOTUmT+rt54sPqOTChL1ifmHeZheaq5lzsIo5pytqwOSL
SI8TNhh5BLZlp5+I1kM0pqir6KDETGiQBchWSRdG4xssjNy5t1yMkckurn4hYH3fx3GLCQTLaDkb
zH9vJwg4QrTfY5SM5jRZ17hHhKsWoD8nG8jvTt0hRtRmGVUU76ONz3L7uOQg8aacB3CgR7yb/nRZ
D/6TZphqh3yrWEYnO2msfWmL6YNbgPK1ssZRjNlk1uMTmZV7h4eolMoCYLMJGo2xnAkVVIEDx2yA
0toMg8Q3Y+WOkThg1euvSbsaFLA2DIPVWeu1/oQ7pU6h8sF6GsA2/ZkvVe7vFHxSkXPwOr9XT/Y3
CZH4KV58fpOnFi1LhC7USTuTG/t/oS2lWDobV1gknCJQAppmNbyQdX8iEBuXgL6VdzLM7h8p91TK
C0hfnsNs0Q+5HqnVQuP19hvZlzjtVgDNNpS0Edufqx9dnHxz7vnQRr93a7OPk3UTwZ+gMR1LnqC4
CaQwIaoisn11zXL9ZnUfqQm/CiIxFeSLsg3oqho6R7KHCxEp2reVSVIjlcqTCc0+X3Cb+vyTb2jc
JmZYxd2NuJ6cI/5M5neT0hAu5ny3OFZt6s1QC9S+829wQhDN4+ixmchxKEBWjnFjYJCYlqmy7pSw
MUNFO5Q8Y3kcs9uAH1G4rACoIb4QCTXLm8t5uwSZ4/GdGAMmte1c4i/1sBzA6ULFlkDsYgBm+391
kPhiGO8K+nPWB9zca/IOhiTm9JxEWeChMZbWvre2tXkFBAiQUCS2liLfeGiGtMzIzR7GrPLVkFcI
La9Wn36gfbgTFdGafhJKBerwsTwwGKohFX8hbD3bL4tkoP0BU/3IEmzhWHI4qvbHk9VUfDF8MMui
qt5tJv6PxV9w+Z0/ERFsAX8n7Zar4vqNp0vTo/LX1psg2ll1KCl2GwGMr3u43JCj8R8Qa+/KkFn2
c1edZOHuXD8GZFnMlIEd/ZAPa+VnEHGzkHSrFFWeWlWoPthzScUb6lH0ONAVIfZO+cNttAXSSd9A
V1q0Dk+CnBk+f5S5PLvyFBKzZOiYALYmt+IiIqTc2Toh+vXwqkNQGjBVr1K38wkZMSZW0Uag+/eu
Ao2JCblrfx5DhemJZsq4V+wboNrvVahL4kvnDs/jMNTwKLSIQKbxRnlMImLrMLIzIZX39RkR3VaF
+8F5YcuQt3NJ97FQTToVgQ/5Kc/AOr/BA7BppDpiRzeLGpw1khtfFteIXIkbJeawM7MDr197148s
z02y6jGX59dPL963SpwCwjWF2T6wgDN23T31Q9iLIeN2vJUq8Ixlr+uBBek67jj3c84Vj+mToO5C
BXwLrk7DLgx1k2kBn8yiLwbQmeoofF5M2v08pUyu2K5tA0BV5cfqC85kJM7Hukx7PTSL5+qJO0LN
ciybg5heW6uuVJrNkgraaNY7Jeb7gCKJSF4OBlZijLfIGP3WgAWTsIgXNm5qU2VtE+yHWY9/mtkS
apiMYbcFz5LT3/0gSGBsYtK3XVJAs9UcSlQgN7sip6XVEOrASqOluJfnq+K7qPxz9GAkeE7t7JYi
Ssr+hqR4nVhGTkMf7+pjm2VBNko997XvSV9fdynkVamCVrei1au/nrpgD96XKLjnSoJULV9uSbQW
gA0Hpv0RH6C6k+nYTV7TBpbRhoSZXnLl2l37IDrN3ybQronE3KMRI4yOuqSpwC+AZ92D4uB4ZTUl
+LItj/H761486GQZBkqImGDxEgTQfKtCDylcUcf4KJiDQKkwto9av2TUN1NvQYcTuNCpfCPyRdpN
sERkI8qdLI9OvSxfWvx3tGcX72OxPNiKwgx+yryo1jI0DA6tp+VdxHVtbnAV47N5yZU8RqSPpYcI
MLFPOhYS2ewwqe5clv/EfqVUaX8mfGdc9CzKVdV/Zmb9EJXLrsKr6xvNQpudjPV9mbKdxp/EI6Zo
d37F0g8zrJwbhzhhzQy7gNDVrfLvYz9+uc9DuhEKdannXtvA8Zarh1l+xpjaKFrNt0p3n5+vgzrh
oIkH5HQSsBobsYzzZKXucrBn9mmTMBmKlTmpBfVzyLu/LN5zLf+bq50QP1eYQNIyPQcKQlZMZ2ML
W4WhjaK5gY416yG7yrIebfSPNoFOiipLtaHl9QRfOtlnn08aTifow7ifdqmwidQ+3+bvAe5b2lDg
+hqXU5DPkS5kTfOpjKK48AalbrUGFp6TBqq1sZJwS+arPE6cRsFsyxrHnnwXJjJwpVZ0gMHt+rGW
cCcNdrYVWWDZl6NaQ6N1Zgu4ffc5m/6Ko2ndRkCeHXVScIE/BZUiF2tIJrDsnZEGwmbklBSsg54t
TuBQAgNiVldzs3HnNbpFVcRAU7sAOk7m5eEiNIvpjsZ57EgtA/uQaL1z6XmGlAEvnw7XYVq4NG2J
yKpu/njiGdOCuD9wf6AXzycVN+bD6FVxbTWjLGXOCYQdHfbZqVxzJFF8iOOKpdVBNXbUs4DifS8o
/wiMHhtT4VyOuGjozpykEKQReoIKOMzRIZophx8wS8wzdvTp9x0cys10u8NfreCxBr3XhX/Zxqi8
oATTNJkozkm+0777RceTrZd1gI2dh9PtY2it9N6fzOd0KZI8FIz497hIZgHhatcCbjj0Bbi+K9XI
n6sGF0LGLXwm7rV3R1mBROM7qaOiv0lDVYL7iriUTW8BeqRds0KxCbvcGkISRYnx0aiLof8CTrF6
cvo3JC6xwlwJWyICQOQ62wa/kbQwkBAbk4ShI8STN7jcmYqKXpUueL5xVQsAmccr/mh4EpqAfnf6
Ey0KbwHfuwpt47Qhk7UOU8OmIZJYBEynRkIIvovQE1ovbN8MKGKR5FH88NhOR7uIJwrIV4a9FWZw
5qwbkO5P6sBjySrmDOHK0YdgIKQgrv1SDEZQrSisY08IUf9c1GiTgNC6gEBBRTkJxIoF0gRmWigV
IIAOipFd5iJ7BtLid7g6yGu1+3Wsm2eBtlybfFKygVf36mpUEt0KyzJrEup+6S9bmrJ9kKZMixdi
NyBTXHEK5RGjaShSf0+gxeKMaWTAwEwe1bNVzllKKMj6jSPl4Xj1V9TDh+3IGoQnmV3yG5ZReut0
q5hid5h8J8gdjVQTQcyUk0pJdMahkQgjbst8sJ7Y/9IBgTmx0IrpmYbcEBLxrMDI+bxH20n0qCcB
I8frtID/cKjhWVjI8aTnVJnQfc+9pUfy3bJsTx2RU//4yXK9DlOW7uB5CbvxqzO2wernHJa0jolH
8W2tOfzHlAgBm0dsNaqzkJTMreQZXzUv9CBALIQ3q6u77EOat3Ic84aVVZr0amGQqD0LSKtLbdif
DWKMVK0Qtr4hnmyRBdGeZJnMMUYOT7xMYDVM61sMA5HKDG+BTgyXvIK1rW4RUBF2SgjQiroPs3bW
hs8lpzxYS2hIojKFX6O0ea7pLSu0/z1OCwEFdE7kwmMMJERYLDY3Pr+JVpREwOyLrGj/pPjcYnOr
ev2RnJ78EfMI1GnPtiXv3zN6Qu0mbl5KmNIGP+WwQ0U3tFOeF8KcSGGjxi2qcrQKfF6FbB/7Y8TR
k6YlPBMI1uIe0gvG0xbHBKqTNON4WJTJQL5xyVTFhMqxLBOw1JCqk0rduRgA9dP0YTrow+FLpW5j
3hZ6njrs+bM/knOlYPtxXx8ZuweWjuesfQftsuH6YtI2y9BcjapPrMBOkt4cuh1NC8hrEXEgx1bS
x6TjXZA5h1UjXyQEwn2VyrzqEoqrD05SbCZpdHEk3lz9xa5+sOFHx5JdSR9BoU6qtluev6ulNKqp
wMvBAl9WufepbDe2DvuGii9JFJewlcSQGWFRmOg9n4katlNp7yFnjz4roa2OD1GjRNH80yGNS6F0
eCOaZBaP8mOe+wwBxW0fP43F+hPZB+jdq6Y09Zmw67Pxx0VY9EOYCVEdmZJR/bZdrwdYSJG4+k7D
ol4yJgC2E6MjsNrsHO/bkrsf56JP589QhxoGUXYwtp1UIGnPeAHcwprsbwpp6E04v8GWT8yW9did
2Lj+4XMBE0ZLro7/SuIJdqfqoMERW2rUhrYZWy/VNZ6S1X180aTh0ClEl8nbGEe3f3SaNfT2F/0X
B5DV9LUBm9eOjwpWxgaODBxKW7qMYgQhNbHezvY2uvsxosQRK6tmcURSPzA8UBNZe8cZEHX5TStl
ORkcfr9iI4i8dYre7ZMflHgjEksYfhLeiFKI3c7xRfMpEe5FG5iYtTvHKZ/vfR5RShRXPtPaKofD
zKLfaX9iAs1lRjcYmZX95Us7OU/QBn4Ou9PtsWtwm5SeTTvmXPO6KUw+9YblIGqEGxNcmbwj0vl1
Lf/pxrYS0iigQxFkiu7QOvH7/iJKeyHL6d5auP5bdJW6kX8X4mSrvMGVN0dj1PHqsZMT/KC80UcE
20PaHIhzyF02hMibf9CE2Jxn53tZUM9cySOpeKH8iVzA6CiSOpeK7hIaDZN1XY1yeUXBJc3M7J/T
KfuDGj5uIQaNOE2VEV9tcYIprfwbIc+qDjgroXbMV7RyCs6vXcD2OlzA3aPTY7A5Bfim5vaF51Bt
Innkljt3nmzRD/ZxKQVzOGIbUXl59wyTXzkbR7HugJX9pnpJxqV44SbUIH6owUJEmggeCc9V/zoG
oK6cU5bm7ccjR3ZILYZb+U2eiGI89Cb7G25MB3h5ubTM9MASxaocwQc2/Xulu2mJTAor3IKL3Cz4
bnF21nAZwjzO826vvH27LlfmdUE1kFXIyJpX026SLR9j27xLNeVpu9IeQdXdclvYeXZ9SeZEVcdY
dHaI0sod+HZmLIt2/7pREXzb8lcjsshOyfZU2KuZ+IpdtFxTvF92g3kBb/4BgPMqlbiXASaviCpc
PSymyrE/GJtgerAZ1ETpn4S207Oxn9De4ab3r0uXdtSWp+RvwWadfVTe6fGwLGl5JFGfSvkqppAb
ogJjI9sP9MXKvdiAvJUhLnDg+pDOG47I6JcNPRodRzAsCTH0SCtpVNtEfuIRfOQOuo3WvR7TVh8S
ZaP8u+YF6z8XW7rMcUZUrAL3ZMoVYKiDxslH0gz0m4rkKZQVwHBmdcrthbHr2BI1NypoHerpaqZF
9HB4ixwd+MUc15gKCSCoxHK8oyAwuGm7J78hAonkSQhq8miPbXFrZTk62a0IXepaESyoFcyz3H/E
ksAUlWkjwzj8yrat8bYWhLvr3FwsUfayddhwJowvdQKDS6h+Et5XXgN9mvOds4Wjh0u3xERnzDVz
L7REf1MszhijNEWyQwGLgRf8lu0Zu//lQ7eUCE9essa1LT8IjTC4gly5iFBdQvxqlYp15W1WH6Gj
N/6dw63yie7p35Y7p9T9orCHVLqmO+1EPQK1uIUgra0WcIZaelj7DuEDbPQJmt6NDXThjklJ4QCV
GFBDuMqK40UlJ6zaXWNFj1Vy7VG/vi3yFD96w1VIxPCrJvRv80a5wqsof6slNHrttnJk5+kAsaLc
pGs9yiUpR6Ashhor6IuKbwQcu1X9FgDnutlZ+423CwYjrO7N4nV3C2WIyM704PjQR07kgf5fsLKr
xtSdGhuKuhE6ITjizZjMD5IhpQvuPMNsch8h8oIVi3fPaZnYXRrziXPdCT2R3XsnHy6yRjbBXQ8q
lYSCWwk5UDLyOJRpIf8JqMQETR6QBnmsHNGACxwigIoepLeKuG5E/Nr5J1vWeEgLXBvQEOt0DhXS
fAEpuvD1YEZDaOtl38WJsOVMIMVlby2Q1EwNf+KA0LpICdsFme5TKs+tjCMjKu96hxRkFjQE2ovI
S3R2EbWqm3jZLfboJNURJO3Otumw2hacLWOW8dZBZMMAjJx+Wn1Tnlxt2uHkxsjwqyn4svJ4QQLU
MBxhKpRmu4lzir3CBvVDprcaS6VIUmFMGX9FJYIsB4MVV8G6FWZirpSU8gpEDCOSYYujCSWPdsaL
dikcdtLNQ42t6QKxzFfM5KRTnMPu3PHgNsLDAnPVUw4OrvIc8X+r7OQOflcSgR80Ont+ygOjzv9O
iUvZFtok2O/ZJWpSR/PKH3a6BfEMgDw7Abu78q9tomiX3xHBtpo6eSUWAIL4SGB43Ne2rcT+Cvbx
Xovo6V++nCaKp7zFqj1q2sWiApo1QH6Z6QiLfFqMJPz6+k7pEGd8fGgR3ztWebyINQMD8zqtFAM8
kFK+EQm128rzb/+30qKs3KtsrVNyA0UveJVOcXeKKDhsSmA1o4GCYJmN6Zil+lDzIV5ZTZWLWVZH
JtG0MnBvg0BIGj+FjuAMvyG6QMqHDU6DlN98u11lq9dUqvAtjdQBdLl2v0ZDKaoBN0RnwHRHmRKT
WSsKMC7YpPYqOAaKUL1CTFy+kngYcopfoc+0g9+0xOKjfdDfV8/0gNwDslMm5jlr8ayrYANY/eHf
gZ/6FVWZ/DCdn+tValAA9gY3T+MlHFOMxbF8wGHcvMzrnT2c+KlaxMxJ17jB4h7kzNsyFTSnVQy0
4+Weh2kzSOMKYE3gVuYnJJVhA/cXsd2N6cwu+LVxcmDHi2IMpNe0M2rpOrv0DvaAmtfEAOim78l8
XOqlZhOT4pNO64rTc9T1XTCjj51rNX3aK6FOAdyD2973kq8RiO6PJajvtk8cKEelqUWpNk4DhTkJ
BzOfg/lzr9YuJXDIMf3ol4vFelqKDKB81GHWrVGFymDOrUbGALbgNoJKgCBfcoEyfN4r12Z/wZmT
BUVCcgGnLn7wnKQIYTw0HXdmoJF2iPqNz7B7aT/kGtRT6XNboDRAgBqymH5nSOrYfvCAenOnAHP5
dTOAQndqEdYEq+EuMHBRenOxmBx/m4vslOfrNui/oKwTuggq3GNDi/Gj+Pqu3gKVqm8y3BxGJRNf
53wXQaVM79uRFW+9+HqtvE6NDKmAop5ZldYwHdgvCJcO+kJbkOSscCJC2whgc7fdadrdpAXYdotf
I/r0svwMo9KwR7oeZ/cFHKHji4e5Nqy6f/W+WfHt7yH7nn0FWH70T7SZsbCJrIuO1y01F3Fq0hVP
0V37qwv6u/sKgvs51u3go7ltcPR/QwbaUcTne+HCq2J3QEQeDrmACn1UI4VpkiEhUbb3F13Mb/KW
HRTlTcTjFGoVh2Qq+gL3QXQP4R4SJ7jXm1jEl2cdgTpcrcT8GrkUe2ZXlx2Gns4adZo03aB2jSEn
GXwLo1YJKK0QqsxHRG5eye/Mgbs5A+QWX94NF2rczc9ItMQgz57rR3aA11it71bwiFyKaoGxBLH/
JkyrXzVz8GXLTCRw28rf+Rrih9QJye3+JlYdcg4a6LAX3kSnHhFXQJ8Ej+Xpx+LtxQ6tQsnV/v3i
67r/OzBurOgAa3xBzWZjTzb+aH6wxETzHtzxolhDDC+8eeGK7WV7THUfKqgyZTmEwCMw4/DsZy8c
euwX8d5C0Ft1YqEIa6kJrdzrBBY/iMs/GqhhDf4d5bhAv6WcAyQtmZoYAptbMdDCdQBD6Jt6DXMw
UBpf5iiGFiJfBliyBZWXnupWpUkdUY7IAtAQPmovixSGvH6rekzzWJNFXnAkgrbHC1b6oq72FXl0
7U4yagRuN8sybNEF4Q==
`protect end_protected

