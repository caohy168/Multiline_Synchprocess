

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pWwQh5Sb5imbFsod2FYQ19gBUkbq7kcbuGVuhUCKd73kDl6k7crelvDRHXtyJRPMw22xkXjbPzIz
X33wqeXDBw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qlvDXwnzOS4Fo1g4u8RA+BsWxVOD8Z+bOGqzcikzQosfyl5m/1mim79P9mPe818H0J4yWRIMhsGq
SkBmM3RvTIsn55U3R93W2/uBtqpvIcHBR63U1fGJNgSraV/6LFdCt8LLL8fKZW4r5oiZkfO4U5YE
KfGUtKuPkCo/6EP8JJ0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNdncZgmymiqRKQmOI62koZcv6zjffzLZZ80+YQSSyz7uVVOD1K75Gwn8ts08JQX8GJ+18XsXOIJ
5wgXIHXuOhXSGvLE6Bpf8L2vopJSNXBgDYhwBbjejyGrRpq3epX2aGeYw8LYhRZh00cWmiQzHt6Q
zG70IV33CBBjC+K8CbbpeoU4gmC+pHB5ET14rH1UACA7iR3RljVIClqA2H3maHbbT4c4lV4pkiyR
mcCMq/Kfoc4vyQhScJd6GJygiMkqFyIVcQGFcO/OM61G2ZeRbfENBv5mcB60EkoG1606iIUuac63
vvdLNcnOtX6XaJR1g6SsFiVLe5KVPVeRPHIlxQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j3/Re3J8S2ThfaQ+KmY+mx+npY8R34n/NUphpBrwlqzP108B4zAoQD4EVtIfKzJPcZbYDaNt3kn6
DSdJEAbVy2HWHXFArqPJUviYuw/7V3ralGwqlnNYcSD/NsdqWpgyvVnSoTjAl7xArDw+Xy9MlUHv
HX+uNq6/q4LlqThnxXIHYjdusmt+b3hGbDFzw8bJmB9TUV+xSYIPrOxuufK+k5NjwRt+mwu3PJqA
lBMh6GgPmEJIN5ufl/L9VOHBaKUUvgOkAiiL9qWQ8nUyKgKWnclKUwGYJ1Cd82JW0Csv35snxm5k
xybZVNQGOTBqWj0gGfUIDS+eISG57QZ6xdetBQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nxw9k33qrlozjJxW+A1s1+W9L3a9RK+/Jhd5ox/5w7+RfvghiyuPUvPZq2F/QV92LGjHESvCyxzI
VoW1FwgDD8F+QSPa50cxVW2tnYueROnBJAs8LMdPM52AQiQe1SxRU4FLNwokqfY47XnfFykdfpBB
iUx6mUCrzJzcX8EGVBE=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BSmYmqPwzZNRr68JzUI2cwjn+LHBvLUjlcEV6OOge2vDmKTF7k6CMdYSOLfpaYmvbaWzxUMxzQny
p17lTMPE07rneL4WfWK2ZA+NbJqILT0vBOdrsnA9aCEJyzDeYNrIwLDHRiheS6bjCkDBzz0cgC0W
SGguBKjr1f5muQ4HiSH6ui/nNaNEV1+PvVjq65zOTyVXwTWDxZJkptYuFqsUbCbm+Qp90nn1pWZo
nGeZ/iEYdIOLom85lROQWSCYOpSAka4eKeZG4XVGb9dVBiVXv3MMUm6NrylKgmdm9+oxzRDF4DIB
oAHdJXmfttMva4jExm3mnQdvyiuRiloy/hdmUQ==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hVzru9wDfsCzjak3N51oQvaoCUyWk5Qiflud6FedVzGNWDmgvIlZxBdqCRodR3lWoZoHAaPe1xFF
c/NGNLUnX08xvGifqvBja5ANDgsWZBJPF/6NHXavV75AqSr/vARvtV/gUdsws7hgxKPPZ+Tiv2xx
wI19CKKYUGdLlC2Hom5krNiJqCf1t9lDYSQoiWRr3Qt5G5JttCbzp5DxZ/GiDy60D9BXGARrrHqE
23hLRMOyE1f0jqpryFdvZkPHkApRsokWTOEFMsAgjoPwLJK+ETh4RcZljZtuKvB22WvEq4wGUfBp
eKjxiX74zqndZvDf6yTg1Lvj8OJpfTb7nasxGw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kZgsIA1bc/jQam3CAD4KP6OHNax5hxPkVUgLyLb8TdnIoufLv8PDtZLw0AguJzFDIYBJzHyqdk3W
WPQH1ZqZbXnFgBJVgw2WH5++U4o/ef08Chz1ENkfOKLWySE6W5xSgwnWA7nvny7zfOnhDRkQXP+9
ytyk6rWVmL4eMba42IDZba9jEdWgSLiEzWrbl0RZeTYMf9SZQ4iVynlJXD2Eo0Pyw+0Qs2JMrJwm
Edtu4AUdbkqYoOkfx5ezdQOgrMUvuhiLm72TljECoxEAvSHJwilRypbnVUH/dc2dKgR2wnsVuKvM
U//MiIX+A+CFR5rcXcw95YOKxJTzk/yTDmQh6w==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
he3U66LNPhflQOtq/OyhlILAo5z6YP2BLZZdK9PuT7AORUgJOECnYt/k9XKn/uC1tQMsWZJ+ksa/
0przddxio3QOS+n8favlM5GugUgHu+MbRbpeg+YMjYaqztihKF7ggtVWoAXLhC5DA7p5ZOsjVlym
Wvoi5O5tIaY87JCNvTU4d9JPMKwaazgzs3JSzY3T5U5WdoYLGsoSYXq7vx8aYFQZhKW421Xo4Rva
Oc4WHvTumSbNTw+dR7DckqnvggPOui1Uc7YLrs5bTNE0r1PTOaY50EfAETGZZ8l7i6hFaOR2gUXx
F38LDeQr5wd+h84RLqwPn42d4E4/3jauNiT5lQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 237728)
`protect data_block
3sRkzkaDOdyxz5MZ3mHSCZBMdrigo9BUXWMDlpTthyfues3gli96VYGugwvW9kc/CzSiORcb9jtL
ar9mdQos8bcu6LeRn6865q0xla00/gG5KjyqSDeuF6izA8M04hXEcAGyuC3e4Ay7HZzinq+sCpwT
MLCpD/Tdhn05Ldjrfjo9ZBRvotqNWZYXX/57FwWItOiZZZ4ozjDp7RMZfeQortU8fm7YyW8YSIcR
BG0DzCpfl27ySNFWXS/7F3tAQkncN9BVdmGUdUDlD1/IDS6HGG62V3knA/mhDwb8ri50YeuD7sSu
LwKqhJKoSV39Ufntw3si6J/rochbGyXGhc2uzDWlFWB5bDftavNZQNgf24xCzS8IWWm4BbMtzUtU
mZO053PE78N9fmshLch/Cg+VLCUBFNfJL0EV34lZ57dH8M139feKJssWcr+6j9bDKM64tRbqA3ok
ZdUPOioeSy0OBjru6EzOsmhqlXlNICh00lzDkBdu/po6dUzOcDmdBw+vod494TR1eSJsNIiEXcqH
ZuF+CTtLm+qGM8jdSD/8sBSLe38453IM7NiwU6Xd3py4t0nqvCL1akPTk/uY6PlV0h8ggR6FqTlC
LkSL/poXZHNNoQ53/s1v2r7f+SZcnDZ3cDcRhP5P+QJaDOMi/9xXcTqmaGJDx0ZF+3vRd2mNGOD5
wd+FxLpHvXDjeCRoZZwRDd5dGx1/thHY9mnRhTJsYKjWrtIvyDaPky3HdLxfky8INKE8/24J2c0y
E0odepVriVxIbO8o0B+McTz+k1DrVgscZc2Wh8l5tP4cML0xre2CNJtFvNfUxEXf9hCwv6XNIoeb
fhKJ1/eynJoLC5+8IqsGLOCWKgI4sPJ8v2cu2NtYzw3OVpimYW6dt4AkoAG5rXEPPXqOSWuhBpnU
zKqgxVNEYUWfjZ2ITIZnTl1ow6YIJCf81HCF1Yw+H3hKuwyBbgeu1jH9WKvnFjNVGcAaTJ9C26Co
u4B80ffzMLkvJJMzr7pJPnQ74A++8lyQbnoxRVBTG6qKM1daE3cOdoNNO5kNG0poPTblcTaNCh6u
yrBxTtFnIZFOwuRqHDmMZ3fV93TmicDR12HvE7waPJy1v5umocS80F07LmsJOyXl6jGHz2ZW5Q4Q
hfN7zxmQElksEWGN73Ge0o73WRQRrZGelB/7+OJoCbR6TMAfhWd4sOgJLvoQm8z3929kH3Cz//ey
mrvVpARGh8KToWucx+Z1HRiMS/GuUyDz4a5S8ZFTMxoIA++U3kBGvZqkb0sIXu7K/unZVCjUPVda
3M95I5Q80Y1BFVCes0qVo/5IC6EuA63f7aUzrpg3B1k6qe2LL6erAC85cHunV39+CmuZSH5Vh0h6
3L1J7cKn1ctcfaBFT/ttmlGdZv3jViq0ARtz5igGa9fcedgeqnHUaHFvjAiwUuPlwubYGDK/J5oU
rwwuhoyz1JZq+hSNQIOgYpODyEXTuck2B2HFX8CPtSE7bfZGpyTOzpgN2+L7aBYvB69x7pcqsgBA
Xb1cOgsmEfNjYM8jYprthc3PXMuOB2EXXTmBaBwZzGl6mIfHHDea9k0P0wKvoB1myQLEzgKLg6qu
ugwo39Mxe0t/aXrwkNhxIxmOPIYQH//a6V3Uv/CsCMBNoJPTgLRHWDVSdNI3UypyI66k9VZqpUwB
pDxkcmXInzZk/Lqz5bQsc2yCSFLS5BrTuF9goHH869GJONRMLbsjAgz9SeS+8OomRQkIdvnnb+0e
mp2JVd7AQEzuXMLPfqR8AYNeyy38t9w9lV6y6t8vCakT4SM8JFSLvoylSDiwk1P9ecrujCYVLXXi
Fbag2GmUO51wwwD60mEcjPENNHRRdVGtVXFhjtb++oTgLrQ1SDqpsd+vJlF5uNQAF2OVgkzJZ03Z
joWiP25robUVlGZY9PfS7gdOfRBQe/UMIGs/qGPAjuZeeGSj8GDmdID486s/4qwdWkXEmwvXenmd
k4OanHRl2bXb8sdkspNFTMyE+wp5PtztocvnrANUAari8bmHUXSOHcREgr5PSoN5qDbJ0s3c/uzj
mfj7WWg2vMsS5pIlztg7tPGA1PcJcidPdV77xsvSv252s0vPOFUrXBuv0A7KqKVDa9adTRG8VZQN
SL8EpiY0gm8fTy+uwWYOht+ESp8YhhJJwvn1+YCb+MCLDg99HbUNvJ4/HD5+7Gv2halKUdfefk8+
Nk0XGGrtNNklor3EqPYH9tWHbN9XqhU0NS6XRefyxQVhraFwCnSD31nEbpTevwGaVHABfIqb40Ls
jF7q1xIj/8rLJnD27Lzv5GBkX3vIgle6+TaFLY97xvHhkKrgcvbKCycBvjLyc+pp6dLU5/oUWVa5
LMhn70HowR2o34+oFtCFeDdDOxbfHEQsBNpO4IO3q3o0XBttis36fuGLgC1Gg3ZElJo9qNsXpDMi
d+fvGgTvvX/xbzIexaJ4vCsdHPiLgT5YLD2J90RWkhRzuUIH1843tLFE0zN3y1BAjf9P7UXt4ety
4Ahc6TNk0fK5YlbbEoO3H3CltPh7cE2B3A9xW63kXiSQrEliqesGEbeI2nl9ik1IVyGPfY0XxkgA
HgOamWO8W8Fj2A5qiJPlhjsrvOez0HCpYVCR9uj1brbkSswiiY7n8k6lkyhb7qna2w4HIEQSZDu2
vTb9l+/sMltuNlBDS/YnFjZ1IHTiy6sY3naAuYrx8/CBCEefWwQMoM+W7r91Lfp4Nh9mI/XTaiZc
cwCYX9+q5NQr+XerFFuA1js1yQGTVKXfCfkLhTZaqudlWgainU7RxgCPy4w2LAg5mephTAdJiYNi
b4oOsrHTG5jwn2aj4+v5zbBYHNgE9gy4aLsu0K42f9JxcFU6AxqXis9BXNMnOMueNbigXPjkdEDl
Bd/LGhVp0tKXIH2qt9ON/1j7FZ+kIr4pYoN9qeltc3K/9ts09Z7ptNYuK+a43FBzbjOvzPkKyykC
MZMIn6zCQkesdjJgsnb11MjfNgAo1JhfLQWKS8Vk7BLAyCb2DM5jji4mEBDh23SJe7Al5VGUxRaj
YL18l5wIHJ+dZGh1mH7uw638ROuh8ImBOXjmfDXca0dXK+nfZkwBVdw4jiuVU+uyPgm2MsaZbqMc
R7U3pBKFPsy7li+r8MX3TNyKgx5PSORTnwbnt9lbIwrLi4r428dugZoGSfL0OfQyqwV0yTHallyZ
dYbvt7eRB+1r7RejP9Y6STWqV20KYTsSP6b2LoyBIvUqtKAd1XDfhhJyUPK+3fbzFFBdXKLXqiy+
LwGZ+e3pW9teG/WVvxbLL5CfXCD7XEKDJIA2Ubc5CtQGCWP5TT7O+BuzrRWp5QxSgi79ArCCdSff
P18qs2qqy4o2Jpvlw8Evtyra7fxomUx44ePgRfp1nVPOqS6xZq50MKu9V+cWd4lShjnDWJgj8t+W
jDpJj5kvt83aivgQW/P71+fC4KOa5AtTwVoE8EaFz53LdaKgPj1D6i+lEfM5HZjhsHmqMnj3LJVp
ds6jR0mPmMldel1TaCcINQljPlkOFILSzPVLO4KF/CKHtB0hnxlzpGuatfj5U2a+LCSn6N1MlLUl
SPHOpSlaIew0imIJH6MFB4KLd1z82i/i1m6GnfvAhTy4scOHD2gzCFnpdq/22wB+2Bj3x8AEhRVY
+7ik2SRMtatFHnWl8pSd/vjcElrNyGZ2eQ6ChKzekkdQCQGbccHQVT61YaKuttom8TfacTldeZK2
Sadm6bA0MqToErnBjmzFlgzUlzERxM/Ee4yt9zl7X/yFXOsku7HzM8Ko6a/oP8mdDHw9Er1HbEl0
L9gHwQW0rdJvZNUOHBXdnrfdHRUUjqvcw66od5VE6eYzpOkMKs4gtR1FUs/eaqfJ35cHQpGU44K7
uZgHU4wmBgr1cifp7l7nBvkCLwFvhYLokqss+8ZUcb1JR2f2LRRWEhiup2SXiBdUMhu5PgJWjh2K
Y3ipGsBVHTHMxF418IDrDYVQv2i/h6DlpPR6rlp1WfiR2MR16p3WLMHypfDRHZgj1grNMGRgGaEJ
iKkA3QXZiRbyOyjiCYpFKqwmQGkjQul61LULgSEcNA4YPy3Fy4Wu8EBAD1RL6bgKN1PlR9Q4Rb0l
1LoSG4qeVEll7neAnXBEjjIjNlfaZiKHqxy9WndWpGr+dz4cLVvsga6jBk0+p/aDj5LXvwVATYeg
EefBAVtXz29CV7we1axVSi0g0tDi9acU+/BpyRQhBvrHTYp+46lzBdptp8svdolHiWTKQchEz5H2
eB+6zvT4qZEVQ1Zu0/QCu5Kbh+9KlpkU3JYLuNCQ7+iETmk3oJm1q8GB3zHI1Sj2cOMev059dYvR
rguUJdCsbLVBj8OcWYgydaEJPNKtBW8b99Q/5S5U15guW8IordZyXd5uOGyEws2CQZpTk1Xa7MmV
N8oVoHQJUjUgp/mP6lTNdscepgIfA7qwg6aA41YrKb2Z8t3I7/ujZWILNDx1JepYwVb8DZzvkLWP
e1c6hMlfxSVT3CB02tj2UdtRZjYuopjVebLPTmaDe6+urdqUhj+KaCTJ72X19cF4z+HT6wpDpPqG
Xc3Gu8LVdNlyo3g4fAQDHKHDJpEGgLCqCEO5zwQGOyfpZEIM2KTcyWiFqMB07lgw20xkdOzrwHU4
KWqoSDp5M2RQ+eBHGHFIL+K37+dAHqF6x+5e5iUzrvVAesdnE2TJDHNPUZMGdl1UdP9kY/+4D3BI
LtH31/CUtorZcGqJ8hbGufAlYO0SiYZIvqV1qEGmCc7KP9CIytHqhdPqpzadGsrIeC6CVm/69U2O
NCsfQo8/Czvpjg+NBe0lxXmJjN1OHYBfqCg8O3djkjtOKO76RV8WjUang3Y5UwOq+CR6G/qV8hew
jGPEVfEEanbjcNIVLRDi/Ip9GGhKmGPc/z996DbESkcobzrZjPG7ZG6s/bygOqZDDoevBlUjqR7P
JullCFMMaVrlS9eH5TGlxzFCFMlkkmagv83NJQyBrNGCP/K4aZ3abwsB4woKdZG2HJNhhDPOu8DV
lhrmhKVQ6/S8AH6IGIoZfb/8UQQyj/Qx6eT5kLG+qPRX8WqxejD2HYtlkm6tfo5tniQtpXOVu+/g
Ig/83O6GC5anw3UBko4qQMBe6LUN3zTD2k+ocp4WzRAfkfN5sx86bFu5aGLbK62NPelUwXxOPoUy
JbuF8rS8xwUcTINyRwpKT1YmL+nzrrURt8Es8IrVM7F+LrPryqUuPTvDeEHOGUvATRt8amv0lSje
u/F4ebLhZOuunkZJt+f8q9A08QDFqKOoDCC63yhQ08mn6xe+fWVRxsmeqlJ4MX0shKLOjWgbbjkP
EdPsh27qnc5sBi29MFS3H95IJQpl9rxFRJGXY04/58FQ5HxIRxwIpr0ltmn2tXkNMxbsNwTWnLW7
MHFz3CJ5715mZKKdbNol4U5XR6tdAz5LGprNe93PMG1/Zt9KcTefYl1lvAvihrmy8diKkz0X0ibH
f5UUx0PiDgZvusHb5Z+rpZNabbqnDKYYAjhyLqZZRk00t/aR3fbIXseEgR4foJIh4duGkSEg3L/z
NqDqcueYAqwwZAcMMxe5iB5IA/X4voQ328opC3MbFEACXUm8PPIRcbrrnIF/TuqxloIX7i/xTfyJ
pUMNin0cwgFz8Vgsjq7NnC/emjXWsxGsO0aUtHlRbF5wytX5I6gYjcrgoPVe4oTEXSkoTlY8FLJj
n0jJN5hN9IbOa7yoSNTrWyVWwt7DAr/RoxDAr+2WcB7W9ZEMMYfKWreT55/LH85H9VT5lZ0QCt91
QawZytZSc1sj6dgk+Ggh3Yn71dZy12tUEIovKHRbrt1FxXZzinYJBx/C5raXZugyfKSIvtxcscFQ
MtCMtX40Br/vVm/eADPMYeYJYbztTVlRNzvUOF+PdRDy9jItGDPKsVOsjkaQaKtOoZzzZDkqakcU
ghYJohF7zSQvdGGo/PTgbtsLVhUpHQ7Kc86AsuC0RSlja5OrDxnN0AbhLY2OMNY0QOh5GN/VRWEA
unobLr8OnV1mnChijBdB0n2o2/ofiJGdYpWQmHWb5SQV6C1Hb0l4B17DoBQSwfuvdC1fiwBGbH38
Nol0JRSToAO+w+ptKentSy59h9LpNu09OOBNNPttqmK3fCY8sQf5yfmCA9SU/ndSEQBkWeVSFE4p
jHI3631CvbNnbtsK0PVze1JhO4RlYLBlr+BdLOMztJlNSw9zbdlLsVXDsfKNbmfJcHSAreuu/Ie3
994R7qi096120Etkg7I7+YuQhINYuJ/hp5h4kHQuk3YnH2bP7NZDByFC8+ccldq1kNK6oQvpz1dp
6ssPa9jRzTFJXggPAjV20PKZuLXQMMZoPBtwU9QWPD+/QmqfJ2PYgRJLx8gmoX0SVAn9rJdzqr1X
BwU63rMYsbisn6tolo20HU6h5anTTfGAUS0Ev37+fFqQC4e9z0dykjyWwo5yGaoNCjMr6JjdFHcI
CAGaQKhtf74mYZ54hYJcblalNG8Dyqylk8FsoNKSN6ca4u/HkTI/TY+1hMQMxTo3G12gN8A91wwt
Nn5X1d++ZYtsQakK32Ozr+iSpE9GB7QO3ra6WE9j9LYBUnUtLNzT56bO0ElRBVtePND9eKh2hEjK
6y1jzwWz+6EhBY0+tgRRbb4zrISHCP0L2xYkE/vzXMbcJFUTtYeMju0gD3prIq8o5t512mMjVTDm
3ivebPVQT2JHqso7jiKlWudPB+we2MCppt16tXuGSD6ZVPpam4p/NBqes+icnd0wsBSBh5DKjU7+
qP0+i/M89TMlToVCZImxgqeTPrdvi6/QZlMeBXeKpl+x9OaiAulz77kYI98AfgA48NaIJc7I5g82
gphjo8B/X9m6tEt4KDXulqSj+flFeyppJIDiw37ebqLCQ3djJXbJxQYmbLfzEkGYFkxlyAOi3/ut
Kf63W3CaxTB1WyIjEUym+kiwqqxv5VK9IhsLztOmE9tIjLGlwIqBf3m22QWLQMFgYTJC8uv5rL0i
D/07gADzayGntNLp1q5nuptXNjKyNSwapCI7xuGsOF25SyIfSqLPWTXXWWuMGFWKqlSZ394o0Gwo
EXHQLxXeSA8MvFRtjUQNdVVWaY8m5i3U9KgTYrIPichExmw9ZQ2+IZNnsKXZeGrr6zIqvr2KliJV
JGIXf4OYFoXeZSdttxN23XX7kulqETOOz8V+UU9V23iRLxoa/AMGoakPCoGRnppeP3/oAm/FpLfd
HskcAjZJJh8fqEggj83fZWNxqmk67SnY8z1evlWvilKyKKhoijYrX/fo6gqb36iTGn/TSefMNG6U
H9rXwVxfm+L4L76XWrhX3OiIyqF9cHYYdA8Ft+92ORfCOc1/c7HrgcyzOfFliv35XcGsm292sb76
mdr15uXnY3O5x1Srt4dJuwsdQtPBpgXd/pW9q3Rf3JgyEbr1LH3Tv+xXUThs93Oz+0SvjVUymF/p
r3I9gt13hR8p8sWimjZ2RaV43UOXbdNwTsPJLO2VJiTmd7MtJgXMoKtNovoJbaf83cuLC3XtV5aL
HAD0pB+Q+oeuLVYqKqaFMYV32mIY0Of6d+2iOEfZZpxeajvQUSvjdiZimne4wBCcQUFeskStw2Yy
QonGGJG0OokLEHBq/8xKm8tVC5VBkd1FVYv1qUnA4fii1WNCQicX5Lrv3EFmwrjoQnc0XWHQ+coZ
qCIT12+DswzNoCtxCAfJCSk0mKk84rLvH0RskyyFu8pdmDGyPj65wdCppNjwwsUf7fMZ3XS8a7y/
Y1HGm0phinoOs5F/rkW21cZRMyb1HvG4QZ/BnOGfYu/HPkUJzNGFMHyhgVuCk2UfDoN2OxO/caun
bVZ2SgfqdEdiWpCVQYRtnU3dTby/Q5XGxDwVow2lfFAtSk0axoCAG2aCOXxJv5pAabMnLO7uyyRJ
6qlfdnRfUsU925FPErzeWHH+MvUdrJtH75t3BI7WKRskJRUZwnf+RSz7KD1Lke6kaNw95BvPsHC/
3Y9zE+2g0QSMtIHCg0NN+MRvhYtBFnQiiMXRiBeW8tVQw6x8BLKaGV8qfF4rXS4pvgsN317DQJOR
X265yVOkzWI95IE9QDAKpGTh17hW1pZqQ9O5zLCWGFGjzbXIgeGsgMhWVxN+kamIr3Cbebo4JvNm
Tbv5iisQ31dEOg5wuZq4ih1DDxmSxzoQulQc6ib+nLIaM0BS8fgOaCOP+x/dOUoekjJ0CHv1yKME
mXPn6RMxABYbHnNynC6zPu5v1iIDRgsdBkrJK5PR9ydmOPvaOdN+/mnmwrldGvR3fqgBuIsl22eN
DADIOHLybfYDI+huYq2pA0h7u0WOnjwAbwqow82J2UQgdE9jwOMCKBZ2hK181SIebqvGE1f1egbT
fYCUM5vggvbIehXjMZurA6VhNVJYW4RBzpkR7fNTGtmLDRcicFN20UX0oMCFSunOFO87xI7K5iPA
FIEW1P+AQGFvSM17fsDhGFXQ/p6QhbIdyxxSFwTKGk1chWRP6BTYsiGFjJ8dMNo1QZzrOckQr4g6
Bu2MqcUMlKnNYp1znwhtEZR4I2NXFduI3T/ETkMPgIn0gbuWqK4PaaJTnFbQzWjgc2Eh5Qm+JImb
0gefte12qpo95om1PnVX9JoEzxwyJTKGDx6lFMo+2iHthOCH5Ha+Oyb4vXsFVJzffcSKGIWVKvSE
HHqkdPUBeBjX525IyioJILvokKuO/IiM8UIA92QWiY+X2RgaYd+FSRzcsD0PrOk6N7jugTFAea+H
VueQmmm2HYe45YQZl0ovnVtL3I6mmIv6JtRUfSC6DBws5L5DuIG9gLohIknTJATITbW1oEGdD5aZ
DWaIYsLOQ2tZSc9y3b1dN668FLym7K2OL7c89XCC0gPMeq5eH4oD377AoAO9fgI842FYUsabfolf
xLoKmINOzy4QAEpIcVcbsO73o9N4gCKiQ1r2xAAe2M/mNZM/q5c63tZlX5up+9p61+TPlz4vjs7g
mYFdP5WcNCMqHBakQSFG2pkESkdHC4RO/KUhLU9zwagv9Opz6h5etuHMBnE00SNaPPmEl9OiuLJC
5nl2x9UHePIxOTvlHsixNxZQa7V2mjh8rc/DwF7ZBsUOmzZpkGawcINa6rT7+ekPqn5Kz/6AB24t
9czV3nwAH73THUqouQSP0FnEpkSgL8CtBVfVf0tZq1XvZEbfc886yrF5Im2VqBlbkUUlBFx06icu
IA+7BuWq8h2RuxgI1cn9asshhKoWHXziS2YomY1Wi27PIW2cNvA25B51ilP90kht8nadOkX6hRDY
kncX/zUMvZLy2P3wFzgY0nAJeR7LnimHDds1oPteY2r9Nu4ORo4Z32UtZfKzDnTW7AAwJ5SZ/m2j
YxHPZwSSi9VIByJ8cIEYAU8/Y24SiQaJPvblz8zK6gR6P6eNxKDSvLcW0YX+fHG9k8KPdsIHtbUJ
9Dpwx4leBn6L9au2HwGE8FEFaypoicSz+OzyRHWrINH6nq7AMY3RH7GOJrGfPieQil+f9qKVw8+I
ZQvUMXCbBs/SatQB10Ruqre7CkCabzbq/9Xz49zmvHFLipUv5XFqWdoYgtvTquxrb2Zjfg4FtVaA
SevIvaWrJyk6YZSx411DQJ6BqrycB3JFqJsE0XOQwzgd0tMNsUgy7GYNCRq6srNAn02THPL6hT7r
3PE8DHAhTIgXHN/VFT2jeLNd1+1Y0c+FUtEvfSmqzAt2+Wiz3ezIREnvCK3WqfkZ0uMfWsWEmH2y
T3gPD/SdhkRw+LvIvD39xDdqEvhx1zj+rXMfqi0c0khsd8LfjzqZjFn8tPnD1eW6Rgg/yeM8DxRS
l9H1/qw6hYimPG9IMobyt4UIHcclqyVV9002mbPIFKKVMeY+I5yDDTAoyL0YdYWFQ27yXtK0l8Mw
nIzh5PnAhNAjNpVmg4osSsMqZ6UEl1h1LmFWYYgthj4WM/G7QQSjWy/C7Ao8gkq0Ku2emv3neHxr
Xxs6Rav+baN9lds6skQXUyNz5ZNOuShrxp6O4pOfF0uxPTi7tBIvvAyUKgAzvrPjpGR6PNCqMqER
ynnLgwDMYIZsZIniTu1hWCdoU/6PSxfpm0dNRLHJCkWEApOluW9GQGu6+Cl2gnE6WeOn58iwYKcr
CfRYq3HcJx4YuqmPtfBRyrr3kkBay03IcVA0RnsW7l7ENMyDcnxXn7eRijr0ZSSlMXDVVV+lnhTW
SvHens6PKZ3nwZaCgLJskhtgElqXsgCyVbZyIS9DbkUEzoG2qL5GdFU/rvDVwMYCsaCg3WMcFAeF
pvkvaT1n4E/oeg5GMXKTUZwyjJs/U3CnCoq3awHC+/rZnTfbnSZ7wx4Rj7H033JH5tOy5uQ0n6cO
nRDh/SIjHLfHXBwTT8z8rsWVjoxQiTT08D8KNo6rXdhSVFI/s+VMU6IxaLeXrbwi752GFwlZIudx
/geuwKaiOM5eGJwT8IU5BO/2Nn2Ix/3kzOoIBZ1xOvDrl1JsFRvGye0sz6xISXUMi8aNbILc6jHO
bEEc2D/V1fxhTFeyEuZnRdhdVasv0fiyhdgfM2nRFJV1LyvwvFdy0BRgKgVchobbTfA7e+rKCkaY
v2WiZ7zRqCCFqThg2uE5nyJmKphCC9bWi9dIZBgJwJNxTxXO3C3z28BUYhF7Icph2f+34xHrJA8q
G5EnjYVllhp+2bUOFkWDYH3xEFvEoV9P5A9jmaJ7BQ0MZjOS7q0vh9/AE9scC5o9wUfduehvLXCx
JcCbEZu3aeplnpt6FYyH9gQTiR5pLZ5tbWpJEqkGoCN1aBC9pvV/e4ZO7ifz/a/Qdh4/liTx4JS2
KKh2RdSy42hLYcS0ViANmH9M8VTE5d8tnABcev3EvBuEueFEDP9zpruCPrVPilTlc/w8iFtU6LwP
NX5lOVOhXBN69PfjqpnyqQ6WgYXM2ZuH0C5ZomuS2bJV6kI7KhRBuOX8Pgaq7nGNEdcP/30eUDLi
oCjgdIZnI/bWDNxx257ExQ5aT7k5FVspSTcFBrnt+vqvDqMdBdJP/bdlRSyLQ7DywIlliy7qdDc9
KdB/Z265UUUSLIJKaegtQkcpK5zCNQTFlTDAIJzHNuuSMyvtWkIUmOMozaZnEpiTSZOkg3rJXuo1
vjtW+xU4gIgErW5JTvw4oB3+l0Fp6C0Ls8taGBfO7byTHI3Ikvy0RPNW2iuGY2bsZxdSUqy/Qp7c
VmsJmNweE1IrBWrvYjXrEJiCRF3VTLJbFVVcb6LNQehG8ayZv7kbTYhWxJcw0JB4yZb9Gklrh1Jt
DshHbUmcdVs+wO3/X4cjzof2nn90XPG5L86knP7Lf6ZUJ12wc2FUADNXUI0aZmWQMCMqSkL10/LN
0xtzy0RXdLrTB92V9imU5DRvnwOq3I8+5syogTA8FMMpUoB98PQf6oT0GI2T3TKzPPfp/q0Nwzfy
YRURbYxk42uMx77uM1r1JkpkPJxEPEUgPFF2ms2fyfllWv7pRkBMtb2wK+juzpoqiSxOJpWLQEZI
0s/52yHnYKDxKsGKNJNK4twEQ3rm6mHKGsHYaXVDUG36PethUnXfS/klzwbnWB8Ik46OTVQWdEAZ
k1C6UGYY+nLwxdwKgG7z19H876wFTuWL1JTtgMIuusj3qE9sUwaQOafsRf1FVcdvm4OSbhR/o14F
GjDmgDBh5QzL7ukmvWd6As/bwMO5ULuB2N3Kit5BW3WYbDFsnfmBY5hwKxAqXSvzbGaD6xbiX5Wf
ChFZ3yRwkYSmjahq7y81d80uxNkM6OsK5b3XupyVA6G05cr43OS7XGgjSU4Ayl/x7hrrH04T7gPD
iY3/PFhYVMpjzM/UmjoCNEl/DCx3i/817GxI1lYlBI4vj2qTmfdCpzjA0k2EEslae6rv1pXUgRP2
4WMNeSZ7bksPohmNa+cB5+GbTydKsOwnektRWp12zsBaqWYU+IEoO+9KPDOHQ6UBfZEZzdobYit1
XWj+yzN4Wq7KTMJ9NC/0wj3mYfZ0pnI0YLgg4jGlEzhxhnZLgzjmtXrprdNmpu8h3jsSF4IGVdMg
99FOpStWS6mWmBb12QkwNDdFgKRXDhKkaQCQr2ywxcxpXLivf7eBFSxIQ7wyl90mS8IsuExqfAAv
LBou0DatrMr/YmTpCAKDM3xltougj9+2dRgsDAHQ3fiXLYA1GxvN07Z0UHge45YUc9ITU58DLvO+
Q8fOTKo8VTXCA2WRrgFwCiwGZ5MAyxO90jSBIK8h3K0iUvAcvIqi5zSsoa8qS7Gq9FCRLmSb/tJz
U+H0BmXlXvhkiy2DEJUYgIhuQcicmwIGvTBuAPiGheV1D/d29B+elx220tpVgyzuA4H6dxZwZ3cn
C95dtRKNigOUfjBXMFBuG0DMXs5kNSCGQ6HzhNS9YwkLtSMkA1nundj9EjIR49rDEgpf6CrzUvCT
QqqnsKHwtfuD+XnV5KXWGn0BX0+Qpk3JBclrMwHbKWvsQsbiE27Na0STCCd4lcdkklMGsn0PAIJH
lyxEbVf76lg4pLkQ17BdO+fAuSLkeBj2rx5cnRG+rlG1XlPsdZ3CbdFHZSlSvFmcrseosLmveFVy
/7SgRZ61ojxFYnyJABY/WexEoSN/SrHrsi3MVXyD3CV041c2m+MEtmMgykRNgaqQ5+B5PBj5T1rP
pGJhSsuLxq4hdCgS6z6tlKKCF5zsB0TTL0SnPeaAw9LPLSiOqM7OU9Wl/8cLlnp9wVYvnQ+lbcga
NW/Tqdk9IvLdKQ0B/eHdZDbzYfHaChjn9oDF0VXuQJo5IgKpjwkwxgwZNJ8mND5fHEyDXFWFaLQI
I/Ry6uCQqpPMgzsmWZ/lcwrbcc6roczUZRp2wnO+hQL/HgkGvRWoDhOjSN6CpfDR7qKr6lZDLNr6
4RoaiS41fxViPt4JLqnCk9as3NLgpuvuw9LJACTDi3t3ryXfR9mGaYb9liMUOMtdTgyZtx8i3vFB
XYF2XUpb8MSAUPSUYEoHrhTFgb22trI6U6tOaVWuHa42NfEzOKilrslywLnVNKiUcJuqk7+TqThz
DrZ3ITOhBITcJEwXcKe35bBv0TlV1AsZWdjtIipsd1Tv1QuP0xQZQG9uAF0NLnoK1jsViOOOYkdP
9J7SnP6uksnYoyqlVjg4LR8pVXKJBR+9wxlpYWKz7FpzAXOxTFB+tqNddLm614Nnq6fuqoAxxxth
Ti4i0Dosv2KfTozCYLeiXhYwiagg2m0m9zMZiv91EIfu7jU8J2GAy7+6mT+zqYOyg8ibl16diLbc
80WK3q2dbhxdSxtqe2pVh9rlnGzHc36A8OcepGrlkyZTbo1o6qLSMzEFb/but6jhhsHtJeMPFysS
7s3AKfFWjRt8SaUMRSYveW3sfHiB8KgMgMh6scBBCM7wC4ilCslYXcD3PeOMbC7emrSO+IkGLme5
P1+EeVUE2HYd62hWWtuHKzjI8HYoiCSZWwWFFPLFMBPjK4fKKzsCa9QvnpUVRx4v3q5I4qIUmWj6
/Svwmz5xJIzZ8gRp8c/tgZ5ta+XbyPE/LxWryNBFe/VwX2xhE5jU08MdeURNVmoAaP1k1EMDTQX/
Q3lH41EgJhHNorkgk6QxjzIcHhQFPbZjLH6bP69/CSiTbP8Y9ZfuDrDLIzPCreL4BDCAkiXK5j+U
dsR+etcDobzWc8H4DxH0F1GXtAf7Eazr2/e0K2ilP2MTVZQ0TiDkgtcL85cUcHBuRy0i3a8atRu+
7/jAkXZhTLiWXnXq8diEd9vhxiiHV9tLdhGsmU6GW527zBfMHW63FElcEFjB6Drv7ISnFhkB2tDe
lHiq53qYn5Xfck4MWssbHGucBi5/SwuEGo8HG/vy0PhdeLuoMayJ3P202wOKhZqGA9RpPmmWeE8k
sbXvjbk7NXkeoDTbekcNUr6GIz1WChv0rUUS8D4px/2j8ZIjhJTMF5j3HK35lpHY2nELj9CKd7Ap
NaNfOdyr73l8TzZQ2715GbtYNciwjmbVp5XC8SdWjN0ozS+HScxZV8huyWc0Jlduq/s25xBoSbGk
KyV0XoLbZ0RvDvHa7Dnn2WkuL84V/wo9osND54ce41+PbrAdBI9KxN1kF+w95SeMDHWSPpfVHg1r
i1HQoFzIojKjiAB1v6kEKdaa0cRDU6o/fFMGM9eTtQgaSLcWcpTCQ1xc2N61HEJLL4SbpQqB//hu
ppRqLMvzzEceRqTx7kujopKsmSN6vZxoZu3jBGA/PQS1RaqfLTOYaHYgTR7PukVixFEG/oISzOol
cec/EAH/EivV+cttHwsR7ugaAgZi1kNoXEuvofb+6ffz0yTTLvk7kqXSLjZRLCVwyXOAqFraRNMh
/bDG94a0XWnR44ieH5QhJUzFRdTX/KBgmdSmqfeR9z5YHNzcpq09s56ICub4X2ekPi1qJz7P9oI5
aAuDBmMs19Z7bu5rW3lyV6ZHqOm8uq3JOQnDnN/A4ubw4cWgjfeMb6jpPFr6q2Zgbhnw3XlboFAi
b6guJQ0J2rI7grx3+jqs9h9yue3sUcBjOXVR9BOfq+FU5LpfCGPgugF1wmvOIwCzVyYcjEXrB7hI
GXHDFg3xBLwWK/QGpZ+jLNStbhMkWqo26UD5XPBdzQVAqG/xGZ8DijpyuJJLkuYBHfh5g1NehS4X
cnhOvMIfmhV8opID/WJjZCjAL3t2tSUoJ4IIRZXd0gZNTEQXtWu91+bzwdiq7/rSBf3THfP3Rdm6
wMIFxt9THr/V6RkxgqtkYADCF1s7HZkMazdwe04r/8boFwTFCaHJrJ5kWv2RCU360TN0sNqDEV2T
jR0omLCtPYMJwWqi0JNRrh2nG+Dnu7TBUdSXI+qmUkXcTmIeZvf71cgFZin6bywPS2OeaYYo8s66
USP1uhhc2vchsQ3sVEaITl660i4o874zDNhraaelfJgap1PQq55w9Ov/v4T8MR6bzSvHDahMAaT+
n2Cjg+Fr2zWlqmMMxLWOK3MYEWUQiCpSDa1BjtHcxexbJ+3gsV1El6IpcnNeSLKWerc7GDV05xg3
MwbZAFlsEAfONqC+aMf+7+cWQftYkGx9eeAJnlUbKNymLi09cmDJINkdPVN7NvY9PHssssKgizw0
63mT6T/6vPwXnFTi5jukArwV03ore87xs+49P7+s7q3mgJTiP3ht7+fIbLFi/dPy8bk+EMqXuTJo
V+klPQX2MUFO36oSWXH/xX1ITfdqTs9/oa8m3//mS5YKMwRPzdPxGznfI1rrWffQRTrnG+zywzUL
wNPloKDqWBPzCp55FjQdQmJML8L4Vd3HCdRdb+fwWSKl7ikCNZQQdkz6wtIvWJHtzoVQCG68tQS2
Td7Yz1GlMFLbaYqbM8hqi1GmlM/PYIEsa4jN3aOo3z58roUaXMKWVXQ953Yb6Y9KKfKc4jkcqnv5
g3DOc+bcx+14isQkUp0qazmXJxwa7Xes4CP6EuV5qmZWq4r7uSbLXHeSWTMQtfDzaKS1oct5R9qF
kzP+7A1d5MqPkQwu9mxqcc2r/qKGYbl20ftpMKKbkznCBS7c3eoso6r3Q77H2kx1+K9ok7Y6MEWC
d0PDU2+Si4Q3W35TbUfpua+y4p4PCxEu6wGURYZZE2bR7UOQmSTmUHXdyTATSR4Z4hSz/IZb5xR7
uEA12aESc2oyzFP8+owzK0oFAGRQkQejBIoUeZCYWFc9Fk1z7+3IApb+qmHD1yfOhkTwqWO1C9FY
cJCkX15KctiCqhK/5Z4XTF9Jj8k8FbjUTn8vmCTsbYyhbHUfWQD8drmZjA03Aiffl8iHpHWM7Sy+
dUfcM+wCvRRLrW5js0yPHrKkJKDelhtbLlSKar7DU/jyngbDpyBhC8ndcufuH7uS4FEN8OeAUaWP
fLtJ36ASSMCcXsmDSJnzSpV0XQtmWOnYXT+v8kGUF/+VmpQJ80Vz2zH8Y9D9RxwAdf8csb/XV0LF
AteCsGBTn99VH5xFJcQ8TdvX4CgBsEn1YfpP+EJoJva8YThc7Epl8XxP9tu19CtCsyPkZVPbY9sp
LYPL8lqFuUxba0MBtNzmof30zf9/7vgRGNRLRWlsgBUsZF86h48rX2v0/PhTPAGkT17EzxfJJHKw
vkK2NOrudqAdPPF8kTt2Z58npPCE1Z7AGzzmgFkLGYtNFnMOyZNbqL3+EACQ1F8QJiXuJQ7PI+Sr
f7JD9LlbWwaB9ObMQSOUr7TP1TYcuIx0uHP7e3dc9CoyID9d091YcCPTkIa6ELLNfFvjlzEbN7xX
mv2YMiSvoGiTR+Lf423WOs2kU8hXMi0DEfbugCGwu5jOHhzapzfWOyFaAhzhbKsqeJmBr3MwFlTC
UmXZjNN7pL6BMBVYIS5jFp/tQUz0OqoRNZBmAS0tJRG+1tqlgb8aGUu8bWuAWPYiY90t+GA81Yoc
v8qOHYBWpA3ucLB1omuI60u6qdZBieYO34MftYU0xfQRZ41+7hRZ9U9f5ogf+yfj7MBkYAAepGIw
u5ZJRms1Ctx12QcOPySDXp2jOGrs6Jt7/si8NEIVSx4JRGDsWpE4GAaQ6x2IgpZ+C7+uCAiSPI4h
Ec/i3P5nj1mvzZzewEX+NAfBu7o2Y261TXkgojBY4uuMuiOvTAEsvpy9YHP+kqm5zUuuxGRPwH67
a3qx/Krhq8RBr3SJCkVeOPvQHW8WA2OH3vsgRBcy93xkEpHuW2gL9JOa6veJsWGrvwUM8PKU+UFi
cs0eM4akBNJCi595/Q/ZYF2O+HfMlOqKMd5NHYS0bDrEAGNazGQl7HN+B/b/zih/Mmab+7P8LTGZ
sHUYL2NuiaBHBDx+7YROCXxwHbgQpyyCQSJHzu6b9Wkd94Vl2Nq1JWW55fSko6Ad5s11nlAsFI58
4XNnqIXdVyC+v39vMUfWiZY3yedvB5im/ssHKT5MjXEVDcKSEyzewRquz5sZMb4/OmiePmoO+qq4
vxMokd340ZfjY7Nh/D47axaDI/5uf7D5MKj0d9tzkDyn+1Qt+uOT30o748fZGjWpg9H10WzCVSRI
FA+z/edu7YUhX+SHkOupr16y+7bseKdeCIUkFqdLAnUWubg8YyRY1VFLglFnmr6bKiBTc3kJ1UwH
P4ailM4do6DnD9huOhMX73Mriq1871EUqMSaBNgdADkgEtIEuWafsQVFkh9jj45DBtRGX8K6wAx1
ARCCT2WxPt2lJz6/OZHPKRXU3h6OFEg3d4dDc9PSrX4M9WVuQse9+KZIoWGrVe85uYJdTI7imLC8
6Jf/5vZjmpdE58E+aUunZgMsd0OW3dFbrz/86krpNq9kKvaPZ381TjYdO4DyglNxCkOyFLomhjZI
HbnghgSOgTisLIloqqbWDx4yJ/vPlbiuYotf0M9TVJgXu/d6rIamcgI3H7dtBJDW2HUvRf4GtjxK
n0T6soPm3ccvrUR/FUXBUWgCs9TVPOS8CmllNi4Qb60cdr8VwqPHxC2aMtU1QCo/7ecHhFL1Jtal
Osd9IOxmaGSryx/5nhTVgOhujVCVlcpzzIn9PcN/oV3Yz4rdTeXMh3frhK9Tm0cvYljazx6uob+i
rQpfLjvmrmr6qlKcdWs8Kt+W+ks1YCse1UlZv95+LGtGUKKOqrzbneNSHUBWeEgUyPe4JxlxxTmN
hceQkGno8r1HdgS5aH9tWO6JBeLtaiyZBbatImBJIrqu97pNYCZWjBhucCNilIxyL/zn2I6VFTmx
jOPP8QMDARwtgYuzF+3qvhRgUFHKpHngl+9wxM/TF8B49xUf7Em55nLdJkXtqex2hN0s7Y2tiG/7
/Rth+dwEKWtcRaRZK5X8Iav998mvQlGD3M0NyFPwPaqyCS+DiBe3CBJfjeahJauj9vqnTxpQr++V
LHgOWQBOaFou4q0pkVOd5OAWVjMZ1zH+V9RyFXYimDJNV/OMhVCCOKJJb8YNJJDewma4ozefN3Bd
QLqd4jMbDQwmLjMv8PHmA96qMQvgfp1iWJl8op5k6T3qCeGl2DiffQgXSzau7bRMAp6I3ArFVc+C
bhPUoq0Dq55Ec2wQ/ihnoJoUT8BmQWEyaT54A5qGkJTCKtl0+fcX73ZAVYZ2zbW4GmMFaRhukCfz
RkyV18aFw3zscwGgGxB66FnSL9qG+8zzlYElwwAiXr3X/PqKJchNU8u0OKAwBPno7vfsh+agvFeI
aqQL2H3J6ldLTsCzjYUU8u/Y6BzHBIRlEStjv0s99Q31d+4xay79IyzAtv1CC+C2ruUcC3P8Tsk7
td2+AOG5gd+V4Nmpe8Psd/CTXMl2kSf+GOHk6jDyGYnucp4PIP/QLGJfhuRt+vCnuqCX5Hc/XwQY
HDDrOr4cdMklLr6iDacUJniy0Xof23Fq6NmthXvkwlWXAigM7dKktl5Z6nmtZYp8lfvjNL5rAj0a
m/rsnI5bAN10Z4LuTuGSUuoEr7gED3k55NZ7a70lUvYPReIU2hyQj+pT9kbfYRoEhOUaA95UTkhn
F5gPAR3vdq/ANszhw9dPHSYyOdzjGoDtybZ3b0ie3yrAayLcCdyVLrngyXQLHO6tWo6ltreW1bdV
nzybxut54i46mcyqim6GNAhYVuUmm9xXByNhnSk3DpiWOWl0JCAZufOee9GAvaMHDCTXXTvhhbPx
upKaaiDpvCi5pM+Y614+DX/6eXq0dj6uwfGIuONStCINzB1yqWkOSoNd6jPikaut866Qdz1ievV/
/Uxwhn8fMBow/+obCii1uattQuWNjNlkJMsZIRaGdB2gkJRhW/UFV47rNyThLIkQB9cdX5bBbEKJ
2h26b+WIQtY27gvKoLoCuH+9aYU+o3LzGHggocbWSmRgvNMLytLVaprz8u5sUjbJ9TA5oPm+PwZR
FTfLtJkpqpMSJF6BulL6tLbLt7tok74rGQpMwEUR47vPCGkeEORlNdN/rK7XfY92jL2Bm8mF5URy
cTDGwIDYj3UDNnUXl4ZctyjST9Ov5+hFSPrlVP9UzRzZN4AjwO/t1IKv+1nvv7cDSrXtfTZabh2W
Iks/hZqCsDHQNVvBmsY7cJ5Zf4wPwHTwdJlJMRW94bUSZNMaWbBKcpdQPSEIta/qO5quhbHqlgLp
OyGiixI/3OpcvrDi857jks+QBDRxg1vy/QZZE9WeYGgeLPvU4AA6C2KEvXnLmywCMO1KGWVeRdhk
Jlq5XQ6berhSc3P/I/ByK7nWBXziPfzWWpM17S4jc/y5s84qks8YbQWAJh8Gh/GUPtY8/IwKTxyL
7G/8UxV1v6/SCeMlJjVbLEb8GCImxqF6+oikgkcPwHU5jKOS9jYO7VYFOEeuXYRip6TJKiX/Zi+Q
omTGYw95DSMLelAxRfCppKMQWzevfqpDsUrOjUEZPdJ/j8ZwMzLez4sDuP4Uc4Z+jhCF7QU0OyCK
+acs7PzGi8GIpFFNHASN4jhUH9MHK9jFzMDoWKnWlYubNDSi3WY4g26eL/f0hO+Rv+GKbA9kxDtT
equ30eJ0lDqBAKTPZ0EtZKHLMGJ0iCbJoKj0OyXpvY9Yxhy6CYfZjS/2ZUojxRZHG7D4api/Gt1L
/98QMHj1tjHS2A3j1xGXaTZBZIKtZQiLUlJAod+Dvi0Q5H+73LCU3/NIlFrmW2ZYJUNcIll5ny6r
kQOd2HTL40gO6q7d/KVwalktlE2fY30cqW1M7zrcUNCLUrw242H561ePxWyhCVH8QL/hxmuItkrH
XEoGTjD2VmMW0teYRVXfAtH8coACYPYAD+036e4ysaTiJwUd80vMz48N/ypbVjDCz5b6iLeCOfFi
fwb1A/g0G8XorcPSNEz0+1fip+y9bpKhHg9vVISx4XJMESz05W5ny6wsoRkwI1AiwgUwIcDtKYA+
LtO32ALPrgC2wUA8s5qOjvNMSwusVsK5EyZ0uyeo8ho8VaFwSoJ6vOT9UM8pLkx5tWwFBqE1+n2b
plume/zagW8VoaEK2Xk2Y8KVZn5Q1hTXHQSqDLopud3aoozwcWFzrnDD67T9XQIk8fe4hIMyClaZ
W80oUf9F/15DEeF6myYuoZXHLM4tdYg3aypdfIyAJ/LI+llpXe9hRvZdSbwh+3BXH23aqf2L1T0x
w6bNHlD86qy4dFJFPQyJJJyO+K6rzXiuILbPP09RrSur+MEPQ7fvMM5ODnsnujBxOtRZY09xMVM8
c5WSi34MIpAZxUxrO4Fsq6vQ4iNVOW93qbzGppyYn9tvJLyBqMItJp3qdv7KCBkpnUGZV7LI2sSj
KFIONPPVfNT+DD8qEkbQSxpuxHST+40EDRcITYeuJThGBZzmJ/oPeFPQiH6HiaW1cWj0M2GvXmni
kUw7JGE+JLiGj4a5+iDt+mohpAlG/dIb7DJrFPl6uKYnq7OABn0brzaK2ML1hFuO749OOkPO2y+S
x5u6jKa1fvZKu2BvGgngTe+gAruR3sWvOPaMxqzgZnYN5+GH1+TGjGCBlsejT9HOerkQh03ZfZ3L
tI24EFd9t/aqflXFl7+ysMflnLTfqZr7/3rxshfK7aiU+1PQCfAsDC+SJIADzhspuzLBwBwZIQOR
d9iY3q9Xm84IFaqdO/6/Hkg+5EYl6qhUvdousa3q7S1o1YWFq/QnI+2ZR1pz6JRG3uQKlZDD5wk3
YznR2oJeF45m9gHSv/EEE0wHGqYWqfpkXtF8noheWMywEUYbeYqm4szAERmkjG8uVUmKgb7Pd/DA
+FlrpAFt1uSl+RJALHztYyZxpmjsPYFx+941kvR8sMpSHAfiqs26jE+7zredPk5Ory4GziptbNhK
6fJR+p7Kk3+JGz5pW+qrwjEfUxl9IqVZYvqIFJGedBLCA+EI2yC67pc+SdMWYupX/dkEv8foQ8Ge
xNbS0sysV5/a22x3cSPUs5Kyiv9Rf92xN7sBqJEnSVxzXI23FYJeYtuLfF2bu7QfWSwgGT00OD7r
Hrkv0yUDd+zZS+CFIqH3/yMwh9sg2yr+1qkiPgw0Hkp4YcKqZGEgiwZPS323VCHvQiaoLTx0LxUk
G6FOef/7Z6zcQNt8RbUh1OIKoSERDGhlR08dGHFQ7iwoTW7Yht1c5W/NZOcezCx9MI4tLT//TteO
kHA3TbGL7k9mNDW8+6J3PEtqdJ3OGEOhIXX7PesWcU95rwstBNIzAd3euYiA9th0v4b5d7Ww0Llu
zM9rV2+Sg69LPyY9Bxmw1q2KHSxcqXYW0YLzdY4LIpGBNc15VVdoCywx8d3TVw9UClgiwUYAwPoo
XFjV1xRpcMWotUTfC/B21QPY9TrOAWDuoMfcxWGGNmItHkh7Pnuzs5QUZkrz76yP5DazgZ1cVJRX
/p3zWpFTNlQMo/0AZLzGWCdm8LRp63kCRB3eY5I/6913RS4VVtvCwqaYvoi2vFu6VTRSdZaAB368
I/Fh06xXiIeFKr3Haa+YInwCepynYiaOzsthGAYhENY7glf4cNLkYzeF5F9Yzfp22EEasL3N7kZ7
sc5A0G73rxx+zGLP4mGMIkG3Kslyqb0n8d8XFM9NX3eWZx5W58Jffd0pGFWey6yUqrIjgTpKGmKs
uZTeffnXNk8PWK1rx3VREVPECC93baejHTPmXEcRoUb8sNge7FlDtYeyfnL5dWx5kVIulLvgp2s5
EifHHOwAVYiM/sRWW/ZEt+EzKMujGqWdqUwh4r0a+DzCWkKOmgOOZ6rPMd7+GjSLqEEBd41p14qb
a0a7jBf0yD+8Dw7WLp7hIIkr0TcivJC+p+Gc4uA51dMVh7tpQ0hmOpgHYkGxhwayCFlf7WDvic4H
L8AMFOuUhUxMLkIfxcFFwuq1rrnRskUlAmt8/SeEJf+ThcO/uZX4fcScCtilqgaUZhJDKiPCwQ1/
syWd9BLBfLwJQJcHOnl+B1JLGdayiX3KUvO2OGUGwO8K7w9QLZ3yfVNsIBaquuL2r34FzWsZ87Yb
EKJ7/nOZf/IZQM2wtfJyr/UILr53GQ9YEQDoYYTlIJkV2RDl+48hgcdXaoAh2boAb9I2X0JkaSQk
7SnQlez2RVLcbw8wUFrSy97nWe+QKu7+HH1Q5Ld88YUQVr6mt3hDXTZcp2iC7gvI6wL6IPcbDXEI
mFuuSDBW3xmakoImZ7Thu/O4Xea06Kp1x7Iz6YUYwKUR7rTg2Brwymkr+iU0ClrURUIKOaf9guXO
8VU1gD1XP8vZWOAQgzlknFNgM+wPM6qVON67/V8AF68HKz2uoVQ83WG/3Iz9e7cb6cBusdkWqRcR
9+eMnut1KIP3Uc7iFUI/SLocj5E9KuUdqwR6AjwS3XMawnsxxrYB59o3r9HDC3PV8aA0zWDDNGYP
hypdxgBtUKjY/V+xYtUQnimo4mVwzfkEJUHM1WRhysBhSs0dhMW+gfWeBPewQyFLKLdMxTFHtcWM
sEnt5eTGn0wuEau/a32e+pX9AXW2bdWK9zAKqrskwEugm3mVO1A4navMGn+O3bVrYROWNuwYB3kw
GPvQy1zrIeHJ5EFwqnnvxD5q7fPNknAocTMQwNPlcmrUvSuRNKdv/j35FaygUPtQ0AgK8ZwrOhNN
MV9wP3PnnQSTkgoEfxs3byfP3fSSv8ghwXUvZ1a3eG/5Z3YUusGs8sVOgUhBrukhkMOHZXfgg/80
86idQMDr9aswxK5tHMgVq4v3BclRiE7/z1rEM2Ar9BXo9iNstTCyM62pdvbvi24cTk/s6SGpPr2q
ZOaKbVcfX/VcYk2as2AGU2ERJl2WADgdo16Uc8K9p++noANHzJyOm2hbInWYhVegSq/UAbquN9wa
L/9IFn+secWjxP2RMd7NGo9Ae4FZkN3u2sL65JstsfbSAvp7ezIQhZ+nDawGPbl648jdBG34bhzv
Xnixwa/nO63vIkx6p6nye60cAPgmV8UH6oNw7JJeZcNEHj9rXBu91N5WzefMgbaz1doSMj9un8gr
SiJ/CTjoRy0zeXztuSQAcN0qqVEm/38YxqvbY7L9oZM1LK44vGRTVfM/2sGVDG/sUowd22qiWbW1
XaTDyyXn8bWgiFSL0oTcasNiDUTR9jVHNB7o0unGDLX017iy4tpN6+ivNKJ89lnLajSvbDGJO1KP
JZtZtG1tLSbXwJs1dWouCx85BLX+95FACDITt5Dj6+q1PcwJ/WBRaD5kfm0RBRL1NjXbJgtXmLkX
HpXWVmMimxBZwTMCVTSBIoRZmCZdkEJJQaORWlvolAWp1G+X1jDyp3IWZNwK2PyrashfvQB6f0ee
/eikp9Hds7LxyzOyzdAbbNZ7lQLMhueR0PT5GIh2il6gS9kIoKjtSfDvtPCDNuNIxUMW3TfJcM4i
a4+OEqPJkpBAtpppBYMGA3u9XGVJtJBbK/MZ3CJJ7Wl6CAedCQ/Fil+msHSfHQ4N99H4LSU8aKi9
2/Uid9JDMapIgx8rVTg8KiAtJydwx8fK6VdufTFix8mCUxUyf68ugQwuhzOfBpuqFaFpRhKDoplf
83SuZGMxzhXOs+cGaFNzWcSQUmWaBdRt7E4jYmGnOMi5mMXSr/429DKv8aR7u3pjm+bi5RU1NCuV
ls1/iBbqcIAPfgp12qoMRFdnufojkStJbL5NwqSX7R9aX7yxIO7sW+6BFxwNTE8xDBDWe9b5pnOM
C1gA/gEQIwMMx7LhNeHAA0WDHh9d6vaTsJ0zi6iQZV0PSc5Pu1areg+653dIA7AWN8lqIWJH415N
SZxxWbcpGWII7mJbBLfDryZ1G4ukoSGOeYbTP7yNdswjaYLQkWhHDEygiSdh0jR3CVx2lb8cDfOO
9Ee6jVh1NZJhOEg5gx31f5J9v0u+m5MPclZE6o72aMWi0pPO+TNvavatbxugzxXT00/5u331KKyi
KRlekBBftkleqCFPIeDg6E86e/eMJvpifsGWANB0ULcAHLpjTEM/iq5qynxUA97YBzu8xjr1GR6K
o9MxD2MRXSUqXMGgaAeJ+udgMF5676ph1SBzJBaur4Z9RZ7ZkSlVDdmQtuuPtEfl5MfOY2x+mufN
yDG11QkaT9nkd5FymAwN0K3SbuwO1FlK54aov2yVHsJDQfN+UPJktFq0oUfdxjfBp8NP5JlNC6HI
3uxUUY72t9JaV+sveOkDDkX89lZC59O5XOczGvxwLAYzI9eoQrW7AFi3O+YcYOFfCWFe0iXiyqOt
NqkNue5V5NcnvsjAVGL40lehNNMYdsPV/R7umljDVgaNhCL+zZXyqEtDoNXU6DsEBDCXVhaQQ8yS
ljhVriuEbRH8aAGAPfFk0dQzsE7ay242IeGJUwgkCJ6hRgRyFHUnlEc7FU1qX6UB8guhDBTri8vx
YiRX1NYc28UGclGzocH20e1PGkDQ0KtCQeTUEbX8ttiAJs8E69ZzGy52YDfd2BIpnAH4J7t147dv
9bbsd5h76Ye49QjSjP/wJQJ2ga3SWq8OMTBxPuheLzrqMZyXAAJfupSzzM+sEjdqbrAaBp2zePYY
RMLlVY6pPIXSwuf1Clju62XjQ8SBYaRYlJMNvLE8k+nrItNWhnAi0GqC7ozRchkqsIx0Q3TCJOC8
KafAV1C39VIamWy3V35i/1rNudADU/ZOTMF3rc7L+wv60kJd4hOo+Ee1TPyV5C6rYyevh8BD/c0c
bg+wcb935kxpIchI13iQLYMz6S7A8Bd3YY27hTSL1L2VK+kmcdmQ+axzIwGwPhclmohOpVvg2WzW
GHa5X+yWzMsJ/bC5D9Q6+oLcVwO3ExI2Q+mUGNthpn3/rDg1VPNeT5aJMkGa3ZL1o8XDTWmC2QFK
lGpTYjelZfS/671Ud0X3CVOcVg+L9WA772uaU8s95rbfpq9/Ce5omARpbDWqbdmtt/aFK5W/KauI
IiS1ReCFgE7g9ERa9X+VG725k1rmLutLID3YJrrz1dcLyPK+28voOog+5QZTH5o4yu99qbbTHZYw
krVlNUaVNPMQCpA0eIqqbOkxNNEWHAkhp2q7g4ZqYQmTpUWXjbMhgHMjc0eqDwCplmnTdDci4R5Y
WhEexv4J1tbWuhmd42KM+vLUe9S4zAyxvWMfuOg/rdlRoFZXrDMr1YahwBIg3DXSFJVHwcMiXpi1
4HEVAAaUf/HnK6nmGJzAxIUDVB7E1bs0sy7k3g6VqwrbE61Om3lQOCTYyD5FyTupro7qceffroV/
ZB6z8TUQCS/21AvYhZNl7m0sl8BK3x6zsC3QyK1wrt5EPap70n2VkrlqcF141pq1rNn/2DzXEVnQ
0IBKJ0OARDX9XscIzzSBOgKkm6h2fkEyHCpMOnWdCk3/YBPz6+NDMkciRM9QR7VVQwekSbVMtFnp
shQbxTjUhhia+XiVA5jz0S42k6nbVdQqL0ol1dE2Gt6INujQno9spJTQbF0T97lt0KwqKb+k2vJp
qYi8uEMMkzbue1de3mR0RtOZg9/iJPyZA5MiPtpqnNZ5iSKD1Aa57lQexApNj64vmg4d6GFlcPCf
IS1uvUD8NI2xjLnmUCOKXpNtEXZ9RQuUHCzD5wPeS7LBSmitg+OMXKPDy9Cx4zZHncJicqahk0x2
KyKuPe88r0KcjYiinJA3djL+W8xoAWJ1T0RaCAeEN1sk2Xy0nRYwVnvZvmA423PnjXEOsnHvUBJz
ne8v74OcWg19kd2ep37Z07LhjHAzUzgf9nyRCyqmiPs1rvD9pKOdPB5PDjs8dzq1ZFVTHTdloBQo
hPeZkw9TgwhsQ98k0jbgNr2PE9qoJCGT+Q5pYiyCqDxGks60vR46NEog9ycTFd5kV60imyTjW2dj
vSXEP6h4HMBcbxTaP0KeuJDyGLElxkQ2fQ9CuDr510VonIQSPSk5/6EauQYMDslQl7cnQExWw/pd
sJzvAhYSdQvfhD7PO4LwkdcWch8h5+7nYkzvrOGj2FOitRAdcmOZIvJp4nEScOhxg7giNwJup4jb
g922ISGC3ZLICmydeWCagrnFRQJRu94BOLqnZfI1N6lqUDjvQIvBWvv5T7LcospfOxlgk5OFnct5
ojba/BGWby4N7qLbPTaNI3EzFYJbNeSv4OeH/txGsn2cZGTH3Nof6ZL5vhSpZ6iVoYgeVLRqB9DU
+jje6Uh5hr2VJn7q2atYpy2ASkoksn+MYlZ95/y9Dldp3zjZ5xNV5L0PfaokzRicGDyXit0so6Ky
DYcW3T6b2L7NVkGgKlZoz6py+87UJ6lzJsB/hLG5faMzsblHO8Pki3kOUzJQ0sLxWDaBOJfpDLiW
WWChHtXpGQ+EvMqvLJRieb/wlS2g2gpbU6PhovBfFtQcXYAQ5D8xK9vLCXf4Iv4N0HDcDRlmvU05
95KXcq5E1yhMdvKfR+dZlxHs9jT+zeLIwFDQ8HaDr/lg4m3whUrLAWrZTyttdrf0b+nDVLlpPc7N
Tpq2JCMA8yrr0890S1cSygn28ps/7WP8dJ57VzrLd1dY/OR0eD3u478CddsTnSOpuAexkD2Ls2G+
FEDX0JSuQwXmN9Qo+C/bmQ1w+U3OSCJsVcDaRiKlrUUZZ9GRgx1RyzZ2fgJCYzYklp2mOJQW2DyK
hRkiWnaEsghaB2U+Ji11mE0EvqNpAGksouXGxFvt8lmXLBINv1oeFeGOJTHzZt8qMXXkmN133+OW
lhwIigrItS6iKoePL24QOcmclaRbqqPEpZbOvCTzdcfqLnvswBoh9c5cunq7sJGhu4MQfz75Pbz1
vkzXeNj+uF0LAL40ZyBtSHUg2MijMOiVD2NqNfhahtiRgDYy+Nfd/wBcqJgO5jbqGrAP85o71iqu
KbvqGgFZwAWykeCu9yGtvtuL3zSHOU/H2cs8gx9Iu8B7YE6x+OlppzGObX/bP6FcA8azzDJVk1Dx
MHia4Yhx7vam+Y3jRqAvFRr2fWRbCyD1GtBNszpLxk7mO2AlZD/ct5U5jXFixxWE5vaM17qJIYRb
11zB5ih8ozmTlMj+vKRkOCaa9qOgkq3mWzI4AfjWHzJ9UfUQdE4dZvkRVA2LQVETtG4sx3oBfqJ4
w9j69nuNVniCHQ1N2PhKLtArlMo5iszH8ep7knNtHiurUY3MeJZxZEmhmKkd96V6GU0SteUhgefz
CnlIei20X9aoEK1sL+C7YF2J9NTATX3gDz7WttRReszFT0x5/GdOt+0PKcJAhHu0h5JRGv1X9X7q
Axw1HyT8LwjKLUX253eRmFnqipc1qDjH6UZEpohyq5Sltp+ZG0hBUB+WAb7U+cvzTQkncHBuMk0/
R7bU5ay9w63859CuMTNdbjAu53OMzpyYe8nRd0zxBwGmAEurlvoN1gtH1WS49tf0nmnSU+nMQJcR
BXxMjFNtoty1qbxOZId3DiHsvcV1GsuugW6Efvx+7d28cyqqTKYx9EFf3osL0L0mToL36Sb4XQB9
OKA8MSDbtluJNrvjjP9n7oJkGhTGJp1LLBKcxVSGKCmF44zfAUaOK8nq9Ujumss3pfSuF0guK8if
NK8XfcMjzsK1k5FGRrVz8NiwWOJDm9MZnRCem68hVfhDPBG5fN9gfZU1IqaaEwnsdIp8s2gQ/OlS
cRbrgBK65iA0wbkeJ+ke5ll+HdTmQgpv3AWuA3wvDEa3ORfMEQ6hJEKFBDrydewSNkEFeiPr7eqR
iFaaHf/fMr9QHO7fZZi2uuql/sfyOKtW3rTFDYqCdZQAY/Xk3aUpHJyEIOhB9yW43Vla50xWM50Y
mqpAeGN21oup2J+hvIX888gcwwh2tJiYSx+gJoTyZE/IaKbOd04rvzXHgcdZzawgibgYR2MoAtkH
9zTAec3TWTF5WNe2Y2fuvm/Y2hCcmnG5QeDpjl+oMX2QVbG4GN8GzBpdZjhSIXREK046yr5RMxTM
hqXlwpzhrWjWtOQlevfrwPU/Y437FswTbEKX2UUQQVo+cDGiYDf6jZN+UoSLnVcAcPQ1QkHRFycw
nr53FT1hgYmO20VXD0EKmh5+jb9qp1zNOd77Q4zl3r+vaTn2YlUzW5dsezkmtGLcIRfPUXACImDQ
m4YCsGsNYzqQjwIoBSwIH93GwdnRSfIzxism1GgLEl1d6p+KP6+ULJV5YyQzq6FJMfBxO9QSeRmc
L2Ksp7tbvJw129NoQlf8n2/UMCT5z7IeXdq/VhjuTUjBHH2VgKG9Y1F0SCsKMXusT84/Cs9TKV8F
idULHRskxXNoR5LeMrM+JnlJG91w81oV7hz+FXbGWIscgFHBE1z7v8FO3OjKltGkWcXWBRlANOcd
PVhZ07JUpsiS6yDLpw2kS5/r0gfOggB2akC+Cr2FwuFaWxoGkrRHuNfS4yjxPYxwi7nvbJ9esLG+
797J15E/u60H96/f7f8EFJCHOpEDVz62M/XUskABTT4+1oFEI5IRmUHKmVw+w0zqvWjMU1P9K7gY
DKO4QRES36jgilB4NSIKrbIHHdntrqHCVlhenLBvFz9XJJ0RALZC4RnCmF1oQ9m2Aa/tInrvbCe3
yccRQ/jgpKMme2bfH8EWH7lbBnzXhFNf6QjXN7DQ+594frB+umqvaUFO5vuuDxlQCAq3AyJ4nQvK
WA51zEwbguj14wGUjt08CsxuBPydcJhQNcODc5S5KR94SzZLd2PzunIH1RjFdNvhdX9yfiy6Audz
TYe8FN3oydkJuRodRUvwG4+bwAZykBYxxqmpyuTRxv8lrxwVTVFbqm/RtgUA17ZPystywDKMxot+
KLEQ+9pNAgAKWv2Mav7W364xOJSjriWul5CHpx7KMYem0FcdmcXdUp9pFKdoylIkOK7ndJE7MtpG
10NxQxVgXjHG8y/7a5l83bHPr/5ob43l+8q9+3EaxNs3eJGudFjGAP3chwFQffdRlMHfMCdCXp7c
U7YcTrAY+jMJRykawW/rv6eSDJYejxTgT0omgOjUzhIW9Z08yOwLlj7pVtv45fUVOVyjr/eV9Rpu
Bn/dfoFahACwG+W6HiIZRkom19ssF3lOQt59lwDY2X2w7jkidN/KyoW4jEqLQ3+fHabs1j8Cccqd
BCoL74xra7ooTphodMo2LnwsCY3VxRn2MJzatGstj3VQkyTe98zrxMTOBioZIzJactZ0Bn4uYWOM
VSopQXUL2Ozd9aHiw39FKyIZsNsWg6TFyl8l8JiwBwgHTqp6U8LKQqlJ17RE36Gex+wXWodGT33G
QWllZjC3VeQtlxaFkxf9rNJvAiWhbQE3fEosYmPo2a1oYWLD+Imq9SJRyeA81tqPOIpvU06Ll0xs
OCnJonovzxNWsTM+eTagyzOSC8YwMJSXJk7cZmxGmOlf4vu3OOxcpMyWukEhYkOs1sVF2YCyT23k
1odbAntk9m0xRbgbzKbxmpS2za5JW34mflSclzWm19UM+SXIfnbU4o+hrFitUochtL1uyUqF//SL
xk9zoGxm7J3D/yTvAv6RztLct5c6Yg7TUcOBoN4AqaoHeyFZF5lM2ztqdAlUbiRF0PHzQA+2WdTw
7BD1kgYuCil1fvlol8rl/HrkIo83HlMqVbQJEyt/EDqBurMnGsAL0sQ6lJuUNh/DvA2CRo5ixmkB
2GCx8t2RGm+1RdFau+rM2IXAzzfOCU3SKJf3/zc45FV+0ta/nrhlOaWpYE3C+QbZNxLpI0cH3Sm+
wcF8rEqg/OgIJJVL47obDo0oxNV4XuijvQF60Lu4XW8UN+X1GSgNh8yXz4Fmguk+FS8fs3X/DrIl
QxieUUfBAmp+7nVNK3hulwy7rcrow9O/NV7l5XTGfaVgcYdi/cGBVBnt/Rxl2P7YbE5GLSg44/d9
w1MhaocLIKfCwBTmckFL8WEdi0WTyEpcp1ke7vPwc1R8ObOwo+/GWSjU+HOd8Yj6jpaXOHAPdMW4
WoZPQZc4w8avfBdOnTraPLevhCzrPWPJ3ccYl5m8tDz2oKTLxXNZOUaKkX5v8FaGbaSGMYfwqq++
aXfCDBYhcZcrvVyD1fy2VugaQrOa0aup1/SxRoA1A+GWxIfLrThjwgswbLa/rp6LzlynwTponJD7
afM+IGknE4xDo+UMvGTGymf6h72/VRYaI9oDTtez/NGJhHzlZmy2xPI/rkZ/wC29LfkOgqyIElaL
OSMjba5jfamw/Lwt4bxt4Em9RLYWvM9i2f92NFNNokozMOaEeAqH6JcQsPHPZalmBq7lFpgisfYD
zQXdUuqxHkVbJ8c/O4IASPPmBTXKwJDRhGc8ra6Ngxm8HO3CjX2CyfMRj6+bCUSnfQnVmRe/OTaa
lhR9Xt3UL1FGOepyYKUzDtoznS8OXrf+fCZRCr3wJq8wVKEv2KaqwTBK3xa186Cf3hlKLah7GLBP
NumElrbsTM1lA62KFHcaZo1kWbDJBrXoobrEC2D0WFL1Rl53pUdOwLVYSSukR9+6L8YjSxybLuQ1
SFoGN2cinndmmtPysYhnHQpLoCvAu79RNh1pp4UXjdFGKROSj+6ZPeV4Q8yTh4/SXS5mA5XMpERV
vih2d0hGRsXhQBDq8pc8f1canmyc4J0Gf2vGnXXYx2LDIX1di4nmjWEtqVCuNV5B/x/Shdr51zY1
JqXOIGESlKcqbNmtRg8pxQjhOJJq955ChCmJz9Gci/Gc7mxeEInAL472ajMKDxoBT4pzLOtOIODc
QrD4jcyzixWg4He6xnkGwlhwwkjWsA1/Lsb09k78539yrpVfA4lPVqX6+8KnLrVE7oUBHRFSHvA+
nDD2Pl5yy+GyJ9CF1ch//B/iKJwAiXeyIwAvHiXX0qfQT5Lh3WDOQetEqzqfyLGnwQTEFw5npPcT
SUf9RfKP9uSIKGH3M51cKawQ3+Kb9l8L6RJjKrpJBnF3AUVoLmrpIn0P89OLHErspkWQjHnUZAD5
sZ7DWcafItSpVimWqGu/iTKylSfBRYljdflwRTZzT5X5RoiM7wFITwqX4B+KGfSV546uEMpvajYu
vOwYpFQihnnpaIbFGwxMXLLtVqj3tzoovlOftL4GuTpMylI7czzngIf2FkXAo30e/j6noX4sO8CY
k9aA/C8A2/W3wxknO8TDLj6bqcQFkZ2mZCP8U2PuWFsBLNEU4b4c+8Z7gm2bmPhA39D40QRzgz4Q
1RT6/Xr2PuhcnE2t8DBaK4YoZzMjj/DvG9+3SDPw11lqzVF3zrz8/7pftGUaw5EKw8HNayuOHC1Q
+gbsu8OIiQboPkYlKykt4O89RpMOZYrTftteuQ/00NrsW1GNkA/+3fADV5DaGXE+ia0RW7WfGseI
Fr7QfLzl9bExXil/V/UoT3FBt5s8DK9hI/7DsatbgtfuBOYOMJ9z9yjwF7IREPx2kMCZY1NXK1iw
tdOm0h8T93vo2971UG6TmXe34irnbNh8BtpQF3ObO4r1cmIcWXanqOoRltGJ+xfm8cFO4UoBooJn
r5TJFfMwLtiP7FcHYqNPQFMuv3nSHa9z8hm0e9bBbcot35EC68/jtSvej0bppkRI+LFt9NaGXYcQ
liEowZNwrD5NnJ/WeOsss5APooRkXD8NRjurCgBKu4GUm1YPdKWd5vh2qgjA0x9MI17IGcNmZGlm
uHHDGfov4XS9Q6dB1P1bqWprm/G9yvAxeG1Wvoq12hmahCnDTwgD3f6E/mCSTvPimyBex/cja/EM
/xwdr9HURD3criZhvzoSAIcpcrxA4wjW05lRzo4XLDjYvgVlR0PJtmXrYZKB1BKQcCjZmBrmvbUm
oAKnwE2MzoexACzCc4sG46gssmiQHj05+TYINbBhmOjmaBEGkhEdD4MH5VE3roIRL5VMQGrloPKV
m3q6Hq/VxV5y9RJzlc0s4sH2/g92gPoSdhCxtxDEF9eeiY8+27o0n96MkrY1VOfhBMlrXOcdG8z9
fi9PGABAKmqJfBOosDH/+qCRBVwrvFI6uRJRDldP8DRr2PE5GmDUzNTZfzHuj5n0bF3FTQ2MXebZ
tqiSR8K8sbfMfvhh2f79RkQsH2ugeIkrI77H+iMaQNY+dYWM1mmhbW0NVUjHCK4C+Cff/bozMzhJ
ThoJNi3Bo6Yguku27rgL/R5V3oA15tmmVtZeLcgOW5vUa5OPNplZ9AfLglJoZyxkdIWG5kq/RH4f
iY3MUBAlBhZD24xJ7hBDqLYr9llkntM3+fjAjqS7qzKA99gvz2C234ly2aFobYZ0S49//NolWI0x
1AjRer5wG6tkukXbGaDiKEf791e6uzgWBMB/MjDZBtJXnTFTScVJgBY7Aq9W3iL/e/OLDPD39Jpc
dLlw2XCCUTr3cDNNGdygShy2py0207kqoIiYYSxGe/+a5iSHXLhJCQHLDRc7uwswlaXOIlejbZw+
KVW9ef7R36kmZuwm6FHh4y/3TNsd8Eh94HAeXhHZsXDOdzn3YjKK9EG7djpEDxkucsSW4z3TPqaG
oM9TMZddZuA/x8kfXYq3FlkFZOxGG5kmcfl7ojo6IdHgzur3Mp9Mym7WmfMR+e4q5nUVK7LFvY8t
3qVYVU4v6xVys2H59quxnS1W012km4X1L3HgCQpsspUBjpl/4PLSB9bfmP0u/jAMBtiZmNOsvYjb
h6iJlH40zJ8iYb2VpClG1HhzYRIQTxIH6V6V9aIZHXZb1STGhErQELaqeTRtc0lwyVkdIAMVLNcw
ehG1kQq1iiuojVTk3wPNK4PUHyANVB4BBbDk41xfKXcj70EYwG3lRIPJv8uSHnrr8zCESmvhrGV4
wwK7BnwYsrzkv1McPZ9XKhfDeM1r1g20ZxhbK87trYc6UhdOre+TNMvnaq+ggt+T4155Ij9BY7yQ
9mwZmRPdD21plYwtjbJNjUDwBRItKbUZq5f/XBR9F7g7KKAF/2rappELrLYHFz2bSD00bpwd0eb1
8F67dzw/OIEuo5m/EjYvINJZ1OwFic1j1bIP0nNEUldxs1NCuhbhtKdrTUhFfDcT/N3TYXDG/cIF
FsSjh22iyHvU8aZg9XBsTT+lSa8CFoPJSxAydSLn90aa7UH5g0yui7IXUtxZALwq1rqXWNejEeLr
7EmjJ8uLwldCkfrw8VaN2ioWpzhO9sISFZS6DOEw1h9kStyMVp/CT8LWwZrc+iSUpTBnO1/1N0xp
LO945b9FxWFi6e0MkuxToxG0AKKv1uCYih+Ph5G5qxo8lodtyIDNAlZbq6ST67dFREdSE2FoGad2
sZFhTBrvq+LNDyW/cqjjtVucpqmWa1k86ADrwVWwehjWRwRF/9H/PZ7W+TerUFt5jaDdzI4i3gmx
hpZhGnWoNbZZNqLzLcQ4u71u2DV1WK5ebYGLZIoLUk8uVQuuMdM05UVG3+gzi4PWT2pU2/0bzU+M
2K3YtxBxwYd/DVFZ4q9+fjl2aDwYTmCvkQn1Zc1qYOhPPQxtPdE2GI4lMGIXi0nfSema5KfZAaBh
TgWz6doda5TI5IRBBlLJ3SsbThdVKiSUD+HxEFxY1b5RuuUUWw5PQJ6HPn4iWxWyUs86fm58hkdZ
c4MuV/M28Kr5v4yOLz86Qop/WNtexJV/YptdX6FPC4ydI8SbFo4Vn50/zW/VZpvSdGh6fAiZisk0
6/UjENUQ0Z0cVj0oaRmA1URlPp6zYcxgfKHOKOqSvOWBd7m7AUVf7SbswuvFyM+jnDyxPAYGp9kE
/qLS34FPae8Q8Tivzmr3RcfntV1ZSOXpN+reiOz8REHRjJZtd9eqXqzpPcH1D90s9qa46+gJ0VzM
1MTSbASJGhHs0Y8quQwLImI0GDhcc88d/mgl3SUgcr+q4mrT6KS17spIazegL7guQpkv4+6e3pAH
MAaYajON8oFa0GVoKKRFuKwBpcMjGTfsHdXQXt7g7P5B8FrzAw42p8Hx6+XqyM+5kVoWO94/ebWc
45CQuaMHJvV8jpc8BlL+rUaOKUnZIDfmy9/FRZtCiIeO2Cb0y1ZsVQhRVBuWVrCMQO+8Ab1v7FIE
4CREXjM4R6AgzoVR1sQ3oVbyP1L1kvpdU/hfeSgWTCkqmqnE33fmaBGXwVO1NzugzBMmMHcfZCcB
Z+T7NyhL4upiKbofOkZEgkECtywoq/9LncQusDhp7Qlbq1KGmAtqdLXCTnXNjDJ/DWrUympnEbfO
BmU6imJLTWxi72X8HSnds0rdTqu7ZDshJSEyuOkeQoI0bLlKdb1X88HyRV+9caOENoNJX2+H8xZE
9k2BwT3urSAfe2ZwRFi0rZtUfJlntpr5MAVwmUm97UCiB5LYTuOIYE4Cz8CvRUvyqzQqUqQqe3fb
IG3plGU+1g4+PMl2SfXxkr4KJiF2S/ZFntbZOkJfb9J//GCHCLJDP3nHFYGQMZZfYGsEcW1T3SsS
/9gx0rL1cZVhqzJnxkfousu96oNUZZEbAqccneUt8jYtE0ysIB91ayujtL/KXLeeWDFnyVFqf0mk
JiLtz6vtdI7qWythT1Ol2AMv6re9FDFXnDJa9ro8RQi/RvetJIcLFIDCrfG+vC3k7G3Ru1DJWF/M
O0TALQiONRqGEBIJa/VCOsT+8DUi/NZXckUrpaSDZ2CYjIxC+OZE+BW1uWfZ9VhJeDJqfVyEUVOO
u7WAN0C/IjwzNwxBp4ODRPgbVmLU6uXoyh0Kh7cRiMXPV321ZClHA8QHCf3Z+3gAkPx9XOC3pK7L
8VYqO33ybZkWcejfyJDqDJ7ybGluTtpL/EaYwEcFgq6hOFEeobzIjVcGKVWWyReYFu1G6pafJBqZ
Kxy5K9KyzvzmRoXYtGF9hY/7E8/TcXm6/QUBmVcLAGcinHoEb09TCvCYcIyJAGMaXa6waC+2G71p
BnZAKYJ1Vxbe25tguTXD1ZRl8Tw7cwa0LfYOOBJSyOmyL5+7OPeUzdH239bvoCI5BRJM1IncHsJu
90Mn5bG7wdUhq/hGEs+R4xtzp5iTeX0I4W5X/BcPaw1dIuimnzDyRfrxYYmJx21sxQSebOV7D5ut
8MEx8ORlZNtSZBg07Mg+4yCrsVMiwzX//odXiSsOkgKTOYC/xp33SHg0sD5S21iqHbnZkeqxP/sB
WbrNEgdWO6oBBgsaDxe258GdYkn9IVcRmd+Y8RpuWB99C18iPwPXEapEB90aHuFbfhep47YUSE4q
e0q74r+5n3pNXE8+fxQ7TdIyLGBL8+zDc3s/VfNAoyZG6ZWeNLAcJKq4cnbqBwcaUgLCOFC32xjc
detUXFMnRXHbewxw/WAjAd+pHatO9hkKBhFt6nYHyemINb2e4Nl/yGmtDQ6w/3X91FO7ArSXXXnv
jhqA7/yxr78Y9vQHTy+Q1puVAiKW1z79Qds6LyhjV0F9xDWZQATonaIlITBRCl1myB3Cud/G4sWI
/bIH9s/C1L1hzSrX/yjlxUg5ck0Fmel9bzBBETXOAO0/sA8qrLKbRerNz8aRt7nfQ/2o0uyrcLOS
d0scJBiRQVQAP7PIYgG7yrWZW5FxGyzBGzPLnPKKGHFuCjrPg2pfaA4E2HDFiGc57StfNDCRnPIG
3OnHqyAche8vnN9y3JxFZWMjDiOT2PFIqrm3Zsb7TPLoGLrHskxTymJQeUO8DuuIwNwpLAFjXBoC
WNeL3eQGO85kmMcJWmKiwl/iH2y1YigtJBhSK+QfAI/S6Kfq0Ptf8quRxORaST5wrBFGn9Vjaklm
CBpcC7fupx9QWoQrvA12NZezsp5pqdh3EkEJVqGtcEuxshmIIkRKrahpYCIce61SQAUyb3eLnShD
fHqv/j9C45Z+tfqLbbEH5ETlsVF/h0ekhyRNZrgr9zh/lprMGDiC9tuz14avEwA2K2bbjK6iyIGB
7MT40KJ4T6tAoBi+OcfLGhM/rNjux05fva6vDcoKW4KVJNtNa35aVF16lMp52+IxPDKG293zjhUo
629JPMOF36fts8HK5cCbZiQ36/WWJDruyKeTpztJUpdn8DWsPsZdlAbISqAiXTamxkZmas5YbjvH
y1lE5uTTpe8BoqY2mMVwClZ9vn/T/3rg/JRdmB/u1/Deuhe+A9Ci120Q7y06H8RQaiglgKpm112z
Ku8N+CX8W+3AiN7dBElIh0pzFLzDJiuW6bQa445ktSdXG4gQYPEDo1se7eK64mhmeSzCm41BWJTD
MHao5nBTnjEON+QkBneErPlLr27idtyWJ2J4CxExCX8OBGJEL699OFCtFG/l1vpepm85oOJ2/2CP
jLaHAEdon2efFZB1Xp3BIx8LO625+BBAH+yFwh2NBvDA0e57BAaKorTdh6LHA8UMw3mwAnNK3DDL
nCP0MDBJUymCLbmoK+vbH5lmulrfmWc2IDIqyf4Kuruvt+/Xxho751ZQvdynfBM7dDMTpf+shNnS
+SlKVKfXoRvP6T8YIg015nKzOkcZrLKoC1m2hT4X/gA25wYxVxs30bZeZQwqihYuZSQ6pFVu3I4e
X2tqqrcq9GnaXWdUW6hx0ff9J16LIbY8SVax26qNDWD4oq9WMArwemerAT4y1RI8Mkdzx26uWEVL
m+CS7haoJKlrpRRTCdESThQCeKwoRNA3ODg7kPHIELJzyIrxANuaX7BgAGWZGd4NfEiUZiz0U7Ph
jCrCEcgvNTm0IJtPAdjxvPlXlnyAhs1/CI8o0Moxwux7G7X3bUheKpx909UTB1XjCDtxJIFH3pjS
v3E0pL5WAekyGGWWdHhVi5yria4PhejqiqQnViuhuFbIBTN20ozODPybdqu2z7DWvqnxFIzQfRe0
2NiUTmylU4wurKLt8M3Wm4AfXZXU2xkcaxb1YwJb4iuT99F1N4jMiV3rPA+W7Ely8GCbdT0cZ48v
WGVKsv1Wf9tnaBSdBuV1xgP3qts24SSiRX+NvSere9ljLV3c95emCEFgnGd/nqJEds4oKDesmlYD
qaqotFtCoAbKJUe26UcqcZTKh2Ot+ii8xpCePWwL6NHktIFPY+Dy9KbElQXa9dfGKqgjm6TzUvZv
aSxevwJaYW4MWYZeGGX86OP58ZlCAfnrXh241TMzjp3BWeK3UvpFuC23tbq/KTagvjbrfzOdm3P2
N7wLmKPcc9wqpFSQypYRHWO79GJkIU+fwFaqlrXk3ybuURLLcVjHZWQf04igO1lx0iH1ZEaMNkiP
km0EXnN9TEAdXBNKgupSv0VCA8qnS8pNBbthvO4+mrK6p69ayDDYtPlfHg7nJZoTJJPMs7gILwGL
dC3llZr7BBEMX1k6mky0739z3w40AYNCyJBhzPslS0T44PP3BzQ92IOkvv61wBMb+bheOR8Zqkrb
GEKdbXSYWYYRfJGWQ7dJtyAPBTlnJRpDX68rFdEHdn4T4zWN/b4NIzs3bigJGun7B0ypvsBCZ7g2
7kc13Bd3+wSw/axfAfX8NIRxH2W+AeoRdHs1m0EKRUcsA7goxCmP4CBzwcG47ng+VwGW2klbcKG7
Tevo0oCza3NrokR1XAluSm/C21Id3uJgb/KfTya6u4xe4ycaEJ7wNxbGcAG0d39o8WL/CjWGISb1
bOVxAiEUkLXf4cfwYZgx4CwqRVvTZyMWg4ZTlgnSBt3vmI9ksFTj/OG5klUkYudhCrE8AdkvfhK6
jpOG0O6xbfsT8swE7spc0Tnn3nWw0/ROYe0ubAnMewyD0RovTcS6V4aoyquZ2V7U24HIZeFRXr2u
ADBGmbEzoJCMZu7aT00CoHEyi4YSmI2JbaMvvA7BkV9vVKc1FlJrGDRTqNVTZvmXapRfeioYfKTa
wSI2jX5EphmbI+sMFlum7XJU0EFvIW0lEC6AImFb4frkE7GB+aAeDsQKsvnKyPm8BQNPzaiToejt
nP3jJb60qCCqlfhr9i2Nile2zmW2Az9Wjvmxikws23Bwpg8/uX9FkgRv+g+P37O7SI5FBUk1ppQQ
UFs1t5g2efy8HP9diDSQjJrw/IjOa9gdhs9fP7XTtPY8v02KdFotC/qH8OMFjLCQMlKYEKSQc2MW
g+1IE5zW5mEvUUOuFhc65etwxkA1yp9KCIXqLii/Ah3tvZ6oUuhpb0W6fKFO65sLNuqUE/6d1fEk
9X8Lf99uF3e33/iLj2v/hoSuEQFHswZhHU96j/gi7mC1WeK/DDQolu06HoObloWgZFYxthq+uMhL
9iLKUnqb4Qd7asA5FT22pE8pp+2NFM9V3bTzqTpmNQAqIAwah47toUcE6YLEbfeVjaxH0wsURgX+
P6Zo8lWXIXG2CYWoomcwaZ7J+3TfFPfuzDg7RVNWPdMuZ3j/i41ZejvZ2Na5pnDxCMpkeafEWV19
GnDnAu1XgkI1EMVFy5KOeGXFVz2n4UL+sHXyRh1oN2WmoasGxI5wNTlFQB/xBiEegXj+Dp9qVF7q
HHCcBs6WFVk+Kj/8ZW1dG5KbzxFAG38dLuw3Lv6NJTE9zZ7TMXGELKIuiAmxkCJJ25js8/6oERwm
BR8BLc11i9g0fk8v/6i8v587Q7wZoDaTnkbkkrQLFvhJqXwwu1XCNwjV5Ww4lpt8+AjXk9fuFStE
X84EZqsA3upvhpS0iykf5eNzyoKfCUnjGDttT7BK55A+1JAsb1hzZpu2fF2yR7BVDEhh9vNa9C8R
nzoBcGHTRQ8C6gvXWrF5W6V+Kh+V3k85Xv/k/v++Gja1ASPbofizy43gHVx15Lr0rUH3nCet7ohk
0/dy2oD6oU3R7NHZAkkpkcS5qlfknetOV/DAMIFXczDPTuEjTyCCMfZBRdnlhGU9yjZ8iqe6K5KR
j/aINMDyRW8gc5yLL1qKE7v6BKh7uw7beLj9xDX2Azkotdv8sl39+IVWtQtLdG1QLxealVLTBwT2
PLoxToKnFUQUYeD7LkOQIzPa1jHPp8hsxLlBKFO7AA3eS82NPqmD+uy7G9B5clu6ihrJNnqi76WQ
a3TalKBlTZf9AmF6gYxF2kDrn3Xvh/Md6TaCtvsxO6mAHz+1ZL2AgUvsXHrLxGJ8HsUY/wd2d6nq
Y4+C1cDDlf5PcddKyzWpBumxJYiCsytaQ/hasd6MKPTIvVwTfW6/VktQw0b+p/BKEb+Iehx7uE9c
a0MizvBV6koA/NGL9AMCxtzKJVAg1YuXamRrlJnAOD/VbldyJrukmXbitbBew6I6ANpCI14zsX10
lznINbUYUza2uDvEqiHC7clvf9GRLlgTkaIoMymlE1XWAQghhbGbhk1Ij5DIIxayYK/fBYYWQs6J
AcPozA1nIV6vRIjuR3pQlCDsM2uVnTJFsvvONF8h++mIQ3WewigeiDo9ZbNCvvl497k45ddCLchi
nsO/l+/LEYFHrthMX530vlibi7GAjXTFyUtLWW8sR7zBbdPPXfBqPRSz+tmU5iTrFPLe1b/j5MhP
ePUAmGI5nNVxukaZTZTnCFAi+0iWke0pyT1cXc9OHkRXMA+pWT3ADHA39ChhAgZ8O18JSStF4EZQ
YuUhEAEzJKEwZl8Pbnf+Ejv0e6FmWYjvyEib2xUGTABX9nEnEoldDSqnb849bBzaYiyq80TX+l0n
VMNi8q9umkRpUs+J68E6lLC7lcN4y4IhBB1tXND7cChPQ3OOAH+6KQzb3jrBK4GtldLgoblqy+yc
A+1ntMuVjAcBYjgJM7uMuqONZIjWgBASqhVC4vZ/vtS3FTo9VilapLqFW4MzGatwOZGFkrcGTRQx
ONVgWUyaROH9yyodq1eHlGxpRlWSD+l4ZdJi8DCMWTuZe8zOv++K8+uBdVjCeF6t0s53c6Tl7acx
5KhEN6a9mP0lCb5TAz2+AAGYkPGoQGHflkrFDVjwJpzgCEXLbOz8CHgcQxZV9SZD0o/e+7kvsc5M
aITqQZahQYwaTMCieHVPUuRh8sRVAGKiBMbjwt8ogomg8LwvOrGd54/r/P+lRS8cBp86+fKKRcny
j5cGdW+Xtlx979lpnZGFqD3DEWW5aEiH/EWHcLD0VRPoe4FN4Q2EBpfJp50Mtp7+MWwXFlFmv9sS
WFuy+GMqXuONEEggHHP7LyG5P3YhwH4TDt1O1nUXUCCnvN/oMd/eg7F7VIvgq4ArFl90awGUVehu
H5N0PDpq8MEzST4jK/BdaluDsqOe2Rv1RU+n3RnXLv6c5l16gKIKZIOuXdW3RmnD5or5E+Etc/Us
nSPiuDzDvzvjsJY8C6WXKYwxeQQaB8Y+7mprJ7f4pwm+YNXENbzyMOtM2LWPJ4LNSdhqqcNYguXO
hMzfhHtwkk+23Njr6ccyvHHeRPn+THMLKUsNZNk+5cJu6f4Y5z9tV3Iq9yCDyJXzUmswbmQX5qCf
fTGNgw2hcqKjiHy8mVRpZUdIhmCyxqbom3vmYd564mREupnHhBYam0CMv9lG0ezwHoh5Pqc8uh/I
EB8QobXVO6fpcOAyseYGe/uFp8pdG7imCa+ZTis9QwpsveQ/R3usyMLHTZVCjPwuAiZR8XOaN1k7
Orf+esphT7NIhHw4awBZjTzznKrUl6FiG4xXI88nPwwe2DEf4cn61WvBHCjgPkdcB8AMqa3tiY0o
ZlEb++xwskGtVweU7XcDlbtRupuozbyFYZ/O1PFkIduLwLxn9g2AeBUXq52oqOjbOAUfN81oGRH4
mOwEjjrQ3WJjx9YIG2G/DlOBF26Ccy4B3z+uUxJUMxFH/BzAFK4+h9EaoSvSFMPRiu8Qcs9K4Zlb
EebGE2jR60q7t8kMtHLmVvofBWE2lOi+c6PA+jDwDT7uaysnXok+5pTxGGVP3V9MCjppfwJkt+/2
FPRxEmmGh74yk3oWvYpbPHQcIR6Hz0LU/esmM7KS+lEhXdVGvCMVjFtelpg9rs9v4TOhfU4OxIE8
gcFYp2GYIS22osmj9+WZdSTOCyrtNoOwfPImVZ0XXukFsVHrGek8sYyEgTI+VQbhLhM4gLVaAIb9
crAA6wlflDtTXKcJcHk5HE51n2ecYt0TlN/tcUoggDkTcb9N3mVtN2I1jRrpr5wdjuLkwEtQtAUN
aLcNJrfMwKR78h1Nx+IQFt2U9RYonbZsNh8y+0GE9aSJjD9XVAhMwYoDAPjA0NnPdfu10aazAJDE
w+g4jCCsr9jDpymkB6xNGYMD8cw7IeV+BfADjr5CGL2dcWqmaPGqJ2ZF0yyNL02Q3IYgRqYFsKrl
MNgFLn92/37Q95O5pLZkORcFdUzLVzo4uLQC0f8Vi5FBrs1rjWvqYRvOppx8AuCv+M5lbEmxvsGQ
zhF970zoXOc8rCrNwSftfX/f9JZMl6YQUOk9TaMFPlK/YYLgk7eOEZnKn3SW2qhGpkvijxyGr6Oy
gJXWIc4TqGTiT99UwfALAh6ValayMa8l0ZzQfqyLQ29EfznhiUmKWhdbUIO1AxQJGv4Jk2y7Du3o
QNpCOSZHv0cQiz8ujgoqJBaVIwD49dXPmnfEfHZ6iqnP1Miqv/ESOLRXWT6WUF87ET863QHIF/fX
rXgy7c/JHqNus3xceqp6ZkM6cm490Ac3b9dbdfD5BnyGSel0V2ENDz8PzQeiDL/34YHvS2Yl7gN3
7GHB6Q7poiy6q64MkgW9xZgOM+R9wfITABZ4Age4wNS3FnSsOVn9mdC/Cj4Qo/CLeEXXH12Peb2o
NzK3V66AkCIZSdJWYlsHZP53ZGeLjF0XW0a3YXzg7fL0N3mAQUTzarBpLIRfCRJM3Sr883uScsI8
WVlmq6/scFYJFnnT8p6bh4+7kPOPSZgNd9bhaj1t/cqmrPQimZ2b9JzQs7QafIrG6hoLway11h/v
Ie2F8UuLDD6wtn6T29uXokD4q3U3exHpMRjgvvT3HaG0/e2PlKVYydLYrcmsU3mY2kS1s9px3a/p
qo+qKrn5sJb/OTn2SJqSFC0UaRIzjDXleMSp7bQ1DwyRZ0UZ06Gk+nrG2zgZxuaEzGv/Ijq7A8Ek
saTdAFBGnz8EJDG1UZYxbAtIF9+fbdF9ZdsxL8eVhq08wheVxpvbqFTURiq6Efy6xx2ttvGzVYmr
VTSnOlCtQmeo5nt/w/tMS0/eJesuHhU0NUZ/STSLXQBcToUs8JLGcRGG5hBN7oqoFP4p3yKpj3Gz
8lyVdviCKNf3ID/yFBPq4STJ5D2g+iUFqBKK6cyWD531At9yz2xEF3LhHMx99Nn1PW/41MzJHE79
gVWqiLxBFEQEiUY5TbEVwV6C/3yX2pQgle3QNGs88SYLXNSK65q7mDZPmuyrbmUzJ0oIovqubCWO
/83HBHGoN9pTu625c1J/V6/Oo4P63zlKAewp/7WsTmvlKEOsUzUuMb/rFuoPpz4lLkMVedpyQaC3
yrN/aJ0lCakuqk7Ya4G+mwDDJEBABksl/pN7tkjF6dK5S8t9zjIEyWK9Rg7os2V+nzwimIB98XPo
53DBoBGDEj9uqqeAxi1Kn21zFlU7BWhezq57fjg7+DMBbvZC8i+6tJ4pUaTEdl9J/mjuqzsMUMzb
UGcPgQ3+HMNFnTPP8xzuQbAekCWowyVXhA5kKhbV6Fhp0idCR9OEz64lWHA+pXPS2ZvRbQJYT2T8
Capp2mLZcwIfZ9V1R193oRI7K4iLgfwf4j87iXPsiFECH05MjKxeqDunbCc1v2gr4Wt8+HdJoX9y
A2+J1XKV+snu+yadqNzrl2pr/pklTvlDQ/Viioate10cGwI/OqHybfEii4wAGVpZM6ZY0gak32Z0
0OwvwszoUGpeo33a5c0DVIalzNi07Kh/urI+IUclgVgfsz3ia2kZKyDmX7uZZuVhgTalSWzLz1/t
2SQZu2bK9tNr0OUbeFuVUeNSbbmesV9FIaNtCWRdeJ/3Ylmm2idjYi3qQt8yLjRPPYpP0kXc8g+o
2CP5EpuZZgFTvr8aXPf+QamRVW0ypmuBWy/1T51KudbgJOV6AieqZ5DqEiROQ3hTuPYzfEhIRy/K
JxmzQJpOPWpCymCKfnn73nnIQh1L6VSGJnsTNUDFk6jDoXZnJuP4rbtkLLeR8a8xMhISTjPbsUYN
XzFlD9jcfvMaN2w/OuYGyUJ0AKgma5vEEX47Tse78HQqRv8u1G51Q2SjwwC+Xox9Y6UYw423Iovf
KsCvPIk1jbW4GLlCYMRRPWZxxeDn8YdWH9/Q1ueYYiawxSo7oqBfK3YQJDyh9l3Xu6yKTz+0qKAc
VHNc2LziL/dinVoOiljafuJi8GCXI1zBtMXuuWctn4MPYR8h82L83lkA8W4TcwN2ilmLeZfXCNuH
8gOKXkhl5AzEy1V3ulw7Xo5+KnKL1O2o5uze1kyJqM2kCcyMflWgtWe0hBXxwaPd2stmKDK9ko1q
IrzLeU8qpq6671jYMtRKcFBDFWlhuSV5S2IJPLXMVhulpQkzRN7ha/ym0VyM+qRbeGWryDmFKevJ
m2e0cSSR5YBn6G3Y5JQOP0Fu9A4Qv8Yc2+TrNDnCM6At9ZyYMtDVhjXTpc2WvRJRXzBfcbQ/XPet
d/cZuAy7pjhwtzNwHKGAdA9sbZtqF9SJJd2fmwy2YZw1sIu/VYHsk0xOp6IkgSVNY3R4cBH9Jxkr
yZvz/5nRglOLl364hRf7qolICSt2u+BgXyCVKnSgbJRRW3Uu9fz95pVAWGCEV93nzDx1zCGy+TEx
kbi7WWR+uNGVYUsSVckWqU/y7w8VJqyCJTsm/S1wWsji5IRhHxIe5KcQU7uZ6v8mLbUenV3sN8qU
hXpy0KIcPUct2HVoPnuepROmY4N5nQEaqXTqInqyuDzM8ZB0+aUeXhWosP0EBBGVZOXcq2kjeT2/
7bCPhcZYfGtozl4KtoAt72UXKi3TVKI9smoLaeUlG5dYsiCYANWxgaV0dypeZgF2fxr53fQvq301
64Uhlv67uQPI0tj3a8EIpt/tHCdA09FSkG2iMJJ90fICp5dG5HYrwHnINelf05mr03Gbg0g6UHa4
uOv7PHzJ8ry9Ezpyjka+7tOshsK4Kl/5wI/uezFyyJP0ZTlHaYurVc76GGIHilvkGuwB0CB2MK5n
IyqIcpJ+Q5C1s7XbgbQWc4cMuhlBMfGq1MLGRp0vtMDvJ2Lb0iWhdUtqqhy4cPsRMDCJBxqUVrub
HZcDgzqs+nIIalUWSSZ++D1bNI+uS7DR1ohRJCCmjoggn6MrvqhonDYgk6Hz2RhjrTfW543ThkkG
AvWpLHd/jEeAs9ptpQWhJrj8g0T/9kc2PezrxBK8yUT3w6bc3ajPLqnX8PLaTHpDkamqaNeytFYz
NEJC0I3STJ3LpvQKl9gYVw4Yvvci3grLxJsVQ4fCxBKP/VcQY0qpibIPKWgFCYsDe6oZ2BFrU0SE
T7ehWhsZ+mJo1qQ7ma+uMzW2fpSA2zCvuXigR5lLbmXY7jinj3k4qiWPgD/vuifoDVXL2xzz8RHE
82tMat6iF93O7jK3D771z3MaqFuor5BUhzxUsXRkPutka9HLy8pSbb7A2T6x53XOnbH0whnyYnsk
tieDqlOk93QKfuXQWpXUerQhNfeY0g8gbQkyhByLjh8qcdduuuBmTAhCNuBSF6ko8dXAxu22oK2o
DU9ve4FtV59pPUwmFD2m58Rr/k+ccHIT5Qilr8mvDmRANxK2Fes/sQdiUOkqI/Zsh39bgU0gB9+f
JQW2BZRKJyE4zj+JJutKveLXL0PTEP7Ibgc2sLAc53zXKidMz++CtjTiO/y8PcVAUyJlJpcSrWWp
8WHTmc3z8wQy38pRBpoBgDLiErSmVUBwIeHZOg1yEIPJbaeNRA4EMP8/qmnLw/dUrDmryfX3ChPo
6WQc5oUfAS6CcQgH6wHpULJwSEVZkz0fvnPwe/rd3Abpzj3pv8V6nRmHGdSnpcvw2Wx1PLHWkzBa
X3laVKg0ajPunqtfBf6CAka3IM5xFRzHejnBedzng2QmsrjlyVv05XvIzYtL67d/EErQWsZ8nhv9
UTKaEPqwYP0QJgYaj3SmQeMbmv3WnsGP7k+yPBXypdm0IKuY565oCliSnGOromAweiqUv4V7oH3r
2TO4J3h5MbutP/S7x92IfQ3q3nd/fdWphgABfhlbLFNApg3GuVbOAU+CH5l0wWe7FwZsZn2k3JM3
Y5Exoopnb0qDmZiXRPZprQH71v20vMLaFTTs+EeB2j1IORnsI46XH3Sv5JD2XyoJ1oU7jzGvZOav
0kuTURQzaEQTzvAGEVldUDNZ2AksQwuTJmLnY22kSLtlali/ISlG1Bf4Ova2IPmnmoJf/mAQOfWG
Y6+YsCzbW6Kq7VKYgiSsXRbJLbGMKyARMKXD9Ba506hcI/NUv9pdzy8eIP0K6D3bKoLonUT1Otxv
ID2mqI+qxLZJk64ppQlfa0AL3QrgVC//GTwVfZPBfD9z8MtI4Ivi4kkJCgP+lbraxIyI1hC4RyYU
r+dLor/dSeGvkfcb0Uw+0KfsZ2PBfel5NGejSwUBH6ewTzfMeJ2iPxP1mzsyzfJO3y4EqoIjr0sk
jgonCsXG7PtiYxAPBncjfO8tIFOdWGQt36u/I44+t5kAksvK2e+LQcQwi8ixBscR+XPhaXDa2bnC
17vU4+9wxBHb8pVksGbcKBcXZMfGmTusXPfROuXynYtuWAdD5G2uYFxf+xnmUIlNaLoeNyEG/925
xUJZmyIfqBsqQEE3Bkz56isF3hSCwxGqSxtSpCkLx5cigGBBRkebW0vXEvnQB9EWyCnsWj77CnEB
xwtH3GYdV9pT06yTk//yXCdOvZVPLcYl1aaDLcZ+uvmh7yiaSlSdGuNoLx7VIFqZnbvc7+zKfXT5
SB4URSE7p0N+ffSxoiaKI3UjBaQKy+u/zIAsjdPsX3b/M0DmhJQ+LLj8oRbwyEWw2VVHkyTCzhn+
E3qtiq/y9eBIVWtIU0qMY7pd/kL629jv0An9Rt9DxxWLovz7SyfrfNsE78rPnCozXWnOZDl8w3z9
Q+p6q6/43YYK8OPipQ4du0CSirf0beCj3Pmh9Rdk4eHZNqG0vuY+dW4di6uoC2XVOUkPmU+gWh9q
tgiChICHDiF5mNCxY52qF/QHB5HtcVBIlbZ4fTD1dgsG7lnVKHG3VgdLXcyqRHSZKX0kNOUJ8g81
Z3iwWaIWau1vAOqt1mIbHM8S+Le5Tt6XiwfYNAnySrS8a4UFbNoVnSQhgdEWAR7mmHiIvmElOEZJ
2AgDLaBlpbfztf7UiVHi3vZBOiMVcKGhspJSFSDMikmdSz8+xSkyJZ4EQPRnXJ7D0E7xFudHe4aC
X3pgiKpbz+A9tXbI7EkhtVM2OlEtqavTLZWZ9RxeCUk0jFjOO4JiiB7+qQrs00PIxWRF7Mv2nns/
yUYveFrE7MKx2PwZLhY9+6ecId9rNSvIZhzhl6SKy7bKq1xMzdc7zvld9IlFewyTrQQNBuQgZMGz
xKoIXw2YL0joB8YDRogWYa2oy4ZLsSJEZjzVZmINiJeBQ1a1Q00hNKhT/8LqtFMJYo83slJpGEPp
+UtyuFxo1VN87UBflqpSmAEjVEuNz7V83FKwZOO2RjJW03PA0Gh1TuzdTr5kxoHFBJlCPQNdIm3m
KHXZUovoBlWyrq6R1Qwyf8TiibzAjM2YmASgxrhlPVUBXkJNSFLJ/aR7xKquk6v3l8beL2tvYWR/
tNX0VXMTqv+Yi1IFOuUIxjvtS5RffmsdTHhneyFOr/IVf6FjXPuOKNJBhWlisKq0DuN0fIAgcqhk
UlIxrSB0pd58apMHj8cI0kwi0U9TdLJ/gWkjrygKalXI5DkHWIVCYjDfwuO1dpVtD9VGhRTquqDI
VuOB1nCOQm7Vdm2TjlUiyoNOIytO2CbPAjKcmvt7q4i2fOdP9QNvW1V0rHRtoUh8cnS9QhiANSAx
0NMz1CvetdZNIPVb6GOHDVUiV4U++Gq9+eWwhWdtO+1sJYGZfUR6cYCzHsLeWcCIw8khflUHS2VV
5MqWSZ3OjGR/NpLwc0Pav2CtYWi7xHRI7NLcD/9rwM4W51G6r6iUMHMhN+mPlAqJdJsSpaR+E2XM
jnnGvZeQLl6Tv9RtdqMgev8Cluc99MJa/jZjAQVVN4A1WDcPYek0uaQqhdA82ZHLjIOluW/d1KRB
v5gDCX8H3cWko2c1xFbboEKAseMO9ajxMvW8Mn8rVfdWZP/N/jCVWMy4Y1Q45M3k/Q310Btpd7t/
RuDG+eFR8o9R64SijMfVNQLXDuzxxsEGKwaGY5xcusRslcu97lHMAQaDzOlE7PcofZhL/FTuJyP6
k1SUL4fZWvTLRy2CYAY7XacpOR+XkQY7YA/GOrb3EJcWPH9t2695E0i1OcUXYciSXpfPKvJYUCD6
KehmEMTvQYeQlsRsHBCfgCMFO0u37iHoHb0Mk+lVQtZCyZxmbHLePMa7L/yDs+pBnfKRPVWNnmKW
T1beWWviRWiiHXUIcVvxNva2mHw/5PUiDSA5gMIbXzpp2T8ogBIEa0Y6Uhbl+e6p7B3Q1GTAsNtc
6pP39e1jHKsusl56ABioJyIuFX8py68t/anM7P0tr1cmUztJ5UMdD1DkjBqSMlB/685Ndk96/mjH
kza1Jh0qJCgNNJAQiuiGeoWR+DB5dH7QJYY5nerTvNda6P1Y7N+22VWW6Xje39s4/uYkaFEkWPml
Lrn7tE0R0NPI0c6A1+ltEIqA4E2DuKE/XWWIVbSyZb0gBHfpIWhAZu3PNh0rELqVCYnfedbrybbd
y9yEpSkxBhSuBIkl28oguOf9dgspkW/raWO3I60JIK3LbTOWgi9aZpHLtAQjipXXRpmIGQgGMWvN
3dgIM6zajQiWG9XhaNScyRBMbBxp2STPL8RRjKoDfI/Q7KwpZqznYBOQGPTWdkHoY85+lSM/cEOB
rQwHojgiak2BPijSkO7xOL5xNJNVnUgZksYAnHQ8u+CWF6yvhCsKqqxAyYPQ8jWuOcTmiqvtGYOj
5Ap6HAEiyNXGVdmHvUqKInE4CCgbPz2AX+83f+M9eRLrio+gehI/S4vsuA5zkfAP9FOEI8AH6arK
fJkW9ym1t+pfXEBWWLWn1EqlbCy6jPFFmTXZRXFonSqm87h1pvhyb8/wUG9Ui5iYmKxj3R45FnD2
7trh7Tes3okN/ydp+a3ywc8llTts16ZdsKb3vdDmC5U5m8daydJ7rV1schnbOJopJ2rTddPuUzQj
e1k6ohHtzQx5rLbxyTv7YKQlzRUipXNChxBa8fl+oIy9FWM70NXusTcWqrONTLBnOYKZU9j0YiGr
NGg4VGGmoVgVSXmHsTpEw4IZUFVFmZuMNELXuaJ7llawVzPm02+TVI2WK1cGn0xOsfYGeWSJ6VPh
UU8arl5mH88kbbzCS9mr/TVAlQujVIGukAXPbwHCgM5COx8iwSSFcyVD0JCkCMA59C14OpZ6i7cw
SL1+HL3AQi2XVPL1Qf2hGzkC2BahSchuR2TDqvmTyV202VoWKLabj1HqPUun2jpIfuxQNh50LCCT
ds5QyrMqq2yRIueg6y0ss7AMn5j8eFy7XWxeujKeRZnJWUHB4rRxCl6gZAJCiBARmv6hd3FZkQPP
1yr8zxUacMPtCH/GmP/D0aqSiAh73LuCoQTkMNHXmEVqchs9K9vHqGuxFNm6NR01HoI9or1nnqRr
Xm8VQFRmtGQr+RnxPV3pLcKSiv6D3CIyW14i35KM5JRv3e4m24HtPPLFORpMVz6B0kNH3orRkPxI
v1dbsYreQfi06cTToem17jndpb9Yomv0iZ99g8Chw8OPsQGtfu2UsMyz2Fh5O5m7aBa4VcNhf6Rw
at1tSKmBKyctvd0sCxg4gRBHdeaghfRRu4rYjhAcL+QoEqTKOZ9LfgmbidcnDJAV5206BsKJDUsi
2NWcSwDNHduAu8/4Jt135pfalRHlZIMO1euz3W82YV65zBpa5QMZ+MU4SzfsGS+cJ35nhqK3K+Y5
iDxjbXSFCesiHi5bDSA7nZalhBxEFpdtN8hQ5Jk9ncf51IANopfw29hnhNO4wtbeWyuGySFyMbz8
y4YXgTZnkG89TFTSg6qUokoC8oKjuDON9os3xRgQXux7Mykgxtg4zj4WCS8pqUsFgP8ylJx4ocwB
irakKrZisFWajy4cu87CsV9CiaVKE+KYIJVl4BF5pVv3vL9ua0kb/NQs9JW3s1jYcliIUyxZQBwf
7Jz9dPIx2spRzP9CaTPC9EIaGIzblophOTs1OFf5s1pUasVti5sSBDMCdcbJbgVutZeJgpLSEpWL
MUNuUBxOQLSZUo2wm82TIdgB6hSA5r6CflzPZj9nG16w506p1ggfHr4pytgMWUpZNxwfIiRmE5Lx
7EebmfUrQaBSRTNC1y1bNk5DZecKNJUDPHTdEoRcmQ2IvnMh0AGWV7TUbx1jCH1n3ICxpTU+cgPT
//f1+MQa3lHc27MugLDuWjk+PY1D5BA41R1xp16sPvCvnxTWHl/DHkcaRCCn7XXoG90iLxQkksgE
6gedjxyT0xm9/eoX7vsF/aiBb3WH2a4zvSWjQA7z7N4+PUD/KlTRvIz/J/F9z+tp4QLz+D0+c/52
j6MoIvMJS/TZFAxP+P5UMOnGK+bOxL+OzQTGeptjjshOUbuLTjpLrYIIRIcYp8fybrKcCBtPum++
nQAw0dIJwN1mtMT3w5HKBEYHpADMLjS2m5wKmFsz4V/Mnc8qAfP/M/mPUHWQrEhPSljWfugWHSlW
oRb1TxyLeKDFmb7xenu74YBZ1VpaqZNa7uiibNekEH3CUu5CImYI3epvGyXfe9X8yej079L/AFHq
8Gdqe0SWair3T3cj0pPODOuyLxBwQvQvM7u422oM1VS5vxJWvTX6NwCMeK7w5rvUpwX/ptr6hrPr
iNQVX65zKg/0GQr5n7+QxAPU9d7aTAOpNTFjybJIJkDYjQ8iesMD1UpZWHHVfzOGOUecnZns57/k
kj7ktcwtFYXDOqG8sM2estYdUbj7c5eLZWMIQXRcOF0ww3jhfTg/+V5ITr50xmkJnOhWLAyBCoaw
1TvLAMc75cHl0GgaQkdb2NaEhJvVg6vAg622ybq6OLvZ9yd2j9MkcSmTHi7UMIGrhm/3ffgYi7Fb
wn3WnsqibzH88YkRtg3gwtObqBDLTFilTLSYR8hm6O+ZGGEH9Dy0hBD/x2uIxR2NPwOCxMCZ0HAJ
5wqHK06V1P4Q+4knK3YNIU7VOeuUtCSFhVK4tIrk6P4RKZYcunVhh8POCqHjkgy3SK9bX2GBX/sU
ov/gNi6VAP5AVoRTv4upour5p2ghMOnIknk4L5MJieF2wmhATRyQIoeY3DhiyIWi5uAG9bzql1kW
Igv1RTwXk9T0iZAC7iwTtMY1sPSinDiESke2Fip7S88iK+Ohh34kmmDk9fHzDbfI06Uf5eDlMCTN
Tn1Juuk1rMm+5+KChr9uXdjjA02LIyecND62vszMu+JSCZYur9l5OxuqF961vo9vJCdQaOpjLBBu
/5eppDTvLloONQDhbcE5XxJyowpiSjdbCE5Vk9gNrn07nKHI17gBzh8QYiD40h5mksmnrbqSEfHf
IMCu8wB37l1hYAvhtTqFn/apX6XP7imF98JL2VEGUcCHqlskl9q/f0yB0rQsqhDvrTch1osZF0Ml
KpnFV2ATFcT+KUL391/ZLXK3kKpByVYLZq1wGqVDs4491YqxcZPi29yL1EyiJWJvZHMWeFanRxjz
/Ga9lB8fGWyngTsDv6KZN8xiQloOcrMcWeESteWIxIQlXGSyP+uw4pj1roRu6Vs2fFIuC9s1gx2Q
+RA/ud/VR2Q1jktPQ08dPlrptLMnFEk38QdTB5rRPBm2XMFy2P34WP3MyfiCYIjUFWCGf8KuNk03
Ar4K77MG3XLnvBup7fPFYDiBDKiYy2skhE45mD5F8c9OLza4cZ9xiMO9leWgYzn5DDvlU6/TzDFm
UrrqdH2WirsC4A+0uNWxkc6Jq8vwxW2EFjMa1V4QDc48uVCm46nN/1tLYdB5dUiHOvuiNLHdAlsX
iO4Tj1brUHU5X96U1CFp8KxBXgrcLCkNIKaQ9SbIrEI+mgZSxxfnxZUSspE07D4aNU7KvFLHAjNW
QdO+M2TqU8UpSCsYZezd5uz41DqUQYR9YBvdE6rKdIGKrOijNnRrVxoIWJPDG48IlKaYDub44XvH
7sBXq7n8o8AbwWZeFVydIKQoiYyRDzj3zAUTWtFN1ZmDTFLIdUiivGuoZdf/mMaEsZApnMDIOVB0
W1U3/eD4+G2tZ20MbDJqTSkJnjYP1r3H8SWgAIrqgTkBtC578mlJQHfdMMJCDgX5ciRkwhO1Ruoo
WTZJTG367LTSFSE1BKaA+bTmT/SsE+YDrh0350CympDM5w7N8TktJUgQiDpTl4iLOMZWLsSv4Cew
hZpXtuFotvtv2vUAeTs/64RoU+ZYORyWUI1r0Llns+x62m+6U0gKWnzM2dwKTAHaxXp7U+zMD7nT
fVWVnxrMwR9/A4BydzmSTm4aJvOt8jR1s/+H/EDyOCmQqNRN3N9TWv8gHyGody//qZGIIIBwpg1X
HjM50LNVX83j74csHmWdPclu7JKl9sdOq+iWuLFHIbjaYGY4kcCv2ktVjsJEXB/aQYIHlfEjU2kX
QxWmcbr0kEeGvwhMrZVecv5fO7dI+Qg/BnfIGcaVQ8Zv+Rv6nrC+Pjle+sZGrzrJV7rEeOHvPAI9
9Beu+VzHcJjkQRKS8ucrqvXR+J2XAhs6OVRs5Yjx2eUgzbakAgntb0H7khkEYfehYTD/4oFHBKs5
j1nlAmcb/9Y/0/+wwNlEBWw72oAokFqKAIIA+trXl78tq04S+ObTHDHwkIHmCc6izVhl+6AEvqGt
3lJVXXLruDKQ0dxAhYO9FI1pnv5md9jPyjJsvSoTKExyu8jpyL7NwquZV0nsk62DD89Fwj9R8TbG
an15oOslHYtpLMo9XusZMBGFBJxQJ7k4dEC3X0HJtwnSIeJoTSZtdPEg0kDeTs32bt3riwNiiZ/A
/wB4UWeRzL+dNIFqPZzeaWIvS/aSiHAdO7pE7P4fKa5J3ECKXGtsLY5pYHOrbpVK66Ku4AHoetJB
mjGvxon58ZSGnGv4WASYgFwbQ5byFMA0gXhsiXB92AmCh3eO9vzN9l3cnnIzfT64+slmqmOgi1Nj
J1fZo2dwikDJ9Ck+KEX5zVs8shUSdFag9K1DTLHL+nDaZ8sanYXWVjf/oGmWLC359qaw1SvSuII9
V2BeYgHCISfwtIfhp4yjwkZinHZu2YmeK3KuFKhgKN1YFa2vhYdUhcB3KJw6cs9BxsOugj8f/jed
U605OspD7C7SpJJdqqNrq/0uSsMvhWt9fVln3fZMjas0hKYJgzd+lY5pIifo1in5N6MBRbG8L0Pb
/7WFGug0YkyyS/lC5FApbujFf0eeqLdL6Lq3bsTpSckmKCJO/Z1Fd5/y8qtMnFpgRHrzERBSpwYL
n6zWJkdonc4RRQ5gfejjotHx3KORgmZzc6FdnDKG1l48e2I8ZtlePYYu0d5ghYBy4x/A2FaGKN+n
+RdLbidj1eDAPa3OpLgQQrQ9YFLwFjPaM2bm0tIMaK00mMnFM++AsdFnqmWUdwrw/Xs0oAm+OnTf
TkGa8idPm1fdCHAtzzXYM5Mp0xisRqQkofRe7I1ZWnEgTbM3r29LYPiGLsU3biIkgqDEcqZSwsJT
UgAMbhBwqrjwzqN8zUCTrDq4/3UhIFHumOrnCQCV+gIiaXQQZklrw5xTqkUTfPxttO96PPjqXjTb
tnlJYxGI+aComHbqLrf4XVZkfWrDjOVQgYS5lZdzHCiaAutQLYpTL/x7IxbXiHFuueN7sAlpn8j0
Ow40511c6REW8U5lUehPmPLdqYGZoYyJtmNQgOgNldFZSIt5yIWIMrhEieDlqVP7YPLOWK8+HAi2
+ImjEaGrz3dI9NSfzSjjh4sMD4CD0tYmP3OXA1WeGhjx4TVVsIrs3bO/UABbWyP8/43NMXgtAt+m
DjPcVjMJNTj73nLureY7hno7WsRa574+Hjs6j7nAlaDloehqSWDyak1upPQEQYKkhnpjbXxcw8HC
RKQ47VT7EcClh70Q7h/IwcV06uKeGK8KdGFn1n+nQU+cFDHjF3CzvwM9Gm+qc8Bsi96T35coq8ju
wss81CLcBYsXUy3/vOzImKrLWI/bCME/HY4y2ZLYO9YQ41aBMpCiV7YYyAn7ds54si5rI8qA/Frb
nzFUi7o5k4Tm3Opkti7ykwmUBtcW8cuuEBajDbvicuncbRiBUtKhetKUvKLg9xOvwlpllExqCTj9
1CzknbiAZk/7IyqphhmLEatR88/RZaqC5PbAqr0KG5BBDOAl/fuX/YU2DblhdBBjCEEwwb39vwkb
4RJSyKZV2xECcwcKN+tiFpiAY8Gjwzkxm65Qsbd0qRvHPbQ93eToUXPDmY49BmgmFV2UJIv/RMk3
Ypw3TrIRPhMhVUVFy29uc8Q6UxycxJmUUtORvUJmwg+bot6P9Ij45ud4KZZDi0dhvKTFRtO5lvoi
xEd6nrKyDAaqvaS8ro+1M+kDD1ytJyJhVr7/geAADtYks13qERBwq/aZF2/3RMmjiDv2rsJTfLsG
rcz0nxunPjrhB1BfE2yOfyBvdn+11R98Gf8QFZ6MAe1E6M1OQVewTMZqlJN3XxIOpOuccabziN8M
9SKquO9zODcL6qssiHIkP1jm/+ZYqGgIWDB4yze4rL/QdbQmPhvy4rLxK2gsDbfSBPJ6dXuyMziT
bg4HUodUqNcwiYduH7itahfIheh1qTVZsuDXjGYwYPmIb3qRhGvBO2/aD84+JtNkDwCM6/gB5Yrj
FERujsyOhK/Rks8GP+eH+xhGU6vIlOHKBibNlC6gvMGLtdrB4WiNmZLCcC6zSBQ0ShLBZXu9jYnT
dKIYfbG0DEEawNWk5rQrzC+mp2RM5hTu/G0g54DuvN5dldQ/9d6ahDhzNeVvzQMG9doy6YYDcH/s
jGTPrYml9bpiYToFH0Uw+G+uMHsEZh42WOFjUAXX81FyCyzQYmMjqJNRnVgXrOm+0zcS31hIv1tZ
CgGBl71oNnIJEkyyQKJGwpLkX4DhrZ6PFD4X4uTEiurNW5KIU+b6dy1uFu20oTSx43EEW6jG6UYZ
89bn1YPZPjRMLT44w9uSb+XBWB49WBs2Qj621cdZ5q+zMjUa5VyWvmVjsRwhX6i9ULwoFyvoP8+S
1eYOajF5FJSCs97IfM7MGtaBcCsLyVgojAMhj+zFXaX+BnBj0w41ISN+xGAzC2B+OY7N6QOrbRJR
1GJO8e00PPJTI+zfXlDdOQwYJSUqVQfoj6jOcS1/IHUniko5rfjhKUY7wpRq0xPyvUtj1iQJumMo
dZh4WllWp6TvwnqdB4R3wpNEIRyveFjix19NX/sFntnvtQ+nTyADXMS0EQ93M6EzTWEflTvQJIoY
nCE64qkAmtSY9eX3uth3CONS34Rcn6X7///JrOrXpUpn0W1DBiZY2xCmfEiHXJq7PjKbvwyy45ju
IyM4zxOyeuJ5eTtwSnVE/urznQA3L9j9TSU41rvIqbNEBBH0vuaIoj8m48kB5g4G64KEQFpICrRT
bf0kdKpNXgiOn1ztc1l5y2m2GuDDxDxnOYks1mGQL26FT0IYm6E1FZf9nRbsgtrGrbzeOs4LJ4u9
zQP7uTaNUAvfrIYQXWWaqSodUGqMePGXvckeseezZ5vRuDvzAX6KAZhu7GEoZh4Ahu+XUFeydiiA
YRRlJ89xPpjsL3wYaxsVdVkbr9oHF9r4HvyMSEF9aQuVHL0Nobf8wC8k+a9FpBjZ2s4mXarKoRrk
ySr/zaa7og2mlOjHlA50RSLG73vGNETE+Tc6fOxwdHUrhVcGzG3Z3bN264q6ngb0iP4aBFxL2ozT
14Bj8Sc+Fd2LdMCYXsEcp4HkStyxvJtXCzhJp9m+OHEOftVPs4+rTmrakouoEIy3/z6QlFN6a6E2
B0H3wFZNeoTA5BusEMySAOb2Uak42t9/vAbntK6suw9cVpyM2DXtpYwYIQLVd5gN6wDLsG9aO9i0
MqTLDj5J+TxBbeNjurlyYGHtIQEPuq/Evjf89MZ50YPpWk3Gq6e3mwGgrbnx1lG55a8sg99F6kK9
SCKwEuzkmCeiYZUR77KrASIEuhzmsggID1poDuLgn2G5cCFWOFBQKb/1P5aaRB5XRutRPtaxbBTJ
v08nL2KqLIlhlEfLZJDqug0Py0xWZZo6uuO+hnQzGW3BDs/rqbYdEv2OL2TIfVEfvFDaLR+o2Pws
EgbOR8lDseHVdQYfHEhYhiBIXCmOY1FmdPrjKQSN4Osja6gTMV8cAiHhVkEfsDfqPqdCYi6t+taE
WC2yaeoqa47kqctwC7FblVxNneRCa238oVJGItVSNgTCb3n1Rf8dqJD2XMU/33+8C0ohIxJM1l2o
IzERDniqt8Py06OpSY6g2RFKDZrh2COf00mVyWn28zxtGF7EODK5yfYocEy2IheEcFys87sx9pBK
OIGM4aGQ83O9kU6+Vqv7ZBVZuiROLdo0cW8SYSBDzZf/FWN0mPJ3A8z9RYqa7hJeLr+wSZLZgWEA
c3ditBpbau0q0M94rCCb8e4MsfeKT8cSQZcCKvW5lxeR5ApL0SQe/HdcIPNCMGbgfRSTDnTWWIiw
8RRTSiSUUQdgzjGlBpqf/Kb5Oar6JvrcILsInO9Iq9xP3vkHWAzbta/rUV43pJoO6RyZPoIkPkRm
ewJA/Sif48BNtSKfBodRGSBjFoAlnQlDknazVJ68RkpFg4BismRTCSJWrzpTzQ0iTGX71ugarodZ
9L6EFk/YsqsiRpmY1saW+slDK4nxBsw2Vg1jCZ/Vqoji7OQ06jSYub3hzCJviLy4zrHRkZmPFuqd
xvDrGYTQg8HNMBnpoAa78DToT3NBqJXV9ntsJJXdAN5OQ/foiLAplJroYAAKscN2O/ySBNFzkoO/
WU7I+e0AeF4WYqAl6FYsl+z9d9YJEZW0/JacJFa5gStd2AN0vgCngZegYBA1Cf9e1RzrLynDv+g+
r4Ce+/AgM+GgVXSF14VRXptQ7hX9xOhO0wBexqzU1CNHkOrSHC72/jn7Q7fz9gmlaPws1lS7BSj9
aTf6rDU2RNVBSt6yzxY1h/Alh9O//Xu4w+2w+rLv9B9ampI0chZSHNYgNME2blDWH7TuObnQNnby
hzqScjZrKKgcvY4Rt+eEqNRFtqo79/Spx1FXCxg9cuocWwvs2BRyn4tL5zOw81B36CiMtKSo4jSX
psBN/HPHq2fuA9DY8ZhIiT7NRXfVDYx69qfRvOE+lbG71YO5JEZG0ThUqWAww4yjWrRLQCNGEn8I
5XGky8KFi0b96Q75y80KYxo+uTww4lVp+JLfZKcln2M2v8l/hfZAhH4U3XjGkBVfCZyLshy5d44E
zvnim4W+B2sSFPWnTiuk7qkDy7713YWbgL9pIKdRaZYL0zpf/GOGAqPSEM5AX/MPem54PHL8aKGc
6rgdQUW8SVICZIAR1uhivmoB3y2M+J19jGgSI1lMsHAAIFWQMGsMTBYtl5oiZszPph6AAWqF5B5n
4nvuujwgC+G2yQ6bcO7v2PwdFYH1u8fVqQUIhoRAmetp1KROrrS2O87++L4rfuwX0/8IOC+HdzHR
y6udi4J1iuxfxCRF/Zw4kESRL2lNHN5K12wPVaHJJwMp+9Vtpjz/yP/SfvmgfvJd041FtwQwmYaL
Vi1Ol4+8GqIRQb8SeiK8tyEqNKrNoFdZo7xRjwb0gJlDfaYAzBtRFUdgDriPgfTOBHHKhNfUp1PS
lNICzZvCRa/r2J8ckSg4a0aLbK1fZ1IHn5dVl3IoUG91vQGA4MEDxz8vGq6Y9CYWOUId3zfMg4tK
QsIqxF4E5TrhXNaWzgl78++yk9Tj1jDavSGMVa5uaZMOs7LrsILNNqF1LsiHMIeLXgN3w6QprGfa
4xLbAeKLGW0AbVYzSPsRngtAD34/n2i1tpLUSioJqnLp0I4emsHAMPoNkY0sAnPsnlSGGHmtgB67
g/Q/yz24o1t0Nc+mtdD6b6jKRfkEA9pA0xSokd67Jao6FORxP+Zka/aoAKs98OBuX1YOSgGKYHjf
Wn4nUEwq31CPXhdwuKYNUDDQF1xuW2D8Vhmg9O/x+yHn6LRb1i8YaooVu0dKJetfdsLbW4Etq85v
pYNSBtMWge5F0G35z6wLtozmY4rGOTtQSwZ53dmHSZ+N5hGVOEymM9ZFxTysJ6WwmsXZzRx65kEK
PzZPZQNwYUbVvwuw/AAuc2YOCcxLyPn4pH140Mjd9uIy6JBB2KnUWK5tLKVSYTw5XF8GqIpaycIc
kTdgkRijmEhyUAK89l8o0EHNe9jX+OXeJ3dAkPbjfAOtIlMfEWbti30OU2sSN+vl+R4RIDaRwqRG
g/giB/JDOpEuoo3MjuP12pAVd9Ki30NZbpmGb12xMlxkw5L9AKmT85cJaAI1Uze3RgQjR9iM8y1s
+MGeaFFAFV07piRAOK0jiIxE6YWzpMV77UYenIUQcpsTRTPHkhUKswPQbP77zKNUpnmw7NJ+pbby
BfzZH4ZNQrUaCYa4JoUvaQKj2f0LDISt99+WdKc4ztU8+EAZvCZqQ3IwQwWEcD+BLMMj2/qUopID
hr64tkzZohVIAEwEBI1catQgA/1Mz1BHxCX9+CXgg+T3fp7VWlkxsOu4zFuHfHRTUJRLvcjWZ1QK
FzpPhnSPv364+3xhUkbPW5G7poUC2YzWIrQ2uFbY2SX1htUvOE6U6KoLzBs3fJj4cUqjJ5ASHnIg
//oHDKQ0VWTig4oHjiuZ14gMdRjxlgIwOa0PJX5Po5BMfn2V4wQDNhdOMtCLoWFx6D9z4ywDCYSg
31aehFIFE6srd8NPj/jhg7mzMIncbYMdVhX/FmEv/rJGp4LswIDfS9Yyx0AQNPi4X5nFbliZnZaO
xvhlrthaawxxZJOo+0XuH0rue28ovDmoISeXoKbBO2e1LHuaOwS8fB9qL7ddGNQ09lu6wW9rcjtw
l6Zeg9gM/V3AgVwdNgWtxmIKdmEQcH0D+FPKU0scl8jOoB1y/IrYRj8+rKJZVLdbnnpYpOWsU9H0
RcGvOfAtRUq6SmYT75oGAZLgU2e/R8EKtk55t8eXlB+JaeFEOKiXzGIP/sCKCb1b6zA/gKvPkiyi
cNp8v5VpLB+QXLuSiYy7gys+5USBFCv0TfFd2ZFrdt8HYcU32e/FDzWhfRr49rypn4PAHyu07XXf
AGGklnUVx9jZh3x4v8hm1br7L65oiWLM36OLVPM7Nq4f7TTvT4jqVefEgIazex0dPueYQhcWqEqX
7ZOnEZoAa+hK+cMMC/SaRMgespP6gGlSW+tlfc3RU+K8JE3LNoh54VuAxHMNfd6M9fUsYEXlXC8v
sF1OO1dBv/Mc1dm0+kKO1qP7R4Nxrm+N1XyGipafP0SbhVrb2pzrduuXc5w00ga7XsJ8D1xTXrKD
tVi1ndi0DyxAUbu1qkpFRRAnzU+6Gyph82kpHrxTdmPRFQ/Sh7YOg1/K4PcgtlL0hSL7W5wSQRA9
+Kb1ozg8JCHyRSOl6aJboYoSx+Xurq+jUGAk5g25kyYDGldalE0XVHYPtbtd7iPXBUbV8J3T/fOr
oavHAscmWtuaH4Ng/PYkrUZggYHqQwR8mUe1mGUi1JX0G/elMNzw3+lxisC5BDRvnekpS8LbJE1a
XDrT4cnm7jRXiLcV6yLy8iARrD+XZrrMbNulB5g2fczQTy2yXC90MrnJIisuVJQA8WbB+ctM0IwP
VJaL3+LniXKVoTQE8VIq3cAvIlXrgN+hkgAsalLNe+pW26T9mMxGu0uVgzgjlytuxe6iwMi2aTDY
wirm5q5nkx3zMnZj/8+FwS9eEkIioQvCvgsMcQkKxkNDeo6qrZUHavdoq6H2hOs/7Cwj74kl2/cb
Tw++LFivys1GXEENMR9Fon3oDx1DgwnZiwUXHne+ZnN5rR2P1HSSFjTD8DZIydihsOLaoW2paTsf
6c8MG+Jz/66lYWJzRUSPYi+1OAFZA++k6KiqLN0itIHYMLalVDtRtG3uw7Npsx2RRN4rUC5fU7es
N4R170Q26Rru94xiApNY68PChaHCEVT8qrfU57HUKlpEdhb8IuLMqj1rxKreXZuogrtpt5u0Drtt
4E/1ffFJ67em8WiFekaJ4iPyZ8mqV8nrTksIoiE8FHjCyGYmwuxvwfUqe8WxQ2l6UKqoNAnoqV4H
uDnjfPLtvBojBhfXR+IH6GSeMWcRBej1Pl2j0D6sO6yxyG+Av577GaiqbyJPhQMkvfSpuyUTYx3E
+N5oGpSPZJrr6FthvGCaYkeClPqgJP5j6Qr8UL2b3AhPFZJ+i5PxifxUvGsokSFsk7kVuyUL5w09
ofDEA+pC5tb2/dAmV5BVSfKXYrdliUiAWdetbM2P6P0XHdbELeUp4ar+jkIhNsNjuA1Cx7wHCMyj
bIxkwQeHR5RZ99YxZh8mni+ZyLTooz2bPqN/v9uYJ693iowPQrtwEx6bkX6rz17QXl3/deLaF2Y/
r38sU0QsTSehUuLf3Jbh3nWWv/ybtCf90WrWwO+XNVvKNrRGh5OYgsuBAUXNzYWaU8qU2XxzpoZA
k4lJMkipn8LJyoix4u/yI0aYdjc1CIlncZ6onvTc5NZMHUF3jS3p0r7J+klE4IjjPc0FpEjElMX+
0qV07p9VZsxLmJtg/oWcMm5wPOIdbPzkIw5bMDjuS4eqgysgq8A1zp/0QGotSCKwIwwdenjuJLeV
5WfZGAalgvl5E+Js93ZsCm8pruJKEG/zvZEbPnU4fPB0eLvyutXkteSb/8a4UWScNOyRvlSzTzXv
oAfNJ1oYsDjcz9whrcOlKp4UezTxofL/7is9Qkgtf+S+AmqhP2Be1OYlEygtOO/ELBid4OVXwTGx
c5foyqijzdH+2ieAXRvQvT9jb71Xdn1leQ+eqpREIjFS+0PSKjJJ3YwmQ6x+SW01MbeT7ESmmA/5
EcwyigwAfYKWBUQ/3Tg7iWxtkypHZOUyt5AOdfZM8/hRWgoMyrhX5YPeRZwjVDfGJ/GLuDZuDWFz
gWm2Hpg6TLuRF07RnXbmhAwKXYBow+a2tCTyRgE5ztJKtvfd4LFgqQout0EOyHVnEkIBeQksFChH
7zbvmZh9N1Dg9l8Voc12Z2UzPeF67nc16pzkUjweX6Ql+s6YspK0NbpqiuGBLzOKTfr/XlCoQCp+
1rdpt3t6D/+LJJBy1KBWUAPWICIsIUMgmTfyr82KmXdHS6I2Zc92B2hKModzpZwRR7g+nFf7+ejV
Eu+zZKq7v4UwQmRii/MKh/zgxa/X6Ehoq8EehAOTWXG3gIE1RB7QXOjxzidwWpzwk6KduQk5Cd7c
6aSR4aVE0r4Iz7vyJRuG6RIUj9SHlZMnVY86U7/6IE+NqJz9L5Jjhu/pk82ZLJnt8D7fC6IRzyuD
XIrsHKNRHs+mqGLybDQsHdBVaWEvhEcZuvzC/KZ6KTF//1oSuO08PJpX6x5/dp2T4PA1Qe2g62sI
ZxkLlw6Z3cmMSO6P1tU/xx8aLF4PChraJkj7wnAY5zhEPhQ8elddE2JEWMZjANRA5Q3FaPheGYDr
mdE6VH/O1cbQjcgkHc0eaQ4u/8gu5WFdcPjYUFWTuavlFObDc/OKuKpGjKTMnQUlXGKc0wE1jsAU
wbkmm1xdddcMrZBSew4CUK3smhxv/wBKUtemvOl5++D2Dba+Kq0pWBX8CSgZA03w5sQeCWo/wFV5
d+TpQQeg0O4m9+Ng8mYMcHBe8VX1pkKTfRZuGX2mFif9Q41geySUDbEJgk9O0Tu5jYjKhsHa/tZP
v7JZd64+BPyAx4TQWeox2yG8HGI+nMvqJ3a6M81EpTnhLRxYubuJwELxlUgr1+hQStrv7zZpgheB
7q2jP7SfIY+szUasWVsM40IVbGKa+mji4KvDqqK2xBNJrKgSTbn8eovxy9bgugiWJeWEm71V3BKL
2P0ZypP28xgJWO80/xo9GJY6JIjXkR5xDTTFYAaHVyWpWm3PVdGzf11oVI6HYefFWjau8vy27CFG
6/e9TmoyjWN5kle8WaOWk2EhnqY/1uOG45mIDBQe7Fbn+ojnOqCZn5EPuGbD0wa4V4a1D/VktPjX
lDF9I4zIRfl1iI7L2+5dBvLc28tjUzs7IfohoEPYeKEmmKiGKNHe9fc4qSK9M99KOIW6BU1/ejdE
rdsqTkbj0RKV6l4o5IyUpgl/3MggzB7ehAQJ5N9TKrAmWMQq5L/DHiclwn4KuS9NqRq13pvPq/ii
68jXCc3UARx3mT9HjEHAvfET/K3V7J9iZQOeD7K5D9U2D7KpR4UrW5E3WaXtwEige5OaIwknaYUo
zyPADxcFc9SNpdSR1r1tw+q2QElYgKoOnDIGTV5ElACpemCJ2+DkAowXtkUIChgBWgVhij/CLoOO
c7rVy2+OwSqdZNLlWIgihccnJLJlKbm3Nzdh4KVqupTcQAu9URhYdSGR5SqQ49ZJEInkFaEnKcMi
L3zCIQpDFsgmdGGtbMwmpMwH53E2hnWP5yT6DrEabouEJF4cNoy+yBHREsHNXLsTaipk/0ZrR3pl
b2tqG2vGWUrPKBfBnDWIzkGKYzeUjEpTTOpmW85H8qfPhfZ7D+oqxw8BotGe6D9riJsbT34LT6ca
FKVR6KFtcLvs+fj78H9oEjNqZISS6LBIddUYHy+s10jAevAYFgEuONR3fHdZt+Sre9QJI6yl+sPY
OD5ULD+tusAfIRoyBLxSWmESVI7g1apYjYNJDqKKqSdMRHu5sPRzJYNt61WmYr2eHYpqpjy9uXhn
uc20thFEnLJfOotOWpkkLsMt3sxMSz4tW7lmeK8fdJb/2i4Vm4rctMtX4AEZO/z7BVmk9q81B0f6
y7C3Ofhkj19ovbUgHTZIoS8uVkQaA5OI3gKvVsO6aIPL74518zvK9QVt0msAPh5IApaqQvYVRaSw
o9pRzBdQBkAM4MuxcJ6ZZJSsNs60EkVQAK5pLPoHprpCT3g7EcYIOnMRfapP+bS7ldXMsuBAhqjb
Un5qWKCaT1C+6L7C9D2/ZavUW76IDF5Pi7PXw8U9Y4I/PK+Q58dWMKzWKgMIG98GCn5R0pRigUSe
0gmylOS9Qhf4KeLx/he1vkWSNrc9TREVcOmsMob4EWPGuiCllyF3nZphW1Xcm/WNIoflHCQ9Wfwz
ImmrmHcMFOOJhQU05E4eFLiU5uCwe0M/E4x7S4yb7RzgSFBrSxsLpzRKTb5CErYFm+eEtcUWog4e
SP8yv6D4cRXHsoEIG5MNBZELqQV5/RBlTPDjCf7qDM+lzTnPe5lfBO7X8Sf3m6IxlnfPXrt1V0pD
u61vAj+SopvGHplYnJQNHWafyiI/FSoFrK+BM7QNFkPxqJ76CTBcv4V1pd1luuYf2Gm6CVbI0Dsk
4187/eIc3M2vHo+aUeDL+AHI2I6r3fJ2oAMThZWiCd6ULpdtFdPY2ISUPYyxKhcOz1ef67W4cIo9
2t4TtXSMo7a1P1qRZWlcYJaX7u2kSRB1g3lPDf/8li0dRWcwTtUqxmjZhE6jLr4p+7iO3ex4QZZZ
lO/OXm8LpGPebBw4D50s0UwTL5E2a2eDEoF7AytGX2kY9PROzcOm7FZSJ2xq1x1k6J/Vxkn9pihg
U+kvBkE33vOzDTmru5bdq/whCkA2PVy246s90uunf04GO9l0fvBcsQcxkhqB9xVptJfwaC13Tz7P
iIKRIiPWf6G5YDh/8NWKOUbsly+dwzu6IFD9D9nS4O8vGMrVKhr/a7+L+VZ+WWWYINvoy7+AC+SH
x2mFlRAATkjkOO+C9gPrv5ycf73l5K9ut2jpsqv5lnktQM/7Nd6F4RAyz/iq8I3zneLy6B3PfpVv
ve8ELQG2cDz2pcS7K7hLEd6R14o5TxQFraMRezTwWgA0pSWdPAA/FAd2I4Ushb9p23+MD/+tBUBU
Y6KM08qIrZmvGFpBx9trojUwEyufk34wbc8W2ob1UuvyrH9wUtNgA/26oXuXupYZ64wAL8XzTJvf
q6H2zpbjE+oq8okx++DQVkaxEE5cXWIU54IlGsDBeDFgJiiHjJjJQfRKG1BeNhY7cTC3tK6gazYG
LPpXEGmlJkFdj0DIJ2fy635kmrcZeGyR9p/T480GDbjJ+rv6u+II4ZHecp2a9CsKjRoi3+nYse5+
Wxcm/2HeBz2TSOUJoQtxq3XV3qqBjQ0eiKH2Oe0n8QhhHYATEMJU+ijwr0vu1jTrFvcsHVt/C4oa
tQrb/RFnMrYBNDHK/5bX1n2Rehtb6+u+hP3rJkxbPoh5/qX7Ee9NyKDEeKmFCJ1CtyVKO7A0UGh3
BSr4Ho8g48Uu++o7TaTSwSi6HSxivnbtXKPSe1B35tI2NAyIrdb8xE4vQtABU964dVz2xgyi9x7r
xsYPAqbFx4K+/UI3H9Zp4DdonATmKI+Jk0IJW7bQffbf+f1rUkm2ewUkmJkmKWLBkMJxRCWk0S/N
jO3TypIBzp7617XH2O4NDMfPy28kgL/UxCUFWqQol7G1eQf9v0AsCapBsa0duXOUas1ywOenhIQs
Y6ulF8BMM3sD1HDahyBSANxm4RyqNz5O9tLEizK26wZmDvoIcXRZ5bRyQpUcJyiCOZV3UPBT+7U5
TFdBK5xYGYz6BfBRKORFZgo/XdVQB9DycXhGtqt2SdivvUvzhkC7N8YLWaYczJASeIYHcTjLoXaI
BFcucuvJHHCR9twk7ljEJWpPK+cisioZGzXqgQp3LhhonteRV+pb0lmqawK2CGR57aA1SUMm9ZY1
aMdte7yv4LOHsehR6n1Cv4HP3oDq3F1gHp/09H+bfYqClUa9NNwhuRDz6MlVZ9H5CmnPyxP4LhmY
RPSNlYysftWV5abCBS/9ldxNDYvPNBSnyneFdudiLKbPxwVqOg+IHeziDP0Kr/Bf9ob18XwvueDZ
Kr/ODlKc1x4fbo7AneQ/aVKg3KFOeXvQq+TJJ1srATgNh9zIIWHPZwtEa5s5oqbY61qCmyGMsYss
wTq00WmlO7IAQMUgkN8ThyCfFBgXxD+eoB++uutV9n1bp+dsS1LbEXVSUpwpw7jE4emjJUXX9WLa
OLOedtgp6FdcciP24kiELTHVacEzorEWS3ijD2P4zkDDt16coubr34ibp9PzJKen7Lr94SPVIW//
KWk5hzpp93rvW61fX7VXLaNnYGUC0GzZqVynsc1rRgn8kaqq4yiVzDXDBXcDlTxKBnZOz+N+MeL7
hdGL+/o74ljstVil8orkPC2OFOQPZj/ZNashIlqqqNPQQ1jjInkDkJ77xI/ITPeuonLSXqLrUIPq
qoDm4oEeyz3woFVlBdC1gWXyjxKSN3PXmKAKVlR7LgYmBttEaJlw1pcoZ823ran8edaPs3zZTwfA
xjXdlms7nb8S9p2PmDMH4qgou2LRGb+wq+tD7hPqpMDH+33hEVBlImEsGQGdeG6VAZp2Lfuas/pw
A1TFvXQHWblml64yaJkAuSlQSRIZLUt8LCL8Lzw87IKxk4JxM+cq1UUlEjVToJUvWQf6WB784tYs
KDamPG0/DQUXATCOMXKUKXU24RcArXY/DZRlvIM3X46/oER2EeifppdtBwAj/0Whv4nZL0boe2uh
D7/0SLgKOVGyAqof/dGlXhTCXgy10DVx+84lE9grD56eKwBP0TZggiMeR3GvhsupYaGa/P5NPeqC
Qd7/rXPA4zq7xYzDp5yVbVWedB/vPDCCbHmHLJDcejiz8giKiha9448dLb7tdfJPrxtU7PeQ4urY
Fom0+1tEXVcTwzRjU1HgCpy+z0pGeGgcQXw1v/lkTdCJUNbf4vV4zHGYXVSSbQR+YaaSGGQJi7HE
vC/y8e+ZneqzYw8EyKsQKlGmuSPDTTW/NUyYCgXemHXHbjRQiZBsxZbC31TLlMlKI8tlfx/4HbVo
9hvYu6tH2aa9gfY20haxf4w3LjmXLtsY2aDekK0q5CJ6G63ELm0CJaOKTMgd096lnmOzS9sABX6J
B2xPZrrSnOKHUtErnuELkhCgkayOyucE3kGnLOZ3h6OqS0OcbvJQzVA14RZTZufsYTzlkcVAGc9P
OWSS4XhFUKfUEoaPkrYRU15pLJsP4/FwiZOEV1ejCd5KvAl+HKHbgfr7UzqEMjb5TB3VFm93JRiJ
rvPSAtYVdPFRa4G4MgGz778AOPfzEoZTNGK3PrCoBItJ/xApE0WuB8993X/FbK7k4EJK0Gro5WKw
tCo0qDzZvU0SB3XsRClaOVr8yCNMlak0jVhSu91tmvUM+vwLohiWvYjwJlGFav+36dR1ZweC/Ukl
4xMHzkkKY40XxCvtSIXu1PosfEyR1Kf/Wrm88F24zHIOSLC2utexOqnlbve0sCYKMfQu/eSS4iwD
eo5jVtz0WNniLcY4r73N7NPBh4LsyRmot6PGs9Sig7gnx4Djb3lkA2BXFwda+wsCumass598IaIF
eNH/OkBWP6DTSMUczppbNCjjGU15Wx/NCniFLKs1BE9c0Ufc3SLCnPox+l6gLNFEMhOObjaTkAL0
nHPdcg7LUxIrMgu7atJo9XSEUCJ/Ktiw3mDNqJiHAkc4mwIr+uF3nx6KTOXSseoqW9yAQvbGB/k2
shHtALnc1zZvlmxoaX5Td9Eox+Ry17qVqGdsEAFo7yFk1z+rarTQoV1qaqUVfQW1VKo5tChVGkMs
/kQD1/Qe6CgtzMMv2G8Ttinjee1F1s2RDU3mXM9DWsdVZBLNBYl0l29NgT+LcVydddVbwEiGTR11
lNqvVnbX6CWCABQW816R8B2LQ0umnQn//2Epl4yQd49kjjGmiCRojcor3oBZxMaktEdUqVM1kax/
sQ4CXAUT0NgmpJ2tP29KZ8EH5+pyiYDOqdZ0cy+9pTy6g48bSlhsReEFbiS/1cU/hmLfedcpiWj2
N3AOEcysXjf/kV/tZwzgvb4RFOkkR09hx45gLhV4Bm+zXcjbt5SWsGkkoiQofQzCEwqP2MCbKO3a
hsv9Sd4JFBMWgiWmoVQReTYkk79Ulk/YJZ+CFnuZGElVCtVf0ml7qThyrg9I3fNt9XgRc25NpLud
Bb5ET0pQaJi8e7NmA0QA5A+Zir0YyyZbs8SDMcUxF1oPT8iHa7Chgvh9SDedPz1BmuSFq/3cQwUa
xLezgrt2Sr2UXB0YiLQZkp1eu2u0eoht+7cOJ5Wzw+Nb5wzA+OEcnW/qSeBZHXCxk3jz+O0pmWsY
01ewNhjmOS2a0nfxRBhApKRMC+n3mS4aA/REwq2YkrcqqQHHcHKI2uWtnHmc9VQzKEqpTelAdVAy
ow5LeOK1eS1qMTYVeI7lsGjEmy05/VeMo4odVkptRbH4oIsu2xapp5KbkowY9LgMrc6MOPkIvEtC
HZUrlmSAnSPQto97NyrZTgrLyP3x2oZ/zii20fXrXFkz7WJ+baYkLF+cehAKRavQXkDfKfQ3xo2H
qoCm02qOVs6RT/NP1Xul/lw90nEeJqrznuMv/HMCvHezIMV5G8n1JRPsX1WO2sTKB51l/19iqdBk
utpqk3SIkZ85vEd7XPkMgNknDr6s+clrzm9txDiIqXXWGD/WFMl01yZc1xeqhDWz8sfhyZCHPPkz
2BzQnshmGwxNdZF41fM01dQRoCIhk6XHadqbn6NLxOrTi7qC2jKEaJWYGuV9t1Ud4ycyWv7bNMH9
BF59r5X0HSfpK5qHgRWmiskIVWjUM9OAnEJffOwJGq0n3n348mfeeTkl1uCT/c80RrCDW7DkN44q
/dQRupmlDfoKxDG9q0sHx0ogGPJ6tbZ/sZfl7uh307BnHgegPB9re4/JZuaMUifrl77BSk7fHJ2k
dTck/ywlMa6CRxu82oXT/fiHlex1L1XdZjJLdC3T6Df96AjUCEeyBCFtPiVOP17QDl6X9//Cc838
xI4NzS9rHCaGJqHQwQ4bPpBblczkqvwz01LaRFjuKO2FbpnmqpNrUGAT/I7VA6xaW/v5AteA0Oax
tO98Gfo3iyRQpA4LQx6OUJz36sKJ0gneJSHUfoSDvUgcSlW2/yXvbfoQuVzkZjWvWFx3hodNEq7r
yKpIq5A0amTEzLLnYT6C/y7S/7IJ3Txodh8H2+sZ6KffAeslHv5U62/pQEHR34FDwqrbAlaCHydy
ll59OqBRuwyLXoWmR92gIJfupVDSjDfm1Qo08+nel4gVAOj+8mj2eh0BQJmn7xj+t+lG3C01X+dx
I665w8MVc3lD17bUq+wTtZcCBX5kt7GxLE+TrRIFeUzYG2y3j97Bv7z3nXHiVqBlcRCMDTB3DXKD
+nd6Msed7uVbTOgxu+64HS12j7alumM4ic7g//9Sr6Ur26XwXYTm32lWb6NKuM6PzFRFUvXWvx+2
XGYtQ0xMSJI0jY3Ct1P9Wyhlf33kRtJS/Q4bsMETO2nlkEdUfIlP4boAFIi0VG8Mj8099gxZ7PlF
7E1DQKj3cgmiTj6V/Yt8Dp9Wnq5cej0uo0yFYZ3AAa/ySVw9V39mE/V0ITil4Pwj9xYjJAHPT/CV
R9thzPNjb4mZ4h4fa8/foPnF1yUxgY4G/1jxVzBO+h9m+6YcxvZAK1zLKesgo3b5VEnGMgF7D7sH
65ePbe2hNyH7I7jIFacZUQHST77bJSRtg3/TU4BiWtVxn8nUp8AgslywnMLdDJcnilDwG+Paie1e
ZVIEZse+W5D1+Vqy58LVB0cjuqlfBVHhpoCiYB2KDALAt4m0kxi7W7lg8VBz+VsuEPFyYF2MTKvi
wuHPyiXt+JlNlFJ6vSiOo/Z912zTQDuiIjxlbIEHGX6qfw39V6l7ZJt8HjwFFI4FPQ46ATw0QKux
WKPNRSytg+FQMB2P7rH+sFg1XYNm2ARGnZxVVKcxZaCym+pV9/ka5BHuGyh5FC4pFM7z3iIor31H
4PUnxBfpWPzypZKbjrrP8ZVw7kUWZef9KiYMk4KQJc7CvTqcy/seSdEE1sLUtkzufuEFgP0A0LL2
x5jnXzb8jeNvl/Lg7wUj6Us5f3YeRqiDACu/ZI0ncRlB4OhNQoosn13wCdIyKc0kzJ47DDE/YP5A
sljpxnBTUuBiDNc4sWls5w4ETAB8Ml25acHFb+LwPzREp0pGDrE8wgAgYvtt1Bl9WlSVCBpw/UE8
U1HHe5E4rL0DwdZuOixFyjAspI0EYSgis0j3w/RmtzPNJn/XorcsSdnMmoTxqn8QJghKBiVZXocB
ZqDLMurX1hpNUya4OxhSQQYUTP/udcASzM1qUU25EGFWXBOk+jNHRbR4IXLaQvrtuvMMtPeLzGrQ
Jt4gSeSj313oEzIg1qXH95YsvN0aZtwrClGavHtU9iJt+9fQFhr+KfilRchVm4wAAEy2KQTu4GlW
7Ke07F9iX9fMkmEXfcFJnzEpizclFj6EM2wOUKoExUhgYURJBByoLRlyTFd86OzIINXMMqFfNsDs
9mU3aAlu0jOBv58EImNYlg2t3O/BXwz0aqAL/7NbdqY37L2oM43SxNK6FrPfpP/JsrHr9F03JiSa
BfLS5pSpEErFPbgt6LbVHWz48BWu+WHOtm5czXxImHiF6thmJ7C97q0ZARj84dG6Ng8CtHVvSbF1
54gj1wJcNk6d+KLzME41dck+xUOdlEJHOzcyKrAuMksw+EkE3u3fBbN5BiaXF66NhNscS99X5/97
/QhOgeTxqjlAna1N2K1QLN4dhuZ0/gC6QO2ENclvOMXC23CCOpiveOQ/ZcuLQ35ND/997H/OaiTC
LXU+BqrbkZ9GX+ktR5XHYeH5fXs9uasKjJNoAOIitRj6ydC7RXFkw/OR9GTuOzSmLc8YY2YTSKpZ
RzCUJAemXd0DCPh3FhsM3noRKcYzKcowaSH5wnj5tm3y5Tb/aU1qdFQPLH5RJXZeZggVkkbcRmpR
KUT2OFU2SBpTL5XBAtKMpFRh5aP+iLmoG+BGASd3jRC8esUoMmABOqHqa3np1jltKTLwJrdbzqy+
zlbuydz9O9D4WlF1WuJ0dG7QgySn9xqyOcV+yGpxyw/THQCTVw01B+k6nA9wifkCmoZXuWi773Fb
HnxSBlIOsfov1ioMz5mM0w+nocE3iAE4UYDLpeNmWJxRxMscRKdFTFs0ZCLnTZ5f04r3SaDM1RYa
+UkWe0eLifMxz+gBwl5b0C8vmXPDM70IockQAsiTCZTNDMD+yL/DlT+gQCDQ/4RUlqESVAbO6hGf
XE0V1JKf47CNOOaB2CcyuHWOHL9UjLGvP0jUs1BEcTFWyqVhxLMN2Y/rIL5eq2+yyL9s06+9ZHzj
plqSUt1tasdyd+Zk8wXMPtnlJBHUQmHirBGtH/o5ziVH/2sbJuJqKTJsRa2Kp+hX2XbV8/vJ/1Oo
JoKufpjruSfSLc9buBayCs2Y5zbghkjDlfWeUs/odTBneDvQlg99+QZZJ1tZW5hr1uMjznDHuYQP
Slte14tw9hW7pdNe4QMwMxCEkYj/6u38vzzyP5kV79mwd7NWeb4kyiDNRRnsbwGOiSnEfjC8PfE/
ISpw9okTZWDhJ3ozaviY3xicymn4kF44X575GuRC4NYIJ2c3Ngt7MOy1ZCbhCSKwfZrX8GL/RbLO
IqlRwBdseE9NdPBt41RzGMWYJB657A5ozonQd4Q8LeZWeZE2/Gv2AiOXaJEPS6+t+LUlpGh99tkw
p+g+SpxIteWCIHNgqADyHdFje/HQmae0g2M5GUNZWtq5kXwq8ES9DciV1mY1ukSma0cVMUiXo6QR
aKUfxHnEtcwrVkxQbDIRN7SEN4HwPQPkkqrzYeDKkZOXVCihyw95zq9Y5Idf8pGtAyUMRXRiJnpU
oNwxot+XCHwZHgDz/6b4HCcT/qdckpKb679hdTErNCJRib50mOzCeblyytx2pZMt8EeipCC4DwZz
E+zhV65RnzPpVefeRwy0soDkgZ5fNW6xTJqOg3BZMClEws7suHOtd2/UP55020vzjHZ7NgAq+Cml
wwA6AVG955L4rKWS1yZr8uyPyY/rn+ldlkSTi5yXn05H54NzjB/lwBk3Bi6RfU6nJHnHV7b78s6H
5s3s+j8ibj+YmkW/XWK+fVYvnfmYwC6GiSMUg9EsnzrZ7PplvmCFpmmyVvIFBWFBA961KpqE88IH
nP5V7OV9dLI7VCiZK/t1gCLfy0rCrsdMqlP0wQYWvP76GbantVJ8sNemPwA0aDv6+goW21MRlG8V
T1r/l32UtKmV68Y5tysofkRFfsp1mTduZmzPddWv2zSK15tvc1RpMa1PKrPeJtLo9jHTGcb6GlzL
CRilkH+X7MP+YYFwhYtEVZGl+wHTsPNn+0wJBOXh20ciY22FJY5CTcQL3xPFATbyiQOq/ma5wtLK
th6kD+5ebGckeZrW7rBEx66EpxnVehQqODxy7t+Ywe2EY+ua/u1u26fHFeAy2fJqigwkePi6IKJQ
i6PniN8tVzZ7vJWrfwTPeM9SHztqKqjgxQFoTNafIpKKinWZjxVcX+M/Qvn5gG8BMETmpAgYSI0K
j+C5Wq8Azz82SAiDZzN9BiF2W1CaxN4rfBRAIBFS+s4ZfAAl/uae4jPIjkjXV1c5btBfTQIBEF7g
+t4AfXQJ6pUzZEYBD+sgCH5aBEz69FvYGf3oRD1kF38PmgYJ0T14+L/nwzUBqsD/JXrrNb9tBkum
6sy4l7v6OOsmwelCb3hVlJm992EVnDgeiRclFzElCPAfu22uPr3nds9dv0muAwhRKGHCpIV9/tce
yLFBv8YjhF2w44DuGJ6Ndrib8pD3ZrTXUFUs40YZPrCZ+3uKowfHxOzeu9W4pHacWyYyTtlPJftM
ikECGarImTQAtuCgNjNsIP6AFxr+MhpQkEX+uefNzkNj2OQCr7ZmZY4hKX1xyC++RopVosEAZNHV
QU2Xxj9+k41P8o52C2sGc5RURZVYe7NX57VVeh7Mbu2P8awSzIYeJTcQ3NT39lEXnPtQHvE8bLZ/
WxYcV8yhLBAwZ7s01H+cEMtA3mjJBQBiXo+0tU6MQMPQaHPo302I1st0DdiJ/UXwdl5CxCTB5AM5
1LsVDqkOqvjkSJAakk8clcgQpWVB9xZzvCwjIxpaG8t0ICkp6lJBiUKS+m8V6QeOg3LrxEhTA0d6
WaPcjXuAYkTOpcB4b7fUqsnk1Bny3XsEDgMX0DbTL03Farq8Vo6xFpMhnTDfbbj7Bk/Of4ayybiK
NGCrD5yBe0vVXmtDxIxcXLUZht6JFBE49DFFG1whhCmN8rvN89ic0ZkksirjRld9evdU1QuuuszK
7bARJ68u9o6HkoNLD9tbYrBW3j9pdooDLQ7Sf2c7qNlU+6Hpou5RvHP+G43rzbGH1i/ApV6k0D25
tDmRgpjs80G9gEoWhvT8jWZPfi7oRx0MlIkkJfSkxTEAnmGb8Tjp1WnXZ3MhUAc4H38WwQcWk/H5
Jk71zagKuliloUxlUuZS6wi6fZW6YJRi3WoJUa3qNapgmjj76vzmfm8Ev6NH+WcIli6ozugUXSoI
tJ2QvOOfEqD6uv7HjYa9rab50sahHuhY6fFHcG5rk5OdeJRqrcGX469XwgaDJtlrwtdxCnNr+a3J
6MeiYRI0fbFLrWelJhsonvO21O46Vx4ZEY6AFPP6fFFm0QPvuRTFgH/q+QUGnANRFEV+WIxYvVxZ
tM6R2BphvQtIna/4IG2CX/ayqKx2OHs50YpU9IE/fTIJ7vxAnJHX5My7QJG3bM3WLfYatILaZpcH
4JXOArlYppFsd71NZJJDb01gP/oq6lnWu98WasxsxNfRvzmwk/JXqzVMkysSJTs1juSg03T6vsic
zJvmwGIL9xvDS8tb055JlzIuvOv2PA5aT5b1lVHbvBUxcm0lb+zbtVsl5ka4UPe3SUrNS1YHYhol
YHngNl0oPVQz9QQA1olXtztDXU5iBSsZINVV3cwXWMF6TbEScW0Rx49+OH7A15AAGnpu9sEHgN4L
L+f9ZT02MBzN1he0/6sr4PES3FEAwR/emtRdmkwBYX7vh+vuAqh48evComwD2h5+xn3DKns3Anas
0FaKamw++ZfZRLcKZsUfpPgTGz0kIdWpXAH76ck0JMFO4yRGSl1CAvYFndfaWplO9Widf6jjovzr
e8B3KedDJZ1W/jZPJNxYw+JFtOxSMWglRkKZ23IoPq1Pt9HZkvs5o/WRgJpqMbcEy4S9OjpE/Y3u
xiLIJ5t6QLneOP0t6H8Fku6uzF/vfhp0pSLMAlUeb+C+NEr/S5Jz+YbcV1i9/O5+kzxu7C3pPXAq
glykh9h2BU/wRV5SE3Yuifm0vwPVaBBsy4ptUOY384ZFUf/efASpC5F2YyaDyug9osVnFH0W9Y35
Ri/MPsAm8Wk+Mf3TTlEBAJtkM137CHVXH5ZdQ4w3N0j6+TyY9Q5CQ4Yu4DznBGAtabaNuIbdHn9v
LxqqT5ec4OQ6Kyh6QDwaGB4GBjHVIRYvN57jgBmxrYQzGhbK/Vg8JXNRClczLztTinPDLJ+h6W6d
w+CBbgtQfBL3cpIsCnNaSyM6FTPwt30cQY2wRp8GQaLF0rssfjzO2JR/ueCnc3+xO5HgEkyl/2q+
+uUzZMV55PN1iJrhpxE4ZUiocJuiW54Rvmq/QpB13pfIT6pGrGASDouorVSzcT8oGA82NLxu/nvA
8FvbGgWlQZjU4I40+HFVaqb4i175PLCq95kdusD63iIRJMcFruth7O+uAqTRf2lmic3cg5NPSMrx
yBXnCOB6fMTD3Qa622QORWO43W/uEJkK2rY5f1WI40CCJYpc75fsBNQlMXJrAWWrBO59dkXDcgS4
qmOzbhnnc8wH2SYF2xGGqK8MRt/xY+ixmym2lCnAtusaEzwbiSxkRSvf9wsOPd+EvHvx2r1z2bUm
zK1M36KSpOkWdMbEygrQviN/3hNkfxZmpS5ZG2KbRu92wwyBE7KZ4MzcFdB/Ai24GFjaRDyCR3+4
sLgESlV3Iu5v/uJiwf9BOGYM7YFEFQInJHzZRDNLsKpbZH1d4e51kZtEomt4CbStKBuzZ3tOOPlM
l4H5+8dYzq6udQeroYOpxBccJ7JsmDchNAnzomrC9tSX4Fa8LhZoThMzcfU1PyiKrbTGQQNt0P/v
y8hMVh8gJoud++AwCqreL9+wJlzTXmPoe3yieDh3RKnm1E1NNJ5umBhPC7exP8AFQYk/5rs2qp4Y
ZiOh5KYJXwhDrVrPnjvya3SbSh+7/Z8hLJNfwNxFNAx+J4S2sdUfwG9FQzU4kWaQF7TmyZKsHsvU
sHA47pqP7SOMwncbqoEKkaFS5CXwbw4I665E/meY6ediAsEdvgNoFCRPhTr/9+SZ/1dCQUr+8Z9G
L4gbONibRnDkg8V0KDOw6Leq0xDdIioPCe67WUUsnSeulSeoowlQZQ9fHASItT5pKUq40FE6BcJ+
4Wm8jrM5iXQC9IMfngM1xJErEyBdrHe6bCEBO4g7oba9mHNH4APvw8+CwhqKoC7MbBcqcCUkWF7J
qaVlpjmHWMarwKt5FiJDlo/R9gIyidMHhfN5mp2Ht6Ex++sIPnsy87dQtPJb5pTw16hs3yuqgLgV
2EKvMIrsZ/elQxicVhVK/Sgs8ryschSKJpGMpG0UuifMAA6xJCrjeM2FbNLA8gcNzVk+dEJt/mxk
qur3MENMug5gBrQeEEGpPzDQDT8PvfK1YpI+Hql8ErASgLOzx8OpIqo/648vCQszChGP96yL2rx+
pt8OF8uMVtoS0R0jT9mIb6svDKpe5Rj4Qwy/huqG+ARYWh/JhyFxNLqRqXgwTGMloaNQOAED+lcf
Bt646ic84MRye84AIengeE9m4KY5RMd5oyVSr2TYnMhY5NmYleGz7Nuth3X+Jhfcv3SGwZDop0r8
2urK8TifLpKhP0fuR55dl9xsqcEx2yRSvXhzbXjrccou4NHTyLnfzwVv4Bw4q+RpJbvcwBpxbUJV
h0Gj+VWKeskOQUVWbDRzNA1h4RTFl5nWmgoDC7+KAON1S6BmUVuPFbf9P4PtG93t9kwX3grW+xaC
DpBuRt4HtTSoeWi5HjQxsXl/P6uJ2V50oeAgp/SgfcjTufIFyY43y90spLvHVDeNGLzdaoAlGBGu
129GTmcHPps6PyclmeQ3Y5xYuYb2Epx1Dv06gyhGG6Sh0m3wbg3P0Dk5kgtlIt2ualI5i7UuP/rp
eP093cjymnnYgtdNsJ69PBtgMjvitZBagCOHSBtKbZOi7Jsraxy7GQ1/Np44OSMYfzJHlXakTNt5
Y1x+IBGbgQ+qyeM16B3j/mczs12vXoO+lf7F9L5XwK26Yg1sTr7o12VKwYfhKTYSXKU6AheceNW2
gGhdlrTbE5+5blXRVbZRj8UABaBjl7lrWZB+Ke5gNbYRGdVr2NJsQe2JjmRPzwvmFgV7YmoNfCPu
do52Tyfjfk8uXQ2FiearmhOxTIl61YU5Jcw6gwgMTHRjKTBjMQZtrhokxuTQ27nD2AScvgVRhpp/
mAXWcS02kfNFx8jDzafA8eNXnHNYt1+5KTFy9Jj9VHDb23zNLfmikT01F95+KQu4fmwGhHirDLFE
efEXvA0L49O5wCDe0qfi5zpL4NzuZqZ1Q5P7h+yh7U6AjwvwAZ+5KsJRafkg8/xagdQqBekdV5IK
QvG+Uo3+J5lf5lzZYEwtluyR6Mcpxqz4NJi8pEeJ88LCSvGBlY8w4ipzbmTTePfTTE7XdG1pZm3a
2Uz62yNb66/U2Gy7UaKakKAaTjkEiohQrFWR8bOjh+vg6vpoNvbPVx2I5aGdPe5uLcvxkyQ9Q5EM
Wypcn/p0fgp+nZ6A7kopHVnIHN05XLyFuHC+BgB77Cmo0/K1WLJ2gKxQFIpnEfzmrt9lm7Vjo0Mr
HcK3OW/7qpbxsJYGquS0SlryHdNSkgpnNTu05C0+sVkbjlSdO+qK1UmW4tn5Jkyob3iGyHw8wA5q
fPH2SeD6uf6q6iMEeYfdoM5mfCJI9p+Z7bI2AzyTn+x2ptaHf6oyIW7uBWqULvxF3g1NZxBibcQu
uV+FWu6s66fZaYlgPlood7mqRdl9QCsuTNGvd2iL/V8rTjQ/wFVxNljJGKnMQ5nllMvY1Z5TTAXD
rugOfA/PuH9Mekmxma80+ZcGwi/frV65uuw/5gSFzFvAj2wMcfJ8hpTs7eyV3REfDnaVEkHjl0YQ
Ei9dWDwc0WMui0S7FL9s7fMsc/+jiTHAKtcjNcDKdvhlTPsqyRP0d1x1VS3OYIVWJQyGpvgtWKB8
F20Jx+yLSTQSopydUnt8yXv1Zzxaw/qxW0DmXCse/f+epMTBI8U9kn9gidg8AgTLy/T6qx3OpbJv
m3s1c4k1NgbACAr87Dd0IdEVdEj5x7p5pNMqb/43YqErbfF67JzJe8nH0Cx0gI93wkmFIj2FRP3t
IxMQX/gPjlnb3andW6ursyCo2dqO+M6s+vTF7aAc27x9t0OrzZVLtov/bcHns/moBOlZL+eDV72w
qFwgiHBtZwJjw0m2YcKojCMOCFuXXYdDgZMphbQEgfYF3mX/uAh4R58rGLKG5uh6Dr7RnGz7b/EE
qs8XAUrc4d7yhnWSXMh0G3ypcFJ78+I9Dofr9G55Fd7B+OU9D77LXJUXbodVDcMM85FMD1BuhGMN
suWUfQRDemWGFMQTbLBmH46Eg3i/tM9mkBA7UWCGvXzdUsJrUlGhvJ7flehPAG5oxPMHMd6rNPSk
nYKwMPNhqhyYC6iEfLMbdySfGF8nNB4ty91oq3Ku2IsPABNFLZilLJdnDlE5BXkCzDAfm5LPwGaS
wywAWSwftuJ88IrrlaYNM+j/cJVolg5muniTBwUmTbvldUu7jTsOZwvi8Z/Z2ZMjwM1G9+tkccrW
QvydgtZVraJs2wumpEzOo3odvsJSnUET//uG5XW3rlcwezaz0nZLRjV/p66FWXIXGxAwAkoSEgUF
jglUrpnGbGRI+KBAtkG8Mm6N5LoAcCc8oifw2/2Mi3D2VyBq2P/TaKLNaseQtqo0W8Hzlp6nAUw8
W8su23cqb25hqHmp5AOgDTsRhv7P7C03kRFVAypkaSPt3qxZwdvh45Jmdw4fdyl7mwydqebXw9xy
YEnzuGN34ZDcxiQ6m9X6pCZMRCiFiWiGrw3873JDvmAwaBPpxH19BxAylnvn8LbC1shNiDOdPSJE
uHjr3DkbAUtoPjIlKJjD1rodO/9+sTvZzfVvzf91hv013P6zC7VKo0EujfQbI7zYkWX67JU7Eh8A
is5fwuQOlEFR1hRWoMvRj098074u2R1yti5pgIGObgSy7IX0UxBURNxXHu2Zp/equqZrigP5L83D
TNhY23/mxM4X6OTpFaG9bQNuMYS4eOiEjXtbmOPiyL3SY1AtBGKRt9dKokkcQ1zE7lnsqqOtIUbe
4C9Aa/NQC53sQL+wEbmhsg8nC6L8oAjK4sWaPr1YA3aFyQQ4u578tte/gvbzf0lwB9yUnMDziVdH
oLBEgARoVU0+7Q6hZpD/LSBesbgzIWDG9uz7OjHX6VUaQRkNretNYMVuVp3JzM6/jtKe+4iwHYFX
QklmkBj4LX9nY7py4kua4jGgk4oQjjgZMTFnrrBNzgWWEF7Dylyum14p+RxveiCppGM+kyZQnfvH
Vgdsr8/VjBC9xPd4zAiuS/JzVKcvky79L/jvZtccrSldYWDu0dcLEbEMlhVC5O/LHZjdPRoRNcOA
S7sSk/hbjA8NAsUuSWBsGM6IBYSzZAS6y2blERJbNaHDdsyeGjSdZiex3S0QoM5xKrga3alEf6OV
FnnZZeOq8LbZPQgfwOhjFdDmMrhcb4lr09QZPsuehIp/4OxqRNqG7Yz/bCP3Piw5cI+7kF7RAX3a
mKWKnUvb6Xj4nZslwRRmri2hljwaaxHsZ/5m1BKrqLrrPU42w62nWDjFx8KG8mW60LP5FBxisN5l
6ypFEk1cXS6eKelqJTyEe4YN2KjTudnbgRn3Nkftqf4rkGERbbQZRkvbDJGWjGOXZco9jnmK6zN4
jq7+HMFZxsgh6scw5KVeZ1ZEbS1psTGJb/nvH4UjxyE8k7VeBUxc26gcwyXDnOqjnZq8eXm3JE/Z
Av2z6hNV8Fu/oYmwfJfzHjVJugTevkiYzFwmqZGI7DhUsAyrzEAx+/eLsEBPxmZPaJb0f6Qv52wF
reJJyWVxmdx3ipvl0EP86PlipIRndQEjzMHom1xoTUWKwvF4aKnwpS+Zn5aIc+ANVORYBre09xPg
3O22+9KHoNCjiuFq7HExOtV/gpTdj+BqtF+K7dziQIjlRi+JsHoQZ8Gl/Kyv9EnQQZ7HHuwkTd1c
l2KSOZFYn/L9xbb3OuqWPfq1MPt3Y1FT0O0mX6vnrqD1lToasUIVF63V+N8UWKvIEkGTpoMyn08S
w7vbleS/VbqKmnWGXqPqxgEGFn7Ehj24AP24f3zbAePHIVnwp2jwBcsExu0z7S8ArSUk6kAudqNr
Id6U/k/ZZAfw06t4ys+sqwdofXHao7XuXFgV76UBbmDQ5P3adX2pa+ksfvThMrubViZUT4B1mODT
QgAByeleoFV3Lnwb4DvvOQS4qMpQ7NJlfMNXw4DcfOn9e4he5HyQKPKPb8pXJosgImow3dQGRv4I
4xwfpLmQF6Qdo6OZW95V9X0t338JMD4Tw1NF8F86H/b7F3REGZFimvV2QDMoKEF9XJ+w6MZEWG4f
MLjXq8WmIgiDKRbcdcniRuZ/IPQ5XGhm9lQmBYQyLPPcxk/hJHWdlyOAX+5sh1UGCZRgEykj5N0Z
PCCHlBZwc8HoIrrJpiVShoKfc0an0PfIRoXtBTQNUxGsbWIjEnU6nuCpL98AkxYjZhs62yr3tYo7
OEm3ICA9XzEqIbfDFdudfl24BHtWsAk5sFnoIG6aHPPLg0Uz5YCq4R4bVQ6LZLCXz2qhaiz/muFi
P6vI36csLE3XO6EBlKTuB4ZWmldlR8xpONqmfNCEdXoaOSDn9aCtfNXWdcdqSS2VpHj1UoSf8cqW
BQDtkratYDD0lI0ZfEn5Tvlqx3bPYrN9TRfNcGR5/uDVVJBQ1k2i0LAJ+lwGUoDsTOhS7GyaD1mS
cpBjKLsqopXya1+RKUQMyPmPjdqUWgm5QKuKN3E1J3uNqbPQaMYRHsQJcDwm/tJXCFH9Qlx9fhKG
PbYmudVapMZpYk50OxI1W9JmEoS+e3XHn28GqUxEIj2vidTtq6dvryQpZcvQraGUOZGJa/2uf5tl
Dk9GdJGQJPOa+EGZvE5rqC+5HbdhNOI96XWDGISWX6MoiWijrib157qssauPtl+ymgLfMLx63M3t
JdN0fhTuOlpgBt7vpN2cqupXcAIvniWkTuIwEyaOdm0bJQZepv2xsz6gaFQa6WWTFoei4QQnHSFw
ZQhGMiFJpGLzl6wd9VUzjM16YG+pSwerwqfwyFMEpsGOzSdInGis8SezmbIlhLYDDiY7ai8Q26Js
g1pCU9wdRqIRZksR648aOJ8EiN4lM9KxkFaDyeeRTuVvYGKtJ2Net9BtRTBFKepolIRtzX58drDl
ySPeDg7rcv0NeCyG9gMnDSDEPev1g8J+YO4oy5XuEhpoEUu9wpgKvKD8zknZt9LbqUoVxW3eifmF
a3AXkFTGwz1onUV6wk2Q00RrH5tr/qvqI+UAJHm3Dz8exa8N1KW6R4L7Pzup791mHR5pUlOlDqBg
PDlSGdxfhVmOUFFFLuKdEb2ULf8832sT7wIsM/cbgB09b1TpXHakhr6lvwbCl3RJ879vbCYpLSBt
2sHyfhzJo39MF3iQHdtTNPJg9gQWF0vZyHyA4AbvAaH4k8FG5EDBLyGPl4pL0zXYMUxjGlF/o4/+
shihgVJUgXr1iDGm4NuBiEnlsUaxIGFljbGHW5ndTMcEH8tOARPs5DWA7Yp+dBpzmQPeU8yirA/y
auWpcZuWSf9M5McyxWzbhqpVR7HvT16B+Psc9rp/4xPPBC3SpTacrWdwNzUeScbQVE8qLAMZPUrW
Pu1Z2ZMUA3AqEMpgUfVSoNMl2IUNgYDfP9FoVMFnomUyCABx4YLsmLAu7s/gVP9gc8idJS/YDwNY
c0Nlxx/QBlN/aO6NVcrshNqF2Pv7r6KcnvPoSV+Ww5JQtJbbhrHSpYlP6w8NHPAUt9dJ23tJ5WPV
3cntmQNw9i0cKcHwt0s9v9InCUkCQC6+TTg5QiH+oGCSZ63o/gIBU5BXIrPZk4OG/49Uwc4yXL1M
hddPWauMFkYTeEW7Zofw9qohd9sp+hq7Szo+Cjpplo2BsWagyfB3pa8ix7Z/AsDOuboIhNUTzN5P
ebuN4D6jXNN7l0B2K+PP65iOaIABgQ6d2rKutMCBE/OsmCArWhAYEyzPBhgHlAYc+9q3W+tx9Sy3
90Wh2H7wpaUgPGfx9xFgQS3ku2RnUU/mSGLN8ovdFQFKk8rU1cnPcuNhzV0qlm1jFRv7srjYNf1i
QB8n+qbWvdI3OerRGsa8ZhK3BwRppGAyZ8JUvvDDnk74Zsp1rWEtKSMgQ7VLF8z3K2XaPuGCr6vf
i+lglTrEUOD9YQWM5x/cce6XAo8rcscN+lqEIUpHffhgN9yTsN0K8N8SFth/OrzRILh6SfgNs3La
uq3216MoiZyQGt9yo0KZwZMlmxrrzsW+MKbbxMu/bxdtQPKe9ikI2RqamXfAyG26XBH1cQfx2T6t
Y08JnMSpF88A83BCcTJYc+d7i8lWiBd2hFaNCRQlmEYKmsUtv7d0wcubXm4hS3CuXzy1c0sHwf62
K0QqfYjTIBx748MUuUjUWs+REp6Z9xJVTUGCaXxy0iYpUEwkhGqykWmcJs7rUn4RlMGRhNdoGN+2
wQqB0VjLvvL0Mzz0GkinUmqxFAldM703XPL3l4E5VE2ixvQEipmjXh2Fbj1j2jiLkXsShBlQQPEf
czopENYvw/OiQGXn2LmKAJOpx+yBCbSietIzsQWfaEBnWu1PbzSGhXe2UOx85gCeRdP712dJn21P
lQrFP043B51oxa77TlRw5YX0VZEBHgtTsnkf8e0bont/XKML+4UYlGT/p0arGk/R3xCvLDY27atL
mphWKpLfEaZEA1rvLRC4JEcjy4m7Tbn3WTYNxktwkIgJZG0skpD7yHrHcOh61e0psCd4f+6mlVMK
iaEaEFB8EYXyb1LHFi71Fj6Vza7fhTeboSLUZwjSIhm+crUC2smYmJpC49F8rw560Ho4QVAR/pbB
WuWe1GZ7uvvbQtybg2tC5/2KhqKkIEGbG610dwX6CWjSoPBYMrZt3Nfp8yA5o1bSTgGj6FImeY09
piMQos6XAPnQqTRuERsuxrULmUnU7wUgRzutLkBmCJwMgDAg92lP8w8hQ/qybSPKyHan/Q+5wGYK
+FUKrGnpUMCL2zKr9IpJJDMisit8ja/g/3jcy0e4R/agWVqHWFU8a9XudeXx7fSjV+joRO6fopRp
SDntEWR0D2iyqHogJbUIJoFAnlRHredRq5sEcXFDZW2plFl6oE2dp/iQSVpMCtjyZRsqKAnl0tgZ
L6zfnwHUuX0amcCjb6UA7HdGzBBxXZI5/HOQdGWhp457NpEsTtf8LUWkYNyCUIAQGtJRXz2fRMVH
lTAMefAmhOFAYzIjna/FbKQbwFOjsCPklePbt/3yr2f0GwmeWUYTj/tICvsdEw+Mx5RG+pUXe/9P
0S/0J34tVwB6IJ3ciSv8SdguCClvBxpl5ffTP3nF75ePKzAfyacVOmYsqTJctIsdesFj2qXR/NK3
sBziPHuIa+ERKVx2EIKcSn8QT9ZXO/Y3GngbECsC8DECEd+4gj4ybMgAh+YC6cnFxiRZXvOfXaGI
aBzCLsNezEfQK5iNj6iz7R6LOtIlkpR+2j2+JldHNDuiudppo3ralAg7agCWfTHRmqkOLDQ8NRr5
x2L00Wi0HD+NYntY4saCB1a87GFulMaNUOAZ6FNYj/Ei6gbfVrkwY78oUMBtgJNQ3CxhuVxWpzKX
mlhY6RXcobdgKhlkpFukuaaihaBU5t8DZFWJEk1+reKxn9DWMwAAGhoilY/kf2rmCjR/MxvEIOOw
/xj1+zEzVecNAJ5ppWt8S9UTDkfPh9w2EZnKpZgpHnmnsbnnJlXQcgEr9Yqrp9QQAM0BuSoiVK0E
7dQX6u9uzIgeaSSNqLz5SZj4HbRMcjG/bzMae82UOZ9zOE203pAo8P7pRp1Y/3e6TOgvmgMrSUeP
8RnvKgmAjEIXZHAslVJ71bEsjGXesnFhfUNNsYky9+D4pZSm3tPIgadNNFOVjb2ysqEcK+GSR5av
REhLc2K79ryitl9BwRC4i0LijosQBVCqYrtMmwitS0Ks33q1grRwuZnvkIa9AvuD4N1stYA5LkEe
sudxi2LePNSwNkNm+g+As6pDuUC0NARf9N9saW04UaZ7Hp3yc0tiBdZz3nxvbMCYIXVdrPpfW5Uq
jMbY9C2cRyIQOJSY1eW9fVFGBhdiTb+tZURkpk8JSRhxIHGBLBtqdZkwtJa4XPATiah9HqD+QPR/
0HBBSeF6tUoTPXtL40wh8gON4dfopOVvMeIwbgCs/PtUvuUpbzrdIak3YlrFnnF6pi9qQFauV2Ee
lkiQjxSCF35NVE5Ub3GIH3qQt17c+z7D8F1n9rchjzA4yTgIXJsnCznhiB8Nw6IsS/LjPfydMy6v
LjjMVJgYTCv8weCbLW2hZw+rpfq+YkKsSe4lJOmDO/BECInJq/k0tpLltw4FoZqqR/0UlhWXKK+K
PF7azF2j9Mnk3rkzFWMj9NuiiwZyLSnQ7Z3hWuzgbz2bhngo0g1JLQf2ffD15YOA8HcTXgg3o3iG
H23lzWk5gEfVtRE0CHhmSWR9hHeR3751lmUXKTcIHxS7DjvvKSj9P8U9xVlC80yeo5muClYs86ZK
xbb4uu44uMo6ji5wbkuwAeosBTiK0+bvRRplN4EIliig4TBjj73YczwYg03EMGdLs+/rfylizz2T
HUbyrchn0XQm/tATzfHgencNurR5Mh9Ut29A6omiv55BjBu/Oc7RKguezSkHlZD/LDm1+xciLbxT
ukVQpvIb7LPH9WSq4mLNsmRR/lCgM0zgFqqr/cFzW8txtoLoG3b9ZtCKH0Y3DvpASNeIZBGeFaDh
vZurVSjAlVtnjGwXrsdRGC8/PYG5qzuQ3SrxxKhDg44D49d1pgoZ6KMBvIcMHefCXUn+6I2KCDE6
tOHw+XXdF6V/9CWj+PjlFOvde0CvLmReOgNUJh8Bnl0VAYrgwQj1mvwP2K22ZMnh0D5MiqSv/Qzo
t7KFf9983pn6O7yNY56DvTB15CZGk5lGXQ1/HDprjyHg6gQ4ZSiURSH9q/sTPBizCumfHNVWovND
0PplMMTQLf3fIRU5alXOMDXohD+vnr5pjJQl6GMTSLCVTEOIQ3ZEXOsmDCSbvZ2wpue/bL+3vOO/
7Pa+fiU/JHrYy4mawuKZwPNEJ75bKJR7qGaleL2EHGE4ndHSBuNqRd2nQMIVaN9q08UocgqTYLYI
sYpaAGxw0Y78qJK1rA9WL3U+qSNVwsNr741v/jgulkUjc3C17M5qI3kEn1O9Q4X03RwGQKFCCjlj
2zRddLPe+xQRz8FL/q2+9SBl9lfOduWBC0FhRV8sYFRyDHSJ7EFbGjaf3CUw+st55kX9UYg4Ehvg
2k/BbpYloqhLm5MRF2sZBMc0r07rTutQ+e19senHenAOW8nsEHSQBJ5ztmxaAsBWXt/WpLPsy0dX
/lmgBi/jHtAwCQdKofD3sNEp0CdSeg5HEc9cspFuIgGzwfVgDwrWJzfS84PU4Tc7n88M697uRHsG
SWixjhAEf/3hvVN9PnugM2ewwqsyX3weX+SvBRrX82FuamYJe6VM4VlJfpQOVuIF9aSqp8NEZQVW
20HaoCxS4PBajiQAJIbFLRNj/eVJb+tRYMjZJmVpb9cRUJ0ufUR9D8q7zx0EeIaBIG+F1KoFQnK7
Uh67IT1sUf995wybNWhiChtQfjIJyC3Wo7XaB658xhuImHJzz8GFrY+3jSxoGhKM+/JsS5S5oo7k
4X4Tt+wENnnbVDOBzY4kmQXJcwmWfkPkMnU3zLK4QsqlQOTVcidB2d7P/xZC1t+Z4Y9Rxedzgz+L
f3buNzUtnkDnAaIMU4fQFecuDcCW8WSzddtPs5VinMlYWTLPYnJ7uuPQyorCporwzHz0NP8KXWeO
452eg7wmODXpLtE/uRQY8a7ZyZJDFxQz4GuPq/smP8FMx923xX5oKBtiu1VojWkxr5DClU8otT7r
2H3X/g0LNVz+uFKGp3TM8LYf25IuLUDXWC1utSqhJNsDqC2kuH2FiktCQ9QJzjcY53gwmNNwKI0y
4ZPfahOciYG220n2FmeYuMAGK7AaeCucGe6kuQypvUKYl+Y2D4brSLWKUT1x8iBxIP/xBOKoKE9z
+23cL0hhP9l3pFplmUEyMFNpslOxKZNoFgFM7yKx/uMbgwoYERcbKK7JeZropRZFZzs6k0Uwm4KH
Sh+DdzyMCPFMxlt01SAqqze80hYn10wQZ9lZ9fNQbI/kRLBCaLd01qRQuqVj/33wFlEDEGjycUzn
UWJgbQ0Ba4U3N+DgBtSXIrK2qT0TkH4l8yzxOQ37i3QEB7D3J/bKHKE5vpoA17q6KgcnBpXDbA57
DWf4UvmCVGYIoZB5IBG9uxslSUDImsCTlWsIXyNpNx0yABG0r4TmNcJQwJMYaS+hRPosuVbMfwdM
i3PEPnxKVEZq2/6iZKijv3iP2brcO9ssZaum9AzfGkw7NFE0TCng3JYh2TUEHfrBzmtBDSUsNy5D
AdsGDmJeHn5fui+sV6ZYdboYhjlu6zw5Znk2Z+3mxeHPiF823QTJgxPWHzWee+/7OqD9yv+1UuY+
B3gKPTCjS3eS3GmnhKG6w18FqL906C1R4EyAk1ZQAYGGLdZyN+w24EWOjKAvQSJgoxj8io72XqRh
eaBUzrSaiiF5Xy6DmfX67t4bwPqYuuAU9M+p5wSUdTmESN51BXW+2PR6Y3Kt3kDlhdtR04aF3UDk
NPLyVQ6okTkYU8SyQWX5ZrWVBYdRkjZwDOCO85eJclukkZ5Xy0ofsDUtPulyK5wkQTXsZBziPhV7
IE97QbBOak30kyZHOFX58z7C+VTOM5isWZ6ulkqWvEK9M0sYs49uvWWo9TiffTpZkSWQlUfa7usi
mkGmDrYFj646CywiRrd4NN4KtVflbgxQsqlggTpJ0jcedUm7HvIv9Z9uaqVAT97TTmmNN17YGuGH
sAUmi+apBxSCYZr+Yxfti3f86piZVMhg3U8qhh246qsgLYsHCFPSP9B1g5s80NbkyE72U3wi80pC
ibr2+d1w2YESBQ/dZXsBMU9aGYgVJD86i8yFyqLaUBJDGl72D2EXOdzwGN19Iko3wQnMuqgR4A38
lMCEB64SPDP36zgf1IYhhSHBnuC01Ko9ImX1tRBvflSdqlIXTCB7DGkAb1tomRdFTJCu1Wg5b7ey
mtYciE2G0fA8g5MfuDghfLApqs6GpIvXZSH2eURR+WxL5tdrWU1nR/LCYQI/UbZGIs88EN0ScOSV
CcIYbJzykcTmNt75HDUZEV7J3McNtP3qJgnhjNV+5vKj8I0BYfYTr//583chWDPkeUryBpmgKuQP
dnNSppP1964G9xaAVDHypPVvj+SgQtHIu/3k3ysHI3A9nxmRE5eWaFvlIeFH2QGrHrZjmvV0q//p
KFBNc0+nwUx7ltwwGQdjTVWTwmVqQapCCHfm25mSeLyi4CB1+1IXWNwTTGZ1MfTuhd+9z68WqLEc
PSSTgVcFQZD52EqGFcRmVj6xvgqW42S35RkCVSvdbG1wQnmrUgKkulZ5qOLNh1TfJxISNcDVOxKD
loJMYSA9886wz3A3SJmmT7Lx0yunzBss6tD6cFoAuzrlHcy5KJtLZYhwHbd+feIyeiXlm1kQtWOr
0TZpLQXSQtFxpPNKeMEJ8roThUif+S06WbJDFPUNpB+NwnmT5pnVcTwVc5luPT3HCVCX4kQ3iEmb
E8RjB9eKtFSWtuodNEmSkKTUWkOYutv67aV2NWcE6b1RfKFrns/HFzeO6US3nb9GHRrDaWiAqf94
mLhXYVHwjCzrTIDDX+MJ1yGFB+Oz7QBTkgb8Qe3IF9cyWbW6kz9pNEeTapWDCVvwCeLtx0PyzHf1
meJQlT0RAJBPEBfeV7q7jNV6AFOsGjuVucmswE1EotRYRPYVftRLgJOEOUNRHqzPQU8oZY5I821K
FvhyQigHKfLYs2CAP6npKoKnmSa6AJAQR+9ru7uEjpcIxtmJb/QulVw1hSnt9dUqGoIZZsIhBp8x
1fP/x0yXWnJq/5d+lSGiXlIOLH05Lt+1Bh0CdT8bBNn7FmiTApm4PNbkEzVE3inoETPQkfC4/gek
ZrJXHx6U+k+R/k5U3au8BOnlz73e3JPpbSCbnl3k0zdt4MgYGTqCYxFkScQ3GsoGMnqY/MRxc7SW
Fx3+SyX9jM9Ib56VEERzYu1fVyykgVFmCYuWDFhaAr98Tw7zcM3twAnbSbSCWAfDwDlOErOwfWuy
VqwCwGQxS1eGG85l+aG4VahAv4Fop1gfr9kKhfjkSYtEpTOr5AIBrFF1kK9Qy3yyT5+9jZ8W2qna
jmPO0tKmcJFWqXic+dmEvPq9hHSqa8sgfzu/1lD+ehIVuCyKY4gAOqoCLPoG/6a+09PedCb0+5+8
LsDUQYU9utTBdYedzBRk5VijOGBITteeywkY9qzBQdAfl5iGfsad3oqbVtfg1oTUvsXuaQ+NTtiT
1YmK4P/OwhZE2T2KLszuze9Uo+Vv4IghPZcSstnQOhtZN26W0VLxJZvJoD+VTok1EzJAkvo1FYmd
h0MpTUUZGEJSy3uCgFzl2QMEy8lui5vu+A+fg6eTH9PN5GFndxTQKcsGfOX1dDOHB4RSkRLJDRkn
u/O1BkKl7yH6ubVGEYozawVwQuuOt0JhrMzmwzsEzQMOJTvrd7q3ibsOH7XEOnjL6FgihO2ssr8J
RSjDsb60z69y52OQx4xhbpwjNZUToiAazLkEcpe7+lmCCWC2jrkgwrIBcU/+swa4o9tNziFc6df3
tBFQf3skAII/+pwoa2wQcfjMZTJ4b9ycF32o5JCxlaVfNrZrakJGgO7hlmtIzZ4K8oLFlXzI7qM8
Q9+c3xX5JYWOcxdczfyhhUSR02GMSiSH54dTdLpzxK8QyPiuN/BIavaA7QAbolbWEwzRmGCiMene
uXtej8V9+9C+12U9HQofWto2lJlpII+4LvMMkAUBERX1BkcKgaSJ5KyKGiZH5Wlx4SHvWyk/XzoA
GnRseNbvLVOpgoOsGOzFK8R6HsNcKeZh0mqxqW37k59BQE61zyh5GayvWOvmZSzNRIIjFchvbICk
9HCdcZNMZnreM6XrQXKtwhZ6Qsa0tQoiQXMEpSKfsdjY/oKz3yl8AMCosLHS7vmXU2Tj6i9c2NdB
zcHD8cTr/r4NL1gRisMuXULbgvI+PWjBhRPu/Nx13IIgHRuGwD7JelUyEoE/Q7YpKyIOc76QI62p
6eoV0Ce2vMCu3eYqgb/S42nsdPyjgalV5eqR/2CsTnoNpbU967bPF/LQrnM97kslO0vMRvMZBo0f
D5wfSIjnKI/lYhK2v1M3OV8y13xzwrTxNNIic0Kvm0T9XYtTE/5LzhLqO9+Z/s8HykSSkF+GzllS
RsB2UYHTVR4Rmte+hT4RvGRgJUaxzn0FO5GoKFd+/kHrYlxx1yyVh168Bueuo7FtflXNJXjZEM2Q
8NXyPNO2+EsibsKW3wBMNFP+GFCN+cfLjg7dHWSOazLFHicYtInOjlx6LaxVZi9S5iUZIkI52eMA
7Mn1V7SqWhWcgbKWyRdlXq7fR8PV/LVSPUSqCavsbapxF17gn3yJrLlI/T9xqHSQPVFz4igJffHA
kSIASqnpfJiou8HgtZg+UtDkttgrsJiXd0HLgXcpmPGJS+yyq2QTWbYtyb0UbPW4sfgSz5zocoxw
H0QIvRWzFL2xc8JFr5rR9jx6VNjQCMnYnoM95QjfxVT6A+BvHi4oFwAa4MoiUEFHnjt+vIDXNSbR
jWGH5YGE+FJLIwwx6LxMGS6tJ/J+MwVd6+4bSZCCm8jfcu1uS/cGXLDba0zhB7eZGTyg1YZZFOAC
Y3vpFOjaZp0c/icKrOe2IPTJ7Nn1nsBlsZhLztaOfpjzj8PpavOFc6r0vmrGAr8FtoOEcHdeUyCZ
ONEwqtYKPCqSfu9WuSBft676fLokXPkgSYhpss9yDQ1aLmJno3f6dzVYIsOLMFEEUb37nPnjOFJ2
IYeb2PgjKzdoekxDSSVxIfjvcoOPo0ELsy7WUjkOGzC3nw/A/YkLbM/1Fcmm/iXRr7HibCDQkuOD
O6Y6YBv6rCzmf1b7N5iT/sv13BokZJ90wCGAIERK522LgzJBZagG0iv37z9h9nTHDpStIBQwcHvA
eABoYHlhdMsY5+7TidoydGYmklS1SAA7wBVc03pV6aSaLIvuBgX2QyEC2qFypT8IOXhRuG56YztL
q1PvLIzDMGMo9VYo2BAXttvD+6w3kCuYPZgABq0i0fa3ysTGp9DwklMVoHxdne9PXuXs1w0qGRu9
S9XyZKVxNkQv4rjF6UKG7A+uRxZJblaIGzLe4slizqog+pfAZTyhLScZPPN0sEfo0+hbIULeqei2
tmCLeJyHylyJMMR/gQD5FuiYZiKejB64+TbEeYS4yo8zM6ODyQSjgUm4E90+co17XbAsiiRICigE
Gvuvd3FCQBFckH3JUN80gtQwZahMzxdhdFJloxFdHN3zxzmgiPhlCQCxuF6gXG+4Rv5rK/y/XRCk
33u+K+UdNKFWv8OZAq4Rt0B1qwyt6Vb/yRVCTXMkq5S+tLhHpQiNDEeQmMwV1iOeAwNMBNJyYXNT
KDwThIE5rYI1RceNqySblPNlKfz+iCnXw+IqIdFZwh71+74EBF6GD399R6Gf8fQbWCRt95o5XefT
G0g94kAu3rGA0lAkndnA5rwT2P2F7Ag1/3UJFU2iVTWDPpCy/7SiGgCjnExbIv+reP5XvRSizgKc
2YZNyPNylxYjyauq0eq2G0DhircMC0VcWupFS/a8cVUBI9/4WfatkeOKmXLqxW+y8KUv0p96Fawq
9kNb4Yo7t9cUzDg8SVSpxcWqD+mEknVNxYbN7qNs8njKOqFambCy3ypkZQDOGQG4QHNF5H7ObTvu
MV3PuPPNky67n18S8IbZwdYSjutvmvfMW8+3Z6oBF/hXqaT4jzZHhvYVimDR/UvV9r4iJojmA4+k
0oMWIUewhqE22teOzfw8e5HVffZGYls3M3gal141gnPmZnIRQ7hw9oVyJcgMPtlJYGywAIMOxf60
5Mynsa1+1miaUyE19dx2ryZB5LobWzH2etSPWDm4bqmFxYthdwqgkcoYbeXXe9mVEPqFCGEexnLz
IKKpvaQQYZ58qZa9V2enCzsr1SLRtBkT3VCFXZXEbSnp3DgSLwstApmymySCvCrbmnSHH2Wlddvr
Uk3/9xsP8+ihYneaKeSqsBVXomkzJRLIhPi0Ljt6rPuVWpXj7yuPAeLXa1U0L87Nt5IRO6mgfzKq
Ppe1D3OC+Pbz0iCWCpC7WNZff9Uxmu8Tqu0zxPY2AWs9mNGdVDrrZB1vZ7tPt3YXXcTWKKAvGUBe
wG5Wk/cZRIjBoUKFDYewk829r6IxhIZHEcmPv2Te5udBRMK0cIFjhnOFx40zTNV4DusCHP+K+4uB
+NjyVlg++7igAt9tBRO2CmouGBwziITwrJWJ5rcCueNrmOXuw87aEYoM2zmkvy3oIAn9ngnKefUF
N03GgaVwSFQ/blLKRoOe8wvqN4NKAbZoPKOHMbAq3uirczgsHyLDASyV6fkBIK46VBxJtNKg/kFn
MrhZxLfCaU6usZQJtnkfiFrcy9ma3Q1OipsgOWHfKsIoAVWD8xRSy4yT85gND5k043xQSUwG8tsy
cxqCtlSuRcj6jKkWO+4FyKG5eP/WaTcsRUeyOVJX8HblhzZeQzV3192G7K/zxBb/hkvlU4IxB6+V
Fjnov62hBm+6AlW+3WnRyf7DvnLK2tuFOFuQdM9cthSdlMjeDtWYHWtgmuRakUii/aoGXOqsqIF2
t2qVrOEy2crDBnbmMsSb377KKkzah3OTW1mCddFQSGoSHiPHkQ6sxEEgOK4nCIlM0lsl9OXDAy/U
ZESdbBkcORbp+w37Dv5auijwwplc9upWbNr73twdY2b8ONrgS3RmnF5GWZ3xM4GEkF0TwngfV6JC
O05tRWyNDUGT2a3iWJB9fqphtYT1eOe0hacz/mR0bID2Omxq8vEeRs3kBWr2T0JqNhhZ22R2ckkt
q1lnGYlWmCv/DbUJML5sLTOOE+44HIS7Y3hYo0ujv2Ew78ns5KvfKXeRvm7TnAxz9rY/A16yBTJQ
TNKr7T/HgOmaNVTBx4lnjygglaJXRWmm9zkUKWXQNMlgypCrjMn4P019LrP0Nf/fdYYvAEqA6saZ
iuAtptxbSnYZjcu0y0PKDv7krS+Tc7S9aXM/T/KTZmb6SGh1GpfM9JP8Xm9W/i8givHbjBUYbQNa
4M0L9hiQmRjQVEibVZJdLiiVcWqHJ3RUqr3kopSSs7G/60VvRXEsHRF3XCzMPc2JZjll+NToihB5
ouh6meQnD+XdrGadSxwfQGr5X0NzFzcGAEcma9nBMf0V0rYSG/8lwI8FqtPuU+8g2pxrGqSZqhm0
DWdYH6Sr1+4RTBsudR5WBlQMrnqQ59gu+LifLsuMJ6hykRTssdvLUgzvzlIbfmxVRbO9KG61+zTe
oc3ORpUTFo3YwrXC1mXzaU3KzippgH7OTXyZd1/g1dduGUCcz5UfZaC6PcRF8ukMRs9NMpZ+PKdd
dFFMZrFx80DK9TwBshZNwARGAwlX9ExOrpG/6LPMCg2SYZ7EWaD5MVbVFZuygKbr2+m5xAkMtyIa
v5Pl+Tmx1jhdF+JpH/W5jDJgcfJJxQCCAyaNKPc7/mP5uOwRsykRYcFQqEFQe7i7+KQhoqIQ7Suo
lAbkU0VNkdOwgTUUBrWftCs3XKSoK+PWW1c2M0MeG83IMfXyLfsMxv98jpA7zV49A23WHGp8tH7V
AXJzPuEtUtQwrT1fYI4ysIhjR7sesiLxwuGdxgEkM3S1WBmW0raOezYAnUDwfqT4t8afrjDn+Rf7
a57AiJ5d/EjNP7Eh11ber7NNXdft3N321oa2fJbux2wRjRCmUn5MUAvZ3yObYiMaH1Ul7drpK/5E
+3II9kb74felyEjZU2Ik1Jldsen1MDDFLz6zNL1xZoxw4GaMd/MnK6qUNMUwL6HimyToCvbyhLnL
EY7qJwmFhirW+3y5YaDugrFjETlnDjnbjiJcRBHlURwydVuO5iJ+vDlzNpPuq167FWnX3YciZpyk
hh1HKGMinb+1N8RBSsG4SFiAKSgdmEPQXWpygGwFIKn3rHUM8REt2llUthscJUPsZz5Imi8MOXdp
L01Ih4QuikPpfD0yDwc/0WHwVNDOipvGEjNOl+bSZI0DjxSjZBuOdUYo77ujCcsmCl8FcY0jIK6N
AR3SX1u399aP+0JmNlwrocAGec7eGUHtE1IF1+BVNJigfaDkb+mJAHxroeXnAMh11UIRK2rH0nUd
J97PaDdNWtSvkKiZAAlgy/akWmiQeuZ387LF6In3N+d9mjeuPj6znaAX5BiulaCW3ofCNhEPhfyC
AJY1Lpr73nQlGl4ECOxfxK4sdyAHIYIG55HMq66j7UEo+jy4pEFyQgYmEcZmRyAFCvDxiZOHvvMg
1IaB5lbVP4JfShppbMzrldi4sMV1jtaFkVMK5WoCSBHlOGNm0ETctZ/yZaMvuFDM7t1DU4HLiKYD
8+1TIubNdP4YfByClofOTFhmyMsYrYg7ZT9lfmq5SSB+DqFKhzJd4GHONrUfjT/vremtTVa4SPQ4
8xnDJBanvRaGwaQqbxP8tXLITq7p56/xmvloqPhkojoFK45OuUzu6K2N4GjcWGm30FLjYLqXJyXU
GYILRp4vNpZvruZaqkV9lShZfjTb8r/YJ0K4qe1KA7Tjx5APmzE+Sl0F1tqSvISf/JTzPP8we7Dg
h9Kjt/qg9SUNInMZQUSlmwry9u4M+lJF7bHvckHaSUd1chZKAGoCVzjPJqgR51SBPmFeJZlSjK9g
Mky4bbRAuKI4yXfxQyXyYsNKFB4P+Pwg+j7jfTPA5DDIH27J42zf8/mK/F7W1FUxbMn15TsaD3Wx
KhBu98+g+yFGKPnT4Xhan0znWiZU92A37pAvLbyuHiBO00Px8pmXVHbRYMp0+fQly90UHD2FkulR
D+/Zvr5Wgu3mXHl0FftvynxVIvoc9XMTDL+nuCXAcCwDWnjl2pTAMGvzz6q3FI1lyYD5C6Dj4cLh
ivGZQoxhj6gI0Bx4i2OEpzcNsy6MhlQoxVCxMnlCODMUPhm8xgiEogquB+I3H8jjGZ6JIa2tZAIO
iNHW/jtcYVN5neqkU5ZrE4EWXrgQ42C334Zpo85MqQpjQuVsZoLvUc75+hF3ZZIB9OcdywNzzKQN
eBX7gErm4MG3i0KXXlNfpmLazQHOza+2L+YmYWoOZTetEhcgYyO/MiuQc9kLNGZa0cy+lWSvskj7
wXuHwY4PBphxX/p3D6mMdJb/Wryma5HgWKjGn8L5iegICXIHZzpY2YuPRSwXMYAFJZvVm74InNwQ
zMMzZoGh8t7/mPbv2HjUye3w8Y+0VlMGmjHKHhtLRzhrPWuT1mRvqSogJLihaouXH7ynXjw/XcoA
iceed+ETarnztdW0GZcsUIgrBylh1RA2cPC0vouJWozJKSXG/11jKs//v07SXgViASzKzXzjixCS
XXWyBuHwMnxhYQP8Ehqb4jrwVhjCrsCnZjQvTBVB13bfpgY0AUEF54I+pIdmX7etFmjpPmPVMOt5
brAsnhIHiwHxJE7/cz5kHCNixwKj359E6pUxHLPQyqHdbndXDpk6+9NWoHx3tQNDir355PdogQPA
f38K6PTDOqs9i1171S7IvLjV8+O3POU+v9uCtNtn1x1UlTGYeO1JC1mXEkYZ85o3OZ2FJ02v1fqJ
hqoXdL/MTIMAFHOZ6Mve7nZ/ewUZWGLcSXf+ZVj8D4NEXAf1T23JDDxoNMcn18J9VKNSOoQnIyYO
+EjcPaSQYvuJhqTv/Ndbi9GgED/KEEyRtrx69+qetykES0/5qSzRftOxdr4+/KItF4JLWXFGNPMv
c01VAHx1qOghl8dYBFGJzaWZCG2BQ+KUc2NZhCq3RGVZStPw8smJD9EJQ6l4QSbgQWLNJI0miLtw
vhNoxYkybMHJYAY76E2SkZM0L3uF+UFsTtA/LlKjlA5oF29R931btkF+NGKT+bdKnRhjxXiP1Biw
GvI97c63BoS4NEjcZNwKXBx9bP302tCa79Ogg4cffvc+i+hswqOdFwng0f4GR/dQWYkN+lHGiN6H
ySgQMnwGxCdEY9/iC007RoN+TfO6aQegmN8+ceVjsQzvQUoFVzfKAJWD8PvA/DrWilrDbS/Cjf8C
/tSVw4YlvFyyMk6mIyCd0FR8jZhRLxTsjxIGpoxLEv6XoFUitp3NiG1uP1kt6KKPr5gJmWknayto
68WyjP81eJBjiiAM4qTBDQ7tpUBiJg9jW2pCXXZg8/bbR60FUsdP/ctXYWQpRSy493AdeQNlRrfs
F7FgvSJBhF3YhBq6b/rr3+Ab6A6GwXncx4kucn3H2pDICD2GWI7NVMXfiMgXvg1AXgWOT6Rv93FL
shRCHSWrxhqQBSpd7/0ImUd8g4TakhEB/MeBThUSNF3pUvRA3+aDG2HRfKRh9cySlZMVwEk7RYfk
uI4PxrKu9PX+Gi+CvnlVELD+nYrZXJQgWmcTCEunTHT+zc3FsEoVmH2FKfHs3CwANKTLMKQ+OyE1
gt4RH/pbVVDQYz/gMXGa5NnGP3LhkrwPVV5nUFvbpe6FYzFLRKd+rWLl4gcAAVNNmogp659avoHa
DcylKJ0Xdw4OLG7wce6d6jxiYED3sC7mtnLnLcmcxNUAMJc5dIMnaXuj6dn1yjE0HJZwi/9PXvTw
Q1ozeWYRo3JjnVW60cKanZ+vI9qgi5fTxFCNYQR12PRFfncUy+1kQ7kZjV1YqbF5GtUPooaP+N01
WirKZMUtGd1vDJT/CR333cuYKvKK/ta6bR7ev7ILmG+BkYKxA84THqfDhZ3lYmfLQLGxDmbBsDY1
+sKXGnKvdl4sND2RDkL9HcU2DEScr+8BzZ6iGMkqy3DdYNg9k2rmMRt5hunN8onf93Yg7aj8jBQ6
ZJ0/2BgPf2S7J0jylvIZTE/zuouBrRQGIUVROz8hOAAkV53dQkvX+uRZLLUE7ANPL29XkQsaSmwF
B+ttjdLUmPmdblNOAMBS0+MTf22sh7Z8TO0Pj3Wzr51julRPIPQZX216iR+qdBzKOCMMstzmKGAp
7TS/3iSjoM8INy60efQrHHEdKGJSyhy+cUVJLYXXE1XATXq+/6O48trtQw3KGTMW1s7L6XZuMYs8
qTrxDsWzMy5TSzrcJas4le11/gF0Pfq8Zc5eEaqYUePfbLz+9/SSEt5hvUnyrdyLbJPsQHBvvoI5
zTQJcFlACNrgbDw/vWOWlCZ3Xff0SqHa/K+vb7XdAe9ZdOtdSrWsIFpecE+6O3g4y+xZiw3l0XW/
QIDX20QPGDCckVNfVzTYlInXqo/VOELT56gNYPWnsPV1bYIAQH+G08Uadl8PcOIGja7W/klAZ6e7
xSBmt5iINmLLEc6G9/qJ9sa1rdONerWZWtxW5hgkKLaUHCbDqz+BzTjEDE4Uj4f6HyRC/jEpqPgW
sZ1JtImiVnRjgfUvzH9GL5WnrvJ0rdekATcb5jJquIboH3I9W2JMnBkPciex72nwXPyyxIggroCI
aZimA4+dEvGqaSYfx3WgKDtJ19uvLCXSlBrp1VrjXWI89zL7TIFuAYRRwLNYAx2v67wRnDX5G7rb
/owgpAItR+tCgd6blNvys9brydNN7U9+L8BzPPcYUJjLxhc77US7YYB6KfDBOJCon3j0/8VnGHdU
zAkJ/i05ZAWy0Gwx7C7wTM0FX2HB89NvalY3L/iIuR9b7d+ecn+8g376TahCoHGSY5WoNePdXoea
UWcj53EsLD/wOqv+WvZd/AFoBIyOP7rUHZjmGepA+OD/qI7ICfyDJYzoGTUJRIEgPTQ1a0/XdwwV
A46/zS+IFepc3ekcgLewxmdoXUz2VT1hquRO56E8f50gyjAsQIX4DRPsr7LgjeoLTdzcNxEIv6lX
wANL12Rdxi0YZvyIbl3x+lwUK3crdoY0kubKNkGG5ws1KAPgxxnjGJE2U/pk6f+8A2mOLqoz25BU
SK+pXyczOcgh8BNDmG9wDQD6rkGgiGFfLzP2OYgFHsCi8/O8cW4M6v/Glno9umtTuvLXCuNbxDf3
/7m5nYI5CgGC4oKYPbhY4x2Pq/T1pWeA6HZHCQBCGOdq9uKuz2vjtgy8oD4d8kz25WxTPPCKDEF9
ZBWpa3VfsVfjiizwEecpb72akK1OCmQtiyMa1m7k3ylXjn9lzngo2NpweSUx1GPORsWoYh7fXvwE
JY6oMaqZpRL/PmFnuZGFENyYljZEKddUIyPPXFj+63UMN+vX9eMd66IrccZs3kF8bbsowgXsjYik
2708K6AnmDXZ9GB5zpcYD7YbiFdFLxmSvIG43Mxmte8s+/sxuZMMlCrYUQ+Rmh0doYUyz1DvOHPm
wk8ikP/x5LZdbNrkfzrtlAp1S4u4bKBAsu/HrwvqkvRBJJIIvpI+qT8NvK57ejIXhhvuD2LwwN9v
hez2jp80vGKcF5aYSO8oPkrKuKdu1qBb8qVAAOk/Fce+mGj+XGiCbEp3JtdkDXpC2OjBva4e2VmR
TbC2GA2taYdcJ9NhNs043Ooj/tKiCn7dBl1aY5hD1gyvKQDtX2YI3SFDGNCFr886MhKb21LFcP++
JHV9NtCrWOs7ZEDxW/EOwfBESjPuiDqsKpQFQ/0QtAlHwyKpLjxduprdCcPU6OBGsSZa2DwI2zRU
EC3MIA8FrAAWJ765PhJZQyaobBe5Im1MKfLh6LCuhckq1jqe+6E/tiIXWyxINguIX1vdjp19bEUl
359PZcw6Vp7NyLoIr4CQVI8ojkWFYI2x31/9g/0HXiJfdDceVm7LHTPUEdV9evPNq967xFi67zYh
8Y3Mq7LJj6WOn41yrHzRr/d1jYNAkLFwDUHi0g5HBRCI1Rs2aZEzp8gYBlU/1vgfh7T5ygmraOKL
h4WdadDZwvu6TbaZBpeQTUz4gfCflAyUmhqvAZcfM5UriigTONp5MLgOJyjZCQQg6AsZRXPECWTh
adtuwB2wEmuTsnnPo+bXHTauSIOsYNAbBruRJZLbyayKsNtdi1MTFXlJxcOQ9W6NvCyMqlsKtco9
g1Mzr7rTHn4/pIMoFAjICvW9aG4wGTHLvPJUdUeAfXdhqMuPxeXm5Q9kT3n7uRIPoS3JqM9aRTB+
kvonlwJ38WyLDJfV6TjocEul63eUUk8QbgAipScW31gqZJ+QG9w1BBxdZnW/9VTLwMV7mzgtwqON
87KGchNMXfjZmciURiD0eFDjUoJBEDlZWVJVo435MFAY0MOCq39mblGyqHHJYA9o2gRyJ5dQc+gE
KAEnvqZ8FZ9qWy26K15mhY4p4Gx14mQk3WxOCGQhr4kfXO0HrsH8LdymI1/eWpU7iGo5nKfsJGDF
1iLtGKezFfc54BrOif2IWn5Qc/BK2g5tQkb5TQdYgl9SDstlxQX7zzdlf7xnU09pAeT9g2LHdLNc
2Uw4LnU8ejGdbLIWS1+du0fuS7YZYg+vHTXcUysmcHDlYsXRgDlLPFPp8gLYr1D4GqNcdbhSDx8m
uNw4IgqGEIW8i5F6KxV2Pf2gPfpTNrTVBOv27mrz7ThQSxjRQgsuU1DPNyDr6Rzvx9XyH0oxyBNy
C9ISXaSVP4quLztcYzmz9ochJ54I6b6qqSvBthT7xTmrilU0BT34LR5k/51TQZHnpoPZP6xitd0K
+P22c8rwkZNLmR2o1gjHLtD7/NxwxI65JDV023ne6mGdiVHdJkst1okzfVGoGbq88gWa3C4PBXWE
Cx1b5f9Kaclb9SEDKKrRuIs3XxNX8m3glE7iMzkBmhm7L6I7dTAFES5av2hw4sikgif55ffdn5iW
TWuEGM0oXnVMAxqnwvhlYxhgSdpbRRlB/dzU0LSIVdJ20ppCmwEDFowimw6a/wfgZe8KrRuCzsZE
csCgzjOdRwZIPUrADT5WfLTD49dCcdpGlh9BODnEjaPAPyZRsZXEuIIp2k+Jft4QOVrwzxuVsxNa
XYLz36J/M2hqS/JV8DW+VWWbmLYvPlWInKYUJovrqz/AFS99iCJGZiS+/g4NiGcLImM7YK71Euo3
+nlnPDe5R/wdcIuwSsh1d8QxYf70enfjQah6CoG0aRkIU4IL6srjGcOFZl3JjFJ0YZE8oFuW000o
g/DrTpe1zZZEs5OonJgmnIaqiyK8R2IghyCZeUYaUemA6L4syZLKmdruq96fNSUIYT9JWcfoK434
/CSgY65gMWLhbOw4lAzjPivfZphpg3r52/+fMKnfPjGRPvVzBKqWMM4DlH2EaeWWGok1dTbRBeyO
kxTZubPWZ8dPUwsOR27CpGzsxDqMXuiMKM9UX17BfqJY7NWj1U+8OzIYu8wCxhKqwwEAnTqyZyMC
gIDxiliVbMQtImyKJWWx0iz+5jmJCRIJ6Di5/5IYjOZDBs8RTq+uOHFOAf/SIhlgE4+xXuBP8WnL
IBaB0z0yazTsf3nG6E7j46YPKpkG9rXBV5ptLkXaiVsYIbDkBUaUv7tS00WGdEEDfXRF9PxRA80+
DRjXz4vmNPsqvMFbUKxnowQOst5U5o2DsuCm6cb0a7jOOsYsXro6ns2nTOiXREb2q8dgTSORo4sF
86WE/lptAQ4GOkp+EyUOUJZmpSPfDmSCHLIG1GXRCM0h0QoaVSui3Zvv+Q0PBKSDobIpDEMsnUdC
XkBmFk82mOHjGiu/9yctJyjp3LABEAJ8jhANW8AZmQtQrmYGwj/LYBMJTJuEFQlvi0hqNXd32yhi
R4OzMY9PlyUpFVL48yVjwEBpcX/n4bK0skNBnh4SinY7OpYaKw1b6YpkyszewwXpDez92zoT4Chk
VJmzcBYa0eY6YW0UT+CI7AimGaWPMMd9p4VChGnL61s1jvLQy+eT2+tWTDv+vakCniKuvKYAOaz2
i3+9kxA4yY+sqrr0AxSx1bcQ9A1Dt1m+lQjDwrA8b6WbbZxBOo5x5d/BF/zPzyTdLzDddpUQa7ql
rBEbqveVC4YuCazQH5vq3M4X1YHag7k0n1XqDwAejA4uaWEoYznrCRxi24wmtnvp4nP42msvronL
qlLQZL4MHxmF8x47GiLCswWOPhQSxTJ7oSHhIIpoGdYAJ8zt2lpmx4cTKsfUmo8IW+K4auiF3ZyY
DTZGvHhces2eEdd6rgwuEguvQmEBCtjymwgJf1Y0bB0xCHFAOw4lDVxf+dy51MhRprjlAHTIBr6E
MaXCh8Wzk/uNjGGj6NFqAziYwzpZ30jNOF0uIYL5nUZ/2grCcpKtMJfoGNkHAiMu2winUHeSVf18
ra4dW05z68qnURzHYUJ7BqMimVt1dK8Cki/kyAyvDp0Pn03jkcc1GQ3MY7Jj7bHqJe0SWqdyRCIn
W98isxyNWzCvMA60iJb4ALYlJl1/FIn7kNGT1eAlwOcm3Jz29M/7z+rbJRJrixOW0wferePALAKE
yfB+YnpdiNj6URklWWjkhKpk8k/PYpYx8IViiiorft668OVMraPCEsXw20uIPOCxBSsv7lMXUilv
On0tD4RgrQcCMDvsI7rTYrMtRMCGyjbK9Z/5EmxtCvm3oL7uA5w4NEhkyqcprn/YaoHN7SziSrEk
i7mFQFwPucMqbsrwvD/GUNlnsAFYPVLJ05Taqs2Q/shFoBXFqOOQNJhnxW0G2HMDIQ+AhL8B/+1d
kuBRET4zAEsf2HvbtD+lW8CGdb6t3DR/CMnjCVwy3sQD1+TW9xX+ffPTriHiSgvFtKJmEIWI1zsY
d0NM2/mohxjZZNzyUloJd7BXqYPLgsvId5xRwZAuqE3x0baDa/odYqvUDUgFEx61r3gDI4IreKmH
IZexlYckDIOOSGQptuFQ10E8L0B/HzFUe/dCYysYGDd46ukxU4zIRatVYGVjeRuNLpwr5YeGdzez
IxbMPMgxQBRjwG5fzMuoE7WBa5EP6MkRusoINqGe4Nn4IGxArMWW5wbX7+jwniy3Isk+WeykVC4c
RWwWvAQtAtc1NhghnwLH1ajHrotmGoY0I5u3D6rqVJz+Jc7yUeHtrBV3hR2Cj2feb7N91kLIUGG0
VHAnDnAsSlA48sMibuqe2NRJGpGOKM41uT7pzBPnzdZIjDCJfeLV6pxpvCJBHqV0DLbWIHYDR3dS
FVLrrcIr5f3c70yz+Kqf8UiDud67fTFo+Pi1rGQjcu1tDRaG2YkRXlFVorkSms31APjpGARNwEdN
tgCBKDLmm7O5xpZkh/150abfd7desnDyTK93SgOH7ygj8dLLT0grKQlXSxmtiAhgysOON7LsCyfH
Vj1YI8q4+jxn3HhzXPy6b7tcV8AbvjHErrhqLrtOGjC2ts54im7r9Fo+jszlGOjQOEcz+dVs3uNB
f3qnDOGrqMnxY2EnhGB6J36DGCfwRvYvCB55ODWr1rimvsdDACGgMeqsjaCvyPv1Bgf5duHudtXD
qa7sDNCL5SjxffXk1O1Q0NW1VhxWhTohQbkLVRAb888t03g6/Ka4+lPpPz+gN+du6tpg2BDVwJPf
PzL3XjpfHUZ9x/k4dPRwBLmeys+66mEh+g3hkVtrxNb6yW0thLFyFeZsD5XctqJdUh4ZBSuLjIzF
ZtBfQQ3oTNxF26kups7SSXXB8BZ/x8PAI5OfE/Sy3uk6qv5mkl86wBgbGHeh0tH4/dlsVCKxczJ2
r4a95fL8494Vxxg0fBzTkdH+xDmvGLQImmBjnoTXjqDExnfdwW4HtQL2oaPaalS/A50b9MnWEc6Q
yMApbZtnNz97tLYBQhaEpsRHM9Lo/3CkOdLr5DAUhBjtnRDnMAn58WAiebc1OIPxVjtPUa3/YtjN
UXD3SlG8HLIURsYXCs9NcmCKyU/6CLjbvx8x7uOXHmHkdBGOS5N4x0bdSXrnbuQyKJSmQEGUUIjx
XY3w1/448SPGIv2R1kDJbUH6joPPOUjw61BkG985ulwU3tAmfqYUUfO1X6JPKV4+BFDgazcc+Ywv
Pvq6R1n2XyHxnNx0ZkGsL65xYxEcYPiqATIqEhYxqXHuucJTvOH09GBFAzr/VMVZxHPaM4//wsSY
GNFwhyZVDWQfmO+lmZHpxj4jE2qBHy2oTUUTapwfXhhF8JojqZXHNG602DNwVSYOUmyZu48eBO09
EqkSKX/0f0RZJs3gND/zS6JVSWokzPSz30yNFIHw3pp8s8GHlm5hSmgSy7B2Z1cYyuzRfl2Fm3wD
ras/eMmn7q+d8YqYy9hDTDrW76FMQNlFZO9mLPdvGg+aYMLtnRABja7lxyOL6IAf0tRlyjTnotZB
+G4p+P6dM0OOBaRYMChwd8aMQjUD1NaN7DR+y3AvRF0tPMlbC1dbhNGMxGsgM+dTjRhSmqsnL9Ea
g3wjMibvX9z/K3/phSww84NUsnVm7Yoq0hqL3Vzd1HAgBmOzr+BBRcRUw5KPZbMAtENZoAzlA4eU
ZdXo5Cas9PEA/bW77i07y7LNY1tP5DreUnzr77XMqbQnEDh1rbQtsOkn9vtHkCOwYC0PrOgpFzOg
eG6kdrw3DJA3k5tgEEXD+OPig2PLg9GdpIWC4G1xoFWgG8V+E9ArahCfCPS1AmqzaVJIrCLYuXVg
9vmwBrO6zYxtvAISwNAD14+ZcUc1rVP3I2bDoTPG2r57p89qUHNVkmzGFP0C9VY2GdNek8Q0XoRG
tsXUcxJe7AOs577JasnwN2hjtVPWxP3yTQJeEKcaZJ/Dztb3iND3b199ddsMyz8pIRTOyGfthjln
mW7i/ngastMMzzlzbpJZ+5YH+n16FOh/d5rFvaLYpmD8dcit8SviBZrfeFL20qUHrOLsUYenPLeJ
RvFpTSyTrXZXcm5I/qVr7Ks09vMhHKPWZkQA9JVTYc8PkIc1t6l7QWyrZKpyGKdxP0kw+SIP1ZPA
zUWzAKnDXiUg7jq4jLlgRDBtfRy9aM5Ee1tkWGyI07vyZZnzfq2sEYCYdeIxfaAGFz38ie9aH/eH
zotyiQ8x5m1fs0Rj759tdz5TyrXeRBVru8t7V2fRCf/hF+dk4By/0+mOfONvev3KUmwqApUCCq+B
wnX1OR1vkEdXtNfhELqtUppdg1Gs6Yi5I5glLIg6m/lSD/m4Zpb77dKf3ix90cReTlLvmtJ0LskI
2RWP5moeiboeIMT8zBN4VD4NvOJ5KDbeX88LOrXQDauLwUh0PSGCNEVHyCcKukT8cCzPOK63J2ME
mNkidTJHDSgqu/UOEb5gEu6azAtfroBBijfWlr/gZryqJ1maE4OD1LitizJsNYYCi7ZH8MGUe9NC
buPTPDiR8tJF2eOcQnEJKmfBOoEF1pLZ+SAQ1XSKX8age++HRycT4nBfNCkWv6n82eVhWr/NECzC
nnX3wGNdkj5TTe3x2/I08kHR2Dqe93RBI3aGApMlJ+hfQaOMi8B+1bI9X17QtOQPKx1BjcSdcWW7
BChNSvimUQAdngvaCEjrziLNu1E4w1yTG0s7IZxOR+6vRtmxatbMxpjD+tuhVNk9FNVO08jLumk8
fIPUWrBCIigZR+WaIotEKo4h744zKJjVf1JKd9Ifdo2AQZsDJ84Oz7TstQludzDPCeGf+wGk968h
aSlwbRIY4o3k+UOFQchQgMMkiz/j/RvucOuHYoO8u72aYJsFRP6ftqmUkS4sDsZLagU8wBVyrWV5
0fwYh3f3wJreTRxXWYvjWTdGcXaktfdz4p6B+ZPVX3SqTn58/vXLX6Vkb7075QblXHzCbYyVk/9h
S+LHJ82+Bq3cdLHJkw3qhlooIg1FHlMuwCuzMijk5OiurqrwDUbwfvjLLjP2wK9hMwE57d+RdW+0
RanHnrxnvig8uKIOVH+pN+2elkwCXPPZcmTcRE0H+Px8/HuopWOauz5cVj7LtnKSp2j2g+LcszPV
YOhUqj9CB1ufJ3FIudXLkbSim9h917ELQXgfB2JNeTUL8xDI6iWyJYVANJiQD9sJdUVYvf2j8Ctb
4WVydflFrEJ8u1IFoxVWf+gwTdHm78394wJgjZNBP8bbYXE7c6iYVFRclhcg738/9Z8fXEGzsHIc
uSIWNEuLO3dnGKkjHgfypT0prRX7K4785yXhYGnTPSbaFGM7PuENIDjErijNWmr2FkeZhgdlF4ir
p77n7cOo+l1tDxidfew4UIbQ9UzOZzIljQH4YwvQPMGatzxySlO49vBB43MVfngUxzKqNzlx/Z6I
vWdMlqXQdmFzhjj52912rTzxuvNK6G1Re8wfNubLNn+E9aQoCX77zEgV46k5G704ylweeQXcApO6
QdYJcol55GdwNqnrOZ+q3Lg565GkGENyVId0sh1JphxgY6Y7v+5vErbo1nSnqm5eHgUsLuAcmYM/
6jGimQLzmj7I4QhlyuoD9T77DBpsIM2Znoodk0knIbF2O4PB6BlQcMo/OJxRyVoArYiHdwk8As8A
u0j4OOxBn///UZvxmnHedhNeGFlNSBuIu+NofFMtqDCYXJCkkhFZGxdTFR64lPn9ByPQFDJ0QwX4
bUAgFRAjvN2VeMJlJ8TojXM8AQoK6JyPsKkZb3hkhLcHwOQJU4Ynz7g5LjK+gdoVweFR9sKe5Nbo
pZfTojKqpy0FXv0e6+VIGVh54We9V0gFr20DErDT1lg1nG/z1jSiHz92tr6VW8PmYpJUtdG+G5fs
+8ftob58TTo01qxuFyDzM8iNsciSlMUP3U2DsIn1bri96lymuD5xPL34Ac+Ct4+zkqECdk0lCD8T
ifCcPvX+XpJsKSQlcq0kBsaFJD43z37GSQgrJoHmVRJSd7wW8/cOpxSscZJQhHrufOwoQ3Re587t
30dn8HUn96MGWPj9feHERp5DbWCCFgU+LvpzAPRAuYCK6QyMMCyLeSGpiuQDtcP1Fv+8tTbi6F5F
kbxqi72QwNZsgdDcLmuZHXhWsRhoQpB0Ytrtg67QwJ32cF3cGL1SbC7C8rRqKVOhSIpA2Gjid5JJ
0PwTn8+Iluckbj47oYSFy+Q6HmnmG3LX7Z891h2KutJmZfgKpLEOVdgESi0xrSu8OM9G42Uxid2L
WQfMNRyR/V3eX/x0d6S/yeMNdaVjeCkzdY0WBSfgvkmrIBzF3X7rPoEfHkTcFlhgCXDOgP3aBymr
f7vsM/uWRBSToniUVSv7QogBQOVqbZ9gfdYFVrQevpUfvm85VdL4BtrIXQ9iDn+8Eq6lmKu9DtW6
GU5zqO2TDf3uQN1e1vfI8pkIgTOd3B2cbj960Ng/b7ax4gSHjg4d7Suuz4oaMQa8RvOY7ReuN74R
zarRx3NNoOI1ptlPEHu1GOg+TNleLTExLv0GLfDBjqzteicpbLzdT3wds9vsWp09NkxD2qbdxzcd
YijQ9BuWe0eA2+hw8jjEEdi/fNUV1eR2HpQ12SOm5DX6mZY9S5vFcWasqCP/UW9bQRs6o/SehBtA
zOSREUE9y2Y1uiNVS66XIZUwUB7nkVMTJ2U8Ajz7GO5eiulNWRdXkGZlOcuVU99LA4yFkjo2EfiV
hW2T6mC5hOhnJ/Jyz8a3ANQ0+nSU/xzzkK1wjH+UUJWPfcqwQewM0CyanuI2hBx1AB3ei8AsGvfV
csctMY3O4K8j+PfvFuWwqQ/DfcQTUNllARfY1Px3s87x30wFR8l44DsGLMMPkAJlyKAGv/14qc7j
bzv2FYR4yCLxHmeFTN+/r4aWY3uriAjgFH7H0H0Eq0vflNR5qe88h4iYXDcJpIYSFttMPY/+S0ev
jJHff57XfEd96zCFr7OvQeDGVcfdWB9vnqhf3YFafHqP6CzK32ujda3Rly4Bj9S/uOQQs5R1+KRE
Y/0rH1dzG+VMPGnbQlQnME1fRcShPx/5Yp0apDUnAqYqaDoqyoXM5f7CMboSqg6j5Ccy5TFR4CwD
cYz8GtWWnCnxFqIPW2WIHFGLODgvjdxTYIN/4//HNY6Nz2Mpr+jkx4DHnFFGEXZBCNAKfGPDnGN5
NJuLZYgKtQeNV/FHaDaXFRsdgauD/4IKrsPQO9f01QdiDjW6g/JEfS//bvt+vU7BeL4BD/5poVUP
oAhl/w1HiywFVnGYtdbVGqU3QunxHruvnUFdFPtbsfgNdYuEh9s7TzFtkjF1mdGNDl4Kv0ap+NQ1
zNX0Vn752gW4oV/gnt8KnV71i8heqoP4edkGP7heXhnHgaZMYbvJQEd+nPTs4TWzbl8K5a3ws7IV
9hnb7wlUmT/tHx6uNMU5ULqs/Z97BA+JDzEyai5acOQzpUz1qculnJsByX7KaaVk0jE8sT8pqH05
+Y6Ek60DbvAvu4DJvJl6q+WdVU2kxAT7Tnm1Xbd7FK/0EVUcywbaCTHUD8wn8tkaGqdsOuEUUPQj
tzC/loqbq86+lmjeEptBbxzzv9jNIxiT7zSzVIvh0vW0821iHikzuXeRJ7pAmPDc5sUR9o39ZD71
GpYXC0NRHktrw/VGxJwlPFNTV7CaWBOQsCC/4vqKyg+szVZG9yJe57uXK4DE2DKG+dEYBmBCg9Dt
fT+kV3ViJlFkoO//zT7JVGCdUAmIGq0QiyptRDLLRigFz0oQ82SCa1P76HS4x9wPvoEy5g1n46gi
6xxutEXPIDmf4YcwRB1bbjLyoKIW/x0sFLFFy6HaX6GoyhUmTBzplgRIc/G74agiCDSqNJGD0vaq
DTVZqo0qqRSJB8H8GJOzjA07368FfuWoVY1KqqtW0d9MOyXOGImuqwAYpd+bxsF57ju18YcHhznT
nPk2EUOvfMMHQ/L6MhKW6rqC49zOaBR5SIaDzWwXq8PgMrjIHmEAdusQNNFWBiYpvD5HOX7vWi7K
mPs4E7o0bNZ+HPlWkpkWrbnMmdlduJWDFtGWWFkSz/BFJeXOS2bVQzPvweg2c+wp7Fe+zGC1psFC
j5DsLR6tztSGjvq2VL5UenO2ZIo8mZxmygjI9pLRyl4HDer7FxecOpiGsHi3VdzQmkVrPLnq8WI+
n3oxc2i8TkXovVYGKTjwuIOtKNSxZs0mmpnZL1I+l1TRWZn8boc16kJYE8LVx3BsOQDagOHxH4W9
qc+0kmc6iCOzovvmoiyOTKSBNG/pc9MzxiFG1mNVB4VJ+l1is6wTXjeJUaVM+QmjM1ivMeJ8qKqk
VBqvoCcRrUHoHxz+HEFnEtSrmZHay/Vr2TTANJCum0J/SVjFLP/f2f18K7VKQIs51GeHuJHVzYEl
IgFJYY64OnVieVSI13BchVzLlws1iX7nam3S2RHcK+GJGDZKVNdnBQ+LgyUxa7AyfFBM1P3HW7FI
kgofLX+lrvyMoL5PdIvHsbvc6M9S52MppYUMpqEodRxNPc7ou5hjH8U4kW7MnVlipE1sSiwbw7wm
xb3aEZraEmURO7Td5qHo2SMg4mF40lE52rUUubS3rKwb9CPNHuBVNDSTdDjDDQs6eREXE84Xgmmn
AaeraVYH8/q2fT3UcXfi0cRYFuJk9mriOqUHX6NPTsnBJ4/MyXXAb8u0QXLPyzABU2Vt0DZ4Tma9
nfGH/nqhSekveoD+bJswF7DMgGn7/TEHOUvgOF4p+JjjMU2+aQ9KZRA56Go7WArgsPYqWYwgMP2L
nTi5BGKOOnb0h4fB3DWWMBY5wslDM3iol/Zt+19a1Ii7QJ2SA8SbV+ZYs9gNrcvjof1fYJ71ix4u
yrGHxlKmaqEmvs0HRdGjfMVzxWqWzOCYmMqklPc3yE0Yc1tx74ULFY1La0ovZFYvk77n+GDSbHs4
V3yMUWXSs5NEHOiVM/gcvLtaUd0B2SA4DqCQ4RaW57VUAPwXJQgU42XQEvI/1n3txQ2b4SVoatay
HCzvU0hfy1OykJfqPRUsp89263Iuj5WEKxDPBDL/Cr5hQg2sXPdXksiHiFXv0svrBQe371uqkJlZ
3du1Wg6QQNrOuSXV8aC/3Bs8W0OBi21KGxpxPWoFF9dlco4nWKv+UZ6dxaQp0yM/LzjBTvJhDePA
pRNm0TE0rwsmSBR4Pd4jDShrtuA/xuYCOTFd1+g3SFFdqyEhBeZvKSq07QZ8AIq3KxSmbKG//EJj
6azBB7GWbRHG0mV5vDsNaQcpSS2wkM7/N7yJFfGOUYhTvur1SfijO4tN1GNKbQmyxXZapiBpGs96
/e19t81r0y2fk1Achvx6VwAYhBDTbn4LfMijQOdCdf2stsmMyBv0T2oxlUf8LlbYkVyoDmNz7bXK
TApL6W8ZX7PK/Oy2oaUPey2SbHyA1dTTyb0auc78VXvO5cy4EN2BNcepVXhW/1D4+FYVTlo8jiHv
4czJQiFdGFqlJTUAYcXYNO0ddpnsx0gKfgkJoD4CONcUGDq2trh6X6ahInszW2QupDc53g4LN11J
J2ct1UHEWQ9q4S1leEmd2YFePCgd9rJk5gydCnzOJBxIQ+SbvaEkgzFSQyAmGkuBzIZtEMqU7bKL
RRlqk81Qpw8t3jrfe4zfFIrDpNSG2uKxa8zeFhvr0rJv3C6ls1oXHTxASrykwqstIWAq+CNhXqrN
Lh9AqXXIfL4AxE0Ac7AVveCLI0rotP/TdAVb7iHYryzJwvCXWcmrdN150pIj6s3UEg1OpNkv/5dk
lq4SJpkAtWo61xxSVaubaSnAa8KQdHt8MCV/LOWNW1gparCE7vYvJNmuN2UaIKym5oG0phb3sNA2
8M/grGykieDUCzXC2OCCCW1Jiu2O8ulrg+TqzPqEQrUVaioofOuxcM2TVmT3dfYGw/J3QYhG4G/M
VCcUqZeXGN2dJ//aWRzgXwp3eigQiBl1wew3qsms1jttF8h1Qy+zdv6So5sWLciqlWrEqUA778xF
yN5uttCmb2phoik/+c0biLEUYHDT4wraE+7E/P+h3kduXulJK3B2dUpv2HLxB4SgbjIFJ+QTyoCF
qHY70lmH/9pcK49t1cRKFhhshJAHfndP1jYNqst1Crp8FDkFYFg99PDG7nNwGKOzzryYmdDAZmHk
ne8EJB2+aJC2/kZBnEaw0Uvxr4h0ABp2qH0oKCiFJUdGCa4DuphWCLn2BnA6FzTgb76dZBPhPJlh
Tv7691CsfcMpzbs4qPBhWJiYXqmIalykAAsphoS0hd0lSEKIV+6jCySH7VI2P7dyxan+3Ai/Ub+l
//1NFBk6z8a0K3LmotIY0ykVzLw+4Dz1smne3wpboD9fRdGbTFoeJZCdJbnol26ArlJRiuPrmJvE
VHNpqE7z9tn7Kew2eHhQkelPZ4fQ4hXDvrYRwsbQZpwDpM9TxIFxd5I28sLQGpRHkZRZZvNov9v3
gKczBp1nKq+zcwWFAbCE72lotBhCceY+N2YbBWIx1UOWJx5jvnbQfxf7rTGcr2Ky/S6L8jGXkA4G
QIsn7BdKsZe/w6fpLPOWEYFGpmx9ucnqkHwnk/AO+tBL0JPZzFEwQ9sGqcHULM1niTbeuDlK2/s4
6TkhV+pk3uiNmKQz/DmtF3s7j1D8OgG44i25P5z80+1VmnrksCLb1YxkXb/ncUUt0u4tAqFLsr0s
LPSr7WUDpUOc0WJ8Pfreq03MTPZQ4JNciFgl2yayA9swKVJ55D2fRgNZtWdQ2b/mOTrzT4drn2tc
q+GjF5LlVH/5ivkQ3IvqtdwmuTx0lG6CijPD6rflRuyzlOAa/gbcAvzDFRFAycwzyYqLt9m6gP6C
K35+Ua9ZTJThqH9WmV8kYkop1MYZAw73EDquDn788YYCkwNyKosvrvmHLJOGME4rPbGRppAy7Gh6
ahqDm62CgpLuFRCxVpES1Z5zcehMv+W0Wfs+jheJLweQulXjBAqCNRCeJRmZ8sIn26hgAem9bnuW
EkuUxMDlUNQfOXHLBz03UjglV9N7cHGe+C8vgRFDO/dhxpiuIBtfMaqSAWPu9e8JjQ/fw42EAPWL
VsN52pN1NPt3Clp3tGJigPvEqXfNgOOlQM85eVaRnbmYOK5kO4eHURMYwbOYuE7pd6f4lwXKRpGg
WN7Cyf5KZFJDQ+NQxyaOKNalPYWAfTWEaYa29kQp9KB/3jldeuL+EEQfZtGPpFzN/Cua9zaD+B6b
yf6m0+vaiiqbWTs1EZu4RbdEWQ9jEOPHh7gTQIkfYRVjgfOp84o55+h6+GpFJpj5Xf+DC1omgfeF
QDrhTdpQr6CG1QkHW8Vypaw9JNLApbpocWMujxb/iINWmlY17RSTeDsW0oENfSyiJEH6fMu8Or7A
pz3ju0Wamqe8nNJVNzHUU0Irp3M9dF1P2iPdGYcvukfoCEjwB4zHMO4xBlBKq0BIuP/dyiKPGzpO
lR9Q96Msvv5DXvvVmQLpKqKf5l4i/Zp8yIsXzsaxxktTaOfiF3mRdzyErD8gDLNWxfjup+pq45Rq
ixLsafqhl7Dhx5AQOwbj+17zDT8crwbcambxTaqWXPoKrOo47PMmMS1nQosL9ZPHYnKo39ymP070
EGJMElzWJZRhVUK0hRmN+ue3/8x72MMuA0GzJOLaEIhcJZ6Iz1yNC1gl5k0jZaTVegJ+0J1rvlq2
hlDEc6z2TumQmkHEuDXof110V3OTPHoPt+xc/UeVbkTpmXtWcYZdBGe8R6X8DfuZMzWfiVmCSrvr
0vu5M1CkczFv1fEPMUX+avEh0Sl4IDXTomCbWqhJDvhrlBZd4nUxBGrhnvAuElhOxV6bWnjQJoTS
E681yQK2Gage0N3JuQWBay+f5Pt0CPHU7ZXmQwe2h5hBAtWKB55c5eFkR7Qx6tU96VZ1fNqGY4yp
dgcptHdkKLMOcd34QeOnN9nRGlAculpy64TRU/pmJqcojxfjqOYVJ2iu+Ge6+u+kATo3vg+AwNAv
yl0vTqpScEI482kLDPsU7ocaYtFOhaZZoxGdjgfuQ4iL9RtEgJUjzGShLZ4q0NmtrblToNuxeJrf
3GKsQqFvEB3HPNO6iKC4/xQ4TCETMNh9INwOAKDiTY0Lj6D4YHHhg2dXqQ6jwwidnDze8+ZaqLk7
GWtgClSE0s/fg6iG9CJNcfF13OSHDwT9k/sHTIsYs2CnJAcYgnfnqeJg0NUzr2ThNdmrWi8F0RIx
tsSX6faT4zwwJ0+rBh2yt79AIhBtsyzG+KzamCAmUUT61KnaHHJKomh4zDf/bRNiK+zG3PZnfu4y
dy2FsX9+c+PAIcie1id6Gt9yAC/12QHk1mnBLlRBmIfQeIyleba8fVBTE5PNm5NcdS6xmzqIGLrY
k+QmqJIbjRLS+08hbPUErnFh68rA/iryuALRC4Smzkt2AzhCZDDIKfO8GzOyb6YqhRHDtp3+yEa/
uyC4icQjDxRtvYsKJztLWv11yr8MVwUtTGz7erhePlgrjFu46IZvuVTXIMYxMKKof8FlZudvlnFP
qm08PZZ/bnyE4vZMveon22RmkBGaJcnl7FACRssQFOmw2l08L2LbT2Wm5igEDs+ykCGZ0HPHQfqc
ZlV1mqfpMIWRxnoL0rU5a8gOCROJCGqSTU2wteVeTfi0hgIKDRPchxgIPrlCkHgbuS0HmWHIDVck
be5+KRnDrokuKNZ/fiigFfCvBO5aFAJzv28SnDuOlJPMsjLVXTr4OR1AD99SN/YxU/i8dno17ify
I32BW5qVeCFYPwRWSpQKm0ZSedQyUZvBplhcarTGmWNwlYmPGZLQcmc9BeyIxXdvN/H+BS+yhWPW
mRkPz7uCFGYymtXcWbo8RD4744t31tu76wF8d3HxGd5as3v2a8migRPsNKNrZR1R6CWs+SXJhFSS
pJvvoMQDer55qS5AHJR9R/SwPNuTtFofXJ8h31bB3msOWMOgpZqOnfgmSCs+nxJl5Clnkj9OJroL
2Kwf/PfTsBn1uGVuUGg2lJCcnBdXNBlycJbeB18fI3KRmzVB6m3T6IZChyysByhf/O+UZ7Hrc7uW
rKez9B8UDUH/DICKdD8qsubSa9Rg+sXsuosqlugIOyFAcHFQQ+tKw3MzrJoQKJe0DjXtBfqvbkHq
61bDMmoIex5UNp3VLk5BL0yWM9VGgKKkRWA/Fa00MqSYH9dwExg7dvLlrV8VOz0h90iCPzlxVRgu
qxMW+BLX+u+dzovkq766APiUxo1qkpoMsvxaS8l5dME2bfQBy21Wc9R8RbNtG4YFmINBvRAzzT9+
giJ7hM6DNyaWQbOvJrT116x7JHC5C/0+UDtrUJsmpj/tCwAVvI5/bhaIRJIOvTsg3Jiq4Egy4E0b
Eb4HzAHYXzlxQ5IkWLazsv+zzwT7vE3UyesrVDZxC4bGef/BwEPMy7IqrMCXTGSQqCaPkLPyADC6
X0f/KZPNzghr3Xhx6ar6kL7BAw0fHKs9Q+vWm01wXVeZhyYu+KZVZlq4aCBB5TtA6P0AQOEUBWGD
rNiIAldYbsbe0QRvXEiE8hxcRW/QTiusDKh28Jldhnu1wGILDFae4FnAIM4XIS/iakeIRXSaXiY/
we0E3s6DRem8DDmRsNOfn+oxM/5Uwy67Rjdg9iYmEM4wL14wBAnqTPCKhpqa/hrIx3MNCqleTvzG
ssbfWoIx8+BjWn5FjTSlxCNBUQaYb1RA1Q4WQmMaEXniettRnVaxmdLjzZn5CTEmPJhG9IwrEVZy
UdgxvxWUl4AVpons42vekJqA5kZ3+bh+UYTtoWl1mNSz4aD4Bydfb6AIpNv3WkO5HBmYGVJDxfx5
x3JNTXtrXrFRqBq8kTRwbAwJPCjB6RgGohZ3GBRgDA2cNCvMzM49xRmW+D4qijlrT6H+JBwDEPWg
IxDr8WKq8wMPbvB2x1ziCDKBcXqQhY6ZZpbqdfyWq3L6ORfX86Zs/oWH/koCBJyxRfLkajBIzly1
SlQ/8Lr65wT7tiHFVp3ef2zUiTeYieFg1joB9hSOvOgRNsKPam4nTRsEcuHqxZU49d+iSKwKaSsc
M0gVQw3+PqEZXtLgeUPaOt6B7mTA+airBvHAfxs352jahxBAxf1DMmSH/7MpGoEIFW5NPzwVJKUb
dZJOa1nJbLCAz9Mkp1TaA1O4lXYCfh6vbn4o85ICjvgtxHmAEUQ5NzDsdyZii1yRliT4pMf6g6qQ
zdqucShUB/oYwU36kbDps5IiIWa81tUO1Df2o3k8ua7YGwR6mBDCu2RZD+tTGU5LmFigO9pOkdAt
Rh8xqKVKmWb7iB36svnRL1QZW9OhFJl8/DCLoknNIX+2MzK5EVtLWj3SnxRCM4Vmj8jnP+jUNT/6
cNUoOR2d+RJpHtqTeoIKVt/pN6iEpZZ9v8zdPZ9jIcYS7suTyyN2xE6nS7pmOoS6SWJoXHFZ3h5n
nVNxTifxdIgnSkYZea0I8JrlNkF58pdmzyx9Lf0F40bWItyudpjGFDRs73SwGsILNhOFwWyFxWra
DS2TWkFvjnqLEQvbmbxOJIiDNlmwVZyIpPrLkDPS2H8+cBasNrCHqXOTQ0Fuzj9QbTRaXmfBnYdG
zkhFmxLC9dn+AG+GfjbWRfwrDHJtJzoCPxBG/Ii+6yBm/Erka8aEAiIQReWdvGECSEQ57tR4x38m
EfAPcrA4XQL3hkMs1Mn8ZCuQ+axYE+H6nbuStiFmum7VXeMr0DMEcAZbogNkNLEv/IGtkbPAE8K+
UQpmFRmGOLdSpzJvkxg0wAYVzXPBDg0AUfjkB2kiZadh+1ZM+9l0zpEz29xxjc9Ize7zd4wkcF8w
IWo9rs4HnAe4KwEXW+miJtXDxTJ8EWpUWSOw5Hnk/SvjIJRhDKusMadksjtkq3alGntuJnuWTmES
aDjcsd1nSkDS1488TCDGGbikCM0ciUyDDRMnc86EvhluX2oIgFnAByJZE5cMjp6IlpLhNJ77tVv4
ERvs8K24q7ixvePU1Jvvrm2kwDUObAuqhZ7fs/joeQlz4nxUM89ZkbGcjfjVZm5S6RYY4rXRwE0o
hQPs84LqNNqC9DHOZgQzrHeRt+ZKFKpiKBOeDOJyBkRcl1xTDUhPOkAVEX7l8+4RA8VWYx3chU8M
Jv2sHxCxbHXYvhP5jlMN5btpwklblkwwc9jHJnQWSC9vK+wqIHflPAe1jONO3YCDHDdXFPes8GkQ
3helPHaBLgEXwcOJoc8IomfzUE9Mm3niznmaoH1Wqv5YY4ZIYoYdJSM5GiBgSv7tu/5VGBNpVj9k
1HEUYZputPLscUthIRO7LSdSJre2cgB92O/p3wb8cwipQVb4CROouZtRs69LrIlcVzeHFR3OGZrl
gAc9HHHNpYYpu0KzXFY3HrUd+JO5thtD84CCt5Wfd+kWVbqESBo7Sw2iGdhLR/RGX9YCt8FZ45d9
ErWRUf217QRJDRvtnI8Ookmk2Zf6oA2cjlPZdnei2xzJ+4q7jWm9Z42GOzERAIHdOTy3cauONIdA
kE/Zd8NJESDNibVg7iTRpELwcGeiCfU6YUDLoVEc3Hy1zASIGbdYietPpyL5fA5eAtCZOlQyMy24
0hORcG/bIpgp54iyG+oBvyRXLRAJtKPUwYT85cqPIZXYuKjtYAUAJEqZKr0IV9TSMPKGrZKEtsmy
opuW5y3N2C1wTQ2fjqcUt1UEyJTCcJDRREiud2oBdqP/dkG6ivHn8h1Zkc/RmY18wsjpZYZd7cM0
uuoE5r8W0U0zQr6jcHUQ33KFch9MObf02HULEqp9xQc0M3LzQQX5eU3vjS5aLUBr70pfdfLqScai
1z614WDMwRPMb/vEccwwqYC9igx77lAkM1Knt+GMObD/8ergk9RK8qhCDXmC8J7CMLEAbl4T4fH/
eWzJ37dO3u5FMRO3GgaFv+GsjFBtGX2pLs75pNK0dDD8dLiKlp9IFMCoITSxaMmGLMa4aHB1bDI5
KCUKTysVpywdNP9Sgkiz0/ifq+aS9ayR86XydNVVrcMtMrWU4dBLq5lbb6qYxr4LXPcO+BLc5pQ4
Zwaq9boZXYH5NReL8pSv1L+1k6EhqUD+r/RsEV0IiRrEITf+oU/920QkqwgLGg4HrnN4yUYGLj1K
Cjc/qFeinjkluYm4YAaPZALarpxodL7GQyn3hT5UwOaqVHe4Lj6ZotuKxJOKrljOxI04ET225YNR
15+mDjX50C+nMPNQyl/E+/GeOzIhv1zW05bKV0skY2S5O9nRvTr9ctOEY5eeAGHXVnbYsQFSCxkv
P7wBXrFXDhWjQJLXfQANuflJkSv7N6VFTVQCFMOUkTz/YsE8O8jyEoZwAwMnsLd7/3aJvxhL1ssh
Lix7SkCxHTKGocoqkLi9EZ7xtDlQj61nioh9HrZ8+u6UkoClQM2A2oKGHBMZzBGstsK3cfmM7JCc
GKLEkfGMEv1xEZAocdktcvxjJ/XFif7yBGD1hM6Z66ILC5X8ZZixdBBWaT+5VhYniu1EgqQA/2K0
b7Hvl7SSjNFGdptDYykpMnSWpkAh3LZo0LFyfF6wYR0S/g43I1QiNdCVgMMeBVPZRoiFZgDIEdLm
eDpw0tc5QgBWqiPz5vRugW0APeNxgHMAt9/1ohqsoVc31AN1AQe62k2Mz92hKzPvGX3WqmobDEJo
3KX44lMG+NzixESsyh7vTjlM2LHC2W2CkiuwNPYJYsDNLJiJ4zm9S7DoSw/DtxYIv6eHGGmat/N9
sglcjfZIviXnoxvTQdTt2y58IU3RlFc+0gm6IGllBWSW9YXI6ah8BjpjKS9cSFkUhLfWSgEkuc/K
mHFwTV493CHtqkm3RxvHDVwt17nEX8PbArk9IuL2WsMC6c04RL1YDJGGGvf+93epu6LoMJZiA9my
+R+GgqplvmqpNWiF91lWGMUGKo9x3KvXPOPgWLbIQxgukKM0uSrITIDyelS4yxk1A797KU9gO21Z
1oYjyvVZbxZWEz7N8Aq2hfErDhS2V4LEimsx+c8wJu0enWWcoIQh6nr7cp9HHlQZbLQAelvROm3L
XGTuobanrH4ygDPN/sZHbQM1q4CZsx2paWuhL1JSB0U9sSbUGXDhGLcd8xmAdYWFbrqysoKdPHtg
86FrstSIQj0j9U3O4ccbl3vMTttMxeE6YpvrUbgEgnKrAyYJRzYLXhoZEzrxzLm5HqMfKOQY03FW
ijuvHcf7AGga9CphpWdE6//n8ZeF4X6SPT69p0VKLYfpqOgOuNxtw965e9UGl0Iz1+AgJ5lGfJEb
xCIjZ/lTvOJL6YR8soa59/h02ydND5q+PrnigXDXtJeqG+zY/TVa+hNXgaHl1yx0evSaULTymPzR
99KoJXyoBOH1sUKvul95GQNq0/0Rc8uBT13VS4rwzojAyJTTe0B/JHs35jgICIUnrkfD32PrrkQP
q0p7tE0jn5ZI5Jb6gpx9d8wnbn2s+xneQmRvmHk9qDy8JirkUeKLNqYXO7vbILWp4QhRNA4xNztA
yBkCvIOabedGUsiQq9kM0Wbzx0+B8pZyslUOlXKQKqAhNfkDbY3EhCiYAw9vwG0Z5OLU0GlUR8ZB
kSZBBf1Ea474qwN1d2kAqtbRkxztOcRiClzibfUPrFLM3RZasgzip+IvbjvhTU2dIGGxQW/N2SRd
BisDBrZ6JrxNjZn/krkgsdIwnUfDhkGQ8WdJF4Q4pkpuSTkPcqmikan4u5E1WE3P2lCspZdg0msm
avZHhAyKVfN5OtWkV/8dbjw6fzUigFZ/7fqANkNqQIhV7zAnjikKcnoNmkqgA3PKKLWsdN/sbV25
hg6IP/uujRG9plCaHWXU6sqPSPlT7ajzaBa3XPEkPrZQRdS4Gf1BhkBfEQ6Bk35hyOkInpKvsFr7
NsIqtYztU1VUjD+NqzNIIfBmXKmUtpk1r6UDa+T9DG4haJpoKolOJ3GOHptDJDnfP1iWfyqHB8yJ
WoRrHJCc30gBjESZhvAu4vYHSjJR+TQj/XjGNVXw2DtFuL0UNBnH+6xAhSwoub3Z5UNGRIs5XtS4
QhPUdKX2TynbczRqDWTcAbBeeyDWQbJr6tRzvsTiyIB3P8lWvbzXyb79RFU+/CsfJFo4jH9TEr5j
c6IMqrPMW+LF7HtXc0tB6HtTBEQe6BDhAkG1b1TwGrCnMiL78/kpm2cFah046XDutibUl50lSWds
fiOswbOXZv4oWCTvpHDbRb+r3iickpZVslCznsyACeDOQL1hSc7/oDWcoYIh4LSYgAnP4PTVS1Iz
/QhyXp70GzklwIiwU1/CY7bPil9VpuqWVa6Y1ctpBnXZ7w7DN3ssOzufxj3QIX6aJvFB7THwp5HY
Jn5BXmPcqiZuRXyKnNML9QT9iIInGaCkI/L7f6TqQP5ev11SfqTNwlANm3a87YoYrHtrKTydE8qx
WiKqsFVmMPXpo9yhc5EChk/H4pIJUtoF/UuX4Q59YvzM6sV9L/VQhBuQjBqthWZIQ5/2nmT+PtqD
A+q0axVqe4gBqwKS++6jzHmYD7uUZKS43SVh9BgWo47yR/GFSYtKZtwnEkqdQO/eg/ifiE1xO6IS
K2qTMKeOL38SUnx2gqN5+faoK8vONgYOFjLvmDQy+71X/BF+Zvj8pBr7HleejVXnRDBmqcddi2DO
cKmUoGZz1N4REV990tZlQbtYfbucwoWakWD7F3l/y8UhAg5/0XEVMjsp5rSpKXRikRmVJBM7+Knc
iyyj5HjxRQt+TDGJXWc1q2ggy7m0cqzTo/nGDNL/gW48zK+xebAAUdz6Fnqs902Jw/QUGLZDOZno
7Egc5RtlWoFEyE4HOtECraSZTMOVYGhb8HJ3dmR7Ze/1zWgXK7RYZ+mEv+YyGyVLsTADfHUQ9PkK
iaSCpUj9eIsRnSqcui4VUuj6JRFIJclZ4laVDe3sj6z6R61SGXqiCYa2UW0Jgt9Spk8knV5uGzo8
AuEfTC1KPzapBvMhpJZ+kL+3Z5BDTwUO4RPY1fm6V/nR/IN1npclFJy2eTfajRcryOD8dbmwDmf4
eDOgDdEqmriB7rrLK44gEBAANLCyvSvtqipDwsjr7MZkosPIA3YRsL4+KESLUNZjyene/KofoZI5
FiWPTMjMT5l9HWVkUn7BDM++LmDipiAO+7O01qaOa82uwR6diPx8dzY9DQyw4Wyo/nf8L79PCaIu
hI1H0VYQ5klQPuZ6KiP6h360uPIQemCh6uEXa+mcJqNjjg6ebzSRIR9qLGmwly/TN0+6ql6ZzJGr
uz7LeNLmmSu+f0Z0SPWQvpuNl/uhcQnIfj1CtVM1G+hidUVWMjpOeXtlmuiyeHYTfbEtdR1Fp9Xm
BdtvjFxl95EFHCkC5B+3GJnh8B7YItVj2a1y78Z6GmGZ06jdDb52TiUdSDBfTcynItAihN0psibo
xu7NfgkErQgf9GL708dkHrA2olGmdPIO+yDhwzHunEdKd0M4k5FUtqXkAW8V9Nmi9wDrVO1lvRDK
JN7VQJOs/3nWpoC0wBCnPhHBATaSsLgREGAh+1rCXWXkRcPWL+XTYKBs/t+sJjdLda4qL/95siZF
3TISXDCjoqdyq/lrk8WkO0DjNxeFL8R1XteAFjmA+JuY5LmNzOf/kmlPBEHZ51Nx/WEO4Fvqorqn
0A35U/ujwiI6vIE4HoHxLN/Z5fbaMkbk1PV0MLtXJVkox4gI7Q/HhvjABEXaGP5y5kgk/yu2AAG2
gmIBeyojhTnkP77p7PsmF0qGf3AOcXUvCS6WjgetmbDmPv5Si6DRx270/qxiLd3WUF5EX64WcoT/
lEgZGNccJc8sO++uOnGRrwZn0WXoBMFc/a4mkCvXbQTebOlQpMMdIMJUNcwpZQxfoYSDcdM8MTUE
JHedXC3oXdSX+KvZfDH+wU5fr4y0MLlcHc+QvQXy12jhrHd+q9Hpfb5yEyvs66JW/CVpswf7xUuE
5GLq2Cphs+mqqq5pdPTqDDU8IduJFT7a8dDG+riHUkifqh4XZZVfQCOS+knqzC4emyk2QIPxOeKs
HJ1/D9ak6jcyu0EmCVfIAl9swtpC29KJQjRgPoGfBkcY+/6iTx6Fx/GHzCj6dTr2HI4OvClyMhU3
uJhjc92qgriPZAE5gsd+bAhRM7ivjcZgCiE5XRJEpN2M/zyY7MGiqQLh8UP6wRqx39gYeTJG1Q/q
4BJqVhSmAtOjPNnI2di+2R16diQBvvkF8Tby/OqzYrcM03bi6F+JNcy/lSxIsTWbaBXe/B+kyM9e
4ufQ7VJbrIMKZ/PRFnEn385Qwxzgkn9ehj0NI2Ce2HEJ+F3v62xbNBYm8SCi1PmbOP52qTj1dCFF
fLILQtg364O0HblLOHpaDGVAC6P/UE62aWafxNtPxs8ybebulvGJSm6KCKX/zXn3OQg6kukpMAsR
POFZX6Vh7tieHn7WQb1lJRKrKUOmimbH6rDJSYRI9xJBPreRwSiTjoQZRW1pGm4XDix/+B/f6yGl
Ee0ha3zqtcFBGmHGRzMFpA491nFhENBK4jXPNzpAC2tzaeHDtIrtFwwTxkLJi2Axr9lpaKvh7AWq
s/mPW9eysC4rcxo3RBCzyIIvN0LNsEXxj4vxEmI1mliPTlSj52xEEZygTdOAvc1O7mY7XPmyo6hP
+EVGWifVu015K0KheHMWR9jE9JhQT/f0ttb2qI9vfvttFf8SqkH6aGoPK2Qag4q23NTOac7CvFaw
QP+xNNLvUVVOoJfQ/PPCmCtYwInXr1PMIyL0x05hGAr8twCZlYmMgO2TTGsMSqNK6ypcLVUgOtE2
8isAneXF3Sg7fWsdyaSw4XMLSQ9CgVuOMyQQvbKoEJJulrWgbHncywWFZgIdNYhkhKxzSUuu1rf+
bIwPfOqVBhqLVV3IvLqxEl3FFLG5TGJTr8Y3Ah6DGclDVoPlgRhFHtxHluSRzli5ksd7mgsFt0uj
lg8jL1m3goDRKTuxMo+rExFRFGTMqbLiPcfemlXP34c5Wan6c43RFNKu7uROfCappoMk1Obf3nVq
byXt3tHeTkm1RxNO1FiUEJcgeCis6ZVqKhGWbX7zFMklvwgQUds11xS/ps+OYA89cxp2OnOOMB/D
STm1nSC5Abey7HcvDseJWTZ9ABH6Ub1KU55Adblvmk7CBO8nIoRir/H+Jb7apnp7PjR3p7BDrZaq
fTBBaO5c7cC9sIavsOE0isn7e6hFIUc844MJoDvITnA8zor2EhbcxLGXTkuim/+j477JEWSszcP9
8M4KaSZFWEBywlfn5Se1Y6Bjc8RILT7bF/C3+TbqTLpcjJm95N9WTPVkaeaOMvl1aUXUC1ptb2YK
hRiiOjlUvd15nt3RnBNCx3qkr4ki3IfIm9bzpNsXNVnuh4kXfGz5b9TFaziZdW8aJqEIuMnt4KIX
dN4u8Lh+Sg67XfxZPnCl8ukmhyxr4sutezxOUfP1WkVGV8gErPOHs2hwdYlwy6pfkBue4tvwHCCN
r6v7cSkw3KXhL225HdahLQM9ta/Js8pKyhIbJkK+q8zVtQX+jTbi6pNby9lx4u32jQDaIAsgJRH/
Rc2UuXI76Pzpm5eN0LVtb1QVYS+1i83wRbEWvaSqGKAh6RGIPU+fXq9S830P2nH9ynfgSKQfXVif
fIi5D40av9W2csXwYaaKiu2he5HY/niXtY4X/nJY0XELL/9ipox0hKcuHykJ7rERzA5cdtN6NZLO
MgYuu4X62u25/3ONhmG2w9m3EzuhzWZgeRVVVTaxWJrl1YSpO3+XFNZqOKY9jnu1bB7Rg9GrAL4a
8J2/gnjCyRmaoCtDdAnFHDH9kC0tv8GkyQ6ZbJ4GKBO0PdGnfrZJcrCzyR4C5AGdHzj9tCCZG/Yj
wOvUbzzLVwK6miSEf12otNWpRD31y+F9IM2EPSo8MfD4KeGle50Fyu8YNtNNKg128NgaWkl8Q1fz
I6s6yKAKmU4eMw11BsN66O1OjFk2lnze8ZI0PgrRhtBA8JaxjY+TP43s6gCy1zTZ/yXswY0BmHzk
4IZB3ajWBMj9g8BjD8ZM9JsIIv/eiYSe/+BIWbrt9pz8gux5Zj3PtWa8ZjHBYktD58G7nrsLscTA
6eqCsUbMYnPIP/QsUKCj261gBOiROeG+NKdv9mSf+TVGell93rkw4K8CDZqg5kglcjIU3iTdJ8v6
/nMEXE3+75ftzvD2nR8IKp7gZywa39WKVdby7G4PZ9OMy129U9xrJuU0jfhAw0Pf5ljSJcDE1OLY
G4+xRK//DNEDNpb7q+0XWUdPCfLysUWKQoXuNhqb4g+4lxdlCeiRAZvzn1kebuBeX9vxGtgRyQih
bU3drLf8CWKFds4/X51RJc/a1PLW4jPy4AKfGrM7V0FRD70rJcAsFprFEfEgnO7b69Y+hIoO/fef
xZ03UqnB5XaaTyJCdkKYiQoKuVsrWJduK7arBc5CNo1+AfKiST6wVC6NegFu5i2Rh65eNuNpmPPS
I62o0Bdo5mijUe6Q9WD5idVeuU+yU55Vhx8yVnXsCsawFrbDoJ3EPs1oRV5EbyLa92n/2ZRkSRmC
iDniyMvOsaYOaPYEVTTkkDGzEDJamcBl3F+YnKfiPeNP08/bSSVmkOeQsyhraEZw5rDOuxrc/SqC
2QkV7VX5qMGTXQ9mEouLKQ7O77TdJow4hdk0KPPqMrHYEz+KXVDELNpfHUbZMFTodUbIUiGINKn/
OyvUXFsJnboz43dKDavN+Ggu485aXrXmjeIpLyP4grg6s5v7lIGRmsndqbS5UNkn0jwclrtsdctk
hgXfQ8q1mdqVPQenxK4GD9XhetFuVVoluKdveadGWDRXURB39ptZgRfYQ3/T6vtVH/qtsBl+NRE1
7OTgLPW7AZ8qUUz6ViNNUt9hyBmKRTz6WOFwiChX5972Ul1v+3oZXZD5QlBoOPNJq9bADN5rB7DA
BQBp3ovaajX7JLXpoSYFn/oASWzPHevPV4fj2MYKwZS07u3Y5cBJJLZZWfqSLo2VHEWGK5o07nH/
aNK7WrEvP24ddKopgmUIk9s9sEeQMYoLQuOyZQUvnNC+8pzViSGzeZyRwqQ/kb6tDwOfy20F1gLS
CMKa9etTCqhHP38TIftWhSxQ7bqTslmXgFMmekCsOT69hyLPRJdSfAMlB5Tr6knZPUmJ2BUNc4Xm
pNsPEdfQTgVFbGJ8pw+gXL8FmTchviF6N8nc6sF3R9JEClH0Kscxov96trgxOLm9peXLte/FIScl
ioqBsUukW+xIt7gTPwtIQe/tcTNfKj+hhMPwTZMrERnoCc3RqLUUhr+X3yGchaTuRJdV4BA7wl9V
+EjEZpJPwqOOxfnH+vjVXa4MaNYh+LhE5N2lY8hgVFumE9sOuH1zGNhGnxLt/+F1K+j+zpGpjwmh
kaLYcrVOUWSo38ancGrr7OEuyWa26AA2IXfbRTwKvefIPy7Cgg2mWw1B5dULD7SiCL6CYMSNEH7K
8iD8SQLvkIPPoFnWa9NBV9pTEauAxGoWkXlPwW0coqUnO6lqnudSJVEA/wOSd9ThSJlJP8Af7S5m
EYUcgczy4QDDlPBJa4Uygel9/jkgsvf2Ge5t3pxe62HwZoBscEcKkUMGJAsrLqlScPen/pB5akdr
BEtU1zKzlwj83PtygJaj+hYjasX/UdcF/SO1NeHi6KPyrleL7pg8L4xBpxfoAPh4LDqOaaugjvEI
mAGMX4K+CThssTrNjTBFQIEbosLaSJ2bNfpYGtzO+7DZW7b1u93bPzBJ2Id77mC9w1vJXeAqFYVe
Bbfl4NGlK6Owa6TCcJgg5bC4WT97P0nssQyAVSBtZQ4ua41B76Km+EC/92igeYz6v4opOcM82bFg
x8+vGzoxZz/oUaOByj0FdGMUUUGcnfwYVkqPzypgZVncUpOcYgugP3G/XM1ybyXJEATsjoR9C9Yx
FMyi48iooqMb0eAoQddzRU926EX8YJgGdpEwQ3EYWXOIv1Q0/+GfsFWmIojR8iakFNGtl/MZOp5s
6hVWJgThJ65Fm06pMQbXhRp/e2WweS5mFA9JBu9VdoLoufPoyk2so+a1sMfHNqi3N7H7eeuqz2NQ
7ndjcHisw8SBKN+zLVDgBTzZDIQZ2nKv6lPs75d3IjapvY2zLaK2H8w9eCT04w2T5mNpAwRd+NuQ
lA8FhNuHcqVcLSLkOWDkg4p3eQdDraIgrL4Fv43WvkFUgpT/xJoEyNYmSXFvngi6E3xY7W92nhfK
9eoyIXa79VccCUL62ma7PLkJebVUYyXBvy0xQ0+u2F92VGCv99taIKmw8LXqE/5QZCZuPiwKpky1
WtdkOECc5bJc/qpeIMaGa64So9gIXKNK6roquQUlHejQRX7FCQxUx6+9BCEX0SGWDS1bgG2k0OLz
DzQs2DVbNuB5QRO9KvReXOQdPG89f0iGvjXm4TThbiMF5DcGeCYM60/UQ3wjhkfJkvoJZppFP9yJ
MyKiiF3ynUZODdHZpecnABN7bVIgiD1LxeDhvMONc8g+Tl0Vu1BV8Gwhg+vUfsrTrm4MSOXfzHvV
U0tadp7vSvfOtA8GAV8ZCJ7DbQ2dV1bgMPX4oxO2IupojZ04kWIMEeQ7568+wC/TKlLtccoEv1r+
X/qLGn7Df3+4FhFJ+Y0LThqEpjpQykrfgjw/8FtC3tkpliYRdrB8MwbdB0bzxTdx9U3rjeAr9z8b
xS+PKPHCHjxwXouTMVSa4IdpDtg87KqNTcOUTn4Hq2+dXpG9x+Nrt1si+qxm1vVlOG9/ldUQlHbF
3hZfbfyZq8fR9mnIDkHseguhaO6xxMYLuOW0e7nUU3u28LcXj6Litpu8Z5ZQQZtp4ykk6YA7YTvI
mJ9itVWmlTyFAr8bMvaT9ZOuchnFvkDiyX09IiXMGAQwqjlwqjLvI410oUHJ1uuEmKmr3nTpaHNY
o2aYf1vshbVSRzU1wfr2J6528vkwHgkMn3uIUnacJCz4geKq/bgdwnn28MoCSCkwj7kjyLPD/9Pw
OrVA/skvW5L7VwY2sTXKr3GpvA5p/Ex3M8BBYSGLMmkCVA6QIlJlG8P4Zm/ggNzJ8JtDO0ymveRu
VqZWU/6pJ+Sg928534hDLk2/04gb6TJ6zgCFkeFxIRl5tD+H6Scp9cN5G/eE+AfyYjUilI9Y2yi3
cmoWbRNVdAUos6hWFVvwYwxSdpmPqaIw5uqBo6b9lwe5hSoY4iE4PKFv1ECRpj7ocYtR0WrTfJ9r
sOFbj/pz9TWAr72XeqdfwgLBLk9pwMW64thrYxedGxKjARZIm30dxpQ9fDt/WUasphXXIi8vGrN0
vGTY6kw3qoyimbw8zvv8i9eaCb8pfGTDue9nzmBzsaUZdqTPQDo+OohQYH3DEoMKhhJozAS9u6z6
76mjyLqD+ymmt37vPu56Fvyn3PTsSCWmxTbkC6fRxc2mfG7EzQ3J9sS9BApD5+2Rxq++Cwe8xiJZ
YxayOYo68nhCRphYwNNxkcXPsEMKJkvC8JnsgwpdpJpARJHiFotD/a4K+Qx183siFOhWUrCjUkDS
PcDPVhJooP+4ceovsKFtnKHrDPrNko6TUFNY6xQ9PvFTJH7XhKlUs+f9bk5sJVnc9ShTRzc7Gpw1
xvpslyYtMoIyeOtrNUi31oV029FbX7M/T+QdouecPVMmoBfwXUTXS1qv0QwjMpvz4iDCEEBq5l01
BNUBCcdzS5IsTExZN9Wpds6Z/nOwNDDqWLSyqJH216VGAty6YfSs/uVCIkERwEOulP2iKHtJqRqs
nRded1H0H/26A2G9KYOPCjZMYhIvh5BZVrfTM1zuiRmOyM7OW4kez0ygxr5l3xvUp4Tm0HfSaW+P
BdtC+1M7IS5OaIDD9P6CMOec/xkMUnueg2nXrPaQVTgwI/5DRX82mZV+LuI8tciwC5t6M6aNIRBV
zklXZRrEJ4bcKy2FhLzCXb3RZMbt9oPUS7ObJLtdMRypsva4vur4NgJg9qgM97ohL7pFRvWnHpIC
IjWzTn1qPnoY5DAJTEsAnPgIM/d06OxyhddtXSDSHZP0YohB8M01KaRdG+l41VsDk7Un2/MJhm7T
SgdDRM7gU7nYyfNEssPcDBDem6vvLmYciAhbzUOiNJqBOU1ZURpznaLBm/xRgzNd7hmJR9xqXZNd
N/3wRjbb6e8uDf5rqrzTP1eJFecUlIdX1GjncFBaT3wowy0snfcfRxg3q5xHmJMwqpIZ6/Y9zNVu
qOjAEPGYzeHofzya0ZoTzF5xxLzRZmuxSUJKj8OhN8gqCfFlrR4PSB5cfUCX7yfYkzBxj+doTbvA
fO3EGsO1HB6AQ+5vzObsfqbThxgKgDaqmjDV9G3rEouiDlLxc/5o1vRHs6XpcHwPkZdUJZwcXILh
X0V+wep7xvtOvJkIazLWf+K6Illjr7+bZA1cqckbYvYWC2Q7YAS+RI+2cA9Qtu7YWiXk55K6XJSp
hNysm3WsJmFjWP0YobAjct2JpbvmoYCLC1V5Ype1Uwf2O+EZ+/v7Vf3lFHOBw7ogjIHBnroIQaOH
dUwkt4TchXyDix7q0eoMIEAH/7Dbe+tkxxB5JWfu1wxCHjcPLZoRf1hU3IRH6utPBVKy6XfK0JIE
ruMHcuSZAeZnFbl7RC06eKzfoD5Ffes0V4gTq/svnk7KjeinWxfD48t19Q84Qqj4SxAd4NzrDv8A
S6r8q+PgsrYfOZFc1Bppj463FCsahRDP1EUq3qaNMkWquy94aGD8pTOxzadCd8IvY8Wp/FzCzxwP
TeDOdAYYzOP1tR5hAckpA5pW1oJvo1lXF6Sa+rwC1NuIKuAr+4OexY/XiupcxGDSYoQPG3YAWxBJ
j/1kfIouMthvNx37KV2pOLdqLNN46jX6M8o/3k6Isc4U3+bSLvZP3BEyvTnHMmUSWhanZH6ISwMd
suhcG97xYKs/+NEx/+DjLgO6whjPk6jwqh+sUyhVI37QbifIlEXHxdtdZddoGWKTJK4dtsOL+RHi
kk5iwdf97eOBlyTpALJEeRGObRYbYUpzx8KpD5ZBK7a8me9K0P7zjM6OPJ2IClDasiTlhxsqC2aM
TAdOBfqwjyJxVC8XlzEEkDDu4LuZsVKgFLJvMWY7NLGKz0Mk/UMK325OqDWWoj7iPXuV+vw/rWjT
cPTcyzG95JiPQToFrib6uo3465Fygtu1QBzHvMGQxhZIMPArzYEK2F6TB2ZOTdzEB2lsYiD1i+pV
UZjjzfAFN41m1f6wtdPPwikuzwzwYcetURAixOWnmlX9SLrmuGh46OlWAkpkKJS8tat65pSywyA+
xi+YxL1E2guVXAmISGNL9/whhXmJv1Lm577gzLPn93pA13clGbAB1fzIcsR2G3kAFDP0ugQFPaIA
6JngSFZiq+PMmJ0bQrgjYegX3cZN852wXCvOEYhk/asnm3AJ9okJhD85rHdiFRHQG0IgXkvuTurN
6NBDxTLrttVinH8D22vaw/zS8n6+OyZsfie/m4F6g38yxg3LNWh/oLBjY0PPI2ZhqCtZk38FTFzS
eImSNAKfM9GKbcnKmnZk5mAKDhsuKn0Mn468hrsDQIx8yJDtCRHr+2d7dEhQnLv/Tn3Z/gnM0qMU
DMKWY4xaDsiYyTeEb4aELNVhYuwCP/Q1rSmx7Wgc8f2Vy7yUXgLNq2FmTpO0BOvcvnx6KrodQbQB
X1yx2Cpy90WhVJcYDglkCOq/hcQb3u4mQguDWvAjAhaqjK0mz0QD9AGonj1s8WGavcMVGPhLLbRV
ldlFcLmCQilJz/3X3Jel11RVmJ1VDNX8b3BHac3kqvjkBQm+Ksx7nAbPBF6StULc94Lgyd+u0kP+
aZaGlfESB3i1VNhDskDeqqpGtg1P/QNKRSuQEwZoswuaDPNAmlJHVVmN0Yg8l9SxbTWsYlEe8OoB
vP0Sa9gwpsmHl97D/Jw39V9I0oHBY/ntzlajXb924NYVGnJNPJQG53e47E2TEjL8heU4IKUW8CWN
rpAL2nnS0ZxGLemuRop6xYqNq571RLYwIyQt676lJU4JAPFmtwwWyOvNCHksUXOxgFaRhCVIr3z/
EYIUdfTzsjhyTEPjeBbgk5otKy5VGgZp9i14R+3EUY5dNxFK05gZl9sx87iyNvUAgPXXqTDVVkwB
YKHVbtsOy8cJwbTGRByQVh/Kxw7ZgJGVDMTnRJz9kv+Dbg4SZ8xIpVOZ6VmzDGxZLH4HgCqoakWL
/9ZGe1Lbp9dNh+SnPoY1s5UNPBi+zANMelmkBQvX7io0BsXwVOlV/X6TeYpPllPibAlw8z4xB1SU
N+3L+9wdFkSgM0/kK5cehEW6Gfr+69xwLh55jzZl641RNI9nwWGr1v27DiWdRdoM0VJ5L/QkB4dX
6ZiKSHz9mh0uKLc0GFnRTZ5X9mUlv1ryWcx/2dNAvu0QjQJQ7vnDT/SilOL5Vc15t35psvncsU6D
GUOfbiJ2GT0lPEkF4ltrECdO6HkW0o4RTKQGL4evmuN8gaSLifw1yxMq4caVxM3awz+7gKUE+AUl
FibCNDvokk29fwTMrA4nwYp7CJlebsJRHNagtuvzvWQ86mEbNDQt+HCJRsuPsYTDGCkion8glTMd
vvxnCeaS3cDGv8EFFy8cc3YMXNMqAlTGTB7o4vuUtddSfHHiq3tfzAPlxdcfsKFtFHjefNuYsrpI
Ng0/K2/pFEbabx4g6xrbbV1A8eDXD+3R96KDhzLrAHaueSuyINUXlEEVRG60UlQj4V49PtvbFBA+
uWV6sz3mOTTDLW9HNs2S2pZTFDHF8QB1R4whe/7Cf0KDmx1vEfl8pLme083pu5bwy1qga+2M4MDR
DkVNkDSFd1zRuUW/J8XOkK5ov0gRcx4DsX7LYj7pebFxjUVR7uCLL5e/DHXnzIepg9TgJdGETjQN
muur2eIVHBuMNE6Z2cS3GFzbq3LajxRkBnuA3TjXEaV4nPx9EumkrIi5Z96vxkKLFJjNGI6G/uUp
zA3/IgzX6Og4oDs/H176CqeaVuAA0hbPqH4Z2ck52ACxZHMeDvYDP1SmvmxQUlZ9BPW6vWGh+PHp
Mlngtsmjbt4gWTZJxedHNKMF/YEklx1QB1zL/PXcVwco0lu89Q2cHtiFnMwAxk2QYgeqEb9/Kxz3
AMUuNuLHZuAfKj6zBhx3wQFr+/7bCvzZUPT2UFcgJQzuhITdEy2iKy+G8lim7GK2c7JSP9fHY73S
75i2yiMF+VHiVJHxEZFRK/vvhdbEHoAoJ3uY49A7C0O/ILI6sJ2x04vfQw2/i3w7aSPg+UB/nt9H
+Plk4j++NKghsZn+PJ2LbqyQ47LzLrdomnLDOY1sj48+e2L+BR+jGQ8jcrUubL3EyAAVZpswn3ZB
0wyEuYTVRF+K6iwS9CzdumC3JC3JuQB/TCnXIF1e7wOjAKYcQ6EVDdmdXZnJgJI2usiERoUKA/Ie
D/Yqh3EK94greXns9WkAuxDHaaMQ1K6e1pFl7zCPNMCLsvfkjSUKnxO6SaHmqdhg/zI5mzeM3aX0
dicx+a6CjkoXLYazOUUBzCkz4mJYlLu9DSqwHMZqIPihQqEpUvHsES8bDmeHzouq5p6uWzAogVw0
i9Txy49N63y+Pn/yAtvNOs7LwN1E+25OLe8iZiZqn+e9BqrsClf3LEkzVCBdKiO9G+2vP5uwYj/j
SK3v1alb5LxdRno9C2S0de9oLiGnwSAU6TtjmEkGew1sPEGVNTsQeQOkPDKWis9C6slFmrOkIjKG
ky9rpYhteTm5Rds8q4DGNI6WXHnp90/ESPQtdPDxRjvwIpUvzxLOGSsn1QodBJY0ec1QvIZFzscU
geRR/77jULe67JqMtDA2WfqkASuiCD8U6nSsiHt8Gg7kb/AjA8Z32064MEsb9IkuSQT63iOlNlll
ccZhWx1uuV9sW+rJq/94Omh/Kppx8yRSXj6RFltAuK/DU8STQd8i5gsOlrGpRIP/i07gnbIIRHbD
Xt4n1t/MEgfXe65CUduwS+iJuLQrlUFFGcxZE71n826k+CC1CJvxww5w0Fn0yt4EOvRe5VjuaGQR
Y3d8C+ox9wkebtf34q6OY4mwyjns6I8BhLFnYozzU3fkDLkaK3wZOfCL3ls+N5KGnQQj5Q1XJQVY
sLQC5uB5zBOc16g97esrYvmS/f5OkS5nRPuy0FE2NHsWI9HWHmP4nIBEKpXWo3doSC06HNCLEVun
xtG+/IT2IHI+Ftv1PrPAM3icJRGPdMxyYO2moQVG+UZKa5fsVg6G8EPebM/Utty0c3P6Z7WGKRYX
YhQE3hDBbFm0YohhGMQvTkYiJrYrhBKFoewIPL7MxQ38Bijqh/wcOTwagV/7577bqfEF+f3uHc/9
8n0aqmUokDoGYh3tyn2VbikzWH8myMonUHbIoNYW25Czk/KTadwMX+nRYZr+u4QfkeMbH4pv1JO1
Ala0N/kd41Cwb9ht/Nbybbdtfq8eLIxsM8qF0mrHCh5zDjObIgRyLuH1Ogn5UfE600aWYLthoD6W
sjKsWKvXJ5aiDKJtHTGW+s0v/x0iXehK9vyfQQ4rKu2BLoiQwx47dRGvhyGCvYKgGw0SSnLr3x+1
6diHQNpuTV3wEy/xdKKOvwS0A40ZqervjMNX4BXkXbAPny3ZJVwMLl55Ktxqie+9K/L03KfQe4Qi
6DJ2BPtT9e/BFgLgJ+kSkoyV9HRQdTqVVM0LuVEM0MAndNkDaviu9YBeHZp1xYFfXBn4MSYLpEru
t5lt2CP/YYFC0BD77a0S90dfU7BrnOqA6qy1JF3KYV6TEqeUZFE5yZ2Jzl+nhNqk3VPMK+xJlS/L
OR1BwxeGy1zoqWwnOAA/5uhNAwAPxLT6RrayyfXQ4Tuo4+epwkkMjwIzdq94+IjLNNxcA2gfe3Vc
zxqWESND6JIvjKTfZW14KBmiYDttXDdK2rXF/a34rCD1YF2Wlv6AzRKsoXNc6FpZL3FqEMtT4iU8
6aGO7O2uXjCN1XgA05t9bBidBuS0UOdY4uzUmvK335bLgJUnAwCs4xJJvBFHOAGMM0wXrLCeig7o
vf28T8enT+22Ev68WDcfJBJOEgshlHRKnILaJGtO4QHuD8IVEbNyw5GFH3+UhBjBF/1OhQ5LQC+R
YHkDR16i0KrXk8uffmADY3J3LZkZeYdaRYmYj8Juz9MzQ+nLLCbrT75hi1Ns/lISjgi285nKnJgE
BMHvCMyIrmHDF0x7QOD0/LRTJEDVjq8Yg/PvIRf1RycbBHLccN+1ngiIgZI0JTySiT7os8/P0uJH
eklRT8pNS7XUlclQIJPgHa971WDm+xtNuibyWNyjTbwb+eZq+0+koFuK3zZO9d5gdG6TYV4UsCjh
5JFVP2yEdP7T23h40FkakpsAXj9fdlNtnJ5jh+96a/MiS2pq5QtkTra0+RnlMIxG5YdgQF/1AzXt
JcOR9ouPLZK6aaOwL3G0iCyJiPVbvKjn4w8az/CDo5U10KqOOhUSWH1O4QqJnhnnkp1NpeI89y49
6WMiXMNsXLgj/fVLWW1YZQ2KE1aeTPZBr4UyXUDUcl1qU+nkKnU9lC7TuuDqS4ZfvFZXSaQmZf6G
2k7k8q5WPoAaXP20aA9LjG6eMisk6BiYsPRgRAF29idQxhsw7tNf5hu4Upd6h4PiaEBP0UCYU3p6
08wNWOWuj1w+km32U/tpLVcm/XSpDQNL8QjTgmVgo9aLJs5wnGtVvU/85N/w7nQ3oZ1OJ173lI4P
WuYp+2GUdMrqbn6QZ4oAMIppgOOCk8j1SdWvUqvdFiaMqEQIkjhbsy+XMDClFKklKaQpYqwP2utX
XnUIkO6D9TCUsiuLwE4PxSmIdoKtWP4UDXyZKRxOEcE6xuMRz36iK3Jbu3uTut+y9tXTKmp4b5wg
CnHejHhbtGOYTMrw+fCnZjo627CHG67+BfEkSwfCG/UfaRsNOYv6etOYV7ED8CKbKsA1ecLD21Zu
b8U2ebF8cdaQaEMtY/kKKLoJzpKorUBerH4AKY97ZMUS2cnJR74KJdibb+PLd5BKxoaesQgzOst0
eMkh6jPwbX9LdMWkXfVRv329a2ScrfDjzyl6v2SavtyVNdkEwUkooeBYh6S/M6yvbSx4i4fncueT
U3F+R5Kt24fVizWdWqdvwllSA6d7G77Nq6Fk6buyrUWWE7yw0D5QEabkVfKj9+K4LBkSy4yOd6lv
AKYsYmUXLwIcq0jHXl0PFkq/OYNev9jMiL0V4HcocRjaH8pJZ4zvsjMiG1XBrqrtqjkUBHLHL4u6
RTbkAqTh6cVNLJRRg6vGhGMkMvwgQu39JA/lFjqp7U0uo9wn81THo7SmRGlqno7tQ7VB4szvtnDa
vFhN8B1tJKaFVEtUbWCGJpanAmdOogHG3nBMtBibAxbWI9QX8h6SA7kYkay2kmJD3t6UYfXFXyAU
KCse/+R/9ORNj2EO6VOIWTLtjJAl5NeOWiGvpwKChytUQz6PtZg/9qOwd0Iqsn6oYjJsqC+S58nx
QiFNLUrZTanXHvyYdkH0m1CuqtRpFipHCGNl1n57Wuqkpzw1Ipi0c02J+PZyOWaHzH024676e/Yz
IBnX/133gIqKCdPLM7CSV5mz0mWoWSorr8xlC5/4cJhZLuNOHZ5ELzggUMFNdE4lwBxj67Z3WQYe
YvFJIJ6VDvDrV5zEg+usgk1h6TOWjgzUJHMvfIU9CrparuYxf00TS4QTolZPgOJ1JA8RYHGe450I
uhOiOpOx8v3lDBdRkwtE4P/Y6MqBAzlIMTooTSuK8nV5PzxUA7qLqSqQhOTWQ/kAwxanFnX/E1pi
ZT5iFH34mX99XgzAJDqa4IdG/EhSS64O1amM/c4parNpms59SpDtQT8QlJMb3Ph3H81ohqGA5Tbl
FFmYVF71AX8jwbu03e0oz14EaA5qQWmG33n+uYDwWbd9MQSPoawD93ZKfpp9BQ0KJqAN77vZbWnG
erXsjl2NOAVRk+LpKzVAzik/s6MJWP5T4XM/JfckZuhhrdFVDXUjALHVu0rcZa8jiu1A1jE8IlZU
0UCYmLkLPYVV7+jt1iJP/J+W8jVhUHo1vE8c5WnzEFhnfPmU/7y9Li6Jt7751UBPIMX8zoXwgwH8
mUFc2ohm1oc4FDfHXauaXoGZciRLGZ3GU1LmibcfK0E9G5z6Y2fRzMYSKeoeg2jSdsix/FYgfQkP
yEQYw8RcB0D3Ivo5dvu/EjpHZnBntChYdelKdVBiNZpCuo5L7kU85S4l0Ro8shu0x4/PwI/mtPT1
TU9cnJwGfXt1lbviW/roYA9ogC/3hP7c51t/FNFvtuBYDwTQywDNiUNbzZoaMUJaSv5Qyj/mM8pZ
TcTGdsQrBoxk7vyteOhwdcOlJAy4LqlefBtCs4duwMqqaHJQC3Aw5EM39nLMrkPm0hidqTwqX9pP
EtpeOJXXG1nN1quniXJxm//J/ReBcWF0spbBgh3ucnMPSPXU605v8QPdvhOZvL1sSQoAdNuhlWgA
3tTVB+WfwG5TGT6tWeHX22AIxB1sAAlViCA8+2jqdOAlz3zRgZUUCRyCxK06/olXdFNWvNYzREIq
48Rpz62fsL3XDf6QXbVKIUTKDQBhW6LG/lALbhRbyyf3MUGatjpeuHAIkapp0Sa/cQovyRxvNx4X
Pkj4KWCK/Sh1yps2xfJjndFgZbv6FZPu1wsTGz0J5Obo4fC4bSJGvb+nOootzPh75LF+SRpiNx0E
vNcOa4KyWWcf3/T9ei/pTWjmVc2MtYvWnUytiJuJqBN8E4DG2W97djNazQxu9b0scwcMCn5MYROx
VwlwMFkMGEetcXBrb05/Cq7Owi8s8ZJDyLhJugdEWdLYOtizPL1th5CxAk6SxGIKG3/PzG896S24
5Kxf6gQfj+1CHhL3g1WsebNOQMqO8K9ZKUPjglk8FfqlQJxn+PIbc8E7GWWKQHB4rNCDeWdM14eg
B3jJRK0Jh9LGtqIUs4+DA+9Rb9zRFOHsgbk3lq0CNoWffJwMU8wcccwn52kz8YRiWmlcznFHbmzG
4NXnIPIKhri0MoZwcP/qusvCz5oNMVw7A4eE9kekXZaMG1+CJMUVxyTf0kzU6OTcLVjXV+CPkiF4
taDO2uIxbtnwL3n9oKfvW+etwUHb7cwASz386k3LdEtr9bIGdWg6AJrZqefApp2WJA+dDdfZ9O92
CGgOHOcEpLeHw5Dyp9vdL5UJbIQDzpMMCsKqHqNoYgS2n/TQzqjp95pa70iKSh//r7j8kevCl7Vt
TU21TSKD31t3YQ+nrB62yTvRP7W0W+DDYL9cDNJDDQx2nz7NFiBqEd0jhLX+nX7nQ49tWNvFvzTR
jycypW+QxpXJuC7/8H0vMXNbKVNaolbWZu1ckP/W5+Z3UKwnGpIqVpH+obghdnqOWafM0wE6H32V
gYNRxbCZhtvXJ9jXm3gvFFBrhYChiM0EdcBnmneV/l+gBVZ0lJHWJzj90R0O3KMhPTf5kb3ftuo5
x+zObJ4ovYoj0KMoFofmhnsgP/gjkeRG7QGkYCPDngTlmW3X9hWmuKNAeDRLW2Ybz9UkSudjY/o1
mv1msZf6U3xnVxfZN7BMtAZxDKlFN2I1BFoqXNTMmUgIx4JJM9sHvjUGeVM0+EmBz3l7LDEZtCIO
G6MCEdx01UzPC47uuhBK2948PrGAZH8yZ5DoSzI0WAtYJ+orxrbl/Oz4G1VPBCxrwszIZTlniZEL
EyHZCLBjbccY0UHMoFQPFFcwHvwWiOCAYF1egiJ6xMEB6LVPFw734XBQzePra//KHcR6U8jiouiV
S1B5Yvjo84oDvyGyRpAKKMOKdl1itJPCccavrZL+QGXKaVjszhYFK6N+D1ki41nm08mnbyf7z/zO
AYyrM6mLgmY9SA60TSsR/NRX9sgR/zFiEM+lbmHcs24XM8eMtSWM3dDoTvBB69zsU7kYS8bZ6p7z
j5rmtN9fJ8dzq3VxWGErqyHCjy1bg51L5wKj8uc31nZ0U42Aq87/LYJhV1NIk0R2GbM/dubR01b1
Q/cwuQyDqPTcx/Lkl40Y4mscwAkdqVJDqxmbPl6SIACwtdN8sFfAuWfc7JJuWw2qfGE19YsBtmOU
11dhop3qMG5/RQJqb/jJirSc+9oEF8RXVzFVRbFOA6Zj6wGNHLdUhiqTy4MuzDzSy7VjezLGWo34
YbxKhMRFYj35f+NUdliJ8oUOvSJUOLtWlWh1n2wJ7FoGI/cPKsszxv+Akcbam3PiyH1J4OHwfxYg
f2G/P5uVsfNc8sOAYWiV1igvkbb1FxfpH60lLennN13JJNol69mIe6sf4UcEBo7WcB2l24F3wOn/
pmXSfJLHuvucRBz9d5xHAJDrBAuMsquPHd7FvTlVH80OssTGONfFxvw01vrGsJws7UXkH5jr8kO6
GC/B4U/fNkDOKQr6yx554y6bVc0anVdGWjR/CL1b/7Hlq9zh6Ol/0OeDLvENmqVxS9jDIBTWDZb0
qnZQtsHCOUWwgRRih39/s0ynz5di0mg/4A7P8hVN1n71Iktc65v7CAfPL+juvxTUwUvJGut4L0qg
BeZWthYCOG6FDiUptzHnCJfedt+EuYcQ6Rg6HcQD7osz3kILt7MmwbXMr5ll/Y9qLc5XX+3qdqGu
wmb/JWV/HNb8vcnTL4NgQ9Yhg3bcOmN1Vffs5FaoMcV9vMdjLqOTcV0cZqO7A6qNRYlDva59JgCp
KwgBuR8yCEMoNt7N+q1uLYtlJJKEx+X9/AjmPr+vr+AMuR1sNLTlnFn2ONh8NbN1eSS9xagLA3He
UVfrXfck5Il/4OxiDoe//5L+6yoS3RMw5H2uwM3PKBKQYwcUM70bBJ52Zf8s1MXbfU9mRw2gN4dc
H2UHTI9UxBJOHb39SPD+x2v7tcQwmJX8FBUSldjHl3G/j4t/dzgMaerumdhwq934So8+wpfEKjcn
EBL7Iz5niJPFBYshVlV6yo3Np5TfiolbFU+6Qi6FmUMC0BN7SN+cPf/82cJI8bkq2OFR62cxg7UN
cr1M0GTf+qc/3ghMyKBK3jpXhwMorp8FpE2UuJrEG8qZaxG5Wh1tDCz0X6kNYwWybCaxZTJPzxCx
i0eb32kAunYKQiDxPvFNVTfE7fTpzWDx+UNnroHMFdzc+ilIl/Ig4xx9CKLJ06lhaOaUBHZ+NsMM
OkcYdOgHF4UYNA5DepeTIKsT/RlQdGQMYZU2IAGIBD1LV8W9l0nIaGfn097WaDMAo+RjnioDr0a1
cy2QcpbCD8K3loPSJOa09KfXb0EJXOJszOotvnhsqwTfVGZ4BmNgNACWL6jHfgKBV8AUyYumIM3l
d552NJ3BukG/xCi5waw630HDcP2Q3zPf0R+GePjHgNAEQXvUNhveEufX7kjsjmv/clxpVAgKhYcT
EMs7o16oo8n3biff8H6nYPT2qPCml7OkVvdNvjS3QVP9GIV7iS4qEq9LJcUqw8paJy+ZnEJBDRlQ
iXnYiixUSJ4Sk9Q8cSr0wUNRlC2dXW2/ptzDZc8sg3dMEAxI8BD62WvVUXbgFbEqAJ7wITRlp7l7
gEVRJPuXikJmUvDgozsNhyxWgWq0y9+FF9z7dH1yD2K8ZzNsHvBerbQQ8OpXRtzRrDTiixck48C7
RJJdVooZp78HNgLWxI+4luXsAhJ7j+drIjX5AGEbxN6/7AFMGZ1+huXNce3J6b3+BIBX2eySPw1r
Qx3uJnoGO2GC34mMPy/VGIfpAteOjSz2NkK4GKqDBgkEJggFuBzqnT5WLvpzsWxmbyOk/Agl9CWj
UfrSUGeYQ6ue8MJLUdf+N6pEu5uZBTkCTI/xiEh5Soiks+2HiWSAtDhDUtKOTr4t+VqcYRExF/x4
IwXMXuvpkmF7DqMdm+heTNW8dWikuzAjcYsMEVRDrBjlwvxlWyBojsr9k2LMYwp7lhgYA5yMndHR
D30FGm1ggTi6Z0r1iHDJripWlcE6xRaTVWlK9XS6B06WMoicCNh1OUcC7yOoBf5ztxiy8K2gS95t
l8kq7+WI43zB55OvHCMoZJY5ytMbid4B88tdGeHxvW1lV5FEoMd32v2qwXiBRCEzqBICKD13Uykh
v5FzqYXyKtrDTD3MoiuV87Eb/QwThcxCPRCcQuWjT7km3vHwhoJwnotTo5Cc2s2ji1RbQ/rnQfSz
9cIPnJHupGa07SVW7gy2G5cNGe5/Yge7w9mJtkMOvKntyroquhBj/l6BfxdbwzL9TVnUpeEyfOxT
AfSl/dpMookcyBAbfCPqDF8OaWWCrOlaSDDy9Y6Fwsit+btCWjpkBPZzKgX+4hhpi2LlsLwatRu5
Wb7+KDSl9CxiCSIxGBQXTjVqBwOxFeM8JIVi42xH7RkH2sIrooqEuSsYK2fguWiZXLV1a1/0haUq
hdUhSHHFQyAK1HqcZ/l0cVn9sStjpE2RI6O6MMFjLkIOug5t8qcc1Sy090KOiysMLhdGnPGBXJdG
DDqOY+DhjmQWdLRVZJye0bJZUuFvOoUTEQPouBshcUT90PWHWz1Ev5/AkvK06FdYaxfB6AW6aIuC
Dwwzk+0jYhnlRaXIN2xzN3vvHdDQUkdPZiLWdDnlNU4ac/GHqpA0bApuICvaB6LxgqD7lmzZVCbz
YWM/Udh3S+vdvgfk+plCGjpgrCZ5e/ufy0LS0Fyo0+4o/TZXvtmghyOTGry0fbsvbQ6yoyVfnyGW
2C4GpGQQ53vNqQkRZzsN+EX9nZS9KsirWz+tVR2yiDvgmqeHxMKf6W/z5/iFMY9YLAq0hMotJvPB
8gKmZ9Kf/COIBbLQll+CTiMWIW22geAOYpCvOG/qhkN+wpprfGYdieM1HavzFMOfetvmfq46IF2w
rFj8eDk6hXcz/SHmD9iIJJhf9zlHvQR8+fx26evoKSqQ0g2S75kqobT3wsxHI+DkC+f+siJIrI70
SwGkn6sGSFg9wk2pi1YqMEjRvaxsSOyzDi+qnHwRSIxQDc0GZn9y+dgn36wC74XLjtowWMgSn8Id
Fj4/QTeTtZggPmoD8ZUvpes16OUI81esqTvxokQeM2S+Ln28dT8lhOglG92YyY/CyZ8146Kcrfqa
4d8GFO6QikKNXEXCvC236/xvzGQRvSpl0JQc1gr9OLloMTMh7spjT6If9QxXqU+Ic9mO2qrGYo51
rDGKhmkAwNue0rR72ry6F45fbRfVwFupwsD4tMdckzuS1h9Xs7BeHCPIItCPbGXsi0aNSq1MuPkE
VVQs4nQR++xsou8mfkhf6TfR+IseYI6E5rOAhpynXo12dbKyaOOaZCMcyHNHgTb2v8ivw417OWvZ
NvkXhZd5yhVYX1DWuyEMdNCPDOr+vB5runjZPsOEEYA1vrxbWxc/uIYogAi8HK0tsP5phYnHPwUy
+7PyqRSrsgZDSFIK7xehzo+Y9bqq26bYSYCtpnu2V8ZMDq4dzC4mhZVKDM/uystkeMaGqYYUCBXQ
eAWfckoqiOKpmwR62qAOb/KLiuBYwAtVSQNmpN43+mfac03jAxztDT8/pEvWXmOxV4w1hvSLeuXL
bgSnYvZISa4W92sWvgrmTCRd2T7RQBNADxoep6RkJ1Pu6pykKJzV5V7sKEM1ROFNr4lIk5mIBwMR
LAlda22go0/HTGN3J2GMAM1PDSKqTyXEni8kAwZifqkoKjkzMXj78H3b1+qelHczUJuaBOF0vjz/
DyWDu5YNqHcqjJC9FgBJ1gpG8PN3gLjfxg3HURiqQfkqQIuHxpdcBOfrz+LdfWVaQwo8FDiQyt4N
E/A+Q1YRnU+HjcXjo23Sbb8tMJvW5HRp6aiGPb2iSMSEsU2Gw64ea8bsCmZUGxfW9RZz1G80IX7X
7VKwYjIhmf7BjZlEg9lde7b1EvaQ1OjKc3OyX4eq1mmCkiKnYeg3lbF4Yh4C1y2ZH6/wX18FgQEA
Wcu4RPMwL7KhLVnkViGis6NKkZ8iecUn6iF/MbnqiqF4ITpgBcORcOEvglRVpHimOjvES3Az7inx
BwQqOZyiOPl5lx5Voh+7gODhBZy0JRGCQulG1alz4ZsFBHWzDDy3b9iXfzFP7sNygaIcXPtSykHQ
7HR7PeZJOOWFAJKjUQboqCDMCr8fM1DV6X0lI/SqaujToVdbt/RqVmShBRYm9EM/Acfp+5K2+aGF
YkIiJ5t4NTla31W59JSiD78DQ5AC0vWgC3uDIyeMdij6QxwF/j7l5bZJ3tl3/ZeM+5bBLmhXeZzW
akaWDF3OR8ovuIDQzduCD6J+jT+qC8bXWfN3AtkmcDED8NyWehaWBjlGIF2IHrf0Dx+Gvy6YkHl0
qb64ZofINkXzgplrG8HNB5OyO1+myc7H56+OZ8otBMAvEkjF40NVeKRvg+H7nTUZkXMGNu/e5FBm
Dr7/X5nMuH50MvV2JuduNtzTp3Hm3Xc9NckUuKHMkI3Ky5VGl3zYHKgCkI+X5bnTG+3SpNN/mJHs
sbSV1onybS3Xp5fG2sxRHJ6C6nVq1CgI0GM2NmMEa+5pzni5B455g7cZamokyd9tmqeEjKGcl+HE
OYFeflU0m0DxZf1udcuiohNDL+IBBQ5dWjsiCbDyZW2pmjS6bdrUWcG64oHjoZJTwoqTsr0dOvIV
2p1mHcLgrEiDQvBkkcRUUVuNL1gBTCKODUoxc9FV5B8EMNFNjBahxTnT8Rcv4OfU0xu5//UtAtu2
dtyEeglfr21sMS/70nuBmXChijtcDo3yW+bpzkhhxfcVsuZBbCWl53Jyh8QYgTzemGbIJRQpvCDi
YIiJZBPEnD8I4DhpUSRm2VhrAnhKzPrNYYq7hYzAZrxQJ5bS9zO6Rx3BlDYJv4qRYwtfLpBSnCXt
yXNsISFvHCPOMb2Fr8h6o4YdYkNyf+s+dxaBNSjzAJ/sNtsL3CAQrU2SiAABaiOApHYyKL5NIdV6
pGZRlTtbY5zTee2DMBWZ+s0lxdwTpKarBOtc012m/i2F5MdHTZI3ujx4KZdcbarX1x11Gpi2ZF1v
yN8yBvf8ndZsSqvT3nvg/1vJLPHuyJoP17EFfizAVsb8WOjlHK2ch/gOionHc0nQCsSdrNYQbSqm
1lEVmm2h7vUMVKdJkNbkN6+VgA80YHtR7FAet/9GvaLM/jCeNYzlE1cYeDJGMKPgFlJ0ySsGcQrE
bKZZckiPDHF2nBiFbXAxoMP2TAa8XDfB6YJTvLGB+YoCaIf9x20h2RcLaa/nzOGCMjQsi5AFqF9b
g/9NYmfp6POqtoHQ2OAX23lXExA2ekOVAukVh3EONsWJFViACFtUA3pc5+5vGC8lIo2uo3gEmNOB
K01tMorpFBjTRHsctT2WWsrQJ1FWENp7CQUk4Dm6RzssnZTJl0+P+kAGSLXJtmL6YE2lBxRitzhL
YzNeMWpCE3nQycxrCk0vqrSYA+dgdp/2Ie7vubSMkXQfObbEe7o8s9fGaPlyKTxt0o5jCpwqBvzI
UNewtlp9R1rLbfUI2LzYQx2ylagk2E19i1x44wh7+PgoorndJOubsyFlAzR1XyEyB/IgqWHIrBzH
kqhdN/KegCbQDf8zL0ag0YvAiwisw1nNELPdWG191OUUqPYLs67BLSSa6nbFRydHU039/Z9n1YnC
nJE/qWs1oe7Fk1H/kNXm3mFNdsO8KWtWtXDFrQFgW6mfg2CyEOEzSBPqqGypwjoqds2uBEQe3dVp
Cb2t8uuz/imP7NCNdQf3wQnfy/zxvMXqE8bSiQwQ4UdQlWO8YM2UGn82vLEz6zp4n30sJb1+nhZ6
BzeaG5FZ8A6fOsGbxlVMF0yg305YuvCoiahKlbiaNbAlSApNYClpG/BCmydwPW0t076Otqxi2xHr
ggnLuoc5a/dDyqIZ+SnHw+IE4TsQV/xwhaQdAUBusObIKZ8/LK5nXfFz68pYNzPh9MgGVlTjBlyJ
OzZUZe00rfcWjs3xFkEzfm1LBlWbqvaLJ+E7lun5+Ce7JyCjpJtfw3I7UV65QX33s3cWABhVfTFo
qmh22Xo+XqrveuxbQ0Mx+LDs+Bah0pKMUdhvOzEtOdgSQEVlN6RDq35Spu7H7nKpyLTpI06o89KX
EMjpd0YEKIu7BU+Dcc3Mc3j3Hxrmn1j086XaLCWK/2e/GDBFKoJPtHW3Jm/TzdqWFrdY+98YDz02
NHYum48D55aiEtDL3u487K4a++r4jfMKIQmK3/0k3inXunNH9clN8YM6FiUk6sBbQfQPC2SzJ04V
A4lML2ld5XkowIzZ9n07fNnnynF5FMNlV8njVYvS/HmVOxUwCdhFXxWIudJwhBFzjT0s0jdeNzUH
uSBsqI+TPw1ilVbwIK7rFr4ZSG25Jrbm63pjdIIeS9YMvG2iiCskd92aKsw8bxj6xyPZph1WfHwo
d6ajNQGFl6BAVCoy9f7/zeWL5engPOiSfEccXqCWOMoalB+EMn+lZIz2GB6tO4YU3Q7MWNcNt5PJ
RM/NGcKFEhbkz2uYbd3kOeH+xEkjXw9ao6OZ8CS/bOQpzSJBe4NDCVgxKt1U6eArSdWDBiVruVcW
3Y0RkAoBG6ZmaS5KtggD8WIQVj0kf5oWol0NVuviR7zi/mZD1m/feG7Ms+e4JO0nC8HJ3O/ei6po
QaJh/qHrBrKW36hvoeroULxAQ6JCIORVcXSY0jw44oiqhCSLRZI5RRRMHz+bErVoLys4SCG5XFkC
sIvq7/HcSCst2zfL4CkuqPajsLKuT+/4Vh090RMPHDtmICoOqL+ax05SthbuHnjPOdVa4i+wAm56
MVfH/bQAYMRnFteyC5iN6NzlyflKyQYTu6babW5rQk3EbifHyIoFhdRShFXTnUlIFs2urZMw4ZPE
nnWES9tIU5wZnyoJJnybazXM7yb+w2wQ53chZOJ/yJ00sw1lEwk/lV2JaIQbgPEMdmJ54Yf2P9It
8zqHuasLIHrzVRsxNN7H1or+9oItGp4uidPmFtiH5VwH5uQQvckNh+hi1WqfvLJuPhgtbTjaVvar
Y0OV0JxgyqyYkVpGGvkHSaSknENqoKH8X8nJr/uMX1cMyvLZJw5glls93ojbMXmhCTZY2DIdUeZk
1ynx+obecI5bam/gtNNKAooP749h/GNb9NJ0bR3AnKiUtM9e52x7WndfBbxFqX/1r63G5CxbuwRR
6myslH8Ho4RWPRentwMVgrVt96ZkJiobI3w1ws1NgWYim/tfBCw4x1qKoJMIJSFF7TDwaObiYeEt
zn3Gvl7d5lJm3wVkSl5fLKaTKCJ6qe82ZCoHM/NDxppJDE47c3Wl3B2a6dZNv6MdIvPf6tSL4uSj
k3DJ6tRY0dv2MzKKHVgmk/SNaTqhdo6k5DR34+8vsExGi5hNrutvKZhsRwlkLZa96B7T/nkEfuw3
ZBpuhk3kzXhdX6SCxyfhSaaZP7Tc911THHs5oNSqz3EXZeGjN0rL53ZKj7hjch3OY5nAzirUjUL1
llLCbL9Ns/93975SpZm9UwWlQJ72x08l/8NuG6Kw76rZrVzSJKelhQgRYNMOpG6LI45RUwabXaz6
vCZVzQMLWPXYQMPKwPOrC7NNfqCq5L1k8WYdpNFAm5aICjPBXE5UAsOl3FeO7CNFaco7bGTfHZMj
updL8lpf27D9EC+CR31dh6zX36D4qnzv9uo1UOwEfd2L3lzh7Vg4avHBLgApBM2LzDB5BEeVTIR/
c/AOhF2nNS2k1s1J0H1/6OE8uPeB69AAjq1Icv6aIxDEPicVY2xiqgByAi18/mYVApNX7CzVJyoS
DHdLfTvtltPj9xav0OuOBranFr1+qLiCbBKeT4QGGCcEDTC1ud9CCr7/Io3aSC3C8gfY+/Lv+9wA
mW0xJyo6NliR6QeCihUpW8CMKxp1CtzbEbcMfb3YfmeBkhti0Wl0+2QL7weysCMX5uumcpzCTdga
pxCtP4xMDkLVy98LpgH9w3srMvNMZU5oOeJLIPpmvHIWWrYZXxxmnNUWy6Hmnz8E6/fBR7oVPY2P
6O2lEh3/DLg3i0LiWTyl9bOAoilOgWXzVP+DE6oDZfU39PNVVt+lrIaDsAHXJdJFNml3CSGoxWtj
hhw0LcI9ikHN6yiyhAHManX0xEJHK3b4EwZCyXiNPLBitJOjM6arCBdI/x7+AhbpEo9mffk5ZZGQ
j/f/pdXdIzuF9Ixk1EMWQ332sCSeRs6CAB5dNCX/LUZGmnaePgnAIxaacqmuvzTQfIe/VTvwQfsB
CQiKIPICyhoTglP1+CDLq8TjWTp/RdQWT+76mpN5WR7LjRetMKwQZ4RS1I/U3ixGfU30A6AmrZoI
z2VqgnT2VORxwwSzz5PBEqXBGs1XRjp4FhzGvRQKnJHv5uYNkcLiNESE+ObRo2ciCLCoPze1gK8Z
NC5Y0UxGEGl5va758rQgSk1d8HZfmYdTO4GyF0pf3+HiItPDHH0SE37Mls8PAPegls9No6AfF4xh
Sxlw/KVDi04eSYwQ7iAlujp0EQT8KViCpwinqvJF5UV/u/gGPMqCdJKVirnx1rVxVMWHcBFod0cR
CgFvZrB1SxtK8xvGcYAhkqhinsjKvoY4vkgPqZvGJ5l9hPiLmxguoyPaG05JvHggt8kNxiIq4/kO
lgZOf9MfSQd2ltoXM9kkvXukj8kDHoCTl7l3L3en+cFxA2AkXIYhnbQVlASeVMLv3xPCmZmcRhuu
mQzKXY3JtXq3xKvhP6ls/MVlNkZPk5AI5xFuTNOyt25EGffZAB4vezcQu2wddwR8cHFhpf+Au4zB
7666t9BPo1UmHfjQQOuY+w6GfJkagGNsbTPt9lU66epGQsI6vc8SHJAYuT+yGNEslANnGcYOjRlC
TpzGzDdJXadIuHhnSvx17ui0PEN/GYuD1yTEEIEGYMkMvO0thNBhSc9tee0A1mPeu3xt44K1Yxu+
sBjPrOfiUWxxgLJl2TlbfDS3pXvfkEJV+9dbmSKHMj1FQQP4SAVuKL6DJanAj6YagEoOUjyPvInU
C0zfnnVnafS7cWdVqB5ntk6//hU+GAmc1Cdm+ejQsPkXflUTHotjgWMUFaHSW5e6JnQDC8axsn7/
71LAP0VcbH2s3o8HTiDjA8OlJVh/+ocwGnX9exRhXqi9U9I8+Hbkr7/ZZJ+uglS0yCU/j0nlrW1O
wDsjIv/NwY4soJbVcoqqMN+S5yQFJ9cVjGW+csGq6LSDVEDYL3lHs37z0vd7ufJNjWt0KwtfDi3R
8YtUMj19xRIT/PSg82LULtxkt05goI6p79XxF37UgTh3kBDAUIKfN281CGeBHfcVLec77sr9TezL
WPB+xCse6EqUaH/kNYGvcSADnK6eij1SRDDVySPLVL4fccssvhaLKnuJB5nRIudGBrV+jtRqLgV1
r0Z3Iizpjf1pb1+qKKqXZS8NNrxF1zvoU0VkZ+IQ9/LvORnChkyz6uEa7P/yiICtnnufISDPLQFI
SoxVk7SylwXdJOfmMnYZ4A29KQrXQ/UcA8sKCSuiAdWxsaX5xGtmWrVboawdF5gz5mnoZZzgzLBY
pHA/JCZbRhk/wZhDbh3GNWlL8C7WZAEKhkyT+3mv9SVnaH3+VjUtk6CG8aDjkw15NuW1oj2Ey6BB
AXNrNxyRU/bamdO3beVN1tMxMr/1ny15t2lN5+ircV6MD0sYUFpzYFEr5OhZDGBSK6OTpLCgSr7b
IgT16dlfTHhQJxqOa51kdCGM8pyRb75Ouxxs5+GySNsRYcPUIXfM2AUyWL1hjzfD6/w5+LBBHi+V
JKFHBj5hA7VYu7pLBvY9L1EsnB4+QCN2JQ6bu+YNyYHLEag+1Wp/z3Clsp22lrWj3cdpIRXeMAjI
hkb56Bwtpf0lKYugLSKhmnXEOKtQN1VbVpqeB/LSFbbxyD19+hLD+sM+sC/19sESeQCTiVVp1Y9H
K8FpbSXXSTjbXjpSgcNbjxf0lRBr0K21ltj+vD/SuMH3+4c2DyKPeDmT5NIcJkp618RMVcXD7Ujk
2FNRPTjWDfk+AWhCAdB1tztS+ZBZ4qrYAUI6lnBS305ZJUG5mXJwIkd1uZVK93J9GUG7Q3hVESEg
lHsOXx5Hmg+tc1l/+1Ic2QEXNi3s/FposwMawyQJcwGnxwNG1Vk2tiGbADxpYQ1vDYT2UOUgftfz
eEh1xKSSS6Bl7UF3IYXsMS6jKXJyzAw2UUn7BcL8RESuGODv1HgxQ5zoWNyCEZanUGYOe2aGOxsW
1ikwHjS/273jyk1Qmbzo2vmjln/hj2dj+n2Zy2g+1sQ7iLm+jlevMyHDBMRpMKzShIaMWriL9yuE
DNnKWUAv/YIZMKvS65wArT2KxA2n9x3Sby6RgyjF+5zOZGFYfFNgpHss4YmdcXGS6FkhH//vPyjM
hERV7bCJdGnKHh8t9Hc0QaCYd9h2bRWdOZ8gKkb39g7iPrvriVNUz7tKvJqJoq5Q1oV8qYCsY8VA
ADPfTTd8hQOaKCDmILjTE1HwdAQTUDb2FJA8KfO3gEBfxUlZYdHPuG0+lAhW1lLDi3TWvZ3R1CAr
aT2sA6gI2srOft4sz4AAuM3TwjQ0tTMQY6itwNnVqFD3UdL2ZO4y9jJrzjgn8hiBP2RVj55gjZGE
m+XAggJrKXzDGYtJ94D+z/WNarXkYg0lVeeLEhhcGGTJNei+znM93OXYFPG7MjMUw/mGhRs5h5Zx
2DASNKzJT8MeoZ8oKtbGg51+5B5/MlCmbqvXON8C1zOSCgH+SpD2ZHEDhidafAMNw/2KtZrC7bA8
fpspDonhewdmaY3L0g/qvDmNZNaThi6gfRhpXSS9vGujp4s+q4HORSA1ao8bjyYRNPC47uZ1MR9P
Ttj4qn23r75Od4rxAv1o0qp8PNH/xtljDV8PMqCMs3VZVm8fBr+WrMGI55f3TU3ANilo42Cce1LA
R+7lLxLhxq2aoHoUOqWtjHHZoXYF8Mp13UUobYJ3g+6GbuJNCmCO/NUhAxYAvUgAdUkCWhUkvbE8
xakcNg4IE8GzkzRZqnDQ2IiQF23e8WjBeEjUKAYp0lQErX3dl6fr2tpdBJasNyXttp64NIZySXv7
/2VnF6TA/oSRxD5yfnCu5byRm+r8xXucpa7fPFLVmdXrw1TM8inQgTrMuet6OwtqlWETHqEcROK1
Fy30wV2fMSxLddiNbkP2IYCXCSihwju1ru/xD0AtHDytWzw1YGzaJFoubk0MrX59k0Tzx63w1NlE
LOxNt+J4Rn3jY+UdIiyhvF37oD0CtS4Fok+sBM+VHzbWKrv2cH+yR9ktRr+gYwN1g0N0Ek2nBAjY
FStOzcUbsDX4nxq3pyg/LKPJShGzM2s2iZwk/UPcPBfp3g/579/zRIpDhlEMaIMyWusJ0emvLJaU
W1WWjZVMfGEz5hd+o7Aeq33BBAR57DheKyQQQT7f/94I5APaCZFWgXMnJUrkK3a8YzR8+yrhvcW+
CLLAlNbk+k4XMPSj7Ssn/9QHtnlhL5pfjzLN6pJGrL6sFup5a4+kWmBBKSxTf2gIVYJLhXpijgEQ
IxXnolbY3riKsQEWbjGkFrJ21og2mLfWY17/CpsZZSLZkK7m+mgcFMwrx62kdz++H23KMT8gwY4E
6U+PtGB3UE/0YKONNBveCQW1IrBDhFsIsaqdk7IxOj8ZWmpZHwJFZrAgvrmBzd9++OFdaYWAZp+c
erZRVdoJNTrYrN/nq87D8LTSaii7bQIMeO+rWd5RaMa50NQpyC9UJQu1/oIUIuPQ+0WBhjSA0PQg
OSh0C45Ty8DRVwTqB5u9gNk9ojIusPsqZfQEH/6hLg38tWA4QDZUXwrnD3gKxVWbDlAuPib5/Iec
mqXoEhgk8KMsHXra3O5YBq0OEGIbuQp2BrlKBbF8bruFOPNeffvhQOH1PNewhesxZohNycLYIf1l
LZdH8Ss1C8U5Xi95W6MKTkuCnbHtGGgad2Rfqbr/P2M1mTvjT6AibmLuLDU+LkxweDQzo3DDI/my
Ru6Am5TfmGGS2K8hZzKJTD9V3H60xtJpNEfYamYXWLQ0CVccW8Etl96cKIicYvQ/ea0AdbcabVxq
ym4DwNdJTr/q5CbpQ5cgURQopi+/Nq4vTr51+Nm2WxEDxCCVDXSGm3pLfT3ZoHMK6ehF/HrliZ80
5X7kvYNucF0sbb/1iJaSu+cfd5wNbnMTm5/CTl+qcBNY0fJv7nIliQmb5kLEyxnRAZau85e+wVmf
jpt4674KSp/mJgu8p1L0ccoUcIzGfTIEPTbhcVC7spXmhk7UBtNvCGQacFllpc687Sxj2A+wCo9Z
jh2jf0N6mI/Kb4qHK7OgSDSmKK0WgDtO+aGAyhW8t6nbRrqsC8MqqXWOdpCXbek7+uiekuWbs35D
GvIxbbt0X37vSN3iag+OizAQ8GlmdPKsxE1kjRN9cg1r2ZuexYSFjSTpssWDWsyhrDB2mS5ZQ9NS
6rBPb8OVtTzzRwJdB5D7M/bjVNlyP3GdCGjFRnLZpihTp7mtvVw397gII+vjvQK4aDdHJpbx4jXT
YQnvAg5f8IYFcCPmXlxkog5E4nUv795kGhcm+eduMUDTnpVgu6c56yab+yo1j1kQhR27bcWBjeev
OKPl7LgYex1qUdmPEfJONAOLNHlR3pHHEkF0IWpEuPJ/afYyvYwT+yLKwY9Qy6PRFAgt0cwqCwCU
XeW4JEDjg0gh3Oup+imrL/FRbbGkIWLN155YCf7EKD0mY3hqsDfNOXWFmj0GZFiMS8XAI3s1BsIV
JMQZg1AQUUknPqF7j4BdIpMjVC4p5NeH2EaHH9M40wLY/poA9zFCdOJZI5PE0RX4vWzSPu/TXI0Y
CoxJxhctCfrtwP9KqeufpJbHbib5qmpF8hMXHN6m44//lp4sKHbEZ3vAV9hI67K7cs7bOdaavnqH
F6P40yUKKwMNInQYqWtAVzJ1tdmKzCdyByGkwr7ZgCkxQafWxEhbiMq23UGTB8Khmp7Y5EpQRSWx
eg72OO3bR1aFs55AT950ApshdnMrLoF0fgDi5gCTZFWruucbQ7Mel+NRCi6N69OAVQPi+6WRLazz
oKiygkOMQtTqFpSvPh8OrjVP5RHc1yTqB902R+UQrCp3OjOSvP/EbfTPkHH0HcNqfkHFL3LxVjN6
hJtlLiO+kRj6AZhoMCSIW9smbw0x2VUAiohx4aP5w+frGHATzHbo0hiX7c59V4YS2K6ccOcIgQpY
oPTLZb7Oz+TLB3nY9h2mX3aI5hLQIs8OdYTC1LJWWE+eXpIAp3ZW8sTnD+lE1ZqCUVpFD22pK2Hj
eEQrjYllOqAcKa6dCq9wTsQMeHghF6dI0eVaolhdMNxXxnkoPoVe7GMJn/2AOh8qbwujkxV0+NMC
i18PRm7VoyW5UsGuIDEtK2uD5UxRLpB1l/yF/3EnL7wDZfjq9Usmua2iIprALxy8Pw+zvZ2nUWkg
++Tio8IGienWTU3kjoIu5UUz2usQSxqL1RSuM+DMfky/kBjLsaBlr8g0hwlhg1ZIgfM7FsifjC+H
eflaikXMFaVYxTGXdYQFpHqTmWxgLlPS1fpsOxvbiGq7UH3/StAcYuoWl38RxgFAK2PANHdP7+8d
tHLao1N+wOVEWblG5eq9JWmPCXjRzU8tG4xhWm8fM6Wk+8E4g5Oq9C1ypETrCf9zYxiSsX1FgCfx
VAw0h5RhhMErxqpHGMXbfzl442Ae9DkUKeEeID0kNkfN8ur8mnuoBIUAbhKl9GCuMLLl8GDdc/aT
K7a8zrwYXknYYzEtWnuw28u9KAEqJ82OGwgOONlQ/ovU55j1vg6MjW9HVZ/VErERtGYpD3adooh3
qug3wxQjnsRnAj7kOxSOsB4eHc2gylU5quwzItpQ9vPs+Ubr6YYBfE7iL9wKWsq63IhjxxIT32tC
3FI2kiDr8st8aZlSqIFhQlInhmmZKmtda2PYLpY376CsPBCR1j7DkWw/bcSQ8WVo+3WcQ9pslXI1
8BF/hNwGhpKBLtYNp63NRlUgc+UWiTcSYrJJND+FXT4YANMMBBDEP++n9xCrESn+uUPGRKk0x1iP
7oK9McMo9luFga7OreqQU8gMFjSVxqTBZpif6mC4j4J85SbB/YLhZjggEtGGI1ddWAopSGAspPFJ
95bQ7E7l60d/a2PGML15JZgo2paTGT2FfGCpVh1OMy/XhFV+M/KfkBrgFDVpUy2VNbzONaiagBux
gOU+Aa6oBhUZxtdJlIAvxIagCcxLjp7GNtHapmmrknXH9NNioCwtMPmNckvln2L44jBOWR6gzF0b
fgAJ63mzcz1qMS8rux48QddFxmBHxN+wO2oWKqDZ9Z/JV+ayAZRxU9bDbOFWtbAXFiT/DQ1//Ut4
Lkw7BPevSLTANNUvJP9T/p8IjM5+Z5MaetqqU4D51+exBaAcya5nq3dEgu8E/euoP5Nkpaa/AjqM
iO5U205aGVoJART6e936wxVKiiB0GPs2eHi1myVyFHlRNxpNTYDqWogpq8ox4S7mgFDIJUl51S2j
JK8/k2XHwL+DJMskLM8MSDZSmTLTPlk6gCabF0TarvDBJDNfARmFXce/0hXDrAr3RhwC4fv1YHfW
mmEz+7uo7YJ8xJsAFpiJEwIBnIMXE/V7AqpSIAYHlLr/UvKrC4D2scrZmV7fEsp+LRv5Qed4hpRE
RiaqFaAZwvHJCYTkQQ+lETkMIWE8eh8NyUsLCmRyMI9wuzS1fHYGPHWPS1Il5QvowKg5U65/jJA9
b7zB3j73uxKhuiTHJa0wUj/JLFyEbiOqO0RlG/JIKtospLjNn90rvmjtSoclt1jT2Ctk1O6N6YCR
M+HNRdEtljCo4zryaLm/gsIoU1U5oXKKHFf3pw8QHd9QEW0gMWLH0y4epvyi8+Mtm9MyObel6YMu
TlfdqvG3VYONjPXpeaLVW5dTyTbrWakBd/ZxmO1XnMbXhvP7Xl2fV3e/9CGxIV12uK03h10MwHm3
H7ePj9as7a5orZGEC++uUQQ7U+YCtiKgVPkZlwg2J+z1JHi19urNgKYJHFDxZZAzsq8+HSK2QSBv
Mpp7O+Kj2+e+wKa8RbKX8gwAlN39NQxVv9O2Z2+ZGHePgccmxnbYKt+o9VPF5dykntz/8eLQjxsf
cFeuUuIxQdo9PnKNDuec1c6fHqaezRuuOBXS3euqogvHS8y3cFJkiD1CuUqf57vO5hAr5h/TevjH
Y19mBFeQpHsxhMSCsnbiw4ngyvWe8vbHvPHQ0vONldDPtqzkl2E4H7rP8Z13IIoeBF8mwP/nSmcw
ZtDW+Qxc9m2FyRNfql1f0l1aPkphWSnYgsRsaL2X4M1XW7bCeQzYs1gnUdsfhQ7JprIM331lYdaU
r4Wu2SHumyLNKIaT0CPC5sTykD/xUe5PRn7ORV85dcISsDZ6Jn2/sxPjSwNPAod4a3GTuAMnxO0y
hraJKfRuvPddMUO29U1Ne/URcJQYBkqswiETi14T7LCFj5A6XclWm2/mS9G1eDBMDe5Ubb4Sd3jL
TSeAowhCZjstKsf3V0VTW2HfkkvuzGN6YQ0tEIhsgl4DPJfePNjjHLPID5xlw86sr6DuFK8rLoSs
aKn+YAE2xwKlyM/Lzoen18MXeBCWpGyanb1dBx/1vW/4+gEkDh8VlbD4LsibJjRfnzdhGz/QBar4
F+dZVMYwgPZb4ynniK6tQBS+/DB7VRl5JYz/mAG2z7f4dBQp6OhvzOjCOVr2DRsYHDnsTjLDuxzY
t3nrFyKfHEEZzz/muRQ0cQdCW5Xy1pVp48+0LndP9RCjM+QbGNW/AlvTB/SmZalBVyp/N5b4B2je
0z75lGEBpdi3gGyUEu6m7nfdQ/1Lp/w9MtqsX4RuSGwtD1WQHgYfgACjAasmG2Rb5M9PxGPvYUh9
N6NYr3dCR2hc20x8wB42nydVZ2MmZtkBgn+ovBGhizJBDuY2hVOx70m8hmRrW5nvYh7nZdw58LQO
b6ockDuGk8tzAi0PZULvirj6sByZRr5GurmgCItHUvFkjvYXC1OPAJPR8PciSJ9HCmWi+gnwdFaO
JE6v6Ljyd1OUxZgA2Z74junFGN1PO57nTFol3+gXuEe4Md1tBHqwbVQhnF0HQt/9YVAi8SyW7c4T
jU+TaKe5D0unPMPNjsMd2OyIOUKsRBjvXVGy96DCwuXXAseKVaX7EjScfKV5TgukBshJ53EeeMUI
m3+v8V/i3Xkmg4eqzF9Gt0Iufl7abEYsETCMiVTHAhEIGiDCQbC93gNlmaAr/gvIzc6wFt7o0Oam
5B/kasFYXT/6AU741p7N1lT1ZSFPbwf6RAOGZ0pnfkkHWGTn9z+edHnwKC+MnPZfcaZslwfWy2wo
cGR+HDpqtz7p9FB4YY8KpUJu7MQuKI0LoNOl5rOqmV2HBvabX4v1u1KKqVUZf+UglY5IraFvt/3y
kQI9i4/NX342dzuXY/xOXHENylbLFLsixJdv5wfYOUHpRdGOcSjlZlTIXH0g521l4k6nYBwPtUCd
UkRonxALoU40sCgmXI7C606PcQ7H5h2Pnid5yCrx13bDGV7yj0gt22gHWsTYJVfrFjc9NPfdFhQr
I8D/SOyhX5735nozgG8cpblSetaahpWg2JSUq025qxee4cFn8c6vk5XUXJG5XuT12DLdjS1mu/4q
ZGfzeuMEakcjISgCVh99+P2aWbZM1J60TxMgXcLqiiyju8NsQhdP5dF7rcr65GNrwOr0ZXVuiy95
YgAwUaBdaKMvE/IEDsjamPNmjS3CiR1osKJKSHPx24CCo4WykZKrMrqADRnVhNNPwGDf0fCF3M2/
0GdT10oSuOU3fTgz5p8SuLVmgoztVOl2SgPtMnjBgiDBG4mkyxRs0qGFBdoLzalASnpaOWQzyW8V
03Gandsnae3CZEpMkfEQ+jYeKVBCy2iQ7xM8+DAdWh5G6BQRP/FIS3IKZmGShlOs3B7k82fSl2J/
LgIcZdnb7S/Fny5hg72btQv2acdBuVECThumq9jhsGRUgoTGAllxmzGth/95Z1vKCcFwX+ahouJQ
DbQvZlauerJxOLjhIgIIEYw8BTl4GEj5xoSqvaIqMpN4QCzhEG9jj4+Cv5yH7R0CBqbSO3q3jNlR
DnlgXXLADQ3/+gKIc9539ybkR/xY/PPBB6orNOFwFFwJsO0xfb0ay1eSUiLwlriXhIiq5laT2y4e
M/VRSgia3xSPbaUactUzZeYcLIjps0oqL8UVRvHVcTNemblL1yOSDtfyE/XqsNExBTYCsi9UPZY0
bMO7HqPwaleKXJ7HRSI9QfGXTXvBYp20VtZ1hfJbq0WN8fs3/lzMTZYyiNj2Iry7o9Tq1WZK335U
NE4eJKu4ez612aBikFLQJhYw/XDbEvRm74YxXb/kBJd4TuSnVrs75l5yPkSa1IDG/j7raEAMy2nV
ONGvOm6tfHMZ3CZOaEykLOxnl/7sNGR6XioUx5vXEbK6QsxXUZJSoVWIOTr+1lsNmmCdl+wvMnUs
nwWtyu5S+TbwRNmN4YbJmh8oNwb9pad3vXVnPP0vTcoz9kdQ6TQ9GxnyUN67nO9en9qywsbKwqto
OtDNo5QBWE9nqPwjqKmXL6TnYWOij+cfVnTwq5x5xQiHH72m+40yj02IxFuo2FLryLxyBMoPGwuZ
Pp1BdE27J/ObcWL00UtqGxD4487KZbksdScDVLrmNkGk+Kbufkrfhaq5KEiELPXt4lXfFBgx9piE
yjKlQyn3kyBdP5fmOgFiDqmvoQuz6KRahtom5HLyjU5oEaR51x2suqZRcczEB+ZSPs4qhSUugNt3
kHM32ycJwvKzSMAgBbuBEuvB3CaUamsb8dofak5ii7ajAjpw4/qn4lazMzWH7UsbdzO++CbP9Wtk
FGlSZo/DoBySotjikSzg+is/YhO3ZGbeuvA82BHhWlYmNDemAxMNa0ASIKB98Hs6bRd52Ce8SHyD
OqOv4Ej/gqRtkZk1GyF9saGi4AHujJG2q98C9Q+Iic8ixlnS1Zl+S5pFiHM2C3XKH0kRfv1d1MHP
YNk4fYJkoBJNQlUBupLd1ldr07rahTsf8fnGu8qTMrN3Lzgwnt2Jxj130kfIlpwvGddx6sSepuPO
SNlxz8p8as0D6LtD0Rgh9V5noCFOtcKcdsqqwJGHiXmU56ibRGJvt7WgKx827+yZ5Zo0j6ZZm9tN
Mw3ueP3ybmNqxViG1THSMu+PQ8YN64lYUly3zlndQd2VYS2+45nN/dBZy78Y9RxvDO3ktIglph7/
yZ6nXpxpfUvJesZzVo+D/PNnsfs6CiijTCArYHYLyM9hc0+1Xri7xA+vIjJkPEAz6hqz+HZsolRt
CyfahzKreIGBQakwKCfrNill/Cb4kjQ7nDyT1kUrhRM1QVU53aojH5p/n4ExlyF2b9dIauJ7G7Sx
gREq2M/wHXzh/uZMN1c98XnBt1l8dMrfqu0X2CpACohSBDCai6+ZMb/kzcAU8/m8o2iwGXT5+DeQ
ipLVZZ4/mWC31GBnM3mbnVUkHQIpItK8MPrFpZXg8xkEqUdVXodOwNiGYE4jgGWmBiLs4qjFRuwD
/vXgIrapdFMTIkCnWplZzc9i7UB6eH8QWoD3oe6aUgut4wdZHq4wx6nYQqF9D2/w4AOp7On5cLMt
rVJkx4uRByvWF27Z/hH9iLemQb6EOZqcQYmevwJoEpN4MrrTMhWVUX1bSqtPzaZdCELemjQMw9QH
lPmzMH2+IQWdG4VMQdwBoAapkWy0ssGRnEsYU2JUVHs6iwTPK4kbwRopfVEBM+R2P9YHqIPPs6GB
mSscEz31IC//IhrKNubKvgweiXPtnZKNQGx+2QGuLhdWZcmdEoY1vG1wlVPDl1pgxr8pXnTG5MlI
liWQHujDvGmcciAjlb6Ilo3i+03nIAc6mp84sjPlxDGqsopxaarlvhlfkCqwoldsN0ddexMnKTJY
o/V9kYjaX+Fx0RwkBceGbJ5h/K12vW4TceICLWSMLOv/BqEmo47QAohoUTedPKBA0G/tx5T003x3
BWBbPGhHO6+HCFGP+JZKTMQSvudPoraVqIkbhkrC+JF4w7jx5su8qyASRLMo6NRXj4JM7F3FDYU9
KXgRjYW6uiHFFG5GT1SISlCFpWd78llde23useW65XJhHUBVQ+p0mx4zt9imf+jm6p39dtdV0b2J
7gDn3sx/OoHeIP3figgHdTerkt5bBOtDfHL1EWXpR+fbDgk7HpoBYrx5moyCdrYuz8hwx6afDZey
JZga0MCMo+4L914hldFVsbUi/4U6eB3FyprEJk6COOdWiwminJ/iBwVqZJXayCLRzsOy/i4kZNIs
k5PIL2enWAZkjrRU9s7rAaQ+MBuitYGvK7Eu9bwHsZvTG5sp6XSSncevrv5RzTWU2Mliw4lNZOLA
7BtelfZMy2x9A4Xi4L578+jUF8K9UwcSFt8Aq1PaBJZnDOumaMxslRuV6sL/0fc88/FysZyqwQL4
/EXq3L6fWGhgmkOH01Ngk6weeHRnTQ0N8G7YtlGoeZn+UXAHaWxXR1UuZdvZSAcGKY5xh7tW3Tts
UUHVaBYnmIEPtN02qidumOzaHawKX28ezW5jeWCZ+c+ononz1cxaTWGYKQk8pH9WuKnmqiXcBPgA
UOPiBwe+SwZ1mAnttQYx+vb3dfmTnTsNR+/QE0o67txa6o9r4pzwDQpvuoWeTYC1e/0WB3B0W9a0
zw6ChvFFQ9hIjJ4nkd3hZuMgnaNzo4QGz+V0yg/7xnjrDt2eHg3Hb1RpZNaDsSkg0GS8tM/Ru9ZP
HhsbEOMCdm3AaLDVk0p70jHIedga0nvDRZNv+QbFL3EHKG7+lDjgt+L6NasIAVANV4GoWsYDHTeu
+085AXYpjlXmwGeRKh8OmURn/2/UHoIx1Qv7pSueI7M/ny78hmtwqyX+oYTicpfXjsXEev0x7xlb
lTXLVO9xk7NmetMPpBPMtxYG3qkXv+hsIupKq3nrfyXc7xGqDUwHqR42lL8832KNU57SeURb6G/G
tcEXyapQT0k4rmrtlozO1089yXIxfWftjvJ4ir07uLlkvHU96lHXGA2vSPQpvYFUes2fuhuCbzUt
1U7S/aP6sX0uGXZYk4TKm0vkOTA1ktUfVhpW6lyootF7TDD/y7xznRo1Ng5xuFm9PD/n8Mc2v4Fv
fHMDdnHT/trj34jc7nd2xBdH9lBTlQd/Qsp3tpeFtX2NPPB46w9DuQo6JdTGC68xokcU77gBAKW+
7O8t19KB/oa98ZpMfNNqgznqP7NeNeVok+GURpIfuZ7pVCiPpCCFxz+R5Q15PAnzg3pXi6VCdw6U
YB8qmC8umKdJXRnvPCne6Py5ooL2MlVLVvE7bZayAgWmJaU0MhxdPOKD+AB6MGpNdmUsGEJivqVH
fZsP1TIWQdzk8kPqovZ3Zo8mQI1AdGjgdv1+iAhuzCndZuY7NrdyzOnCoMvFN531V3ep/gc1h+rg
/9b8wdpq8JbrQ+uJy7JR6qYF7OuuhPRkA7jffEFTcUxPnFwJPwqmnE/QLGgNLuahKcMUVXkWNahy
1K71/m1dUzlbjzPTbh0BR0WOxEBL2I4RoZ83SkW9Dy0TYBF3ZiuDim4OVT4mijckyucnHLXHoSmT
tDnmGgnXxxHIvQ0+MZNswyz5U89atiXdx9nydH9AaseDHJM6UHqfX9BqmWx7ELS9ban3fTLXDOjm
ncGXu60mbuKoWLhSQ59Iz5d+7GrK4OZpfoZJ5Ytmmhde/R3t3HVaaJ1GIrgS7Y1RbOEEkzSc0qNg
LpZHf3mISunK/bH+c0hVGZwN6RBASKoR2qblw8LL66eNehaBA/stLg7kwH88kXYcInoCag3Cl/cI
Zhl2OwhFm9iMoPNtc/lWBmshTD/+UGBMcBatyAQWVKTsoLyCI632Wwv3B9QLZ+hrApQ57CW8oPTB
3UJUCrTo60EtjzYY2RW5zAsOH3X+aQ+aYRu1S2uE/WoY00oxDQtpa/gUMGyI58qnT3wkFQ1KltmR
3v0cwunPZfRXN6GotSOy0c12/Dnf1GQz0g3u+e20H0RsTxx5B4jVpOnPoQTYxrq8EcX4HMFAIbhN
X4iz5B7Jwlg2IA1Pyhhk7oQLdf89fDx8ooIlBsBdva84cKGedZH2obvYx/DzPXFIWrMmy6nA8bSf
4ZjE1/Fk+TaH9tOLmGox6sxnGzeacSgQ5ccyiCK7Gf8FQmK4nviYXx49U7ejs3ySC4HKWfhmPWJN
Bs6khoL8EiBa8b8sK2VpDxNp3qs3k2c0upZUvizAfodNs0X932MS61C7lNpBRTBzxRCaCJZozFbd
7jnmiq0rSmvkBvu0M64fTlTqg+kj7CI//24s5AyMg70B4fW/xWC8mb5UmfHx80l/HpSlbQg5QWZ7
PtxkHAmcX/m0AklJPqBZoOJHD2GvaH7SW8H0ZJ9cMIhKiNJ0BryR8pQTSJBuH1BygAyFeQh9o4Vb
15aAVyR9d1w//fiSAOW6SY5oZDOlRzXjsW1RARxJh+vTknq5alUUgETNOETi3l0OO3FOHASYY7ir
iWdu357QJIcGYKeKXqkXF41qaTulw4kbUSFo1TaxwWs9oxsFuXRfD2rwhOPApagrfKWo/wJjyEqx
dgg6orl8FYKOOlA4jWYMcALCJWfJOoCL2kQvHOaNhNAj1OlOgH5B4S6+SQzfQ7Kw9haA4HtziOxx
x/0a268rrY9ofmmOXqEqRsyx9LY5Py5i4Ne+NgJzbkANndRsO8J205HzVnA5rD9hoYDqOREdqSmM
aarQlWlAf9z9YMn4xHAyf1SLXwhca8rvfi/BnDiUvhBi6Hz4+YBjkO81m7oRpld7JkStEFCfKdxd
vm2XsJ0OFP7biqIADxitBcBwpTByedDb4pwxFSkgwNvt3JwEW0WbLeC9vy0xJhN8CfYpyHs88ozM
hlrZJhL+y/HEgbAoSIx+Sg/KFNhjLp65NHEKDwuWqycqHY/kGTFYBBDWW04pRthCE1TuMPnFayyo
Xi/NDoi6X1xm0Ul26DIKdgQ1oOkZFKkXiqW2FXsT2xFrqFeUCi+MhfAal5CfEUHwtWZx/LC4HgR3
s3vfA/0y/vaisGxK3qGtNq42ARnMoq4shTvWx54kSzzHDMIjLr8KWVYcYLC6ZsFwn0dZ6fnjSTxq
VmpyOZ1OauVLlh4SflX3YggaNoqwP9V93FWTdmIFUJ5wbO08py++P597u0MT/ilGrf4fR3seQvDe
VcOOXvUEAS4YF02/WS/4vSCIag4bNJlHpTDLUwB6CxR12DE/7DhycyIf34+adkgozuU7eaHGp5s9
tFGg12GHhWALlnsGdUM75k+ydi7mWDGNhx0tyDEjPQBSmrpRumvVWt9v+UnutLcEvbNDrB6w7RTV
MzXCqxG+Jm9N16EQy8p6Pe11RwK/mGNZYM0KxHDLhRAPkCyvb873zOkK/WC4wGKDS6yp9hptrHJk
rGLgx6kgIGt4y7Hb5l4xUhc+5TElUMgz6t12DUB59UKBKF7QHF81Iz9JQQxOhSDQ3J8ia+JF7plS
XjpZdttvy84bRzQ0Xdg/Y4yJyTaRdDhrYBx5PUGiCyfm/D656bo7UKxPGSDh3KCa5iucNZaZbnxk
KEu3uF3s0aTgYmilVBVd78XrIUfHxXsYFaFYaWy0OV13DCQF/vXlMYWKzux0OzrfUc+kTnDn6yKH
FjXPz0dy9+I6l3qDk3ZO8Lc9Yonj211vYkVlaY8Rk4K64Q472T1isPL6JD4bH+G2X0/WeirzVU1e
q+rlmbuBzPmj+romAO5V1QsnlCjFKayGyZunDD9eCEJAXZU8RziismMM/nXJ/Xq3YJuIuKKlLuZq
Gpjz1dtgR+CiR5SGFW0sOrB2qZDsisgNJWZMiNzjCkNKM++GgnJ+PYwQJ+D8BcPujjNSIfEgWuBk
rJh0kaCC5W0wKPjWTV/rfKB4F+jAk9gtGEuMY0iB+DVAQL0QKXcV56zZAkteZ5lmhRrcjAJdasX6
sCblxbsHxpzpQ/M4F+1/P2TasKIwf3i2jxq36PGLOB5gC8f0q65opkqNXyjecFmhEX6TuTi8/pCw
iTHrehpzSLIjqgYhM36QZWmB20UyYT7/bsJpSlCd1PwoTNV3QSZlh2TQsl48qkdr7cpvdtUNvrw8
1uGjQguBccizwfs7fneNgpJJjOzDvMVw9KoH68sZ/Rft3fv7b4qV8Qzs4UeXdXsKgCXLi9pV74Kp
YN6TFJwAAHQ2PjtStD2XOSwDgsShwJZowTFHfi6+0APh/1r1UfGts9xjF6+VjGoJLZc7F6CEpltY
o7GUknpUlahITa7rvrmUADdmyQilwygTzpoOTbvmd+qG04dfwHzzAkc7DAAvCx/a0cDBVhTKwxCl
sUQTivXW1TgKIsNtaD8TDcvxNsdWVr7UQYJyTyl8EnML5On9HW46zoJmeu7f1Z5ShdCjq9J8j0WG
8xbTX4RjldnrUPgfrallzqwHiIlY0LFjZ/bwz7Yi8JmoqoS2GlO+D0UEHJjb8tcIpEDs2PVEFwOM
S0q1W01j/f8KCmsr0bP2MGGLxTo6Y1Nrq8aVzH4GvijfooNhoRuZfCSqGteqryiZxyCrfCjpwZqd
NBnBdmmYbIXMx+/oKAR4Qw2O3BRCQKj2IvrfJhvhQDskwP394gy1YYl0OMf9kfw66zEp83pob0f6
ta++n3OYW2RYOjCn4aFlY73QO/4ymQROenO+PWUWHAFEwZ7sl8e/sZj+Gf4toU8guSW3eUNx7bCZ
Qcp7GI2CFglgl5JeQOlKjyTr9u+m+fMVpohJ9mBbaqDY02WcvA5Q9HNZcV5Mp7eq9+UkRsqEOXjH
A+1fm9/0G8t+BPbKjutricm4Xe241DiPSQ3Zpr1jhwUfcO21Iglte9A0DZS/8iaXTMepBH0A7yJM
AbWQJCkW39+lYYstKOtt/lxNRD2rFeYDTWaxf4aM1WBvQ0+jv13wuB3UVs0wQZaiwUFfbgMzjhuf
SdPKG2ZsOVgAHfDtLvWgtmgOeFSghvjOensi7WlPxeT38t1WXGRmwt5vDRzb10ax8gwvMQwDoJ42
C3Gn0VOdYS5nAKHi31ecjlMtqBqkZk7Q7+ZQbzYCATZB1Dz6IPJmz9ZVYeJB5tcBLA62VhCiVAXS
yNJ8h9viHXQtvMNTzhnhYstLxc+bMD6f67xOMAWS4RnwFV8NQl42tyvC+e64zMMaVN0qhcdsXziR
lr0uuGSuItVYSef2BHBr2XIK1INnaWBKGu606XdDtkzQVcxmJg4eTKXnLUOu683mn9KAziqB9lWJ
WThum3wc8pBs27q9QU++3b6oq/jK1CQtwKyFph025oO/5Q3vK5ksZA8TC26Qi+lk+2Yc+y/aJKt7
5sh3wTRd4FQvBD38aRs55Kr0BSTO4ivoVliyuyDmzcWJ/xaLf3XlIP+sKAUoJrvfLg/FMNLXfNSH
2rImFkfapFokryr8YX6ctw2UM5uao/jIaov5fimbRd7tNXKWwUroIeZghUs2Tas4fD3jGC6hrr3I
IqoNnsv/dNm+9lzuqFTDdKIsTyFdyfR5OiXEIM9HAsYJ+w2enGYj/Kh6+NQZU0XqZX/q1NAZFWcx
q2MjMPM560NAgL3KUg6OnHwvp7mFPhSjv8SJ9CTkfrVyGwdjKmkf9KpKyuljZDuMQEi1yjeax2d3
yKk8Oos1v4CPcjMhB2Po2PwoZu9PSxWeyLeVXVXJplGwuoff80BJm7c51EiOEDmzjP3DrsV8+b9C
plEP4OMIHs0rTZlAOS37JAoLDeevbD4yuQKez+1VQJ7xPty0SHRP09F+oHFL1rRRyfgLYiDSyiOb
DHGV5mNGSi2hdxsy40OVlPGEzQ4ZbtaDsaJQWWhn+/r7+cqm488iY2hhWbD6gmpaNW+jgDc9F4NE
WnU14IQPABSvTH7NI1wicSMUrhZ3m5e+Pb1aNr9Vy8KYmzh84wpUoqP7mKJFSqkW44/810EFL8js
bB2WzZR4L1twddGBtiOJ1kdNZRzn+skCVNbM07fbUNujPW218fWvooSaZb/B09/I048mEashyEvR
CQ7Fi9ODebxAsnNZbMeIF25ZrFNwzaCZ1+x89DBJJr5Z0m8bDPBOhHi0cJrjbXJsWPYMtt6raGBd
qqDsLRVavScFwUwSgZtRF0EuKSYCNnh2TQXra+GLEmfsrtiYYTRhMVOafgwC1tK5gc3nE42PYi5S
Fg91ZLQhCf+Zv0vv0RWOW5v/I0qHG5cO67+q5W+ldIxZ0piqfY1trY5QQnKo+BkiWJR7r0nDYTAM
9FW9O+59NyEKmm/T5n5c2ZkeVFzwzQCauTtXEiLU7g3Nf/gV4TZC6Q3htj1Nkt/hiHLCSx29WZf2
N1CScZa8dc76wcDE7WMfQH0NsQKGsP2t8IHrBl7srljwzyqcIeyXMsIOrBsER5W4siktTor7KdVA
Zlh/owKYZlgrvTqrgx3jgEh4ANsxxq7U61+VfCMMVvMh0e5Juq9QoE5OXk5XR3958+FnLPzo1tFR
+QR2kUrwgNmspH/S7xVxOJZdU3UwKOAxUkD/N/PlZeoqZM32wF2Yhp7JLVJrOe4+irJfhZfo1kV4
cRaV5qgPAUSpVeWQ8SdXf92k9jWI8+LnTSeKK79LGVKMp0+e43PR5LVO5VvIGKvr1flL+yPS+8Hx
hQHU7rvnsplZlNIo8nAES+h+PzLfYF+PwPZe8hY32nqq9afYMShfrEoaa2Ozqnk9enACc/hILItf
ot5tWP9tTfhnTXt/eQapkv0wxfP9k8J4ue9k5Nc76qhPdsWAbvJnzlwcgj8ehQByiqkrYB4PIdV+
4pF9mkkGrxL2NJg3fEQ45QYo7Swoi66U75Y49GDt94F/NkCxAsxL1KC65YQmLtxykanDspDMRkkm
3cy8LH79YtUkIxVuvHK6YLQ46kMGgIDcKZ5NkM72/uU4xQPTJJL3ix/hX+IWX80a5O4YxS4COnl2
XXZFFCVgWw8pNqty3Ah4r/k9zq8JzjLdXt0SDFhS4xRFV5UDJFYHcNL166e4eUHzXQ+vEDW70o4t
DfaN/19hcO/R0MtzkYD716xcs2+zTuXqQ9jEk4V+KEcQfq4oOuoNiUHbrnqHzZAypFafoAx+WEg1
HggBBPVLGkEtkTJLiUoDhEu7HNTQxsHbhvlmcjftCz4Z0IpfEg6FaJnuSsIWpSj79qZuQ2jmuqdQ
m4HXVar3gSUvLfQkbXAFfW0t+J2J2VcFLFhospQIyJK4wznWnwH1GWw2dqeGwmB0HbJ0++Urmy4W
u6pIKr+WekhoiQfnq9PNE4jaKVuJLifR8uiGQA6P1GebM3c5HygpivkhugdzVA61b61pAubPYtAj
7HgJqrFat2j692JE20Kzj3lGz6Bzmou3tH4DCGf8LkoyD20fTVQR6XJhMt4WcgRJLLSHZ7ralYTz
c24Ik0rupQoOv7HHM13l6wtQmk3e6wIRmPaAIujf+ay+2jqPUId557v3wCP0tivQ7/D26FhcaJU1
FxuxeUW/CNzZbF1ZgKay2dpDJRuAQQivjP0l+XagCG2XVN7wvlakwT90AEw8CiRaZMMnGjDo9puj
+AluyV35Wt04IQUY/EB4WtvaytQHBk2PCfTD/n+9yJWjG9bvhV3fP/g1R75Eyq97UIc+MRPxSVFo
En2YaeRoQ+OCu/FJJgGDZf7DA6Nqyc3uInBVthJ+uvcoYtRgrkk/IWmVZdnECaaoEPSXSTk/b/b8
SPjGuq0ESag/RD0AKewCmZC9OKFwi+rJz3mE8l3YtIv/xfoU497NrQ4oRDSRPB3dhxw7fBL+GZdZ
jiLMZSDtI1nluEzexSN1D6bM71wFl6u6rjZZt/P92vINHbgGSR4W8oQRcNV/rHpOXEK5SVZ2t2ON
6c2uWseAH7AcuQSoBhuyeq4hZchqbstkBUDkaeN1+KPJxdSwQ8ZO1axbobJZvjAN1TWvi3I2k9nY
lmBED3hVb7M9kM1k/uKJ8ZOeRth1RCpmFQJ55DBJKtkdOkRX0hMridG2zvxi0GC8uXJ90IGXqmUX
jwXI50mW1JVd9ub4NQEw2lKLbUN2o9ucuUxNT2Sdj0MYf/pi98AOEVH20TxHtkF3DBpR/ZyPZB8F
1ZiPfqZSBFtuhCXkvh4eJsLcusr0GAXPaThhN5M697L7+hf2IEpRD5XXzPyb6hp+x8HlRdJFGKnm
XZMlhWzaGeLfM1o4C7UZ3NqSDvnRxvZtLujpf8O93T7TftS710G32C+LO+eUkqg0xzpntf1p4CZh
ov8b0cILrGhHTkJlozX2hIIgJ3hC2JfuxNxX23iTVbR+BxZX2y1ptFqcWBq5Cn3B5IPjct1SgyQN
L4XiDDNcn+Ip3bVnQOo39PJoGfphqof/hVZLVBB2u/yYyKSb7TSIDKC6vsDtF7mkt3Gq7rURm1HR
o9U/FQM5OvZyFFTn6fqJp83ak6bicjQgSirV9qGnJqrqX8nCugIrUIbBJTWsXF6Tp/c6rSSK3dmF
dgK+OsyrThsHg2ehLXbYCZ9wUgafhD+/vVK4hf+LkEj/FnGOePvuYlHvQFXgYR6B92eyKDLq2Idg
25Q7tAkZprCQmpCQ9p7xmmCXn7gaRqDSAjntD0yx/EM36hWMsJaH0E5tE79jlaj0+fV9dVu8xk8f
RNeEZwlA8yIlAzOFdH9Tw3hwcSfboBjAVCvcJxHpv0BD0oN9ceTfzu2xBDsoIgQefoL6rVhHNprI
TAu0Hp1661XoCXQyCKjA8DUNqW3uZJCuGLTu3x8a836qPYT35OYShV1P5o+pxQ3etBp7dpU6xTT1
rF1bhS1BxYECWCHqAhbOnQCbI8bQWqdBD2t751FZ56tGDlRHIamiFPc3zZxiZjCSRo1Q99s8t05T
j2ViGKjJnom2PJG6BM5xA5bCRfd7uS1IaYlSq046aeQfAdaxSXHDrlFaJX0iAiID7oCAaut2waLO
LtuA87ELc517Ej/TKvkSVJ5XVq25sFti77PLNANufWf1cxH0LCrkcqPk+JMA+xj8OOTUdGVLNA4w
3xY4dLLGSvpSWfLkZsFNRgwpxxEsQo39btN+J2M//SpDLYNfD2u4E4h5T4tHrnH+Do7XWTbY/rVv
ZPgaYRh7ZtpaEoWVW8kZEdxuSMGlGtlt00IEzzuGkFDzdkQkjgQym4mZFPcpNGXMfre41XlgH3DL
suxUv3epfw+7QPVo7FovdkRGY49RfhoFJbmO+mbp2NDvXOUmMuVM7S+XCg5qqlvDMc49RuhH6YBQ
TghQAPJ5Y4nC1+prD3cWWqlxMyUKV6vALpzBGFAJgcsP/5Jz2whcRlNF8EKn71muL29kQKhkzKUt
2IXKJEgxiS5RJEu2zko51mhCvmv4h5n3t3i/x4DCMcYS7rlRY9IDwjaBxfwfGyVE4D/QQpes4XEn
J7bS7kQiyYdXf5WQ7a4QHNGHtNJudI1BJZ/DYR77GWPEZSxKSW/FmGfYLIehHdM5s8SsmRThV0jM
t1GXFwj3y3XzO3ulqioc6leRm4qME0I3kGWcMeA+HBv6zUQHWJanH1nQJ10F5j9fkLxHUf+QIHyI
oql4PN/Ym0PQduHxfCsFjak7iYIU1K4ymioF5sVaBvWt6xt9xrnaPlYjtd8NeoJCRRB0w0qFsFZY
WCucBCWvLd49EIsavc2OQ7UWif+QyrER7inn5MXjpoIxTzKJaRNn4Aqnisj2OaHP3hrDPTSmoj1Z
/dSj+gpWGfrMjKNAzca05aOnv2s69s4IYZ28UPLuBtwptWyXfI2fwRZtN+eXzS/GB/x5p67J1EbP
y1NomqaMPD1RFNbPPATyYRcaUivSnbffevIMan+NHLISDVtfGFZi/YW597IT0ZXaIDLUbCE9mNJb
xYTQa1YBsC9nwtVvUbrT/kn2DLoSUaPmAx6cdL2A0vwRXPa8WgXHEJhKaNR6H8XEEWNe6SDqXuta
wg9gqG05CnhJvZJZ8UOxJxIVFEmW/2WUdFxMciBRp2OA7lVjYab7bovCUpxMdaXkYGvxquDrZU24
EO7dY/ePPQ63wUZybTnR3tmjPDKHLABaNkKmg/IVqblpEsjJ0B0uUxtyyanuRdRB41y0uCoj910S
uJt/pV6wLjKx9qPVfpKMSMF25rgrWTIVP5MzjLgRBMGrNv9I5pVSZmRR8NQb7QADtZpafe0/Kiv8
47JEq6spehtmQGujebM/5NikMGW3/5o0FUKi3SOaR3AikTWdXDBdLIZKGxWokNwsmaOAoTBf6Pe/
3ZwLdvMZLIqfrXlJjqqbGRrQ0OQVON2BcvPjPIlYo4clpxTEVkZeoE4BqGY5BaBlAV9YxdbC4cv9
tY2b2cINcpAmTM+Z02H0GgvFdxgXJXIaDIpdYQfwJc7C5AXDHWdFUw8Hg20bhXyx9lO6//EvDvy0
h5HKFjoUx/Pi6Brlg/saiw7GJUIGlq0G+l7bB71d3iWb5s7w68tXebAL5tUkW5ygrFqr1D69f7vK
AyYFflbQtsvDdC52XGOoMGa+5ZDi2FcN1fUEQB0rVBw+pUocNxY35BgheYdKsd7ri/PxVfNVVwUZ
8QK+Pm3OOQi5ZupO/ehDRPiclaRZfd309KfYe0iDmhGy5mlyq5+twDxCiMn4b0bMogbvb9G7AFWz
uMOPTTCmfh92aOjnVEt2Lk99pmUJBpYADnz7yT7Ma6mUBscDLcwPMnEseGP01UkUM63X9sewWSp+
NPhIi774q5JHfQzRpEFLZiOAfw9/dGtFD2n6dwFmma2VdTNXukByD1dxp+zv2kXGkFGrXyEAv93x
9FuxQftdGMy5xA6wLg9JTzAT+uscg/d7nbCPvUe8Nz1W8zNK/lS5x6Ypte23aWt1NLplSMY//9l+
b9iDoqoVqo/Alq7RmEa9VYJWqGw0PxrEZ4eS3L6QwXejwHiUg02i5dFrkn94R8I8Mb47K+QwNIBa
k0oplvAHUpwF2a7dz9Ok+fdZCR8i9El0NW+YKoWZHYLNZD/0oH+BsE/s3bNXEEa3wYbKwcL2r6lW
lk8GgO3UQMwloHAzE0+qJOlGeS4d0LOd0yotOdRgLT+DduiPRb4IyRK7pRtEI1hXObi8sbhb1xrZ
i+IfaCarzeKYwWzxeiybdsN27TrlfIIXEIlNWUVYKskTypr7v2NOeTgreCuY7gzxkZVVuz3orRxB
ApjwcKPGk4eZ4rW++Cv6YJOKiwWVqw4QOQrggLJMIuCkG/VIGl+REJy0/GkQ/1xtE6G8HpUGUYWx
jeEv+/eV3Jn1yfDUEud666qiAyCizr7sM0fFdnfqntfhGdyhXVl4Fo4OutmoCfgeNsAv0AKU4CYm
egXp0h8RlofxgLh+ugCkTyxJU562jysQRWAX9cuwH0Buf0DgdCrxnrK28stZ5Oz8/MayjRc4JMKM
9W0VxDqwIWD9UsIhF08hVZiZ3CSLdrgm1zzdER3SLNZwuCYVHYwLTk19jFXWZbQHwPPyrCDz7GUO
mebDBLecrXw8dq96y40V0AOdvQmQsGclaos7he1x315jlbqFjbVn3FbwjT9P/9v4Bd/UFqsFyeto
j8pfbAuPnfnTIp4GRGcVC3N2EQ52AE30vXx32u4t+P9obkH14d0nBa4+JEEJrUIfGWwA7vQQ33Y8
x4nNunXo0tXIAowBcu7F9ZEAg5QS4dKExVH23stKqUca3sAVeKBKovZpzP4FXAL5GH86mM0vD4ja
izeRCzJWYJZ1vO6WmCbYZD66r954Z0fCXz5BTtZqtElw7b9/DAyXHIo4aKnqA5BMY4ABJPQ+d3Dt
xTnNr6Nx8r1RchkYbfODdfBTLOhW+58o9dHNXjX2L3p4qVopHJf2qsm5RXRBzliVxWKtJIW3qq57
U84huxjLoeuqZ5xSWJi8kYd7QSUMf56wnPGzoiom62jedSQztvNd4St18FsEgzA7C87FXAERAee1
TJc3TM0PmcowXQ4IA/fb5k+/6A4Tf0ap4Dbmc9wIC7YnjdxKi0E2hgd3ApgZva2FLoKPm6XmCGiF
IgoVLAvM6Lt9j1EGD0rmrF6x/GAYOisKBt6vhaxLCApWPTYLuVUkgF5of8yRb/0wnWvIoUKl4etS
qbOUZ2PniR1zBfqwXqlK6ivoUOKHeTKR+xPWLr2y4HI6KBVpW8HqLcy6SjYFXqpgsamx00xZGpxK
96fg9ysUJhK1s5pWZvlfzEKDWdLub3IFrHJ2eb5xfMDu7Lsqo0fX/pn9A4chHyy2NV3hw2WWLF/N
YhgCd2lkBSDr/bAVP+sfXZwd/SQABpslYkSZ4ewK7YV32Phu4UbUiK7vEHnTwl6UjvweChfUB7Dd
6bMtG4mpuc/G/0QjLeK+OeSBC7c0Uusy8Q5sm39Oj1CynsaRCJa3uCFGHT8oA7ZAm1FDUc2CM4Jo
Kebd7wgcKX88Kx+11ew3ZBIotGt6gMBIrIQk/NEK9NEMMt9iBkOINxlBgIUQBmekvftkhof8j0rU
yUx2egMORQ1NIT6TMo+6u1Uv9uCQive710+GpCg1Xaiu2yy1Z15KDN9M2y/E+lvn2N0BV6QUx963
IXspmSS4PI8AJmlwic9vBkaxGv4SSUJlxcofNMLVwL7Ou6VXjb4yvHkReIA9g/LRFjsk0T5e/8nf
DYbTEfFq/gxpNTSmgKs6H9YTuJimClrePk0+FpD7zyeCBNaT3u3vYOT/qdLbzVsd98BtL4eyQjTE
c91cBToQTUZOKjALFxz+CkFmhmmaN0Bz96oZWv+G7qJ8LHXhCX8P2JX8FbyoEQNJcUf3H4boUBq+
jrIwQ/DJDFsWMnJ4OPZ/7/YxFGB1qk3Mu9BV5UdhHVWqnZ86S65VIDvEXq5Ec3B1ODPFs8p4QjGg
gcf51e1UUlEfBiJ8f5kR7ScH3gIz04pW3OpUJui/4296BdXop6An8prybkc2esfFnrhad392TzZH
umwj52c3skSY1e3LqLhqs2ThGmSSs2WaOfGgNRz56W7P9OMyKl2vcaO6y7WsHn8PN1qhJZmv/cCw
25plWKRfG1O/U+WWPl3jtyb2q9auzh92HA26llNCiaR9JBVWRdiAfLiOOUZVnn5hPAP7SYE2QWSp
bCraPpgMQ2TqaPGUfVoFHg09dvvNTUn7gPHQ/cHBx591ZGvAZlmGDu0+JyLTvjVRua4n8k6+wNxZ
ytbnYzAuSf1qnT7iQFgWsydxuGpLdLJXXUdqxHlZkmPnBsjZwISzfBQwV+TQ0+eyHbXAlaJVqL8L
P2LsMFl5O4YTF67pBVVPjZEXa4JMULLuiUGl5CBXOUlCg79tQefBethePf6iDnbXl2TxyIqdNz6v
ehXtQktYEyhCR+06qYtgT9gD5YyfzDkIeAPoUYXW+MlTRIaOEb/z6PUijCqUyyg1UALi9AgeKSgq
dTO7gMlDNWylfMVBz0AvHq6Xifv77adr6GpxPDaGEAOujAaGc31J9Mupb7n0nwQ2GRgOFoCmFONN
dA7mk6VGjz1YsDPgtOM+BBgJLSE93Rawjva7G7bKetTPYIrJ2al4kjTyfy1QdY4qZkfuG7yluEva
T6RPCg7IGGYjQHN6vanMiB/7zRtyG4LCZkRSj+5k4otR/Mgx6tUo+wPJnQevze5BKksUdaMyeyEu
CgqlxNym4j1TWLmkr/a3BRjTsc/CLYL9TRfQrSGCzPQarJRVjNaWURrV2BuBOt1DryKVkmNXxz75
XBiX6JeViVdZjOLUDw4hsWBsoPk0Cc4hw4XOeIibv6V+zfH9WXaGupwnKwJ2N4TAKjt7KOmsQAGJ
HNBmBM3UzSRt82LCXOt6QP0QUuybOyEfwthiBp2PKg3wUJtHEhI7bWXZNONEcBEqAqm1MrwpLqa3
aFvdJZOuM9LiTqFdg9tZ3tTszh1pPv8iShI+XclCMajtDSrGZDnO4BHNEDp+Ym0ZlWunt/vsjAZy
rUyO/JL8RNLLzvxQT6jjjOYH153BfXA/x7okLqpQ1pQhHeS3rUXpp9S8Fccq2/AEKEQ0U2CZ12kK
5RU852nJdxY1Xdzr+3Nr3YMAsZ4zGvCjvcP8bzh8uCYO7RaTzRflq68sQBQKSnu1mudoa4jOQzid
+V72NEzHr553dxPYnm0KhY1FZRBzb7/2Nyt3LZ2BI3sTJWV9Tvn/d4beYw0VQlccoj5NZcU823Sy
HniniFK2GW8klyqDaujBvZFmrsJg6WGmxUyuJkU+Skym801pQageYmdDIoORbCZLtBlhE9Tj3sD4
1MnFtNRbtz+iPUEGQWTAysqgnsGdKVWdiYlSiZ0CKIEAGLCNTb/+YOCkCQlixUIh26Y1AbcJIor4
teXYoveCw1VlWKWJH5zvdUNVci9VEube2jQslK8h69tfTjuxpmPrF6+D6W+Un0QmU0HEoqYPesKK
8q7su4ykwQIEww5p62PQBE12KZFFZbYrChyoVPgy90JTFeqV+SDr/VfUJRsMtis+LK1kh0XDV7Q5
oui3B7wtylamAxXHFbajS+fV0gkODZuHF/XoN2Gr4SN+OK5gRDagJmH+QO8TnCJVcXfKurlKe9bs
M7fF3FjmvtSm77e1gXF3CaZ4vyPex4SwAXIcMYB0HtYfBufioWPvZsy7U7QU3npDuua8d4q4+NNZ
41pDLl5wDXPNqn5Bc/0vu5tpzapq3HNokgW/sRCvTp2R6jc2oyKj1zuKPIebcoNjpW3Ntj5EXBlN
lcLbdIgNyjIkPr6Tc0+5S0T9XYMR565jh3r2RobJ2l5FL93L9JmuFLRH6rPg4fKwpXKu4x+i1l25
UF50DDEAaWQtN52Qx5q/ULPufiBHmflcHxq80CCk9YN8YjZVvoBKNLTiLo9szuzf0kF8sbgPBefd
wTlVKMQyAb5DwKKzkbNkB500hyaI9qsUEp6LBQ9r/s0xhyAOhkKNcbd0PqzHFM7AYS0mbQdLk+0o
VCZsWLdLeVsbAR1c8N126vv02KE0p67eGCq125xRdnQn04GFVphHSYqjGR88r7tUgWFvwBPKDaQx
UgHiYRhptnQGtPKUpJa3soqXLCrhxP2G4zO9RLg8wPEh36/AUmb+6zMbRcPXkZWm7CRhycGifaYp
y8jN8lCfepxYtnltJzNe6e/syMifiMVPcjhHmMFxd7XLH+hjoGqQPsqHn8mpkFBtcQ9aTMRb2P6o
UMfdoe5yXfv9qnptrHCgCHlQ9pqc3Q+i/u8rHz8gdzO+qI8haOngHUhfNE/7aXpJuO88rvy8bY+V
gxI9epu72CYhBmFoqjlM5LxgDwa5ekgAseJbxfXNHQ6TaDgI2ClQy/lrN4K0VdD19LfdMopmEMJZ
O4aBFlmj4MP/hMxHjWyZDJIqvl6gH4Ne++zXUNrkc5nfcC66MXBk9jfr62tPtCgoitczQzVClK7x
L5HQrif6uDimStTXviz2PZtLOIO7zs1Lw49NtZNBR7cbbkh98h5TXaNLs7xsl2+HokD5uBXqWYcR
H8bTDOTFptxO5qga2WjpSDjAjewzE8T0bxR5qMyZ8lrNSl2bA1akEV/1BreRJijBqzWao7yG7jAz
XALoltI5CSHYKX4q0+C6qc3MYPY6i0tArlq4hbpmETrDWGJqVeudPdYImcc+w6bBFNrYklzmS16Y
zcmkF1SrbBoMROZ/sIliVFdS5wsdBzx9Ne2N9J1h7N5ySvgXzMMOvywbWa8vyY0ncSJtsLQH4CRc
3IMsEJu/XnQBSPe4j8kJ4NOorxnyJUj4Pb5tZdD1OTt6fG2QBO8eUZ5My2RErdGuqN9YR19ppncH
7jb1b2FUFZRDa1NzhVSSl4zd9ZIU5rBblhWUrqZq2l5VpGP/9FqcCq++W29GAyjvxIGffMaN8pKe
G0AFZhC19OkMidjTmPXRAU5Kyrrug5cJT9jGeV3n7VwKv/JvK812jh+qim1ISopx3heRvBMW7NtU
nnaQ7yZ2ZTKRQWwo4dtKUy7ywqQ7DGn8+sRZqBb+kR94tSlMcWgYaCWqpTSkofAQjqUjcu1nhjgz
YvDLr1YADUZKgKpfbH5dM7DeTA0wj60bVrvF+ttauBAGyXNcmxO7bwZWGLLYs5Jsuc6zrbYeZm+w
dPUyDf6HmoAtbIUi70GmqIc64ecJ3KdtydosJbH7SZ6rESyRbXoscYB2cyACl3KdFWb4qV/YFcdg
pXdXGd4s6GxYneCFCIkLqiUCEae0OaVKWCJdr9F4krigKb/BucimJmL5mBwp5al9YwBLMTWMRAmf
Tgvlvk7SDEDjH0OnoCfdAoFN6nWSAPYmRDMICIU+25Dr/CUhPo/b947C1rACwKzBBK2bnbpzL7Bg
o2h4oiEMzg4qdE8vZxlDfN+2m8nmtIkKtizKeRsS9KbDMwd65P2qDz4CTXSw30Pa5EbbBDhfHaWI
8RWPybM2rcFC8ehEE56jjQCdoI6lR+S6IB4aIoihyzgtuNR0CgR5BbE09aOR3KTve6OS9MaWZJOD
qnfc/RycehFr/XRJwgdavUR2/B2p7GFu3pkbP5cNr7MOmraZz069TtMR6bYajTUl4ez+kuX6h4OD
SEsOVcA2pjBsQOmIOdfJziQo7vg78DNo6qK5noHtDAF0WsI3KjL1EIex3qnYwjYlxpF6JjVYVKLs
NDBhMtBQA1TDUbbsXibr7s3laiBfOFGY+AVIDMitrBenTciRKPcTOGDiNxWcXvvT+Nt7o19JmGOX
wP+x0snyz8ADV1RmRlvrDe4RI0rcy6UJk+7J6ArQQmWyzRwflEc39WKJ2gL1CS1km3c4m6hZVX91
qFs4rIgKJwuX1kVd282HxfTIlqAPJ/laOFpk4bSD9k6yhCghTFsvqhxXJeQGj0N0dHjxGaM7v9+P
ZxIJNOTZKVeLNnaH3OmGsMvJ14xEpPkSD5JunElktI0DCRzhmirqmQPq4c4PsP+Dsijlg8lOiumE
Ny5fv7/dbzO0pXnFiToQbsGWWVvXA3rEuepYC3Jcz+CcX6FJNMt5BAFsPm82yT0i+UnQFX2HiD5h
pIs2/XjiiyQ66aSGrTDkVAZRMpd6xsGgLjt3MSty9/NcVrV0sFUuII21an8jIcH8GQO0YDemHa2X
YqNbSix9SQaFjOiKIaS2A7PKb5E2Bl7SB30KeqwGHg6B9m2gt18NGLbIoGHYylarpe97FZJYZOFQ
arFbVf6Hlu8FYx3ihKD6l4tO1aRAbdoXctZ9C1haMD8Vfg/+NQELXJYM1uggHR2MPO5iXtDOr9Ap
7YOszUY2I/zNDXMvs9Incpmjq0AUW3lWR89fwdg+bmjX6aVJTLk6+pgsiMZh8lR9qmp2FiBFmj9u
fkqUn66FO0TPVgKs3usekDPQEJ3+OPNH8FjnrO3OOHeuXVHvgsRumn3HPyMR/3CBJfRrwqjXa0Kk
QE8Bj9eny1BlhB4gYPuA6KUzzG9Nk5wq72GiTDzqWGW3PjeNLqHpuwh3mQFbU5gz4RMUczaaapB0
1lGVLyWoPZ9OGBkIv+iNICGwQSmd77JNUYtOyroEHwU/4n+9QeQWwatu0v8gPrR2Pz/jZpw4931z
hU9nydjixRUHm6Bprnzh1ZPo9q48/sjAxcrA3nu6GXU/TNfxFaEAwz/YIK/oMod3IkXI2DcCwwKM
QJGsCC41Yshbaa5PzTfdU6868u3n8P8dm12k1G4uhqH+abHV0rvTHEj1H7H0XQPY5rfrnf+BNR3b
ogAYqVfsBAQLwAG2AZAoKUOwxUCoA5gFDZSwvUJol7itV2fGcK4OmuBimI0NCyjkeKIN7kBJN5rc
XYY428UJ5BUDKeZ/h8agIZYlHRrMHznBaTpKTwuMbwCmGXTfZ2alPfrgFjmwFZdDL3D6Tl7I9rW3
q3qWqrNk5wUMajHZTGSkROsustHgpLkasrlXE86OhCjq32txJCS9iXRK884zZ3wtFlUD+VmVHe2M
4OTZr6Hu7FTY+XTkzUfKpFPa4fRuMqaC9bDLNS2+fPBKHI5DtFaGzYk4h3IBpsM2PdGmUkHoOymB
pl1kGUdN0JpGsrGQLumSwlvbzWTTAvY8a9nITXfLuw0iw52V0VUAZE9e/za9f/2r2P2aLSvfillz
fNxgyudD8kPIM9W+/TIaawpaGx0aJFPgwZUfCUF/dgqsuOdMxhU6bLPTN60wD7qNLakpaS5phNqT
+MHnAl0mMBmcFdQSXfNqq78UlZa3qUmbooKYd+4DpkH5usyPlxxY3Ef1V3LlGtmh1164rYFVoZqn
OeqQ4TsIAmXqq/tlQACgXTKw/YHSFiBhihjpFymCZHtIhWtjtNvsPqVbsGjif96ggoPwc/w9Cguz
olnjMc+GAWI2F35+1dwsuSBoY5pQupFePSNhzmDD9ZiEBt1So79amVSZbHix9VbJlFYmlUIMjLAC
icUzwh6myzkQd6khixO5WPQdhPnzjiWG+m7MgalqmMikhxrFt8xZ8WE69wt+rZajOqc1XsG+tJ2d
F88UGkCLOaxKS8XEPH392QXSqyODpKR/LO7QZKT8BmozBZI1ZV/qpx06L8Re/I1rfnKJRdIAdzJj
vMy+3lO9BVTZElMKWhyAua9pcV3iLG2EogwHc92ASqPmZdNTSyyS/s2pneQbaJE0kP37JUdtMuNH
FBNx2zFA6LrazQEsZMCOxPRRg2YrdkAWPEUJzT/O8I/FrH54CjRq/UcNVBHR49JCni2I93KXA+qX
AiEJQO+ORsQGyeqHW08fiKqvlAPjlr94WUBQoshbRY2NIPVc2rEsVx2kFIdpwqZ1iCcmA/PDIuWT
ihV3yy3nYLIBpvUt0Hoc8wPrbUuaRe8DZtHm2bX37N+1CjzSyZcG9YKzSU0autfFQpthSrXqVZBA
UVTG3yQUuWzlWmDuDt5zuOQOZlOdX8npQTafuaXZK+R+sJ9aevB4LIkFgdDZ4GI8H7vJYddg3BMm
2a+/G5FWpQmEDC5ynwTWOgiWhGG8wgS/yf/SpfPvVVwAkb3vRhaIKPEKwvx1aUZF0p1P90b/ViMb
OaYS/v0l+WGZHcPzf+vVx/SYSuMR0kEW0xOAjO4NqkgATVWOUi7khkXIA246AlfTvcLAemU27maw
d/ByiMDX2KG0cNKt7nABaavAchIkuS7Jl+UB6AZ6jQCzpqDYiz2X1NgFnJEQPjunS/usfRrZXfw5
ol7Lgyk/04GEM988WwIW9Pnm+LKrrmuZimIKTdsr0F0QYrPhpNeHYTXEo0nvUrqNPEPs1uMoOCQN
GTeED/+bLHb6uKNZLN+vXI6DNsAMcppbNCJ0vTgvPtoH60dceYl2XqUR4VJfKXvHwMreJ0U5m8NC
rEeUZfUpKDphWcouUVUXOsDq6fkZjdkBbOKPvpq3c49xzm0IHyPucgFIttIo5US35LOKvaR6L7zO
QpO9XflxLzBvn6LUcs+cSimVwKt87gAgIV1Q9hekiquassxWKBabUmPmUacj1dMQvXijhOaQNup9
uh22jivVR2lgEbc2WH7JQYzJuRHdMIc75hw+WkJuBRBaJkgLRz57dmD6NLoefJpI1CWnMY174RWq
UQUKVj2pUWHPVHLRUTdAxssQX98DSkrUhm+bLS1cG5ukceAW0KHuJ1451dZ/zXRKSolfLj9/BhAi
GwDzwi+HBLIDOoa7CZ1bXKmDLFsvr91u5S/StQhhlXTD4y0DZlKSj6sCZKY3CPzu/vcBrbMDHF0m
iDTMNmDgZXV14zsaK2BUqKl0w6eaGgloyre/SYKmwi1vv/+DMjXilORdGDo4vwfthE+GnsOounbL
KCKHcPeLbrus6OeqlyOx51/UMX6SdEF+4iii31gK+qxWwmWipquygV9DkyQy9iG3Vf951XWy+HVu
99LVrQlMZz1+Pyu4kBIHBWwDsuAEIfK64T4nhPLplIeRRaoP9CilbQJ5Y133DomviDeki/JEVbCh
RTeCUVoynut8GHduCKypubgyok5tIL02n6STpaXAblkkfofHeLQtxiiU/BDPVSoHb87s1pD9BbdI
JUwpxIJ+N+tbyIaZs7uuZTXHy2ZOEIicUjMYT/No4f8Xxm8XCVm5TrmAErPDlJ5Ywx6LeftoX14Q
aLqNHe2CUzPkWe2UQzNmO/M4IV3YEE1D/CGLuq8AfMTTPZUz4gIhWzmWKuayQxqrqhiNn5D4nGKk
sNkS2hGh6Zg+cH9+IYR67gt2wlkilRdfOxXOswxaak6MaBVVXOdeZCHxZq100VR+VbG00Sn1TYOY
xYAQBqgZoIl5lJZfrxMOPAW8XC7ryEnQ1ixPQQBXmrQv5Y9+vvF2Ac9HSyB27RB3QFVeXo6c8uNz
Ah2hAT4lNzf903xjmKu6QiQFQDD4cpymMw06ZNLvctV8MFAp2EefuWXkvnydb9mqO2ALKyn9fZVC
oxRWnxLm32ILmKGo4osp8CB5w6fnC67Hw1jGRqm+ypZtiKbORELJvGFtqFgJ50LFlfjwiWMCqab4
hfrEDOBgpUnXyyUZD51I8/MOoeV9JrqnG0gqlSmqujphyXE5kZfT1klzd+o/jj2yJlF8HqOSvmPT
A73PmeUnxyoEdDXsTlhSdIYtbnKoVfiEkmVlVnI234NrJotbfYksxsYKokydywmRMoypPOxf8TmZ
655uUVuba2eFMhrH5sfLL+gM9wZZE+446wbeEV23mWjeRkN2afcjuiogN0Jp9qorzxLpQQ2ofAj2
5DHBbKcpAcIlDf/i4zhS/e5dMaSFHiHZQn+lhYzUrd9q5nGSEiS7ETI6mqUSvG+9MMI0RZI5tNDl
QEgDZJBZnnCghvcg6rNFcyGohQ7NOyiE1w6HY20d1NayKS+3vjAAobEtZLePrPulJsM0jyst5vVC
CeQVpQ4uGocR+SRixMikMNNDaRQmAeIEqWX13Ib0V+m3xlVT/UJERjhxsZwdLsylVMicduKKJoyv
b/l/4FU4aM1mpqwrvdIpBWc7PvX6r2PIJfGXWZ+5w++5DsR4iEHY/BEy6Kz6hG2jCGTcQ4+F3y8z
dO69VbJmlCPrgNb9A2ClK2RtpCsBPt7rsI3D5emlcEW+G340KFy+Ij3Y4NsvAceiIbDemb7oOykA
bEL98Njdx2TPg1WVXJoIoAv5YceGrXMOzCopwXWrokPq7LwIi4faqcjndrzyq1yVwdFg/rtFDz6R
OgriZ8rO/CppPu88MPtf0I25Uu9l1Mpc7cV320115hzuvZUlH2sY8jBaH5sh5ED9iV/luZVjTfGr
toVuKeZ//unyiyLQLekAC94c0q6yn15qTW4+uliqr3sVonH6iaRQa6BpndCc5ayBwoHNDkZ4XcOB
hojy3h5pGsEBTqJym2O6L5JOdnrjT/0FFwwdqGchc5PsRBAdcNQBX/SKGdATGhoTA+3k3P7qxuqe
9FZgtagr4dQtcDPnR7ywMBPkfSNgtilM95AdIXuhue6n/dt3nUExtUMzuskFcljFr044q2y9wyr3
brtOBOX6+DSxp9psuGKAVNaAhqib9kYbhGcgI2uYfeshIZiIiyRhLRz2tiAS6aaQDVU+lmrs+8QZ
W0s4kSmAOMlYMeD+FBDcTLj2T4gW69axbee5P6s7M/pgPDWaQe4O79TMGVGfWyJBgnBaOjrsOm3A
4PQmYq+swEqHc1mOPECLkF7zkkLoHklNz5yCV8/UXUQiUEQW6Uq2CVyp8u2DItswBAyE7uanzfuM
dm48GGfYwji1Wb65RWba6DgWousjZM1XZSeA3UbuqD4IczL+9+f4W7TDt1vNC78hqxP2NEAsovwp
KHlMktXDzPcswLudvRTcfm+hCjAR47pOCUHpwec8SB0Ey/hssHnEkiKnzKCJd1GoSpXhTSi0qr6G
p5z4IsZ3+XVIX5R9m1Jwuuv7/3GjEFXKqk+mjlguKsNH6LF2GZdAnufsMyLcoUiYwwZcF0oGswQs
CHFpMuidacTc8iLGKKM3SVbqhVEy5t+BKRfocducgXDQVZs3Uwgdk/tNkCJtSQBPVZJSFPmrHRxf
S3E4ImzE31mzC/ClpMOtzBROBCOXoht875FPdYIFDrCbGGj1M6tCEYxCvHMP0Ojt0W8GXj518/Kr
VD99MS5papVmvEXLX4yHboiHmPVFM6Wmn1M+Qamxg9lEsG/BIuiLlv+5biLk6YKTgeuW3kRrYqx9
erwdKEkTSvO1sxkTU+txEEvFygt4vBPyRZEiwWqfWNuBtsDD+rmOTXhV+yfUlf5Qn0Y9MILT73ci
xdhCo/kZzH7tVSSx6rIrM/6UrVsmTvkr0ry80fSZblhV0mYrV6hcLvJU5MaRS+Twepp/Nfqy01B/
Ep73be8YDKxgJ6itEoLFXzrbpy6PrVs3BfmN1/eMPXOJ/3AK335LYZWu5SCBx5SE69o1rJV5JLp5
ILW3FJIfCQLbt/GwY/kUbhPeZD47/hbUfiwDjAFbHES84hYWFcVRSbSEUf623/xG/ZTiAIqMovIH
5tjjL3iqQqk2qwQl3adaTVLSNT4RpVhIBcJqZLsjwdCnwFyZ60qmzMy+JydGofN35gW+k2kMc6hV
mcfBYf3vKy3Lqdy+AdFkWDyD8G2qcoPBtATwKz3jIGQvlLA+7/qzf+/hrI+pXxuiRz7bQgt6Nl/+
nmYVAny62T65QeVEWjsVn6zA+sayVuzZfcd7yy0bPO5n2ORbxEF3a51uw+L871fR0J0nHA207qWg
EZvx3pU22rDHgKxD1GqVOtSpbmapxLEQ+4Dt4MtoBCO9ZweXDKTiwJN3tNH0qskqxGjGk9iTdAOk
DIs3bZxZuAVcbeuQgqXlOq2eyLMW+3LO/C7f125EJDZaDrBcgi9TcarGH7ajJEAr7yBfgjSdVjBY
KBuQnWScv8azRrB6UQnRNxKRpJb/AlZnwIrbMGWPDXEn23uZteuXMA224+Nu/K40ghUqwvrPsQ8i
tkeJzowBgzDpr+lY3ukpXbT4AbpNFjAqBC5iDfL50PbKuCnpVtEGaGYOwVwcLqoPXpoYRFRsR1gb
a9NtC1I57PryGGEDb+iA4REH6RRSGw5sT2dt90F0ct+kNy4rgbyJwoGbvBuZXI8TAO3RKpREPHKN
nGVvaTDUEpAbyFvJvN+RqYybUZJJ2CghvPH2GebHw8HKw1Q11SzHubzZEQgAB5KaGjzJE6x2Wa44
db/k9Sx7BfuRWeMhwUmE0Q1WVwEZYElBLGoBEd2/3TikBmP+Ju7sbzJkZKx5ub4rhPsMmG89QtCo
KdbyzxQlw0zS7i/AhunqBPBRHAyijnU84H+Yix0+MsTKJt5EryQSDTHwIiTht4NCPYoESqJKoCov
i2vegj1sWVPoL/NETVtlbK6ozqGZu6GDyZXPuoQl1j052wHgjuJ2pJPsfyKfNpWl3sDXkO9Up9T3
rUML4hDYLubu2LMcDJk7FA9tjFxz04HioyXyy8K02Ft557A/c78o9BKn4r9WcbITMdcfaP1wTUAM
/vCU0qyYKAgJ3hkiCXL0dAPaS7JfZ5Pe1Ix9y32Zr8K9sM2iXn4XoqNqJcKcMpIHFGWHBRYwZkfr
+ZuKq9n/8g4TGKrOb1RxalRcjsE5W0t4PK3tSpy06U5N0p3FeAS1hYrIKKWdYjcW4q8WefzSl7z3
jUwXJNuFA2U5WZwa3HTd23RPWnpT9TV5eK5UV+tl7OkuNChnnI0/WB82eej8vGw+dqnOgY0bq3Rm
uwf23sNcdSUK8uRdZp5KpD4CHfECM7T3CVMDoWlP63wzvi4Bo6GtRVU70kEy12X45SPtwrkkmnza
c9qnwsG9ao63p0OQggFDBkW536BRGwXvRdHfFniC4JBKwwjJaATn8q3G1WCHclzNX0DGIUG8FUmO
x3kVoxjeY432woiT576Qln3cHzchCG2asNgKErPnf2bfNKNj6wCx9vjyVHUG8Hb6zOtjCFboFBLg
pD872Hp8ZDXulaDlqDmwX9JBt6JmJiwIF4FjeUa74BzRKUH+jj4fYUUWLDo0qOrMRxwtzxT7zNFU
7e9KLc5z0vSBJ38Xi0ifOaNuLUFtlSSHFzxVKCr3ywp5pbzhO0CxUfMYNeAqsAAbVuY9IrV0Ey7a
8xN+IrdJ3CekoO5mfkY8om0BSyoeYW1RI/3c3jUIn0BM7rhibss1jr63+RuyiuUvNhqdijV5Vd79
7d82Tq23/yQILD3fUKbw6kpkb2SCF0HU93kqUna+gTl5jxnUf+3uMqI51oMKtFRC8G1EVn/9bnx/
4gjnjhdFeGjQfs12vyFsKZ9GMFdjCyGjZd6x9Nt2OghkTCkPGHQd28iExUWCC9lzCqbk3FLvYuGm
VQzqSR/aiwcF5ZVkMQabIuvvc6fcAhGBRZzW+q+W3GLgGPl4i2cMowaKP2KCW+AITYrR7PH1KjwF
qAGRJWidJ/5uLNJRKLDUQVVWLU4VulH5HZHStnDwwiZkWkBp6t7ndX7vp+UkLIFS0Fd/rR8qdaqe
fTuiDfsXb1kcNzuKufix49F+tfOcDdRTCLMCP0cMk++anrBwE/uwgWObyM+RPgMi0Iv5m8lxU5fd
5SFdXd93K9G5955UxX/lZLXaI+E7JhaZnadmpBctuKLvBBv2+eNbk8dnSwPOPPmuWRuzFY4V3tH4
NrSQvhaRbXsLecjctenG5Uh4SXe4rP5KCNzzJdhnaGk8S/9EkdAOMgLkNCdqfLZpXW9x7WAO3g82
ovYrmqBw9nV1gWHPUkHGNUVC5c8Rh5l2JI9X4Wy2ZGwhVoj5o71HZuQe0dpgAFqnCWTeK/oATG4p
JfPw5a5CsJacB4STnhs1jSPjvW0yKxurnPUjQsJux+QQyDobn77aW92y1MkuDiPyQDW70prQA7/L
AM1doQfUK8WYpAA9+tbG1KYDWgnp8usClOQ6MahIe0lukZBrRpIgc0ogbHDdnLCDJXBIlG+FGLMF
Jx5GJY7kQZDA92VC41Oerp50FrghDHsjOvKobywdINeyM6MNAICIjRv0BQJqxvltNW/Gf7U/21b1
3fp64RtBHGW0gVgAVrg8XDMxrLq791Sx4X5BZgKPD6XP7TKIw2OGZUFFxfE8d9oBU5uPzYiN0g2Q
CAMv3/mVWdx7NNk2pZ5t6DojyI5YXsbamqgymkmknM/fgNvmSWYb0YsycMGGVA+q6uB8cx6DyYFv
y0Ebf8yW0+TCqTeyHdKJaDH3DqLyX73cnsduVCUkCedCoX+os0MlR4wceGV0bPrsXu9C8XZbUUqV
tzJzt/tZDs+eQJll0xe6KLDYfpZnXS2TNuugVM13WvNtz+RUqHfPXNhwTp64Cwf8PJ1X343Pe28R
Ktx/3svZhI3Q7ChJF8QjMP7+j+VDQEFL/yxJtqJawudxrZVzr4mXvZh3RT3iy6/7n6KNDruOUnlh
5g2ecEK/FBTMR7gkaTSsxy6KL2OKhfzjYv4xRoCP5rKfOYaLULnqNFTqPH9P3PkaX9l77+5Y8D6b
yMtVdBpuMPFLn5IXxFKRrVDP4i8Od/8ZF3/e36JAVrSA69bdRUmaMIwi0xxR9paz6tn6tZDeGxFm
OekJ6W6iNhRCS21eX1ZXPtzyFFY5VqvFK7+Mjy0ET1QxCcafyrdKA+Nc5LRJt1prcuUux4iQd7W8
Y8Le42GdkY+3ikDCwxmi748+A4QF4w2PtrPccSq/tx88nfFWbHMBSepLcjy7uwix2QSsmQwshVYM
FY9gEdQB0hTbkbDwXdjjhS6W79fxHZMljimoli3BokhOG+V8n1vbd7QMccRP+FyuXLOKF3D/j0i+
0p4R3W2ngL0aGcitZFIPEKg7ENxjXXItmjAFxzp8q4XikIliHkIm2je0/r+mNHnvY6sqmQjXrwLx
b29aCP7bQ1ATSk16GgSkcFLPXgFPIxc+zw/WklDdS3+cKfqF+Iq/ZVoggK1zT9L4XT5qK6M4st4+
/z9ZI73u9SHqK62XWHiDI18c4JbyuPI4KCu/CcCa8o6GEcDAl1N4GHyfnwwoj9PeFpRm0cmbGmWt
L6jkuGxCmj/cg4tFrR1l/7XPEH5ofj+dgKYA0n1dfGL73tDIubr7AysE7TbSmrSogYNFAyJLQ0Ny
a0HnJuXZTzb1JNjl1c5ALqGGMwU51xRNC1yXLXC26aprZsRM8cW5VkJZoTAXUPlb4TCydG8UjqN3
r8hXyy/f8LXy6aRctG4rWG5znRUEHk04Yar6V8SbkubaHWNjfFDS1mCI7bbHwiMsKU6lfujZtn0F
QuRtGkTCcf1pZ6YSwJepSMVij5hPWm97orYEw7D2T0BZ4QxBD+goXF6I8SjANzCtio3l8KhIFJsR
4qSt5yR0YKkHHTJhczUA7JKTos6YgdnQhL+e5w5ucgkh0jEXC4ly14YrX7QLslQ5O4IzLp6khkrR
WJ3aFNKFBZu8lxazZZkzrespAH9E0RbIaLLJmi6zoMAqxo/yFUF+8lovx3G1667NyjmcLV1yDON1
pJxRZ3y11oXyOP4bhDFmWUAEamyhKafZCe4oA1K1J7X7hWvmWn4tkoCCmSYkoDNNmhf7Vhxw2zEl
JdO9Ox8+V4c5NHta3JKXjKUpHW2lVWhznBVt30uQCWM91kOHKE6sw1yAfk01D3wXWWOvWguUX/zX
w/C7FlyOQwh5Di219ZMwgUGzb33xR3zm3P2jrXjsNPZIaypwGbkHWYIcMSN5xuu9GIyAG/GL0AlO
he1eq4LfAZQ2hb97s0GeaIp1VupPMWUhmnCUbXiNeBZU4LKbvNiaxErR18+Hm0VYjik+liBPJSkC
7sCqLNiTvH1rKNiQMtZ61JmGiS47+xlEhccFqvEIBnx6Fx/xKQtNpEVQwGvdLm+UqfM/vcXTQ95/
+NEXZEMNnWf8cUQkfgDw94l3uI8ZhWfrm/OltCBASC2nwE4A7IzHK6hiE4vvmIaJ3WiggzTSzjvz
y+gk+JVwojsuA0EheQxqNlXN8okHxQF7EkY7EXs79BDg7srbRk15FCLgKrtpbg26v0aEk9RZb9E2
K7Ph2h57/samMRc3+KXaIDzb+SXRmCeB+GaLDvuzs5GS6K8zCzmGQgICNAA15DPsDGz7QVXGTekM
YQRCyXEMiELkP/9o7LXjyTG1CwY18dmPOUjuQk7qCZWRUkopG0kcpZVF8a3KS1nzsqNEO7umwlFK
NlmOv3NBqfWu/74LhlOlnFdlOpJexDODtL1O1Oy5bD8jGuIQi2QgCB7SrcK8+JNR+SUEYdvmrUcN
4kt/UdEpLskwHAmfpKHBindWP60tUv6BIpnHRNmdydO4Jn2gVY0JIfZuDaCbvBDqgwhOMKY6Owsa
B0IpCN1ZVIx6bcwvOx6hjUc6QGQ4Hs9QN88y+AOFJcunLNrTatfOc1rT0WvjYiwTXxBbPtvoSZaP
hx6ucNDfy9cL/Bk/cMyqGrqUYmV1Thbu3afvn6pjTPO41w4d1dsr66tfWJdOYS4S4+/5ncf4aUQo
KTIgEp97tLDDzbBweOVXLKy6iGxoQVzQHqXycFlUN/Xn6UQ4dg4BAXe43sRGz2pu+bqc1vPCPgwV
inCAq7FyAuIN2SLvAzO/5g1Tkp8DGOZispg1inHrZrROZOff3TEEtwd1Km71p5sdWbpTja9Jch8W
FcCZbB4r7dk6Pv8Oxj3xMGhaBC2C39SisCnICIf7wWH8rbQ+/qt6h8DwJ5Y4XOj1MgO0lhmQXSKL
LhUezqeGqoUJDB050rOG0h8LhkxgBaxl6CUdJShhK9FtYCUfcXjaSXBB/cgxyLS9uu8IJBZhxHIF
jiVLogHzna30OP+LcKj/Wh4d6mPvFqVUfsVyzCpejqsVq8p7x0T0vzSgddM85hhFL/kyhRyTF6Pn
OoUxs5APja6jP4y3wixqLh7OhLEv6dODTJ6bjuwcIpFD4aiRRNhvNoVQmNBDTLnA53RbY2K92x8Z
RCat7A20hO8v14hirGeF4Hg7ej+avWZuaa367GA4Qp9eldyUC3jsmk7ceN4895vqzseA0WDThGTO
sstWEXne45eTMdnGFXxO+Nue93OKLFPFBjHlMS8+QGxFsOOTENDRXRVmBZReQ44aMmOixtfTkXr0
RIEU0GMHFM10WqlLeRdoBrY7rdWLPtAx/g/bTzpQWRvhKpI1zxa5b0DRxAs3Z97DvkTgAjIaGqjY
cgzTAGXeBdd44ydvpsc2u4wWjmBsA5sHrCcyPm6YtuUisd3V1PHAiFinHvRrcDS010FbYUujPNMa
dyu4wcwXAk2EckeEgVPljxXwPiKJN6/16Jk3mR4ZUGwYY6QWNqYUuVpXtLcOI7jdMsoRk8qtAaFQ
Ax4ynBy2JAV8YP+LCdX47rm6V2M1bfN3D8fhsg9bcuaf1Q8l9xyILmVI8CE0cE6QOhcAHt2sztCW
4CWk6sa0rFVIEwuNCsvZmdpDCJ9pJT+44mBCpDovs1Bg/cNumlEFLsZIdchH073AN35fR7k2XTD2
wcl5Bj6hGq8SAIYtsQLncZG/bilomLWLmlVWsk8pQcCWJvW4TIVtCIXiHZ5UXZjCtOTQrwAAGAnp
n5Oe9CU6jAPNWkRcp2aFbFfRAhCYeHHEu0i5BL4oPfSyywfoskduY6NIv2S4PUbJqw+E4C1yNrVd
339gs6X/6q+uNso5BITgYC6PIDsusr05eoK9bVi2/7SXtpyL5rhRlbIPM14lpEBhSQ6+BbQk4rzF
IS7W5v3PW9fCAIdEPMoMUB+LvzOezV8H1uxukTnQanlQEH9eJIFVKYsY9Viz8eu8BZeononV/Tm8
1kojKGW1Pz6uDO/Nikr5F1Dcdif3lu6b1L3kIYbQKpOXxbi74yOyMe4ToJtNDObx1zkEEySjiJxA
gHt8tACNzRa4XJzUqbWguCqGw4qgKBRWidq8kSlqmT5M9t07g5HHOP+U0yduTkk8qEuFuvLDmbZc
YzRZiaWtxtgYeSTnEfOiFzxBcQv25Ujoz3yR2VeAwwTshoHj2kqdZcpgDfmZGgpYg2H1elf2H3cH
+gpMBpXrVuZKQutYB6u/wYut07BqJycfbVraj8PJixFanAJ4uBSshNgdQRp7trtNeDiEF+qbRFy3
4x6z1Z85BVVSmPuap13XccWhveww/XDLV2jYNxSjlVoVqCzVTPe+CTLUkpsa9ik9/WBIjzY4f+uV
vITSJTBjER3R/y6xC+iz3yZFXJnucecsk99IkHlOnmtxOkMOixWLejzhPLgtvi0vf27SUIYY6Zse
byoAgVlwGJSAvj2bQ8/6YDWzLs/1LZ22JOcsrmxrKXgF0nMqLYvtDgmzLHw26pVqSxlreeHv5O7w
gRQqZaboPZtnkr+PAVJx5C0ItEouxUqGKsyY1QBWivio582wWFcvNAnN8CVdK/SqST5auRuJxo2Q
oHY4dOxsBXjMRfyVjp04y3dRh9wfJZTsWwZfjyed+ToGVqmFGPqGyvtUTWArl/Y5eNe73aX2qo/H
DAy6Ni0anP5NPHHw6V3KDJCv+siqJlSoOaxPSPWIJcz3IipdIpMJRs7Kb1JpbSiX7yRu5CY5M5Yt
PMnm8TJ0Xse4CpPavFykEBUZ9HiU8eGc8Wuu6ozuRbwdYsawSkWpEusNKZlhpCi6kF1J1mNUW6Mk
+pJUnf52+V/GusfQmS6uQpeS6pwuG0qTsa4FdyW8neFNJmF//TamuWmxMYFZg0JmgruuHPRzUwB4
WfXksYGv7p0Rd/vtHuh+Rw72YjHlTJH8dNaZQKabOSAPug3JgRs6jU4uBp3PgCE66TH2LnCCUw7H
A0UH+evHNY8h388FLi+p/kk1lmKoE/2I69tESTt2JSequfufcEATe2qxmr/SZTVG3tH8D3U9Ti4c
76zcJ2SK5vjRVrN4031a3TCq+4kf1J2dxugU5Ad03VB/EbMqzLEj6YPQyBYi/SOlQIUcrUoF3srF
d37F7dwnRWBuwWDHskGqiVHqxljCZLpUCxFdpV4CbrhVhl8wGEecBTqU8tpRysffpFrTr6px1dUq
jPqiKA4EFeYxpIIKgr/fLvqO3rJzLY72CV+plJEK0DsFOLwMK9+L0pE6wsQQ3yOjGUGXTku7ionJ
yYeWy6QCnZ/RuR79dBfwF2jTeguum0JbIypM/L4++JjqOKEsF/odEH2gbsK4cnUYugu0OAeLLE6K
mqYlGkfwjxQrH4tFoGTGPf3ZKPgkUbM9fkuUm2ZSchGNqqT7QD1xE8nxoit95CxoHBrEtI9tZkeZ
lYzjaxK3DwyISj93PBdmoWE1Xlh53lhjycP8mlBkYURMpmsLpVdaijwczIpXwTOsj6kxrhWWqIYK
HlHD/NuGBwWHKMu6+CvzZNql81havCJOuQ6gwmKb5Wfr2QlNfF/KBRPwZqmNA8mWMKEyL0wL0E2T
J6JZ2SXv+p0Uj42yTVKLvOtmy0B75XBCLxVbmC2HVSebwWHP0/mOnYvRb9B/Z7FpvtbuBXxBdx62
U5vW5Ay0NrXEfEhih688BYlEfzwR/TCfJ12WDSZzoCdmbOJP9/VmlPSvHpX4TakSHawasDTVYvq7
91CYhogve61zAwMhT8CB7U6cJeFZeeh60Oyoc+eTYQ7vxjKCRqCQbwD25bqt/JosSVr4QwzENRdY
QQ228suTbXo6M4byLFHOlmEZ4sWHqbDCengbuac3iQHyaUYF7Qk/93bELzY8EpiJybSef95hHD22
ZhcCIi69HKQo6S2Nd950OBRTpdTMpzYmZm5+57XwADFZUC4fnr/qAv6oauqR02D58+VU6IgzCznV
ExLjSb/N4gvSfOHIbApOicn9TaeEzHqwLlqIBsR0axiDXgeRci2OicxVg3tnzzZHBlikbpk1eu+D
4hpnWUUmc7QttJ0w0u53Hc4ZhQSKX1fTtKahIFnuaa6gqg2rPfgC9r12O+JLeNjZvEZOV3xO8U8S
yxJcg6pjWN+byUnS61dKnyuxtBMFbICW7+3/OGyvWphZPjRBHF6RHJmZ+CsbImHGfnwGMqnhaUTj
kH9g+jtNpZI6gwPMgC6KwfRfvQc7ctf0jsjOTBYvV4JDxGx+6Z5yce+gp6iJbfxKrFvvavDheTxb
L4XJZ30Bxw4aZuHgeg+2vjMYqBI5BhQubVGV4dUp5RlJqyWaneVeWoGh7VFXLg6spzYJhms18LbK
a7J2R2qF4mNtbHFWFNaXgHRfBl0i7V/1549PTfh+C/XArpdTuaFnOtkif36TJeG6uJgEHdbK5YVK
/Vw1ldqfwvvw/vcLZzIb5Ekn53AS80bqtKJqfIGA5SHrV3R2w0+6rDp2SbbAPIOKOTV9iZ1T4VQr
t9dAzHq9MQp0pi37KlP7c9k0YvnAsHIv3/hvARsf+6d1/rO3iCNo5Nuj9c/a4RxGnLESBqcageyB
1PxgMY0JeTSVvNL/ynfwDRcjY8losSGjFIeejz5N8uDZjM1VJ5t74RbgTUH4eBEUFd7iPY4kVa60
Ra7TFPYf6tIVsmhuaL66cgeka+MG9T6bUIgjuCwGXh1HqC9rFSlIuyIv3oeTZyWs985+6GM6mKmn
nFuaO/xN1ezaNXsMUHEK9KhW1ABLi5JXi/e1hxpeFNwKhbFXuXULKmRJ6AIwJzWPNY9QBD/jwLMR
FDQ1KTiLRJk7g35WnEjcG4KBAfqv6mESotIzhITO2yarOzgGiX1jTG38tPnUKkND56oYD4TbXsK1
PYJ0ldlONKImrXv0TFaIjhXegMsmYYW2r07fykNOMqjIXATYsc0f1GfHikBniP2pRUmDhJx/Wodb
aCqO4HMoD3RM07G91DE7LppHp0EIk5aQBT7Yv4a9zu8cBKcx4O7Z0wNu3VDfCzZyNgxNU9tK4yfF
+J15RvYYFZQF3Y7keNAPkMDvuFcBimbiDZZY5h+h+ujv+D+dduyD3VbPk1Y8rYTnezykc6cFyz+t
ZCNuJ+dgVE9HRRgkK36zKteAuxWFf5e6Iojiou9CRKSYO40GpzB2KXQXFdAS8ci4yawwSrtcb1RW
CrX5AR+D1U7ayCtX76CL2bEn2EMMe3UByG8naLCa7ljtcGUKY8k12EZDZAtaPqANEg+AoyOMfCyi
y9ZVntgUSq8LsFSHOCU1nDvnq/ObKrgkSr6Qcf5ILPzaZ9a8vh6C9jkVvIY3KVHPrDdYuRx3WLgF
nO/85oCxkN6SeriXCDjwNqGVnXjOZgz2Pa68UBxb9RSsyNnpbDuRK9mpISrJNlHsLCZ/EqEUPtaq
ZVglql4LnCZ8a0nnRxYy0iDUDUiMlzwFRQpDVv7hywPoqcWbyPFuK0mJpssjGyf9WuzO+qZGEwap
CRMUdts4m6VVIT5GoJmABxnLSewxW3DK8jZacmHOjBf6AlbIDTvQmM1K/mkv2HYxXYndk8owCXgG
3fKVpGyoxnYzttLJ+XJRyU9CrHM06HB4mDk/pCHFLiKYZJabejQb6rm7Unr3rhP60vTkLOxK5rg7
VY6nwgHmivGrDhdlfTWrWCllvjs+Vdspxq04HPeFjL7f+cKWhZYGXcVoEWlt5TxYorSX+pthhZiW
WDhT/uJcVa5UsDll48IBqmW3gRQMSxeK3lRJcVos59VL5N1zu+P6ueuOC8npuKaE+sOgnsKHlD8D
7BdGKYUbHIuXjjwvbZviNZESSuGePXRnVxdg7kBYgQU9aDT+c85n8CKDJSaIdmVq8HOirlSDOC47
7s3gtHan4VxnWFdPEusXvdpxgoGUnpoqiMfC0zahou30MXsQEIfdp2nK1SNUs9auOjSLNUk6EZ3l
AR+O5taUonagAGXEC7C9afr/gl7xEh2SCAqU4RGVcEkaDCYq8oM0iTCqSQI/lneCsHNNiFSI+ImT
7nbcX6oZ56cb9HZpuAj2/ZrhjjBJX/KWMcWpxFSar755wFGy2tYTD2/VOXFwNtwAh9NLsWYs/shm
z+0MJhY9MZFHuXIw+zvZDHeFKMs8W8mc8vXkyz8bGblN5/rNeeGeZ10e8NgtPXbkeyMQuGnjfbRG
2mvus2XwbUNZ3e3KsGRVxPqTiY6u6BTzjiFIaY5/q/VbSTdLwetchv0A/SY57AlR5cOl3Le2p45M
MX3xti+s709tz0twR5wgefuEOotCEcYHhUMeHoseVHyy0DmDilo70Jxbm03CSvatyz0fwOzRZ+BX
xxWCy/BbLsifjTfnKKXSWPAf4ZylDNiBfw3+I6saQne9nRkKd+h5AFSIas2WcxclXQFpQCxvwsRs
aI5xFtFAcUDTEDeRCObNuVsN8IuY9ky3iF0ThCmsHRbEyzhV0O1aWHvLkmFrTzDCYlb1AWZCPXFX
eUrRSOudeFJw2qCRbCIkdzIOmxEyRrkUo0uKfl9/+RKYZmrhd9LVLeYFiv5TPpVHcPKj6tt2NFPh
qBi+ES+GtiPG9HU4gVjp3fOKvg7bDVYJQwTj9rsDeBdtKz/HYVj48pQD4BHW2Sei5NCAbAvOOFcG
espLTZ7bWkym80qcQ0pPKuQp9bpnlABXM5SaOG9QLTpGo0/Kq7x1zVgfa6SUMO+53evbZvrztY8U
qafBKdjGLO36WpehkLhPMaA5ZQZpjaf+qKt54R/3/Dmei8DTAOX1C75eav4Nyh608va58A+D8hX6
WWjzw+2KJeb9uRR/KEXZFihzC1c29kB1PU015S2Ph6zaIUogGWIKOAMDa5ipCmMROhFiKuEDOwch
sTR5XlQpwhkhMf72zPyG4J6vPbYf3FPWX3itPA7/hx2eUSFOwAJjAMcMz/5WOWHdATMk/Rkzmypu
GD2zTNbuyTY/rNru3+mrJRCa5iSnzqRlPITYxfY4w98YatccuQKmpAjVAM0ulxKBWgXAyhy/o3Vb
YzDE01IrX37iSGB1Lc31smPD/HvUAaxztiyWYcVxfKpPcSZUgUkUQoUTnYDGypr2QyOiDMdOsnEp
ha6/fx/R7J2BPmbqUL/MP6e7rqjVw1HykhbXdbPS/5dYbZj69iEALRUNztkiwXyZGTZxJO6ecQVn
2USwdPLyZslz+8XP1di2+dmyyxgcld3zGyD7YWRAR1JBG392vIDgutzvBEbczXHS4yizy/hIpcoK
9VBXb7zVfZgAHvIpg9TJQCVSUXkV3VYWPWDFwtTGHyaLvO9KGBCGcbuCTYob4mzefHGkbGIMc7pf
YdfbRbOIOMkhHTAYhYwg8yo9u1ERvodqtGw6/CPLYHqktt2BnsH8hplORguCpSgKNmkQ8g31Lc0S
RgKOATt9XoabZfqLzmvRNSnpA+DHdKVkHzKT/0+XjIHy1HTTrmEA8G2ab/jdW6UsVEdwT48cfHC9
O+vHoT0cICqHKAFtbxyKaYQUYnb4nij3lcUGm6aLhuOpiyNW9Qs8LcwRaNHS94nHZXjDSz0rdNbq
NwZ+zmJ2JHTfRM8E1/9fhshAm9yEkMVD4SSqRfFOAV+2mHo9xANTt4uQDI1V5DN2Z3HDkSCYEy27
i5FAhIgDUNiCqe/rBF6DddL7OsKYJLxv8dM1t4GF2OANeXzUogcg+EVpjSjUBU1yTFzxQjp9KXri
tXjgHyYrICOF1LRXDHVjfL53lRE9DF9kTWGc4C5v/Y/HNd4vrgAASOjUygVzmZhP+wF5hQngEfNQ
Yb1IP6KhJL3pbAKVqn4DK+zokpeL1rFAoAatGDAYqNTUChq01jJjc2L0ApsJbOFtDGCE4ymJNnA+
fRSn5AKEJdLZNdH7HEgTa3dINOZtgwyCtapJKQzqGFWkes96nG7jtmchWNi/xDODVaHvVyDCN+J4
ZaaG877QLYxWhEHVfpnC1QhnoJplMJcWlRh0VL2JmGPszf8yjMNiF/KjY8OL0Jdo+7aK57x7Rhhp
5exDOjbf2uG6ZaG7eV0cAyDrUnYPW6UTB2Tgcc8ewzt1ULpsS/kbB0kjMvdDrymhhcftZ/15ALPd
QOLAaPWuvrEGrE99PL7l2ah1RJ4oZ4vp5tn6O7oKCSYkjNWbVIaXblIqU0HpJ4T86qAPCGb/X1Du
6Mb2SxEz+el4a1yhfdLyaOlJQwvHypDuXV1hjGaaZ2YIJcmQpB2Ly8ZopznVVirKgSO4PablB8DH
c0fjN3l9ZG7kCVpFeE05hvSRGlloFFq2g58ze4thLAQqVejcsXyBXztnTEonZpFB0KEyl966L4+h
7BiXhLsnn5LVa+qPQfQrC7AuDmhIQeJ6NLBgotQ3FpoIQTLK/X5q1OuH37BqPJ4ohZPRBbNE4qwK
/WLHV/y7olGTaXwwS8fuBsrYgBvA91kiCajAEH8/fSDpF6TM62OOggRWdB1blxEO72rTaOE96Za6
AUKjtzloI/q71b7fX9EH0/KfSg1mRsCX+Cc3a7UeIxf53sLqJC1oyxaKoN6S/y6xHuPO30sTiydF
uf6JFtcYOdp1Re3Gs7KWtNSEiOwKL6Sq/GL+SKZXmscDZEPJhTwOtnr5wOETTkb92t7ioA4T//fc
9OnD1RX7v/u8RhewRg+K/4q6asMhV5+2N9u5zelwzDPY3VfzNXpixYhLy4lxTzu7F4J++pSAUtPL
ALvZDmcwHD+COVW9mUH9MmBuVImMctyPBIq/s+1GEcKLMIMoiQu7DLznpE9Mj9WVoLOFV8YhNbrS
cg4aMR7Bt2yEry/ROnmylynhp4i8zhze4cx+bo1714MZ7Z48ZYkZRIjz8fa8LrmGHDIGQnzEjDH+
sTL+OXlGlpYsk6leeV2jXma7mLLzdCA2YTuwk/2BmHmV+UN/WFjBy4kQAhSmYP/3pzkEsqDMf019
jEcCORZW5tIzLSILBTYkfKvJXFDSsYomO6nBzCXvyn+pxPYyfpiLknfu2g0sroReochBrn28dc5Y
E9E9iPY6Yw4GxCT4SRPe2kAD75VuwnsvJhBHtfUWdGEWc5N0Z0uoHROeIhAatBIDtQoeRNBPqw1n
dqNcJeKZq9KwlSelBsRZJ2liNjlOqr0TGZz3A/PQoN+vH99FyO3YPvMqlppgRTWEbaxRH0GnzJLD
JhNVwuXYmRseO2wCVBj1TUweaLwf3BGVLhkULRQq9hIOLcu82nMrfCWFWWg09ZFE1Km/8B6N75cR
4nHqhRFBxGSUuEq0bbA9FMzt5nnGs4RjgNCaLaSiabbsQooDBc3G/nddacIABVawNzWu7LCZr2SA
b9gD9GLaeFgFkgpkDa5+aNObqdVFDCXvcCiXtNTchAgP0CRA3RjjcV5LBeirifSchnlyErZjnaFa
N73UTB6DMf9FgfGfbtb570yoSGoaG8ZVQlBFnyK8K9GDE+cytmMULT+1nNOWwVj4yb4884S/R2pY
uGRpj+4PcQM1BHtljwDLXgyJBUHdHBtaw7CqWDg0QQFdbB7NZZrg1lUIk9EhejbLEIejAg7X0WIR
MsJQ+PFvRNmRFllINxQuuUqtdeIEyak0LL2cTZ23xfRQZ1xdTMVE3LJ2kktSnl3+3UZMbZTXTE3y
HZLuAsy2vlAJ5K/FbVqZ8aZ+GK0geuXK2eDNMCzDdGcIf3L10b2wgBHCHexoIBReg3L/e4iLsQye
CBKVjike8sDuYSTszYndUDDxYn/t8Lwq0oU3r55EndUeiJK+NefyiYvNGmWSROkuiLOSpsAxFC7j
inCKasE04rJfLD2iRJ2Urw7HMLkzI2yDAnTVjc1g+eyMgQNCaDXpuITxVO1z69iTenLdi41m7Rm6
R+V/hnekRkSe8PdGsXib7TYEkLqpNX+fKcJ7AvboqirgvAbDQkRgii3STBWb+oRqlBLnmGBQo2Hg
XfFCkmn+0z2hmTvaLBt7caNEpObVYlhyOkA1dCLfb1RjbgJpWoJvZTn22FG7ZLzE9/soeLizEo/p
gUKPoOBbZK1QKHJNp/Os/04Pzhkk8gcbRE/4Mt7bX6mUhUvDjooZecmTbZFjq+fOdg5EfFP2Ly5j
zTuMfGJXMFpl0OZuyOx2TWj2q0RI0PZS4PmipqGtMjJT+7nFLM1oOaqpPfl1CSoeKTMA1+feCMeF
427VCPrmXuozBC/ZCmjwBOwPSa4Tuv7GYV2bfPgy+m6hE7td2uixQLGLt7nO6RyGKPsRTqv7KiTm
ENET2RSpDrOjzkFsktfjZNoc8B79ttzSMRCvOUHh7JI+fVEZP+xItHDTAi02bdOxxd/4hIwGeVUZ
WIAFCljNiwst8t6zd8+/kRkgokiU/lwEKkpzwvsg6BVdPk83bLb9rqkXHortfHSBSca/Q0jyebwY
bOLEODOIIgGcXlsJV8ENviBZz/XgomXPR9MmyoU6eWSFmoANeJlCHY3YIiAQTrvWwTpZRFKPCnx7
4b5SkoZOxQqkc0rlHGgplxlEPaG1h2kNasRN5PLccvjpq6/YNq1okkyhnL6IwtZeowXYApcR5su3
feegDF03aY7oxswcype4rfp/qn3S0pig333HKS7dfA38gpY/6wUCVVezpEo0aaAf4QlD3Ypre8uT
P2bGxXK+YtmqGsB21n9nIR7XHHOS3/kf3czs2akmM197vJxA13Hx4L/EWjPuaebccAakAsk3urIF
apKV9vqt+65Az4YiJGONbgVtXjM2El7wy4E/ubV4SdSoXNZ5x3NUUWzzNpipIxWuvvhAs6RtnQm2
sr+p9piuHhFmin0dB8JRbzJx2J/HiwtGRd1ILybtT+Pa2QPFWd6sis/ijR6MvNx87HA7xcFD9BZ0
b6xDj5vsz3yI1MyJlFEHP6PTqeqLwkD1ClALSKVwl2TDOVmHrUAJbbZ2T6s3iaAxi3jOOdstK7ue
UmdRBSfve9mMI27HFogDTMCuIe/28AC4Vw7lJI3BcslfIvcafhvdbBNeNYJXI+tzYhFeqBgNpfTr
wTPSDrGMKDoq3SzCDkAWkPWqofBp4vZ9UINvIHVTvgZulMD1NHwE7+sa+wPXHBPD8m3nZFgl1Z54
kSxV8iNDMzNnue6vGTuH57XY9brS5kC1OvWMdtM9PUnYYBubStUMQArRaMY/qcYgyY7q6HgdHtPh
QoVebYamVJUmWQjxn5R3tnZY0PiHxXcwJiKpsObffe5o7wjQCiFhCPOSeIMo+YXOePLZ0YiNzGxs
Kr3+fotffTT16yUwwEmoZd8SxCKqa1nSKtT+npENxc4xDoD3eoqGejNJeJWgp8x8Xp9fjvTp904H
voHSRBgoySxsyxplQP43Qd614153MMakyLIOdMShq/LtZlIXHGt4qBs5U4hHdaOI64NHlPr9LoHy
x+HWb5630qcxBhwiGKWnu1q0CgLbQ9TpTojvcGNTkLDF2NPTd3XvM0I35qnWta3VjF0s30bqmsIL
XWwPnSbFRNuh1bsNVUrpH1BjpfNB+4l3AYOyfrauRX24iBBXnbquinSdUytxNdaycnPUlHzJp6DD
Y5MAkUE0rdUc1Qp33kw42g9e6IEZCvjBSnff4bnPZGf5Qw+tNx21YPUZUtlamqxqRRMLoRdEodhj
toA/u6V2MP1dVNm0mJc/DaKaHOKIJ1ZgLf0Wl7PmGB8gHLmxeSj3JkMClwmUwGRVza75LTuhSduO
6MaED87ns9wdfVV9ZEDeDkHigSSC1ZdHfdXkyFmXiRXk6ugGcVsM1K4/P+FZtkmGliKse0L2TtjT
1ktcTL1fT2CeSatuqGQpZY1gKa1RAv65kNbPHOc7ojQgPTjIlOKRRORJIebUOXUk68fZ8Oe2Kwe7
aJGZ8uLk+Zc7wqY07BAwVI+rdQsmGeDg2d23pFDxuRUy9BkeLtfgKp/QWBWcGF3bd/sHrQjk/Kz7
U/0k2pxszBbiH22Vdz20689Vbd/+A1r1SL7PVcQMZi0MkGJtxYcxhDjwZ3Ox0v5WffbHyWLwSc0c
4IjkdiKnUPs9yByMXeDvrYDU3p8fR0sAOJerW3p2+lYkydRMW1zA5ydrylJBVDAqA1HSQDevkIOE
+jOwrwjb8qn5S1fJP5j4yLt/cPqXq1lV7Mh2gEgQHX7CL0QhT56v1LJ/c3AnfJFYXNfiliM8AeUr
PaqvTCNMGNa2no3PrRVE0daI6qaZ3DeTjupo7pEtV1p054x5cH6JCtcAvroqEiUVWSBmbxXzQbVq
Q1y7+jHVEPl+XkWu5NL8FIyjrSxiLoEXeNh3m2MTyLNjYsoaO9vDKb/Dkt/mc9tBbI5Nicsf482C
RdmutFe35KwDPQEjyZcV6xz7aQQwb0T2+gFqpqioToZaYA9O5jLpsLsOQcLXTcIsQnZdALT0i4Fp
oKW3CKY+v6400f4BGg23YyJOpoI0drY7eht2zH6X7uaWtjEXVaDPG20BLPWpjl4DqhEz0NIMasCE
HaenzowlGhsrQUTLJDrCW6dcabE96dp6PrUH9URJM8ebizV+VqkukoJH2m00sY9Qvn1iz247KT+m
nO1GIc8yqu8bU1OvUtnnHvqLUTXqp5LWBmRDxvKJQTDBdeCU672h13DjWZKvc3T4k1+022OOm+TV
8R4IZUXhkfKNSI+rB/cfIWwqP8ZhGKnz3+M7EZiNq9ZbrZaBPjxl5s25H8zJUXz+UnvKK7E9RSjj
e7dF7r9qk7plowgYy3zBtFcXkLVRdj7qT0F14KR1nVIoohX2Enz9PWZvyINzAIRk89GzPBSYGCA5
QUh5/ZkzFgnCzlnsufpb1eyNsKrh4jvqPcoi29vrXIYVbCryVuInZ9jw2a1HFdgDLRuV2igoXaAO
ME7dmKW2LUoITMxpFOSUrBTV8NbsAwsSSDAByEe959GkCri6jUE5CF8TXWeCe+UtiFx8Igpq1dW9
+QG61R0Ai7h/twR6TK05dQi4gcxJHubCQd2W5xKfn+/zVm73b+fL8NHSTnP13Ec3oWMMkywxqzda
LV88pq2Fd5qnQnYFLtxfKoSJBb91mKvuTRAsDk1Ui+/KMl8n6jBtc04OfxYO5C3cnIxZmjn5iMw8
CKvEbg9U9IaGnJje2dnO0sT4FVQ2eqeGwWd5eVG08EgHDXFa2E7Q9slpm2oK1JdxDDGq3wPbsINd
fcmY0eYt3lRo1mTm2vuC4NydxyTP3aAJFiIDKMY0fIFA4HPL+ncwVTs3ReKFJBaI4+2T1xa6J5q/
irbbF9DpQPQZQxZ9c5IAvel8wPnWQCDwA5aLrVrv6CQ3AQD9dv9LcnEiBYBNd7p+k40JLSd+ZqjI
HA3LC8O0npCKePR6BNjSwDkoxuMdMEE8Hbp0ymncl41k92hys08nhsA0LKa0PQkU/QBnnGfbGUHp
PpD1Jy8yU5088gm4b2d8HKRgrqwWpQuhgnFtXj6GJ06EiYpOH9dZZ9M7jv/mh5JNxzlXAoe8WEgx
ZoiNvW2jv66El3EPDJuyfCb+MTbJXIeYG0G0rUVqClGmJ6DloP1iFzHdSMIxTijrRoOyBEdiW57/
TegOUYIQ1HzHZdZf0h2sKneEescbweCljxEd/8QS/4WmvcLm0DniySabcYIMH4oVPAsGRzSKV+Gq
10UNgq9jqYwMh4+aWgScjQ/CVycrx2K4x1gPf2aVlO/w7Yl6zF5AVzx1lJBTGodTQ0lXzVRa2Ove
ZEs4UG2nK8i/UqEq6NmiiOLPTrWNswcm4ejAFuQs8Rh8ttDeLhxR6J+Vip4/VjJyTVPTXdOSiOCI
A7PyPYSvov2hAxuUbTBCYfAP77L3kdlC49uB0Yf3K9vtzgtHguJcSw75jBhfjIkI+4BEnj8Je/Hy
86GjhO0RQ6xlY7VhUuIFzE7rsjjW0cgICsecDgc8XyyitNGFWHdedU8xBrWqyIkY121jzA33x9/B
vDFj3Oa4Hk73LnPlFvYQ/kqzIJs7UDhDvtxHtkW10tQbgtBesj9TSFBwcgo+3qhW5jHebSPBwiGa
FwOpRLpcQlROKv9yMpG2kU8+/H+5eHjO+KX5fmyvL5eOqhBcz1t4+hCn4ZbUiluczbdrT7C8xYBP
Ei33YvOHk4l2KeNdX/Cqpbg1eTkPim+Qzee5FIDL/5wqO8QD90yvYNJ+rZkrrihksJBKE6Jt4eaD
274oNma/9rCeQRsBXkRgWIzRCd7OVt2PExRW3x4TaNI2BZzwRraLwybNYwwDxurtYLE+yi8f7ZOf
Mrj9/H3t4xD0fTY95vfEetMDpf215EyvZujMKfmqZkjYzQxlcyEvDAJE8YcajKAWw5ynAmZpFU+3
+9FHWimuNEUKliZ9XgurtnpFf5ZifeTaI2smFZqOvA/XsTfenpZU6bNprfPCVWnsFIqM81PJaScg
o9D8+HkuJ4Twc+48Geux/AiYrL8PHWxxggahvbhQf3cONaEkPXayotgPQqQMUJtCZ/cmiQNkCLoo
PuQwCYNdm5Fj9JqH5ee5/yc9HIgJEzLwzJ34dyAp+JqhgdEEa0tZ36SbLGS1JcG9VyHUTT2FH+ph
UBXPyTCAEQnzIDNkujadzx8IYDJjQGgnY9zFd3OFt3vHPH3iSOPYgarDR6HotJ3IalewlvppGV9U
vbWFMGyVAIjj/lHoAIbjtV4pTwSgQQIUgF1uGhBce4oKoB7VFxPx9wjWONT1NYzXFGocq5j8ghA3
PdeDFbr6v7SAzuqDkkHROQZkkUXXzMFVsNnhHxjNYO5Azp6VmTehIqIm+9BNxBN4fiuMFyJeZGNl
Yqb+73GfKHujlGtMb/OcFdY46qs8IFZhTiVamxv7NQhSUyfGTRnrkJZCmAFqM8uescupKHeYtMmn
++8+zQKa2KTyAFuWulvOrkNKarjxVZsYAjhotsbqGe8NxGbOUTNWtzqgezwKwqG1ZCXMud2vs3fK
aVKM1kdNweD8KZXw86Fi/kDoNQMgtGLKiu6KUSrtNhEeHef7uanNIwDxHrcweJ967T+QlIraZho/
j0PEDinUdgvGRJupO0BxZ/bYUvEBTtcIkVxNt3pCFSLDfZQHNKjI4HFznmGxdtv8jXrFgQvz5ujH
hrdoRi2I7pTjIGHVut/3+DIBJY5834qgvM6Ivm79d1SWhibANmObGhgGy9AxQarxi7K/9B/gbt2J
uoWoY91CWS2oXO1Ex299ThYvwk9hTuFrd0q/frab+1qJL3lVY9bfP0b+cnSbjDieP6mn1fWYw0ml
rZ75HV3WdnJLsCy+gIOugwZUdpRuDufSStk+TGraMlbJV34ZNZqWjcUrTDfi4gjQj8ZG337JszR7
ZwOAfDD85TkDydrxx4MMaEWfwutzWpXMda5arnj97v+B/IvfafjRPn1tTe+Tfnb8HzFIpEOg6QXO
pRrjLelsFoaIr2mqom5/5B56vQkL6zD7u1mV5ii6kOVMlV5uMH9z+YQh6Xchh36H+TRvdOtTKkfM
irTTQ0svcKcFTqQutmK72l/N3ifgHbMtK7vY05ZIazugq05aRxa66CoQJbfsXC7PhnEN5xUBfFiJ
BGUhCUI1+fhaum2g+zYq+matKm2Clznb9mnXikG3NLC6+v9nRRvOyEUGhgwjbnqVW4HwJ4jITbCT
t+OhMdjL22EqRAYUtTdsAC0MyQu3U0d4QF17W3Qsq79ELB5b3juX6vA4H8QwiRmfrw//2VnEQ7gr
OecgrA1hAYBuCOegVpEkQniW4P3dLOpbHPZej9k7Ojv3/jvDjUYiunxxZrQrAlrFvOFqHvgr2ciK
V50ZidMkQHheMIvjPXe3/2Uxq5qmWxdXMkuVlEEg6bksrUGwAXEy8xtofvS5YEXBW6edP76jM536
euzl9rlKf1BPsmDPWEJWJZ3w8QgDRwlwXvxA5jIkasj51ihHSumtpVTAleHHNUPzWdPeKx7pVnhX
TMlRcnvEDowD42byPoJY3vVripgvUdASvm4WlArkrRm+9nkfRUTQLWtoO4aD7BVKELzpoROius67
8IR99IBogkPb7b1cTr2o2ai6BmUE7KrxwBBgGI52q4wWBBfNcpCWs9Gij9t+RyIPMVCNpTfLA75W
hFhH/RiC7Mho0GBTHFFFfZYQOdMVzvaiRgkMVDe/Kh5tTTz086+pJvEBqm4XvdGhqILh4WVWG/BF
kT6Salm9eeSBxJQ6pIvhKAUiIDtXFf1KPuiBC2E97y79D/VagCBsilBqnSe6kwB279qh0hIFZJsS
I/QP3lg0Tv0xCsEToi6nEQhzB5y7A0BXYGQQW/xyDW5z2iTfvw7Ro4lgi73PXw4bSxFiPV37Pivy
d2aqN8YMPlcpDJeAk/TTtv8ke2WJBlivg9oZmFjk5pIxjaN+jtkqY248dnz3Qk6ZLr4J8GgDLJwL
16TqWnFmlSx22z12fyZ/8LSD2o45HRgG7xPgn+KyKg5FAypfhN2zgTJ1M+wVQwCp83n3csXLjO/c
9jaxrz+EJXgeAKnyHm7eh/j69r5XHqbLtQ3oaVp1Hp7o76r2pCM/ej3TZbv84AXK5Klr1sSBIAdH
qTlKKljMZcJ6m9hdIPni1rledpfQ2GDoX/U1uo7KeiKWEaS7aTdHbaAGJUxUG+85zJ7BA9ps6Pwf
8dO1qMn7vjzy4Uee3Es5D5XqLHipjWR52mW5w/xOYj81EyoJt1PiJhZUG6GAOCreSRL9AWyD8OEz
jZ7LQ1oj8UABFIVy2nAeFjDazDmN/mRV6aYhcuPemob9Zpamc3Y4AWKShI7XHFoM6a5hB/Mx46yE
9lh/GTy1wM3k9qUdT3WGAqZG3N+T2QlGEFZwxBoGND9AfhCXs33qsgeC7NdmmasjUA6HZDN4eWXK
95eZIMYvNvYm7teYCcYkGHiV5We8BPD4tW9ZZEGmVkHbJvbmNVGF3/bbFGCspM8tXhZlardKmRwO
TLLypps5+30PSlsgqt0M4TufCK7tHWaQcDoGi1Vj4jReR5ayT0qs+SGBM05h+O0facMQ6gHqcOuw
iBaS63BHy6yfKBTHwskdGJdp7lx0xuRMNpL9Nd5EXHLFn7+Ohy0wvvJfqGijlOsDKxgc7uIGQWcR
aO5S/WQxvnttj1pOQBLLZzCpImrknuTHNSBnHRLu0Om5CbUNluqysOCsN+2wJIe190vl86jcFj9E
0QUbOqyNCeJcvcRBzFzs6/VGTwD2CuqCx7v6oRKr0Cx+OepRcVTXj4w9RHICD6qUdK260r6IRDLk
6zXHPk8FK/X6y76toA8LJmjfCSQIhVmrS0UGO7/h3tC7D2zQqEcOBcq9Toj+8FkUvmcvEemA3OXy
JXgIfgxFmY8QpvMGLUkv/l49rmLO+zmtQlT/wA4HHXYIyLSMQ5m0MHOuJ1K169Af0uKmhR3Jov0R
16UbzZUM7Kd37P8DHjqo51D7ezgm2/kDsIkMm+uTGj9/2t3Ye9t9xRz2ZZH7raIlrcREkaDSXdnX
MMu4GznzgjbxnzHwUAoOmjBkwenB2tDAzPDGbwJI4fx0a1KBnL/JQQ7eOmKBmKlKAnb1mINb3AP0
tk2HZFLwiKxxKoRYsV4UjUejgBafX7j2aJ/5/LAvHwxqWShc5eCeNRuDSj3d8KE29tEZDRV0aUs8
CBJNpdl7aBaWDw/Pb9idt5TbKC5/myCZu8B9UE25BlsuGmVKArqdASmro/tQn8t+5ti9QuJjbmiZ
GbAT0Qty0N6EKo7MXMvhGBeMrv0moh9ABKN33F87I+1PBPeZPEeil7fQb/r/E/NnxPRn2c8umhN6
5EXqXmLkCAcjDoZ9gw1Uajb7H4GnLr8YysGmx8Ya94FxB/2z1zSdXfcC/krp3M/M5cwwDWf3DxPn
kuT5J5WayjKCzvOjfGidiWTwXRZeMnMQ+qJeePCvuP3Ko3CvxTNaBXo1whNYga8PVvoxfRkjKSUg
GSW9+1TAwZzxioPFihd7RMtFDl3TWNtVccOlNCRHmzzZd2GnH/Uyp9FboE3LaxkcqKZYsNf+3KDM
HPuO0oanCwmXhc5KXkZoSr9NTQ8yEEDeEBOTUZmr4hBTxqWEXa4NMdJ1qzRQp8+R7ez9D9Dl0jAG
Zy2qktrbfPsFroOZqSpRwI93X3q08XIGk2jskJQunp6HDedNF9FktbBZLI/j3gSo8W7RuXZFUsrV
f6ZNG5T+TK0NP4WnITm746iMPJwqoqYkfKLNxLPRWhLTRcOnaBT3fetWfNjI9tgtv0lftpQgsJB1
HfUs9GKv/fgmFaHyGqNpqfW59pCTIjHihoGLTWodR8cHcvqHT3KhFsFu1magWB088RgJF0iKPsBn
mb2nCyNHWqj4jqgNmfc3bsVAAatfHVU5W4JPeDO6dzITgpMC6a6kh5wMDWogolSgKxXnVNPoJc2Z
2I4g84DsmWRHstSMfFJyHG/MPI/vXmMvgHNnijX87uCH1bTFXQJ3cSxyP6DzdMZ66zNSIBpva3mB
SoePdV0T4rM3eW1xLwFai6wkdKs6AEo5/JpBSGiBW9nEIZ/qDtKE9r4j1fZQgHuQU8v/MtOJ5Ub2
gv4ozUzHoksNiVvWHPc/CoFe9cbWz3kuoPqb/NaOw9u2EfZlFgmAUKeBAYOEHrJeDjDY2RaXesIZ
SjChuCexgxSJyfANp61JAlnkzFcN75GVq9PyBZ0L4bDMpkj17jo9IOAZ/H0z5l8/arw5XydrsWy1
jigl6dGlOcnDdQnV1TcZ5kAcbzAMXqvS4Ruku5z2GL5C6ET8ooUA1xkKgC8/B26E5T4ZkqBdwDCj
+Tvyiko4I3OabFrT3QJVEkGppQNZ31+qs9OXj4kA/49fWiRbuuxxjPDOjE+sxJ8loOhsP2IQ5T9p
JzqvJe/cA7C0aCSQ6yB3admOb8at4PYaviMGnf7hlIaDjQsdjgnEK8fGM8YOXJIVGaBkrjdVT63t
vSRPsBNg2YexuDfUKo8W7Z3SCx3TdulgKtaUr57eVXRV9nLYA7hudYepZDi1tuYMMoBlNvA3H79/
nFcSbEicfYaDkB5V6W3GkPv4ug9OZn7XZDvfuJqDaApuyeB401DWeYDdoF8toGSLfguxp2aBoSrZ
laY3lSpQjTCRRtWJpovy6npENC4MthINKmHPLLYXJrXMh3SUEih24K0Kc0XJQoqR9AZsbMa2Rqem
9hJHelN7KYK7fm3s6b78rdxOPct3AXCgjrIw51AUZvBOEx9fpS86kENJNlOjopeet4OqVWRMG7ps
8heg8mYqwO31qHGJAzPRPfpgmgPfbqdHI2s9X7p6DBEOXZyr8m3x9TOjOgxsdQQnPsZuphX59DQd
qtN/tEY3hlrYPCC56gdB4k4EQP5rvyLIVnMRVZoDuympa4jbNY3cdJtcz6mhze2JK5awBBekI7YC
XkGmUJ5fmENM98iO4mVBCJjxsdPDwl1N6fTScNouvCtta3IgXd2sbHGhfLjH47BlTk5ft1bvseV6
ZUzGH+/RtlGCLUPMXp3hR1WwoOj3ZpcnVU4JhVbvoFMNJrLb6sKcRvhMwCGgG84myGrNDyhHtRFg
zVrBuTZXiApX4LVLq2C/hEAtFM7L58B9sSPzQ2s8dKt1svuMjMWW3nUfFhOJs+RwJq/QMYG7nHi7
MTfR+9UYMkTWEsS/8s2VoxR8EN+X6fDQoAOw8BuY3zEwuhd2wguXvZHlD+3sCE4nzdNkICuxheun
zZw+5OLk4oD+BgC2Xz8zo6fOuG5y+SJzEh10j9hmI4cFuPWB0NqboVCsNxj/lnPTyiLmbBLxTVUW
PhL8aX+N5gRXwjvRvv9FHFQ5wU+Tl8QSOoX6gnldPi30e6LbvrvVJfZYbRKXF+R6Lf2C/oNCuhfI
ugCLWzPkRc0oCns7RjZryQsEoJKx0Iv7LZGxU3r2e2WWb+cSy2c3KioO6KXtQ9WvnpyvhWmZMbhf
XPC3SV6x2W0HasOh94oYk1Sz4hv2r3PGPKQA17R1KGxdwwCk0LveMHWsY2XpkMDlgLlWAT3bo9NE
klNJxFSWwb8lTRTRdr8psCQ8x6DISVAuCgCSGneDRU0f25bv0KFBiSHtfNKSVigsrtsKTNUQVwkh
S96jYoAuN0ughQuS83qURbmFBpWhLCClVGhnZO6tuj+DvECDvEcr0eslqr7XQFJj19fzSYJvBSKj
4SUH7MQ5yj2CehQv7PYR2pn/9VbT6S06u/IRI3zA5PxWI8Izw7c966ATsMj5QDC5JGSQm42Oermn
XSXIAPqDKw2br0fab2noMdKoz/moq65x0Fr6HJzyWsosm7lbBFA0FtaqkLXOOiT/yPSt0WUzyvXs
x7KK9XCL3xD7kICmDOnIp1DxS0H7vTNrdZhajFm2vGQrXdMPvAUmaxd0XHuGQaG9pOh/Zus+XW2+
cwDZWScdHWOdwz4SBV2MobsUKNPxK61Iz19SPE3q2ZyNxe0P8YM6aKH8qjK9U0s2nb/gkSOYCl7q
N0B8bwC0dYFhUDt9RN3pfMTLWfEwu5WuwIoAFselIjX1BN4ibK/zPczOmX5BBivxLMCMg47G4nAr
18xpcX95pdqOSBVCNw2RAhZU+w7j4w+BiPhjTyUISYG+DeRfPOtEreTP6TsYCMHmr01VGDoWxKR0
0cH2+rA64Aqh3BNK79aasRRJ4HcUdVYOhc75zbu2tCGthNlF40QX3pnrbWpkuEty0EaQ3riHwFuA
sf4rLknOPsyBUW8WFEfh+iyxrhcFCnkqZ16ydEryw2omrbRY3qOjoEauot1DaIncCbeWFz0SCn4R
g1ijOkM/zyl04dlpXyQevW3lDXMAPtYksL03/l9jjPMi1mlbdKeMJjM3RwOjPN4zVXHrSjSO/yDz
LjvOMeMLZLR9PoJGNEHSYZ8ni7YvbQoa3LT1uW7lf0cntiN0QOoHRGT/xJLJlZe3fcbPMdRgil/k
WK6IRClRjF3aZRnzjE0xxJuusBCPmb6B7E0CasncABBUKC4kNMqAN747UprtvO2h8paqPwjuFPPu
flo2UMkR0hvbKxWuzacvFVbjiF0FtWzvb/ohwm04Awi0Y1ahAuwHHzOEM0+vzNxr0IDwxKoxhtyo
hkCVk7bY+4uUtC6KIgSgcGUjzfx6ahSm1LPQVdj2Yr95LGjzHrwwBoiW1LzzF+piF1GOTVVusVx6
AxGaq/0qt1ayFX2Y9kJr4LNEKYmBVik58YYlvgT2FlVpha5eOerb+DQ5lSgQRqvWaFaFauh3A1jE
EyqF8hlekMOKszH3K/4mczh+I5oUVNk+LMuiSF0tTewWrBWL0uLMungbvxOrQMI4kxyZljoLUJ18
WXjqG5qMcj/viOAOFJPVDhheqXEgaWN6UaAfIrCxr3pGtJpGUVGMT39OFOmrF9s7H6YSxIzw4vLt
yBF8wAwJ8IX+yVE46wOgomG60phfI8AfJSqky2YipvTcOTEggalnMwlelRDwFS1GWrblgNlH7HHW
5maV9lBnd6uW+9nkxg6GUhWwhwoQRDgqgwBcJVN8AhesiZ9+9aKWsVfNE7AuzUJkCdFtXKAftwlI
AbiqjZq5Bak5jZijLPgAXCxTESlZYJLBv+Z8iOjL5h0sOzc5dwBMizU++oTPpsTwijMah9XC2XAD
ZG/LYGBi+qmTFbuzOK163zxqujStOjwJqVFZKSSV9kVbvkKk4l0HXa+LbtI9MbwuNd+vrNjN32/5
BQ3ok3YC8BcSsm000pPURwgO3C0hbBdFHmXlaqwyioKmCmIuM8xvvLKUt5aiihLquEpVRkSAq7Mx
xKstt2DtLRyoxXsmHt9aARGZRYJdOmtuoe2Ng3mPFcmraU21CyA7m1tL5zHGTg52OraQGYZ74LfB
NlAgFBUi3OFz+w/OlpDRjQsx+mohJlkm3l53I5h/tvpGFlo/d+goWnZ8wpc6NQdkSp7f/Uy2N2/t
7M5boIgEZYyHPu7t/d81et1Q3P6/DxwCzpyXOuwDom3K8Vww/LXyRhN8dJkdHfyFUamfO3KmNu4E
VP/yU50LyJ3kTHuLMDbz4pXvki8jZWXdW90YPtwRx15bWABIPTy30zGmopwcPZEDlbzeRaDIUF9B
/ZSXzOZuDixRRbB4kakKQXo33eA0o2zvFwNJ7w5r4l2x0qLIi3uQx0SiDuR2mSU1PvfEb3jOCnLn
k1rUQsj5pFS4ZYiQ3juWgQuQB5O+gFfn0lHzwnX9+X3oZnMWlUgziT9nHubmjcCgJlpzJa0qsw22
x7fRsj3kJgpeAJa9e6j84p3I7ATx8u0C3kDzF3gv4CbM8n7jWVh9OpEpsnH67tlhjZGIbbFT40Py
v3HnFZklH9nxcyz8bWaQB7QFplqcqqh6RnGGA7UuxUPzBgmEOaxGIS7zRmUv36QuivhPBYsD1qWj
EUVvWuLMcG2Cz6h6cuY9gBqABvSjXze4rDqAUG/ZpyDmL4PBPjAePR87hgmLfl4Jj5jBmK2Oz31E
oJ3yjeolh1UVFf/xg1XnJiXO1ll7B+KEuArYwBBGnzZUTqflnDTppvfiKooWab1lkxxWcASmJo1E
DS4uSvWQ3ngqwQek78x+PD5n/MYwHcBho7pa94kSrK+mYJXl1hb3bYzTFEkaYbJIFUMphUzgl6g0
ibSoY2T0Gn5G890axw/J7YN+GYgA7pFpF90NGQ36u9MtGl3uw77rgCkfQEkpRIjcdgsdcXy8RBh4
lq8XAavgFVpUq4REQIQL0RQo+vSkuIt3yhV3E3lq13t6HNqdCwj+XwxovSCeYeCnuffvRTAAZ2P+
rx5KIpYAHSMMLh4Q82k9jdwUquZLWH29dc6vxc+LS63MQ2mXsnh1RiDAs2EUJwXpgN22vD0t+7RK
uLrG9acYuqRyEwQMsEj3E2SpG+MGg7P99Jejrpl6THdCUUNOyAmH6QkEFENTbshVKAiYgVArI2j7
7Zbz276P/Mf9lU33k+OEeh157d2dWxeJ+//aeHzho1f05w5icvB0OoNZw8pLlMWTUpJAN7heANMm
Im3GL/DN9BCi2ru7a4g5tgaAlaqZvYu5oV1AjaSzgJw4ckrm/6RzE+Ngk/4mwtYZGfaRrmmCOJJT
zmNu/xo8hY5z/yJZnxwVRUk766d9SLmAD/5QHSBm4OvMedidN5pHAGcrJJjipFx9Ws8PoKx0Bugw
l85bVi/DrSO1Cj13kwjQ3nP2hrLQg+KEE3r9iLW3XuxMjaYpvbq/LIDdo0k6NRSVuFxo86+QLI0K
a2wV3S+GqhMZexEMU9zQp4DdLb09QFyifBNBMVcevrZ2JJNj6HV/MXcmhCBc/11khTn0tmY1zjLp
0ULKJtP9cL+SiG/miN7YFFI7t7dQlg54nymnmAfkhuKSWpxEQ4H9TutotA48vPaL0+YcJ/GlmaSK
tALdYCKZqVogGmSwz8Q4BBH22zPlM8lYlTurM79mAlDczU1d2JtW2UrAH+h2OIGmcmcVoR0blXDf
MB4ePCDCCHUQE3tW3rZw78qPvqEwSXpizvTqJHs4fSunzoTaHwvpUl8tj5ywEK41ZIdD95h1b2jA
FPz9ImfaAcyJpGrJznBEZUDdDKv1NfjmQL2cuxf3iDfXDu3J0emrMoPo7+WjKqvE6+3CaV2XZ7zK
SrZ48XCt5sBoNhyBWjsFIZz+oImgzSHzylZLDfGeYhxiOnpArsfgUUwnsB4JBXSoqNBo5uFDa40n
crwydSDie9Te6QOOpoYMphIlFJh3sZI8DwLcKaByfWYVO9XLMHYuRfXz8Sri6cEQCLskygRaaYzV
rqJe23WycwRdReM05Hvh8+BK2GacsuRovFDr4TTRroVHL6mYSHjPkRPNl6b7ng35yvhtpCW+PDaQ
lOYdMUDKlRWk3PdmpcN9+65WTqNkcePIz93RnAFbE09HNfw3xfSN73ezcIs8zYA3ZHYc/ddZrjO+
tM/KKh1XCBGBr+jlt6GcRehFV0miwL8Uh5xxJYJbnDBLzYwqujKE37FAXXqtXAX+8HjDM+1KIXU9
Umx4MEk4h758oqNTE+jRnMQkvy9kvS7SFaBBfNj+rc6tIl8a5xaNwYjO8r4MIdN5/j8hIaL/+GUf
N6pE5/EWyxeGab46hRYoD0Qt+MOdWJuVzHDJQa41Qzfhm3v5i+xFuPMDmlaMTgnxDETwlJaXTroy
vWcTNoK3NfRv89v016/ogiSVSM78t+/0fhke6rdVy43Q5eXrQKfvRi7inOCYt8RCRAUG31sEn1J8
OJamj6m2NvivQCs1SyHsigu0LpO5b2Pg+sFI5q7oUz3dy/0fc61dVNkDPLZzlPefWmLp/OGmbiH3
F638jz785emeMTlbSuLLFbyKSkcb5AW0CjrYui/MG9brxtq6e2MBGqV8/UewEitawJlwZC6Ij5or
PwKpmJtzVveuaTECSuB0gBG4429rjoMM3X/xBMUq7pHISDDzlWVV99KwIQpmBRkV16kKV/QzV8cy
/mKM26ocIflWrlit4qwhLMxFsBtusAZ1eirOgRFTS4RSKgl3PDbkJ+RIbw9MJAi6sPiALKk/78Ck
K3UDrAvLbG23gEWbRAXJ4emwm5BoJBvt9B5zy90Pi8QuMoiNoA3a2qJid/MiAbAsPBoY9c2oSsVQ
C7OVRMP0/7Mlty+UXOGJWu/3XkMe7NZHOsARsA/40SkCtOswUuwQe88UlWGEtlz4e7WlkT0KWpyf
X3lNYJlyulf3XL/BdH6xBlbD1AvE4E/BepkXW0hMnzqNN7T4Z5urHJVnpGdzvrEX9pPbEmGi3xMG
1i1cxN/WzrNWoQIj94LV9WbaVzYHC3nAt31X887AJ5HeLBmole4chemQuJ8m8+W/p89h8kw2a0SZ
75zYJe4FiY6iYvaC1N+ZoIC0aGpzYKsDP/R0e+s1Z2NwH+int+sGPycIW8fpgPEm3oNdd6bcKynn
AbFwckTugOEIUxH9ljAMqK/HBd29zIpyl5r0Nyhj1k4rlXPVDYhI7KcoylwwjClzlRYdtwq0ewAr
f0wQx1p5RYbDRWm6nTKC82fiteSGerv5f66Lr/v1fzMqWxFsyJ9dHzmNrC3VrEpDS1WuDfIX3JWb
hK5CL8t0W66wNOK7e3CSmfgPw61s0vSqk8WAJr8p4ppPIVaIhmQkTYncKsPkc6EeE+gH8hbS4iV8
yAJ3RvwJQkcPU42U6QkEblNYvkERBa+Cfa5/bta+gAsqMuLAUzLS/N3DFTNmoiQ88SYbDSpmz4mR
dcliyhUiojRyg56ExH5EIFMknN7bYCNN46FiRe/vrAaJEEkmHZmlJxT8p3GnfodBNRpoLKrtCjj7
aoceWKFr036kMHXowO8nqk2seQLxH1JRoGwrbBpGr/StNJv9ZRi+J2HgC97CuK2Wj9Y2wdOOEqtp
NZ/GThGgryPerZpSQHSoYDXKA3NdpGxCdc/jfxhq4fVTFDD8CQUyES5IEV93r5mMVKrGvu4QRvt6
dz32Togqh1LChBF6x4MgILZoCzc2/og+l2q5EAydcseEHUgZpjjBGArPUHCr2Z7xY51Jyv2YXSa2
Htonobgx54CFcEwGyEWNfpHqhttCXd5QIK0vdrqOtnJGZgaMJWVB0taKoPbv7VqTsd1j/dIsurQg
CF2CixwC9qcUkrpMJA/hzsF7guO1AyUTK/eJqWXd4y63+UiRdv93oCQYBMwV66OsfICLEfsyAxf/
SMpC5z+nZqrrn53JFrR4MOamc13omrfkKcjp6FiPGUfaysGDdVuz/B/m4vppuMRDobQruqi/TQO2
MOdJlRKR/STg+xrrz4vgRFziAftnO553FcA9r3ZNwuVvcDi+VkKzOZgLeFUVgifiC5NzAiVSCcmx
XjApgva31sRzGDB6ugcZofHN3x3BXFWU7XiHVRTZpIgI2lF/V6Cohk0+ZVt6xQ5N8a/hrPoz/xcD
fLcpd/mw/Yyjz3A3PowIrkSBsCF/YS6Ydlw/mALbjbOvuQNcVaOkyUm53HFARgpPh+wJtUf6f0Qh
/NW4bn+H28ZwdM1sln911Lp4gbKRcqEAwZnZiVYRJYKLaAGCcS+mC6PVtavo0VOzEfpHYc7lzj7U
f3p92fUza+nSGj4OCsTIG9FnQkZHaztUxfxU1aN0ehZaWlkNKchkm8XbIDqtwJjq4Qg0wctjYZHt
VYSXHrswy7Aor4Wvxdiz3puMY47Ru0qGBGAH3bCec7Xe07gg6lmybB+T4K+FBPpICAJKtHnSTEDa
BFCng2UFvsdOUWX1pgIbwiOCyLEtitfemJZGouYwLBwidsE4kL3UgUT60LIJQdV+CyvySMnSQjFX
QNsDeYfuwXPNFw8SeO423jbBBDCrbUWqW75nCqkuPAVsr722jPcjwfwmgxjoTAlOgyK4PJHiA5p1
VJ7YpnrOhdAp7uKAK2+YNit3N6qFaKvPh4noPLyckKC9Vvos4Bff2t8X1uLQdPWLyxWEK04JwJYe
xEdIPNmv3mX70UlO4VHO2E1eQUJn4IcsbszQSNP4+IHRZSJr7rL4KsxBYlr2dyfxEPcGThcN89Df
s3q4RH4kg9u+wZ/p/0gmFfvKbebdbdT8+5pmXtAKzmpFExwa3dBxwWLvohQNx/bC3F0nnA09L265
QFNbqP5cCbj4fl7nkz7nmWn4RjEARURWXg878kDMBlWxz6Uwtro/sI6PKTwwig4Uta+tcciUGRY6
j3hlT0nzv56a5+zmRMxNw9gGzkR7f6QA9WbX2ppEqWLLjlmso55rroTggDbtU3+nGKGBLgsflizh
6ykWCLNO8AyEF6JeHRuqaWcU0yNs6hsl/p/2/OIlS4T+9T0zPLC1XOZjIo/9hyYvOWp/pBuCdSb5
SZDEQr14iXPdHCAppTFydvjlOzuuPtY4+OynOUNDbaIMiM1cspa08xGoEaVeUeNuEdKFXROBfg5I
pOaLLoaHEUn6Yx+YDNALg9edCEO5mEVihmAFTZY3J3z+xg2HDnZVbfUJeSNdyXdpGZjsP3nIXEEw
19qEboYvdSXTkrqiEz9cdTiekHiaeLAaNx/32KzDrDMoZiga0WwM/Tbkz4dwK2P2WTgj6ZkmECrM
bqCSgVVK1PoKDCA3u7blFzlIZBfw/9Az42jhjLhMpocyPwxTMme/ResBDHQbbyXsFHWDiwsFsrOr
1s86penSeVah+vDI20QeDj+r3MobstUHwxlpbpuaiMqEycgJFN8PecqX32j1V8onFdEUzA3ssuBu
TseGSD5/W/pX1NxQtNRFXnSA1WwIENsuIu94gzdi7Qlrn2ZVzVhAGpdzhr9K/wlIqe2xRBeo0IQf
DvynFAGMvxovvZZZLHdZtzAeSZ2PG2+0GveUSuGEOJXAbYrnfB/eHbrzW32nSezpUH+uNO/Oyu+/
tA2aim+7oy6J5TeOMsCFAbWBqw1IHoOQ0pP1/4OTqbUTi9+3eUBUkARyL6+XoC6jPkhckLQkISF2
IqLTZT+ih5jsLeX/+vU//OH0a79NV3ZX1WJkY+DHHS+N78LZ/U7uKt5lAu+ketobSFclc3jKmoFc
h+hEHcMAvFmQhgCdSuz3UvbccsHPEDlXEAof7htRX0oDKWpRM00imrDMoP+v+D8j8nBG8SoQqLOn
+dAOd138KYpWyDy0y6Xfd5X9SeYfEe/dtY54ZwZhJOwVLPCbdKjAFYoyfR1cnq/r2Jyp29Ufq02N
rljeFK3Q0TX3EhskjrdNGxXSwKUaN5Fy9k/4n2NBXHqb4Id7910HIGg86UvvNdge33dOCABiPkUk
nGVIqLZF6E9vpU95wRKKmAZfjkX0fHLQeUwsUik0PRS8ApJESDaJmFMHBv+kPoNP+laPqUzaJmYu
OfCyljUtKid9u/bAkCwLfj4q3VZISJHAD4VME5KgB2C7dBophROg0X8zioTO9lfvVUye0F7Cauk3
xopWf45Vq4KF++iOOMNoViq/s1jsfE3GgCQ0J/Cxw5k1ry4uGX1S0gAibo9UQIwMjDG7QHcsID6/
bsX69VKLnRrJbcJvxDoKD5uTgNSuaAKaQNyLOlkEg5iCe8MJ4l5gtf3XYOOVFnpRVtLefNY6Qr7+
MVldvcZZjlhvlUwxg8l6Qt25PmuFAasBvssyNO4osvs+4zUKk3Q/0TmlIrfw7wZZ/+J4lkLBXzan
Q8ygGV0/mH/XmKkTXf1u9IAn0epJIIgzgFM1ute4Vvq4wZaRYJP7V6FQLumKv8ooGHRyWdXjNcDu
0VZ2Ma3PS++TwYXSWLA1Oz8BBZ6eddZaxTgWJNxwgVr5h5fg4kbLCIVv7RZgNm2B+AQ379D0zkgz
O0ZdaumudIeCB17chSLC2Z2smB0q4TAfbu69QH5z+fTtK8WHz80V77ndhLo8EZgPNtBJj1PyteCp
uuysYlMoE8c+4awGc0Qt1Gd4RZRluCZJZ3pXmeQx2AxnC5hsZZaSlYmSEdCv2eslieuyBU9e8q2X
AV1nWrKwoYboJDlT3Y+y9lc8ozlUwxHCrCwyiHsZe8nqyEL+xMhSuh9yUniXvnmP9r6azDpo3DQh
zpSel5Bo+nkdLLupkKkp7IUOkWNMeY8FrA4CADNhTk8PRjosI+i/YxjL5mrT4ufe5qBK+xbqyYD7
1rgCBgKVVU78LnKvg3+PAf3Co9QBwa+qkZjnU0HCu9crQdnwb+epHdkW7YRDUzckkGcxYIUctto2
4ApWQT60d/XAJPFuxiwG40LAPr/z4sIxwWaupFhjSMyTGpkwRK9zZ9f7qiu0Eb1BCK8w8XWENYiM
iRp99FPsCDBekCmdY746FWaYRiKPQQIAicJiajOaHrcOV67M3tZtsxVJS6ho6g59YS2Q1OffXm2a
NI83OrHC0ZLihj2cxBP3Xrxz3a3KCzsA2xzc/xm+J4e5ZaIsNCTSYUfQ+EbvrIpqELOe97lPAgsc
sipIUmuJWedTYeRUX2aWb3xLm7Jy/2tlmY4qRmv74KRJ2sfUFfdTSuwbrkOuk4YSGOUqDv1V5ZQw
eBkwuPziivRf8z7ylf0sYUtN8PjO73MA6FPMTSRKgbWjCzeEgpKWlE6yYzt8Vq0xf7o89H9XU3CR
o3AXWdwTmrR/QpYOkRgEQ7boqg2h9eTjHZx2xbzhE09yenINorpSwh6XPBKqVIFZqv1nrVg9rPK9
sxH1HZFpqjDYAUGIfhZCwEnrUFtyGPLxyFAgw5nuoZGy9s82tFtmNEcbR0nGnZ+9s/xO4f2VXCUi
YEVoZJt5f0PeVGzIva5dGsxr9rdRhzRfiAVYzv2dwadL7FQO1GCB7JU3Bql3grTawbja4H4mD/vR
tImKsXjh8wp/N0mXnfMO6FnqcQL0dNbm2eHl3UrgU2qAptXAqQlPdV9s480YOsdqoCBP3hUWVqxJ
MJicJrmu5UnGHXSeLTXpMXzldBMemdBrTiAXuv5PFjIDABlp50MR4ZmHdzJ9k31UcADg4U9Ab8f8
6xfG2yPUml7wNr2d091C1Mh2VIwyHysaQ2kKXJbHUE3+85OVyjV6uQkbOme51wOFGqYg3C/RP9lP
Iz5RaF31DsNNjHPNft6wjlhgxyX5wOXnoxfoEPWuOhIQwRq5yb9vT1RVGAr3lxbZ1eojVobQPRqQ
GhNO3r5Pq9+EiKD2mqXWMgpNGEF4NYv32CMZ+T+bsDcU+pPO7jN5nJQ+LvXgFQA1GbKnCW1QfR+j
keVBZjlCLt4bhzGYCE6xuFicbJeUJzHUz6jQtnV1aDAtFUFMg/bDdA0GgJD/DGeDI/h5M5bTX+CI
7/SOh/cms6s+n9wGgtQ5I9DUtgD+xKP0z6ZvPTq9r/OnJRba9TUwMK9iohPGxQB4XhE3wxEfHxPk
ryDBdfBS/Xq0jPqoksYOUvQtyg6OUuWzqNOsV8x4RzfzPLdhWFZJt3lVIfRmpHeueMmf20jSR1MA
jvjs7fwruUyzk0polsBYbBOPn6YuPAJwztWXwz+K6adXGs/hHgGjFSlx+KkTSwmh3IpVgacyXtzw
9k0QncTKgVvowYenZAhLZJAt7pFoccKs0xLjUS6s8C5iZLiODwZVFLPwyHL2UpVZgrCcuhjrs7h0
cwX8Vij6zj1WNQFaeRe1SUKamx2Gtlt7Er8j7dig+bZSJDKf08do/8CaqztscD72vOEvgyDBQEUe
aBR375C/85XM4iOdBNVXhR3Z/HSO6u8C8rRu0pAETJxhzOytgUri/zGvTnPRGQA70B9cXyukjvtO
qFAlN7wpgY/WjRQdNIBcOYvl3yqgOvtX182fb4F+JteCGKbTADUL4TDNL31aAqX1sXVm//fYTY+w
U4jlPpEXM0oepbbX52SlV7Ww3GctKIklymx9qp6EMnmmOHL3If3KTDqz1QARVIQtujkBt5cJGM42
cVCurlFzfNUxDv/6n4tALGwmD1vesn15f/OfPJLphRJQcEgLjeqtO9jkJWc75xbdksnchS/ITU/2
SPpzqNnbD0lrdeLMaZAppBRkK2gupFn34gyJYoBQB7YJxJOu8otoYu3jbBuN/VYI5rCUvE3I3wOw
dhV6Mm+Wqmn3hbOAL9Wuc4hq5L899PPTkvhr5d/RLH5rQ/JLgwr8s3v7qg3F3cFd/6VQ6d3LxoA0
Zde8bWIsOKEH4W5NPfZXhuHrmWMOGI9uEob2WHpS9ZNzh/WG7q35LYBiqif3AiuP3OW81/wvAEDj
6LZ5O8VJfAONKlVc2ZkQgwkQnUQTdqcIYmh2j2LmrEJA7Bh/rINHrhQ97Jik7Do5F34hp7usQTkZ
1/HJem4omCsktWKmq0mLZ2T+BkTBTNCncbDXcr46MpIscRFoPQy5ZyXPijKgdhXJthkOaD/VKAKT
LikYl8EsWoQPjH8mnwfTWkbEXdMGy0mw2ZS1kUqOzbwr3yidKOY7rLNcK1VHcIO+EaRq6X4YniMl
wUkfkVC6r7BRVPiDaA3H7DxYqQF5ESXo8Kik+jbeVDlY8b9sCy2Tq3C19gTSvYwVfBK5DIb9/RPS
M9QY6573zRfCN/L02ZHPgFVk/xBsSPuE89fPMdalv0x+bRCQ2xXm/bOLO9jtJC/Jafyi/o9y8bTZ
wMUgrEUNzpDlRW4nWsOVo/nMBd1XDjcVUbpGPhA3PWW2+PaYQCnl5Zb0YCEHEqSOFuLjnVSBXw5M
7ymS2e8gxBx7J1ehw0jupEW6ySpNJuXN1DqTfOJsmw8PGw+eaHUTJXqxMVhg/Xt5GLP1z8TBByNf
urWNIF/d6FVcq91YS6bFaMUIt2guz2YLew0gtE+clnC9iSKWzF6u4lw0mNEqLtheBcGCi/MTtrlI
G36i/CrwN12JNXwwrfdQdbPVDKfzAAtwv0rH6hojfBhM+h3e87W9jYlp361XdMCYC72rFsOlKXOQ
ZXM0e25efFI9eiXdPnLpqdXhd/nYOWqaLxrBqfL4X4a8O9L/SGurWVAG9dhyc6T64X2vh9G61ZpH
DY2hJfbheYdESxICLhRMKUdGs8WXhzNTsTSCkRWuObwN7f9ESqY9+qSaCORqqvleqapDM91lwzzZ
U3gUo6j3RNC0T0l7us+p9zJgUPs1regkLEAEp7wC+po4uWV3WHLW+hXYZfgoCXVWFiS9webBtdS5
zH9vLH6Mh+Q0yDKs5N9MGA6cJCLJsyyPSOVbkWH0wvrdc1+nNV9yRAdKWSKBDAVBjwG/VMlYvYgm
dGEACLvDdmb12DTjrL6/5vV/+0Wn9391v7fLtmnc0Tl5FliCtdJgnsauYVM2fp+v6jz3xoCgAzJh
zwvKJF/+5vPJ6KQBaFxrdh628KY5i86OlAfHMmI73R54mcJ+aRuGuaw6IXABF/uTxWqgRwp4pYYe
V2OFCtpeTtpPod7OGyONYzlXOXbpACnNkdjYERNFeL9RxsRiYz5VOuSnAwOq1Gu/D2109VttfJ2G
hCWKf5WP2NsGHHNbkQG7BCKDm49UUV38ErRO2B5gdOnMNoITuJEqgQ1A9wCa5RpYAOMdGFrmR46W
zzHoH2olmAQPJe9wOQvWNbC/4Xa7eJVbC0oPtuzOzkyok3fa2V+Us3XtZI2wnGXXkyYOCkEsKK0C
xSlWXi45yZOJAjF35eOWdL5p5zOPlo65hrKJFB9oxr0txZ0iUAYy9i/HYaXgQOQUaYAQyZii1xMe
wfDzHei/+o9XXELfg+b5Z42dINjNPSzVAjVd73H1L1Au8rdHq7JI3tmNRzxVxW0UqIDPwG23xRSH
gjuIpq9WmBXjlLzScze8tOUe8cQXrxp9AIaN/upgAkG1bn8O+XfTQLUv2uW61nQ0NOZrKZNAKupt
w90lGLAidjClVI5EQWu4py/j6W03OEEfFSBiVjvG3Hk8TcAiR2l7ZHmDf+zKiVVpqbCDiXotBzOx
ox44kLzMIqf11YunXUZWpQ5zZoJ/Wd4NvagPvwfy4svZHx5nw1I8pXjlcK97PS0Y7/sZyU9T3Aii
8HZRVaBwpIRV8vwBrVnoNImk0VZvve3VmiNeCdSnHt/yjSRLRSf+LZwF2Xq5MF2wFBxzBa2AQVX/
4SH4QW+iZ/8Wvfnj1XpiHFxoq+YSuMZeq3eXZi186yudYdxHfPshv9/tXiQs2DV1wF5ZCHoxnaC3
eVouz1Dd6RvbB4Q8zGXOpTbjjyJ4oZFJ0KyT5lnv+bsU+MVwMUyAFwLjecWJbvoduTk+R2/R15Hf
GJ1ZAZiVp22o7nbfBXDRxEpPqwFSOrIu2AMvqyQND4nxKSIybWUuD1y1HH7WgZLyzcLfuPpaUoRI
0ge2/wwF1qN+GMsdnH15/a1OijGdDwR4kZvm9tzNUwVBTZQeNtpU707Q+YH175nF5Naguplv5Dsk
/53VczH0CVe/I0cpPpGB5edXrjDJVfrHd+AFC/E1zeFs0lIJ40Z4a2mB8WCNOtjx7vWRp1te6m6/
OgBYaZWS7FvFl3TAFIemSEtrAVBzcIX07X2HBwCvu3MdMKL8/np75USjKP77TSPRGXHNWCXnK8+i
PpGey5ifOWqJb+ayn2aTu3dZr8/YInYHFtm41DZMQFsJMNHiofNsgk+k9x9/ZlAw5KEpkwPiKlCx
8RvxfKujEc8STOb+OG8XNJEO3gYSO+p5uzWN4mg6JTfP9Q2trWl8L5trQXq/nCoUVqKO5FiThR8I
Xo+DOIdXgrESZEGmg2sWqPXb9vgmH6y0mI2kEcIqo1+UvR6xRRGneaDzAsRFbx5jGDnIihaGgj/1
PveJNrQmJZmN9CUcYWA9XSIGtdQp9spm+zo4WvlICLu23loYCd+BZl9i/h05DVypKPPNa+ct+3hK
jltp2TD1CMAt0hsC9bKwFqkUFFaofOtJdg1+oZGHJb4HQ4xiLo0DWkZl1Vmrt3de7zOAo5NcFwdl
Oz3awlG1+7VGDbuCeMTsn95kAUgXcTqxZ779w8HB68CQkvZxrqiHVd9ER510uNGfcxa6yZLhAuad
O6tdMcTjNkAuGl/ne8+y7PHuPbuCJoPAcz8AzZqqTS8m9bPct3FEk2SQhb8rEXfKutdQzyVsD+xh
5mE2TN8N8fefKHVdnlkj+be0oSJkILvDM0yN4a7fAB2NPY38XRpPof88qv8fUoqUKVCUTrX5ClZT
uwwudK8q7M0aUmOJAq8XCeg5YlhaRVDYh3hWvN01Mjx8zj2aHOFGIemb5yXFVdTlZxxXEZRtHXhU
uLDT9cGETniPtYNCRcR0CpVXSnO1FPdgkTVeEBWvJT6Cd7wbBpaEodlQ0/wcRp5j9oShgPRA4IF8
kOEZ7YCCi7tyR5AtIJ1Weoq0Y7grT+teUp2xGlWbkcfR1LOB6wmcauRUd0qTNVLH7J/GblD1vfob
xse7QlYAcw+uNrnKoHdR/PfrWySpP+/NLDo+FATLTvo+E3ht11C+BdRX5wijNBZvqahhwOIHdS5S
7wQMO2YSPp2Kkn854KfLZ+LLrJsdIheKoujUt9hOrbbEGaouc/uGsSPzYFrcO3Cdbs7MeKPHGLK4
HIHv9QUId+1Wm91pGB/jbQfk174yJBBxtrhSjle66lYz67tu994/46+H5W3xJUSBuslu5vCT2VOU
jzPBGZQsodvxx9dgEvVaylydVdNiVqJz5LueUGy0EpNx3cSCZ7twzsZh4bon5sLT/0kNCq5DZ8Tz
x5uyIXe5gs9DQlyzACNmaHa80p2JF/MAhfYjQaoOjh6jNvjd+2Sy7RoKWpBvuyQH2F4gWNHLA7z0
v55dkV5BgwAP4aq5haD0+lR8oW3sI5ulVxWmanEq/O0dIJG64HwT6bUZV9zP1C3U8RH0TiwgFIq+
5cm3rTuRq6PmghBoDP+aFKBvmeOUeiXC2bijmbMbE7Ux5GjR2zCNQBVhU9XzgzblG3tMj08/gyOg
6ozYQIHR8F1W3jkU2sKBb5zHVBlqx5ppgKW1Jvx0MhM6jEclZmTxHYBOJeFTo2QnyiRPhCZ/nMn2
0Jgh1hIwtAG11vKV7H46pD6t9i47IAn3LQqwYmyltrPPWzrgYnrfYLJXoR3xzaGhzQePcz8iU3Cl
33kR5LIIWR+91RospBVGeIiBo82qwCA3UBeFAIJjFB3ieVkQcs6Yf3n/mRHw+Ox9AWRN2dfIV2Or
P31rchtj5ZYsgb5im2QQS7SK4l7A61xoDxeNlRoy782Of3V2ukarvit3+54SogxZbJGjZdTCiDw5
qztVhpBwwdbqK5muLxJVKMTnu7GrBSp/GOlZVmG8gAG3cxqoQH4bPv2pN2b2goNG5T2+c5KvPUoR
413Rmj3bihxGZhR+wrqL5Fron2LbC60FmTXTyySnANpwdQzm5SwopXTY/KkDRERYNk8GinMWbhfv
ioLK3S2x/EPA0w5XNz15/NOB1dAqKMR8l5/vrpzLr1LICEm3KlQo8l0ABc/zeVPNYwGznCvrKg0F
D/Ua7/XalayxV/00Jg6G1NILDsZ3o4HzDeNtwhrbiyDwYd5oqL8zrdwmmOh5E6Ks2dRJH78KjcDy
bDCVBDOCRlVQujFJbNT7d4jS+QpbNBAtsbu6O8R/HVy7jnEEK01ty8wKIbTHBHWFzKbgDChdRQ6G
5Ua5E7Bagq2KewwwwqRcCvTEnQmAIjNUhrBB/GBqyMmb9ArdTnUWyJtYC0uxx9ymmGqRrrlkSKH7
aXfHIQT53pzfEwlculY6JoyozuNCa1tsV/kcm1jWxHTcehi6jwt+Q7OYPSeAT+lSkrs8zEgtHUJ5
XqWnDKViN2zE0QcWDptwjmZ58L+C/Ju02ftGthll/4aceGOGeJYLUB0wfvpSD6uCDeI5mB6pyqeV
dlIHu8V7USGQFitapgglnokWd/uG6WQfhGqNcclt3+UUFaG2p5h7wcAxMTwTwYA75GP5ZDGYiyMM
fKPSatIIicV8wNvY84KD22X0qjieyigGk3KbaRI2G2TKs0MR8U+hSpeCnKMapmZ6ekNRcLUrlSvK
EzKL1Hnkt9FkFqtl1VYjPXclM4lMEJm4fGs/ZlA68R1vaZH1tCCGlHgUQ8a7ErLTBmAXHk0odpxs
ODYbXwEUWDwqxjmVGaPxPnTI7+GZhMp195CH/NGEiZDrws5AbucPZ08qrCWcgENUNrZlaMhKBuW7
TIHgTrPZSo+20Cf+wBLpwwvZKVQXgcHDmkKL2VfCP5QjXfZizpuTK3LOpqWqxalkYuee7HmLC2gW
RArzz2hI/+mMtRjjrSFDzX6iADTF9MVKhq5RDllzM8YSaEjyT5vPsi8fjSAo7W6KNVp+3DF+Js2c
+w0smek+3aOqYtsAqF5usogcJk9U+T30Dy1qbaDHK8G8UJ+hGzfoyI01V58HrLPbLFDUzoKDUUh8
Wg/EkMImBIAA/1MldJw/afpR1Jseic6pPYCQNmeoA0SivWYtckqnyalb+J4nCjz9aleuvYeyUV26
EHO4+GBJE9HvUIcJir7IYchwgO2TZv67OdDQrWCQkRcPY+BPINS70LN0nvHC+4L9Lo3zbNYtSmG0
AZATfpBWmspzqfEM2P2SywXJafZJqhNTZcNUm70niK5oDQdISUKs7XltIEnMufxLo53wiv7nxCh3
YZDjpL2oJif0+e3O++FeNs+TfHJW4gNpZ1JqVXNdaj4rR1rg4bbO7lDNZo87ZvHxjXjS/++CJAUU
FW4O5zH/NN1VFfSU12d/b430umpJTpjY0CPUCa3PZ50sVz9N+H2PUmHlP67+5t9BJwQswMvd3ZbH
AM/SCk0S6Hy3eyjBIP/ivOr9ORQ7RzezgozabnTFVkCxmUZzBVcsi6gY64e804OkERyRx94kW4Ao
2DDcxgOSER9c72UwVkeMDGY7CZfp0vhZng4ha7afABfaXTzaBfLkt7Kw6+tPUQKV1YapNEr0+MiD
273XX/xivsJ2+tjRn7KX6EcZXhRpmypV0sF9U7gRNKuRLu2gQG9CJfe5g12OBaZ7SuQe1+CGe6g6
UH4wR2qlM9IE+udlJFcYkU4PshtmX4/UVlMMzWKjn/Rc34tqonYCuO9I3vkvfOuapMcRpuVlUEU/
gK6+UQC5bYYDXtRzoFavGHoyj+0F6nP6OsK/qTXBBmoq4BQvWjvcKn4/rkeoy9YGmv0gd6AOljvb
0IKgj7jlDt0NfaNBd0BRq0E4BPp3AQNPKGzQZ8t5QaYuL569KezrZV5eltAZEm/pwVBBihJO/4vA
J+68VlqoIuasX6ce6CotsLvHCM9kzo8XtftDaQaDJra3Uj6c7zLzxKT7tkRC3K2NARHalrpENRd1
Fdn71h3tAvGh5B8vr3SqhfTBOCyDYViSXzg47atcpiXOBaXjEU67SB9Ie5shPMy6CeLvuls8pQvj
iRFkY1M0xmHb2QmG8AFScp4geNqpwrWVRrlu6J4wgLIsm9CAyXbMB0rQUANR+ic3XEYaifgud/7Q
hThvjL3QfyS+tl4ET3/5DMf0gXNGpdme1n9Vs8KtYKn4J956k6o7hYUP4jFxVAYhQxgoJnd+PAjd
cGE4PF/9IMYyq6W7SJn/ck0d094SFI+4tX5+398/w+pPDaJ1abpzGKSdd8aZTmIsp3hkB+hI2So+
MDPjzpoO0g8cdQsVzPBJpa8sp1QWD3tr8fYirofhI/8haXQhUZ7B+N+PvwwKE6rzescHb4zlZbtH
c9TOdD2bxcneTkUclL/iA4g9oeIBIkZVfLMcDFdx0WUDtmGUqlMSm8tLujz3wabhNIOTXx0N94wY
q/Ey0mx1kPjYMk+Lo77j1NebBDh6cnuL7r7NCSMttG4ri76Xpn8nBxd4QL2Ve/njFZrZ2bp5e1Xo
317le+lHp2fJHPid08bSU+xeuMSXnP/IHsJ3KzW2BldN2uK+Pmk0ETFpK1PVQQc7BgPEOVOr679U
kfEONJZz9ga5fHq3QnBoZf62ygEPWoYQTPb6L9Bx5dM0yll/qOyCAXB8dUxgipPjWrYJGYBrKgZx
dBP3I9c0/z/YQlLTlptjr7Tdt09I2B0DrJIs2Vp87kQHuq13hoaSMnMOhk8jM6IUsiLOfWHBiLM/
pyQC0XPyhJLF3kbzNndIEjHh1uAKzMWyvua9FoeqNSYudPY1WFItgpQFAUu7zDqnHa6OKLTTbv83
Va3LPMsRiGiQAD5tQOV3mWD1x0iaoI5yC00Z5iqRPk/iNCdPuApqItd5Erv8tBY1WBGmg6vNT+41
eAnFR529hESMlXfidDP+d+oh7HKi/4UVwJNKqVsyoiwC+zO2cpae3t7gH9AWEp1CRxcOWka9e62V
jdMPae/6ox/DfpM5VXshq5dbo+AGzqRFXoSpzKevxZjdk3Y/gi1ErC5sr7odwvNoR9EdLGdmzgS6
kvO707vkFCzMS14wFnaHEUgyG6n8Hz2A9ZUsHlYLGnG/pJE6C5TJjtp3MVyuD3GkvHBpYUWziQC4
+5f6skxFj9tlH1S3dPppO35buJpcBg9ZJDdPIL1sTYleugTVhEcZo/yseQIFAjcqwrxyGw/pHJVi
lMFKnN/FJQHWnKdJX+ql79Qppnzl7npY7mbShDt1DwlP26Oc9SHlvDTysvpK5M0HyToaDn2uqvBa
mljvs+kuEX5RwUmt07hegc74yrGL0QLPkAtxZhIPHDhX7F3x4rUmVezzO+/gfHOdm61DOCGKmdcu
jFshrJmHDnNV5ozSZVdGcRb9Pm3e53OC+tUoHgmkaquA4tzzBjXbRTFH+EHB9RCtioETUP46Dvq9
vyr1cG9icSEz1eaOtBmn1zzL6OcwucFZOHHq7/aMwKa7tvPh9ClRt7rCtalblIVNXnc067awDIfm
gsSWO9sMgom9J8oKCe2r4wXQJduZ+Bgj4x6g7zBY+JGx+ae99IyoLgQSEfsXNHlM92kGNaFSv+70
bdHjokEPG1QYx3k6/jPYihCeqH/JZVFQGp/gMNDGapLkVE4xS/5i17Dc2f9xHi6j5B29wH2E9rYE
2iSKpUqZiKzrlwhXyXJ1QMhE4PRPqimrCwe9R4fD8jKtmMBXI6kweNUi3HQ8zXN4vR3ZKt14CIn9
MWvnhd0P8rvo6/G32VomcE+o1PCbCOo17KzSpetyhFxFeB6GtNkrsESybTkIJKmwEJ0jI7f5Lodb
3jbFTGMwgja3nJPNqbyf2kW+ImmJHLTd3ew2yLWum7FUH6M7hKpES6GPficdbsdGcTYjYr6tibO2
HMTuWarhKGbOvmTkKFmsF0FFX53E5X54wcn6B9HUXBUpS1Bx7euL7z0HQhp6U5w5JLFzny/knuWk
VOAGeTtSEfAb8L4FzT4AKbXNZ2OxEs7mCeCCQdlMkBy3iHSIt0QoGx9UzD/PW9dyZtmkXuDuKW1O
coAiwuS0o/DNgcEFpGeEn1vJ0B1pp1zPR57NbatxeOv13yXpdKc2v6gtiO6UI58QCs8UoFrdgT14
fztuoXkx6sKxDSyepDG7kjx0xHCASk9kPl0uivVXxjQMPxJogBgvCH1puRfXgL/jGtm7h9U/1bV6
BqxIsR7JDT8RiIe6xeYVOHBGBhPvKVX10roJ88ZvdHSn1ov4RiinB8g4zDWnJ6phrr4NJ1cBcbiS
xu0Ky4cH/oe/2LIIOCYfkePnzYqA0mFsJihc4qbtf5tSP81pUZSI9CJJZ44pzmo+m9JqoY22BTOI
YDmEnLC6A7CJY5wHenkDFUaxiUn+C+b37khkiTWB5sZQXjJrK49rnmcWsc9MU5NIw/1wsHHyh7Dh
QtiXNi7qn5jEp/Q7ARfoVQtTC10AYMLme9Wvy5CTBGmts8Qlnpoe/cweEZQUik7kJICKibdSvM7j
qg5bEUd8L9PzzNQjwy8jaj4e9VKLpSmMyhQS8bOCrSdqCHcTt1eSh/SbuQhNH7s5AkWPHiL5CuEp
hP2XEztEWD5sb1k70nT/Rsz9eRiEhHo7g8I51GNpl1agtoggeB5OzNO2rQPz/oaIII0vq21MIeAJ
07yy9FwfTBmRZtdMTVei0kRVhma/0YHm2epDlC6EO8aCKuiSFa43aJuMihEfJjzzYVVfrjkmcZKx
GFWILrMulLmtyWKXQ667Uw79jIwc5RdxLn0H1p7rIRt5u6IVzEU/TltMT8OajotyDIZz1XF2H4vr
taRX2QjiFbeXpcvA0fZJ4InqYM+fzpUc9xUq5tj6o1UJ/EuK+zkOqp7D8VPhzB37y0C79s8a27Mt
gge2jxa86Ifjv5IDBCgptJ5QxQBMI2JElNjVRYnEx3hlUB1BIMU3CfB7TS83CvT6KoRQI4D8JuhQ
nqe7ozM9SS6k5IV9hVhHksZkVtboT30LLLLwtfcIGPx9XEsusRW+OME3fw62d7FBIaB+SsPOax32
w985VFMV9QdD5ANOqRdDuWEfsIlsTaUMrOx8iAsX59YeNJ6Gq6je1p45MnOiHwkJiEugD6Iq+vea
xfzH+76XtytuRGlQsyr5kBM8f2T6zdwQZ5Sm0Y8CfuYxhonYsF6oSg7XvtgZ6PFrnMyeliUMbWHE
s7rqNCbZY4hkFnIIbrbmxviN3g2yCfBeI2Pbug+XriHtyQU55bV8gexst4vBIXfQeZS0Dj6/NhXx
75WNwM5N0yGPrwtJ+FKJH4nAHUTenXEGN6jRN9KxDKStJ0Gd8CfRgDpDHX6N/D4rU9FLYdPSCu44
X/Wgykrr5lLpi0wWGk2jF+dXSlYyLekB9APzZimk+BlGX1M8h8Vafxna0Tet/ApFTSqceUhFH5WE
1VLxN8Vt6Rf3QBpC3aUKKe4zhe09cjnaKmrl1i6BVN0jU9G9k8aFDtVe0bveOPNyuj3hDFl2Edwx
GzLBjm7qnG+jLvJtel9Pgx0prkM827hUnKR6wT2Oi5fVZdJbPdy/0zOfEhh1aj4Fnp9tzlucpXhQ
R3uo3fscZOQz4O2/YTRcqETyaCOSdzyd6LcwYthcpvq9d062seDU44+SjRiXVwm1HJnVhArDscVZ
j1v84AkanbYhIW7lZjIuXSBiK/QR166qiRq3LMEAuXhoyOnuTqWYlMulMQ2AoWWJNGotDEYZT9qD
NOgBNYGPbuYMtwxGkbuyH8YkO9EGPQ0p4datSwDbTc+/e9MezMpeXePTMVl+VZuCq5W6GvdD98m6
PVjz2SqK1O64z1FeydI9TJHWxv5MENPZm/yXVmxUVqWBLML/yFkR4XnWpebNqYEU6pi1so0nDfPq
ds++VXf8S0fmTH6bUhWV17uvL87LkEwKldJs31gxNViHEdo+QLZwncVMUIihCiT5GTe7giBvA3fA
L2sWRrAXRkHT7pVWRENVzXnXRlf6k1J07fuHZLgoEzx4la1Ho2u5/hoeubLpapGdScwE0LJuReJW
DepRZMd6pmZEiQ+rvvMg91OtsiP+b7VKs3hbdr1tPl+rAoVs1fTmNkNaCACTDQRiywfudbeci3dk
U6u0HTnbP+AOZwgHiWcwXrsQ1NcFqLBQK/ePBxFC3a+zM2U1rBD1y9SImLOPH8gdUUPN5WFLTNrX
JVwFcAYLuOXRx6i8ShdYK7BYCkmxQ+z67QCLVYOGOng1UmeNUtU2pkgwDyjq5d8Tvh/QfFbzJAy+
c4lR+7qjyvbFdHx8jkpimhXOikx3HjDdmnMA9X+q51yJqNrqVfiVlIFQJOHZEUKJOPJZLdAgR/nm
Kuqyb/Oiehd6FxDNgpQTQOIT9qH6BIAWS0H5qIqD8EeDsDFdauNcZhkHqzyhl864DrBzdDzvmfy6
0/G+xmMP9AM32cxrokxT6pWn9JmDz6lxd+mLZHh6HjKtaXHQGMcvzPkuSD3g2ajl+Ft1eCsp4yGU
m7LSs7i91nUe05Ybm/s3+MTowqdNlbAXQooyCKrkKaAqcV4ti+MCiTtny6c8rpl5wmCT/f74M/sp
oSAHW8ukhmsaENFzZphmaSljDiNk/WBLNbXQj8hUHhgFyPdBcdsxTJY6Paq9g+iI5huvFpmx2CW4
XVGtD7pVmuLeYdk6YZH0Vb6WRd2DBM1ovrT7hWu0Zt1RSqOu+6dt8OMnN+obf1duFLraxOyjWtTm
V6VXy9JvaVenjySe8tvfiCBvUeN+BfZ/RjvfhnUourtMIZM8JEIxm16nOXOQomgjnLTQgeIg1Ma4
EReluMdvQI4YcdcuAFFqQhGHJ5IGb3sFvshdIiZUZ5BOa1XpBJARzMECPJW9wILlQaUjhALZhoQ3
q9kSCtkOH6QIWLF1Zf9heT/9Jxqpmw5pqQ2UQJ9vpKqcMIgeeMMEaWyUCjLSXXRucRAtqijyVdyg
uz2KYuKkvsbFbIAlNypaUSfN838vNvF/hiJXf9Tc+hNxuMB2YHhOBmSxmksNKWxxsYdjSdTEaq0U
Ms2oTIsgGqqryfOuc5WCdwnWnGqu9AW9DBHs2m7HZuYX/at+4CHHWDJiSXtKf3n89IZRYCLaMb7s
Bwn1H4o4hN0uZVuM1xeAVJEuSD0J1RkSlWHOhQh3tSfIgaUGuRZF2OrzabzUFudA+qH1DZY02ASo
8l+1Z6cRSpxTWDHNOzsSvfNNJ5tJ7n7fOW/cjxevAV8FTefmKblPmlHZdTu6w1ZOqRA2Pa7HldWt
MQgvbKQD0TX9m41KdYHO8DcZoB0wFQJMwDTPOhqe3/jM2Wb416qKwKu3uBzaJg8fW4kU7jExOPOu
3ryf/lLnNzh2KKln0Rp8LFvarXuZP9m4i9wR1720YZvgFRa69NQQSM/Nsw2Mdp9/MAyspGBjlCrX
h8tGtxIcxLaertYr3Vlw060z3tHEhLbPVMu7Jj/CA2OknZf0Zn5dPyzcnRt4YBOYU/loyPmA+GJq
TPGJKjfLDT/6e1X9qzskxQhR//TqoUnrLwxis/a6rfkv6aqS52sBPUmf2rffn4A21bfaQ1xFl6mR
nEyDV040d7KXx1BzS/tXoa8K1miiezLGaY1/6U8bCIclEFZed/k7o7G4DHlpiKKXWWsVAYWM9TR8
inXSFUGh4ghMPG7Ov6zH5rys3coWGQVVM0widedoWXIS0sw4z65b/yRQSdeO6WH789j3ERtT47jv
ZBSaq+bwa7thOZ3vOrATvTmyE1ITqZhTBYX6TCI7/e/BrTQkmenENiz9thBbCBa8oIRws6sKkc4R
+zi/zRaWloketCs03UvhEpuT7dHqFGFTu22+EHoh0GasmrzLcp1JK83/iCXGneCkihW8wfwIpD08
LlkMy64WPqShHpKSz631/EQpT8BTAU1hV4Rd+64fZ4eEqFkZ4hJvsJV5baDzK+lFoGTrBR4Lsjw3
404DB+0DuOY7PibVwElg/GkePnWi7NYkp5NHarWkmX6gWpB43zAx9rf+59qGvpNQl+e0k/q6Ssjm
tyNqeu7F5B87xd11+51P9qBGi8jycTQo8kKm2hhaXoSlJ70ChheU3kRYxXYY5vCiQOKKRJ2WJYla
3xCdQdTAahpZ2ndPqv+gePZeK5jqY5+M1BUvIUa/+50oPYv0pqcQeHwEfoALyTFZRIYapqM36vkB
R24Slhfuf3mNq3Qq9/lSpbIPYJjOGWMSuaFGHcUPmDOpoa333DBsGxqM89uLD7eySVDYZPuntVjM
DqyrAzQL4DnQg42ci2bjAhDQ54/J2F00Q8a2k1ToHmthtq6QNRZEwHF0EV567Hnn1xepOoeuou6X
CIssS9xgz1JXy82bTvUP0ZRGhXDSbI617Gh4/5gFzdZRcUJGZtnXeIyurvwcFzziGMPBUBmaTFl2
G9OOODIFNgTUSEunzdaSHn+r0P48tn240/GNvr0jU0piBstX8fP7mu33cRi6J5voWuZCIAegcbaI
4llY+hdNV9qWPdwuWXHOxBpQtK4UID1w+ZAxp4aNKZuDb4fSZVFQRLwQIblnvYXtvkxprpV6fERi
Lm5tFom54AKrMvdyqYT1lzaw9l86u+rydAu1rziF4gGPhQtFrmLe2b0dxWZi2OgMkl/26D3BGozS
nPg3NHqmH4pbqz/xnLodZjefE/IvNhpeIxwQAJTTxxI1/F4bNYL2kcOjQfT/xRjtiqZ8YNzgbw+H
2VJIs+yNjpXfRbbrs9kxi3HOetO92jveym9Ow+e1NRKil5Ek6O3TXNXfmqUFlKC8wHLqa6/+/7c3
hOETC3CM3E7Q3ywqdFhepTPBrYYOyXZ/pEomB30drt1JVMF12Um3frfNTG55mpsBbphIXh+WsryJ
qf5420VRzhpMOIRmqaKVs5lbMr8+qILXQX5A8I4DomeNAOltTcX5Ismmj8nJ1BZACfU9PlBcb6dd
jktwOAue5V6kbNhdktPDDQYloNgs8bCQnjfX7YOvaGgRI4rlYfRifGSwBU1iOYUQr6L353VGoLIq
Xv2hSMLfIcAWbsrnGChyxRkkE00m3edHK49Uq7cAE2olQbUyOY7zHaZJ32hsH2Re5cBb2+I8/dwU
IIgmybpSmyt/jDh/Lfrd69Bx2aXx0iSSj8V/G3Vuy+wz9Yg4L8Mfy5L0wAqKl1GEXNhMoFbRmKYR
bPc9LzGYZX8q9iZexAFgMmQzLXuOIysBU6b/l9ui7mJuDUGm1FSz2JXDB8r1lf23uiu9tJ1I6hsW
+HbODANzGa5Y+hrBXRZfupGlVadSDtrZzadqnP8yEte5RWUIABMGcQpI+GEQas2PNpIdNdJYCzCf
swbdXzkHk6I4c9Witylhe4rHAvJXUcW+kL39WNSa9blSy3SgE8RBiUfFwXSpLwW2ZNep5QLdb4Xb
m73WgKlrk62EBjDtqj2/Erfbn6BzyPc7GHK3ibXI9hdJ+l2PeUIa2pj0QL4uPbja8E6OtZRyptGW
CheXW5VFznl8JE7j0Qlh4qcZrp8GIFzxOqJY2rP3nvzMNFOuFaKk2l9EqNIDQQCqpfjN6mmsgwil
eC2o/ORVD8taY8x+xYl9x0ZG9aYeamNBtagXAZs+eToPri9gr7cfyzA44k2yDrpDZW9breiB+HhS
PbSBPD+bgrLKReD38iLSgNnmGAhHvGRmvxzH7F2aSmhGdxi8VHiFmNwuBdsa9sE3/0u8tFy/FUmy
XGc7aywpYNYpKAp1+mC0Z5ltN6DrXAtUx0au7b7Mcf3Ac5HcPEqgMud39aq20BaKZVsUD5yGpo7J
dNgMp+n3oZwr/JHCWLWRSupDkvpPyvJhp3nhYuE8kXPSgoL1DFMZelInCYjwQ+qZMmq0OSJGJbFm
nQccBYODlzmhTQmcVLBQJjYBFCFR89Rbb3HSjzlcub+qJZdbNJ/sBdBs2A+9xa7YU3XZQcZDn0Qg
1eoUNkuIEvtWC1NXpCIpUCydH+rr/QOXql3+7MyOr2jODXU6uumdDQ8VZrZDDVQ6e3bWXg6hD69m
Co2JzP0wrM4B5tn1ktxD1lGLWKVYQQafmIEjY0P4vnFid4xL+gI2dfZYs/705AcqxBV6Aod9WzPD
J5FokqyMECi6PwJMf2WH7wngIySlansQApzgqVlLrtCVdht72R3eI74Q8Y+0mxa8ml7Ix1Jy7S5K
WnAGranZgPOMfIG8S/L5THNwGljBEQpREI4b3+koVDUyKpo8iYZ6ssFwQGXffYP0okj4/Nirj8To
+HxB+tb/Bcz6tROSCnhjw7ViEqNmw4f7VC1ub6z7HzZQu4+d1W/aBlFpO0xJrCHkx0WWzoTga9qO
i/N+rmJexKYdNrskMWVFTUMyxOp2qf+rdea2eEDoLLschdps8lfleHgcCYnS5TYxWMYRndx1uxD2
E4F9Pzir3FITuS0J9rTT3AtYoD5+pmqaViemtTAZOnBb7CKevJkSNuuZBXgr+mbAUefgq31+nHKZ
ZJzGMQcyyxMidTIDbpvht7XsXCI7YnklG8opFLOH3RJS/fZNlVBWQ8Or13Vze8td2TjvTGR+v0R0
foU5Idgnz+R1D1tNnau7Y3P9x/Vo5VhondjPxu+wtFAwV4I0VjY1qTQQ5hdpYnbnHFqeSeCLT8xo
616SjWlpIwax/UwQYhlHdkF1qKN7u66eVk7QeXYKqhrsI33mfh1w0mg1QsIL+BDfKrOzbEs1/IAt
zovQnTmyVuNq81w6Qe6yT+wjyY+AOEUUEak2A5B0qmZEkkOObArmGyecUGiMBuTbbl9h4kikRxXw
zk/Qpmlo+bSicA+SQdDvU8K6rYHUN4jBq2VEfHNN7tobMdmDnmXXALFggzlq6xQwfykzxAdz7zux
NRZzwa7fg5cTcm4PS75fM28SCy23JkMSzD7MdRbfitIOTkELAO0BPFjy5IJf3pESaMEFdguFpqKV
Gr0j7r7/gdn1t7n+8coJeERSAWw9pjdRqttIQLzobQwApLjpFqYlDa1XIX3cylZSXN+Wt3ZB7hFK
gkZat4CRbEVucjmlAJVZXVYjlanM3H51PxnphOJ3xXJS9w09lFBCgO9uxFUbfzGw3Q5M4/baL6NT
w3L42TGtBNZpWkWYSKm9Idr+F8O5yEsmL3DRhWZ6NUm8WWVfqer/M8mO2b9kipao6CVvXSoto7Tr
r10vZXGFm5h4THIv/6SQWXeU4mqiRjonxEWppxss2gCdOOcRJVcVzaaXUUyC+sHBp9NkHHHjt/L7
Okvz/kRfWaWdEn8k1TRhJ0WGSbA/fRDqkTPRhM7j7ukzklnDrt11bW5r1QAqlEspiJg4Ro+Py4h0
mqJP/D4eIlkJ7Vt28ORoD+qwyqghyANfjGwkQKpRumIVWwNZm4d+rJY91XlxMJcWhhUtuabn5865
AJP53MlcoBFNugkQT3sd/BQ4qEZPwPSPHx/7RJD8nYOCfmj6Tdkm2iq+9ZNUN3Wuaw/sgt738ZXZ
Hk1dYZhuZc20Qo502KEs1kCbeoiZ9qZH8EfV9DVWbvYRFiy+7DLXLwJBOCk/4LqVe/LoK4eqMkD+
aj+luAwOfpTgA4cYZ9pTQQoBIKVPiQWFf6RC0nc0S9y4stG0JgtEUlsQBEmDZvtx4RdPYxoATLq6
SM8tXgu8bBsa4oVF3HYQDi4yBjkmBK43We3eBWvnbCE0M/hlkKs4IA74dU9PjmGBaoKaLJTodHPt
H7M3oOgWX6uNbBJ2tR3Y2GwEFlanHONdIfIs3blufQdxlhJ8cye2VCPrs0SOL8d+tCOSA0dFfnpZ
3d0/i/qj0oWcWh/2CjBQ078jvjP4WJcdzxp5S8Rfc2XlocDzvqRCSHJ/CtpJUsmuiEmyPKxJHpEz
JJGwHr1cCBPWeiZ9RGcdPI3LDPk2Ep+JNm4ceITczaL26tHAbW8358G6vR2q476kHtreL+XDX+A0
5VeZxWVphKsnvh29JxSAdFDVRN3ctq2+M7zfQ/YR+Rh8FR+4SnwjkU5fxry8X2pSZOL2hcgBQiM0
LW9qIJHMmivMTNxDoQ1+LqoTJQgzDDXsA1Dn6bR8AGcyDw/SNU995B2SBw2LIgsiMDdceKfeb1H+
M8vgXsoFfXAcqLo5voki6b8zic9FSiSVZgJpLVx64Gos/JQ4MsdAJyX6Kg9DETBzuS93axgn7Qps
HrLQPkOHOd/XRHBmgmL3hk4HH30ifVqyGrF6vdyG38wbQ5nVnWv8oDZxP+a7mJvfGxXpQcKK7yt2
J7EyyykKIFlzQuNMZFPbXl4u/HQt+zzbe2afQoD+gtzNHrZ862GtIKPerq8GoNC7NIppY7LtVqbn
0mchjz7Lw5c1ZPiw+nEuLk5V7T2TYh37BKAN5DddDIkZFLE7yl38FGxhp4Yha0qrgNeOrIFZhYBP
6WODQgWqwBPS4ru4e6bZAeKr0xIwPDPNAC1gNccSq6wjDcx3bsD50gvE5ijT7wLbdSej9qg2n1iV
X8H9tmGzGmp37wLZOoT7p0HTmJqotW6U4LDFBfmL+0Y2y9f8h8cGWXvmjlkhJ7dJSsZCnPvDiBTL
Xmx6yW/LM6OTRF1gYK2vSI+/PsnPx73MnSDSKpftW4AewPZU15P7e3ut4qiy5CEVA5e37JQpjIJL
Sl1DP5K9Pvu+xFKEbt2e1rVfDA361s56hOr0EC4gKn2ZZlPZvbp11axYUMlvVRiTbUdJ8f590my4
pusXFtXbfi87/ABM18D0c45XbojNs10MxagqooPTJK+1C8Fo/uPT1/XdCgO6R3tzxGeu0zx+WnEw
Y/4e+SAvdTJUlMdLWqL9uvLPaR7h0daYO8sh9fReo5kYLOBMOUFKFAVqYTDPrfaEhlmlMVm0xepi
EbrDaluYYnLDuta6Wh7nfQtR4FXRDEiMOvu9feDSBtYqQ2+jylfRUXDC93+DUT1Jq5PNJ5Iieq4l
sUKobxuA218q7/MyyrTxaCquieX+A8L9Rypumt5RQWq2gixsNoBF3kXO3Nb87nJ/9SZzNNeSXdzg
rz9Y7PfcgIozqKnn0NZS3G7LMnr6k9FnYohBMWMTFBTUdlHkOikiyKy6ctsz5yr1OJYHtkk/2sbN
3o2LyhbSn8QFZc3zOKPOjcidSm09BIwZLgZzZExwZ22gqn/dyocxycVu/iQazgPJywqrXoS3MGs3
7dNGsKLWEDcy1Z8YRfZSWfgl8+QHYbUQrnYHwaywjM+v2vw6zpOqcj8aUi7j+Vso2Jm5jEYiHB5g
T/xHDLSY+HdibA3IjRDWphYvSJE3EP61rQgnphGyOhTf1IqqDX9Og16mNSXh89KTi+TcQ4+ZKMaC
3d1lLQMXMUaHyXtC7/ZVQFUI6HQnINcFoWEH8Y8H8ImpdHaGORcJFvwkrBbtGCX3rXw39vSlPPsT
iF9aSkLqEdv/irQovymOqUQ8lbIr/hHa7RrMsC7+3fU2f9zuRtf4TFo8cV/9KjKeorViXj7J6Fle
bzmHE2xWK/XSYEhik/NZcgyUUSh6K5xpsm3JOlgJ2YJAIF6BNFGcb+W5t2YEUqZ9bg9hR9+TjWlN
sw9UnLU367kBvrWKtM89xDOju9DzB4iWneeMvzYS6t/prWmPgp5heltqZ0vM1nJ+gVC8ocpfS89x
DzDs/ZkjlDbWAQ+O34g9J7vOofwfbQgpqrPBd7Esou1Hlr1Qp5yUV5wsV49fUmRdOKr+J2t1gsIk
glZQp42emVzNuF+oGsFzltQmxwwiGVVOjVjD3mpvb30qV3zLMf9XPEJGU2Fj+8AtQQnWlX5adx3a
XljS4rCei39nnnHsgUdPlCRerjmL49tN9ipq5L3FALVLrqbEJixlpGaoGRzMYZDIcT9rRgsmjp+C
zAi2jPb8dnLr2QaorDAQ4gvf8nwFs0e0NPjCSEu1a1B9utGh+FL7BNV4AigOPTWlt/sOUokOUqS3
788lgM9wkWxbOJ+b/HajarStxS/VbrrDqQEAwelNABYUxjqQqaVXCpdH3Zinw7cHYQRrMKPLv6Pe
/mgy1ORo4JAo1xDyQhmYRwzOIb/lFEBOQIzPLm+qaJ0mxaXUmnXQdJXXUATTWjUOkvLpbC6M+NIF
Jzi3w+vZt2ZRB7s06B+o3+EQlxQd/2KJsAVKPdoxPCOL6Mrdnunj4aB9VRRS2hePA1Sz+5Y4GLkJ
erSOgF/Vdy1oYfv6tJXYAfw/dcs59jc7pCU3a5dTWpXNJDY4T+aCnNsF5uC8H+0LRe09JZyD5Abu
9VSoNZJvSjz44dj9O/YrtN5zjs8O/+C7gTyID7G9Q5gRsmBczOVVx4wxLmi/4WVr5ed+uMRkxeEK
t0Frp1TrHYnB2L+mXmcNV7tcLgm/Ah3PIOX0/xT3zSrsirYVzUdmieqAuqHQLwlMjZW8kNDjn6/y
bIbPKrCaZ32rQTzlViwG4Q33LhRz4ZVME8lLEfpbi9X5cGOGLx/MfqsIAmLs2+Zons0g8C1Ymesx
LnCfVWxu7EMP8ZJZ6PtWEPAH7dIB2iF7kUChNJFThhVsje2N96fjQk1RT9dgEIkkjcmnNxF8sRNr
RZY8tFEpUh7uov2jNNL8kwjn3uk/c7P+o5KdBvsE9KwX/9ZvcYCISZuKLNq7tAKmUHMwEdXaF4yo
uOY9S0Vk8n2pnA0vER99vgUiZ1EEoRPtaAiJFTLQNPXIFBNykNl5r3BXeBqHW9Tm2wpDf2zowmzH
ATjQLhgXcCRilLG2ch2v7jcb9saPwL3d9S4nDnaX29JCnOGIfqYyrTrJKVqB8tfOMZiF/Qu9qTDt
UR/+r+ZC+4osRxc/b2zqwovueH1ouGjPtFtWPGmZT+NHxm1lTEjYcbYZ+e4I3HDdPh+ixDZxvUUq
+PoklSGa1mI2VTc6Wv9kuPin3C7mrxnwNDTyqjinKyJeYNwmHC7/7a5q3Oj8/U7ksLD1Z6W/DIbs
rg6pRIhWI7PQhf5dGtTe/cZkonuw020KikQy0KqKHuD1RKqOVyLDiZMHe171Ipu4748XFw5L4mr1
iG4rqjhnCu53gJ2z2tn85ftbvjATU1m1pkUzoDNceBHcfd/Ih7VZQLgyRCPxdDdw23A8C7ZFWTJv
G7Jwb390yo/pyUrhaAh2tfquH3aD2yWO3wx+XwIp+bQrZBNhlir1GqjSpJnWrW8aRtZ2wfDySbk8
i/gHXxmocC/zSf74y4sFCLv6SkYqYv2N/0mK6KjGpYwTdIvK/jGmaLY41FMf3lnTLZI8gbrDFGQa
3FBvh4jRAag7JTpSin3SYzxT6DO9qHiaczSUBPSeZiT67a1wBmkicM+8dp2ZmNO8ibiRvYfxShg5
Xqf8M7wrDo20wQYeEfc6SKlAm/XK8JB/MfzCYM4YqayxZJ7GARUZeFCaUc0F/Y6UXoe1voJ6XwKv
QT1YHTl3Pwty7pj4oAq/W2i/ElansiTrgyshc/Hvqs/0/GJ5dI8WaZqfG9TB5kgcW56PT0GErXfv
PFfZ6rBp3aiN2YlFaZGMexKerlBBaDNc3rxTyOQjRObAG3y9dvz5wR5w78DPadRqratOGSY5T24x
LDF/oRGwyGr3Pv0dsgT/lfBbUhya7uTE/HxQg5DsW5knxgzCUYsUr5I5jgViIRp5pITPxxat5Hus
e/GlFqIyxqFhrUJb6BqtLaUm/fBlR4fNIxveAlE4HW6mGUL5PpP7B2qjZf2dR3BrJywbHgGaQRLz
84RXiCbCOP2Wa5AK6ZT3gmXnx8On97eiJdndBO1fuhj9N23GlBEDSfVlkt3x6p0s/EizbSjLm1IK
z+4GFQgeUX5gamJYGsQIKhsMCEsHvret0uTg+W6aFG3SzKGRfCCOeLCtKsiQztbJPVcuNYIYN08e
fXtspUl0K1tMLlnFScxg6ZI/gsQUPG0C+9qVTpTIKbcdbgCqlkKWT/X10Y8ZcbJECrntNzlWOaAf
vlBfHgM2Zrtd+43J4GagcjtKW+cxum5KJy8nE9RtaiKT798eSC1lADk2j642CeZafZv/iw3EtSab
AWO130Zsl8qHmmaOcwApblmi9RX0A4M7+iXEjMxsZEx4uFaJGjNcaG9zdYglmRuY9QbR0ArknPHL
f3LDJnAoodq40kEOtJmtUI0LIcrAFvFlUCzzlxAD2bJ57tngiPnnJMiDy9vHHLlsSAU5bwaIvWSz
pqbdKnKrUkjhzU4DXEo2pGMLmS45tgyHc0fAKU+ZBht84eUTNv+lhEE2vVEPjw/ShvmIX0ksKnOb
J/wcOA7/QIHeCsbAJyyArrEixBnq/x7XCKy3LbhoKYRAWykIT6z7aqOKztzJpCGO3gYVoQPXuSAU
eq8xfhdw/L7y2GtyE33U1kmjd5IWJGIpWnlrOApBnBRLVxMKmPNU0ObQR/xuBOx1OGGaRSp8eiAe
zGlKkqni8S7P4FFBquV03zFFDMVpEuD55z4EVlz29UAX+lQ2O/WKffUmNa5RAc6ZnjiT2zER1xqG
KMoKqIdqnp0JSiBV/tNE/1uFM7ooz6MKvA0V28nuYBRnI4OhWqTtf/x9y7TOiIGhjjoUsugxmXQu
G6Y3m/kje3nUIs7JS9C4qRWBAbrzVYNUxLuJe07TPrYQR9NbLdtWw1M8iipFmA4FLSJNEwIGqEdp
OsCxuhqHuTlpjj0cGCKOBNyE3WILM/LJYkhH3hZX0AWv3BMyL8431iebT3igarBImrOD0KdUoMX5
2wH1jtmM6NngNw5xInVd7My4nvjvgEpFYbBH3eFyShVCFIpM7mrb0AOJ9vooZeOSvQd3BubaZL4B
S3Q6+xnDVMk34LX3cmBP3g6Ze9aCEp+uiNksXmEa0hWfsb7IBiHoREWfLPm4UTADVcpER58EFTyY
RaQw4QgGv7TNyMJ1M6J9kT2rFuoTC7CtCCZ5L6Ym+wHJFQ+i7kIhXszKVaE8MXpEG4U22NB+1FsN
FnKYWjKjhHpLgetn7z4PP3kaPVOsSSJb0CTIbJaOVVqJLG3lqJFwCWkBBJnNkQQibeYWyyxAMzad
rfnQyaQUyNhPRib9C+tCnHZLZ1RZA7Xou6vJ1LiZFNPI4Ptlwn3e836wTtpeKR0v6XTQOzR4bwZ5
QZ4feHz53jWsF/8s/ceTA6JvZXokMV7eoNQEgqwQWe7pZ83hQKdqbvoy9z9no0uwjFlf1SHREeT7
7J9lNcby6PuTCl9qm04NotykoIbE0SUPMne2EYv8N3HFcQ2vUKxbeRYKC45IvwL5bKWzapOuJbhL
q9NA6VGph0zMfQ0nmqOtYcvvK0tqmJsTwPu/5dnZ/BTwmKeYQtu+aMAnLbTN0YMj5wIPqnmWPjTT
1le2SUwIWL8xFl0jNrcmCvBf/6cQMhH5UjkU32cz8mNOJamhpBZqZvHR4KY0gBZNq7nDvd9kmXPU
5J5zKtgLFWxTD53iByRb/RHvcvvpp8NdQfR0JCBGTfF8V83Wjm23+3YeH/+ZcjxKaF6bagUHDliD
qjpQlDe1cEjaoxCVz2XZE+R1UwgAc3vLUJ/P1MEZdHD7pft/D2VeJelYgxKW8qQrDEZJqJA8fZld
P+a9HUbyL75IQ2rRsmp3YUDDChLhVUspGjUv4RhuXZOrHKh6A3g/TtrxqRCWGx21sap6vtg3Q2SV
O2q/BhnzS6wTqabJidJMMlMZByDc0sC9nhiapkN00kTPzA1ghK7nL2nph+wEHqiMAduKFY35enlp
j28nyoCjiBX4+jLQgQ2omZPwwlQJE2NvO7PZr8FJFMAsHg2OIwNNmPXFqEfcLEmHV5KywxGV3qi9
vse0R5jkTpBFui1pW3eutuy+WPXLxi0Vlj3IXJkkGRFgrG1K6Bx2miB89YSLQ8gFK535eRWOb4qT
Z5TXG28nz0/KUI8hRd5QQl5ASmhBY69yqaeRvgMbjpPH7xiOxFUv6pA5QU/PBMJrgOV0OY78z2V3
N+0/bfSDJeIbUjd8Jtyl17PcWY3QCXCu4Dv7bffev2VXPoh7IzsQy0NHv2hQheXB2tOlW5qfGpBR
3KF+c3DJ7QGoqivQy5NJKke4K3OmLNZyGe/OnDDuuJ2r/bSVV3Uplvf3BdVhNsRHXsCpC6zSe9MI
CxIKJ16SkFii7125AOGqzizxBcGc1so/WeW908T4Sq2st+KEITEuoDUdueOy9SNTpoAACc9mHsXU
05RKoAdlwD1ka3G+rL5p4Yj2rLp4q+R5BdG9Puy+WwM3mel7q4nGrelEFeOBmnVGiyoUkAKC+fe1
0m9v/DbqVXkY0CzjUaRQGojaaw4v3M5+SW7bzEL929GURd6/x/28i4PDR/m8kN5AGAQ3DISJ3xSK
LGl0lU0QymZw90O6TqvyRQBHimxl5FqnjCycsKziri0oKOvHkWKQlnAEYTlivWta0rFTAObDJiUu
yir9kwXha+M2KK6sJqZNXEW2p4jPD2VaKobwEPVihO2qhCqzEoCmsC/vppnAfAdkZ/F+8EBK+L08
THUI6/a2Dtl00V4pEqH+ib7j64gTv0b09bsz4dt8/Us8G9vcRJeQxT6+TFgs1xM5G6AdJvgevLO/
fye8Xw0IG+7/hjFVLrALdcO0hr+y2fqYKGXRfXobrby4RFFWngfDB3ETZp6xGBdrhotZwqLNrc7g
KzI7hOlC9FpZZRwD2/uqzKZN0igaXM+vRYhuC67w3r+j0uozumth9UgyGhlSKVMOLHM7iStHzQxQ
e46QiOV9KsdyUhmI4ZtwD9+51t6O+zxuFr7jHggOlGiohDL/iSfi1KcFqDCtx8x5yBErswpAEMLM
yvXhiZj7XCK3XrSxuK7JaHnWkGPHvP3x8ylncFKwPMKY9H6iSw+sDeZIa6ZCkfiwl6cUkiES9Ewo
vyYWbcO1RTndyiLbq3h6HVlR++VCNojm39KERfTEUG4feUgC1h4uggnMiYQq+EUqGcn0Hyi7ofMk
0SugxY2IeRqlabuSPktDt6WtF7vycJiZzG0M+mNKoeYz8yCEJhtLQco1UayhHiepL9dRXNYy3WNo
7DlE7p7+U/twuiNfOEih0ut9osBJjXcSG12sJCn3m1JUtB9cKDpnS3VuxeGO0Uz0zl00Hs63tWi5
J+ezTT9pcOIYnOCnp/Lb2sJNSU9rtk2Vl/jCHCb6w8CJgYuYWupM2UEmOMK3D8OjbU2uKlEczTAZ
WpxQ/mf8QfoSdPjoftiHBocKYnGOLHV8oolqXBroXODKfwOIqqBeZkyOJqhIqD2taKAT/pM4hxTf
PsGYG78iE0r5MVjhlYkCgm6uDDfzX/H5SsV+OcEGoChe47oig1HXZeCpUX8VyFA808N6YNSgVKPM
TcjWeqgHysPe0VZZ6RoMG6GwlKzC30QikgVWqins9BP4iy/nPCp1IA5YKaKzrJWFlfQ6Nm/JO7zM
KEUvUj8tcwH7t2FLErKRA7DIcigsvF8NECQevZx80t3PuY7guQlfRrDBaqgiDRmfTtUZe+K301k5
o08sN2ooaU7HLhMRsFR44dyn8wa/FnOY4XnuFguIzDa3r5S06DfQCrZfeEtJLTn3iDJnQWxeKZIl
5OOJR1GBejo1pFNLfVnfsyYDwrluUan9Em2RtoVstP4LzHhXtIBRVpJAhBIowi7y0jZM14Z4Q5f/
w0CqjLxnM4Q9d8C8Oq80U/cIDAOi8fz4VV8SjNyM9fC1MRVqxPOt/qexAuTlt8EfV+PP4H/9rh/1
srhCv+3U+fQbQ9sxW1Cpu+FoDedgz8/6qa1sLivnTMpcBGGn0bFayDqWRjm5RxIzBAzvwcEHsEtJ
+5vuT4W0l+M0cOEKKhIaJTixCyR5G5e9Hk9J8G82gM6FUZdvLci4wTsihTjIRki9wF5eSQouSXXT
1oXRFUmcmOyFFDiYyHsgsAkAv/Em8ONh4Vp8GF66hjSf4zkHJz7l0POKsIT9IHvwx+1mugq7HR6h
f0ktP9v8EoYjT9K+/dNZ+7JpwM8QkM9e0FndcZnD47YGYOKWozctkTbMGvwq/PPhbRFBZrNkjS5w
2T05FxbuStOp3+PXuljvhF2JZ2/d04dKDT4zQeZGVXJmIJAHa12WX/X2N0Frek3BAnN30O+sGhjy
ho3VqXXj1oERU4E2DYvA1LyohNe+JrFMPpUby5FwFq9iN33Qvr7SXzj5P2Twmh3gZYm/0gvjno3q
AJyiWBo7pSnJh/FrURidEROMOXdcVVbX9hQEtV6o4anZUSeqtign4MtQoaBM0tANDdOJwGQ92MKa
uUaR6NnaYiz/YO4RBoL9sMiuZ7SjhHcqmIUeMRunQBjX+SsNWckAeLsFwJ78fyRTJolgKWGAno+R
mHCef/0xsvygYaJMIx1LqhrDnrFu5CGGwjor25nwM8jfkjJFnybiLUMOL+1jDaSMttr0a9FNdTZG
2lvfJwLesZq8roE/axSQP1NiuoOAhh8BSKW6vJe/vIBc0MWlBB4rlPc/RBkkVAGzt6abt70leOpd
fdKliYdS7PR/fcOyNQQZSQG3k6sew+AC0AKIpbtfg0b+QKlcNQmn8rxdH6zzARRzD9enpdpB6yre
T/TZ1RAF+eD3By90M0tSaXiZL1hFPDT3NwjBWXjIT1/cUbh0+fO4VJDDuWP3ErWlu8z7wS8OORjP
nOxzU8XyIw8WxObnicyFLdcEi30k9Ymi2RrTH1NA8yfyAY+MtdwqQu8z+O7PfM/nBpaXXOE7JkMz
Mb8iJQ/KDmGXbUuOF6IMPsay4/KOBtmi1Yu8m/Oz5+9cdPi5+itGk2GMhedScroAjCSJRGIBlOFh
7swFFh5kBVh8s8mVf0zHeAVidQlsZ87d7L4Mdeef3617I1XKEbk3GslXtLCLHp5wCBCtnUmYux9e
nE6Mv/5uxdEocopNFpBMAhdfqEh4pXMxzzvZgqlLMmiUm64Fmev9Dx6XkU/MW4cmzCDi7oH0MgeV
gQCsXPG5WQVBUaVqjyt7ACXXGRATb2Wxqc7ovW9cg61DsgDzg7MrjSqZfAaxSu/8hgZpNFQAEtT2
8xfab1n+Rt21S34slsgbUGOQmtHJX/WNAtFPb2RAGm0QBZtVme5U6Rao6vItyndIaKGs6kd3jzwE
4ocIwn3TczG0qAnecviWBu1gJunMX6tZZfjZiwKvNBYzpz4dAsf5G6tZL1dPcIfuYGnLsjBT/AfJ
Gc+ZlMSGNM4P60iwCPqLPaueLEFtStYo+civLpgBnU21koS593/u8qDopuVPBvUxX581lZz/+10u
mzBlHdYKOPI8UNkm1LGw7zMd6qLc1Qto2xQ0dpEPOrF+i4ulQ9zRZuSitmdDbR7SYGzZp/mSEBsR
eliKTr0es2pn5z4JDVPuWkRnVHgtD9ER0f3viraBZNSBzip2nsq1d/XjRYMgYjXRkrmkwNOsqpSh
EZYW91CfZX9PLu4ESt2E0W18cmFZOt3M5AC8Wn41FzDJW3tr1fJqxQWKsW3iGvXXGUAh12NJ8fRg
+iF+vuZl+6agx9+OWP55SZxoXL74hhNl2sWugz7lM24pvhPU63nxMFlIdmmadK826tg39rOKsBSL
pJYhV6DJUZs+BK9cqjXicGKdaSjqjhLXDg7IKKZOF2ROqaOi/NZ+oVHaPfNIL4DCv6NbJ0TKwJ3T
BmouJWnmowGjNPZzibJmer2M2TJoPxFp8CPPy7SSatIyFIT68FsBikcOvJQ4FNwPP3DV/cEaxtDk
eiP7W/yuc0Nc1xy83SFrcXz1cysxJgll/63bCDfrS2a2sYFlf/919aY1KxmRoO1Yg5AVCCLud5qs
RbjAkRu6ovcQIVEASR3gWqqXspeA8jA5nkaBJEx4YWCYsop8B+1y2tkWlPwCjsGr9bkAoh3xQ72d
htQ5nX/kPXnNBV0h7j+9025og74d0crhLZxUr6Snl7ky0QnTrG1ifcbZoXCcszV3dQ6cI5LwHIvX
8x86XvXs5cax19mum9CsfIIfAZTvKSQtL06tbx/uCoD6g4HR6sOTY/Ftv9Aziy4GaF8S01rQuUnY
X5RN58IEX4BT9dXJ/8x2th83wFHA9LdccA4zfmY4wHX+fz00nw8LXFsXBTgU4xisv504xrxCT0eS
8YujJrKr5JY5LRswICj1wX17Yxcr5qMHwXhfJBCvq7OqqYXyU6K4NVCBXCSy5E3HEhYKMcjyhASs
DEdJE8go1S3ly2rjgcdbsClswLMlkixUjtQX/1HCsbJw4ENPchkhSS71shhYAlVzMwXEx5sH9/eD
m57Q29tnDLGm5al9h1c/Q3IYl0nUanCkxQOrN/f8Cgw11FlUUYJtTZsCuNMe79dEHOZqlEL/S6oF
MUmsGmK88ENXPEZSM7BBsqDOpGKql89GgcSYRURRUT9axX5reff2emUb7mD1+bqh1Xin4d1JfIXN
Wt9ESd56U1tGlMXGphiHQjNtelwkRTJHm2WQPYLCGzZIoV/zLlnoSb49UaKOv0/z1gud6TQUK1TH
MLeHVnF+fyjBlQ/VkcqtYCvds+Jl6y7aWHPv0OIcMgv4+64+CtTMAWEIKxp70nNCX6vXCyH/vAl7
xm6RYU1bNEpRe0EjEVb1lfxK0eFzqTD7kfuhSharCWNOcdiROz6Xs5P6YMDcAIydSqFYqNULR1cL
JelKcvFI1KKsO5TE1fKefLUlkKjsQ8YfP6Dfu5nDUQzgrF0m6UziVeedZUK4t3igHmRk1Lk6sAYq
8LWJUjnDdErE1CJMGQdiVerggKsViRkkZ8CSxp075rGEkWy/IoSOqRwYidlz32Eyj+Q+e//9mYGz
zuDOLQkbSWDwsqKR7zqAMYvZv624qLBCtD5gmfjndf/lf3voVlzJzIxsPfGdqBh+qpYjsZUvdAUI
wefDva0ppgVqUw3QM9SS6HDkALdOvuVc/euAgmiEC7laFVDDsaYzDNpW2ABuIAbRkXNd/Juy6nkm
6+v6z13myzQYn6FRKbLPsdaAr/Q4kIBYpSlVsSNnsEfqvY1Ry+7LLehgvy2fsaGdRlyAuVjfQxM8
7njEuDcyOUQnC9SwUFMPBcdKb4u4BYalfKlHp5by7999b0O4SsLVZUovD9XCe1B72YuubZNSJXlV
+kGg5u+QsMAORKIhoD7fHrBZ6ly8HjpBF5Z3ISiHmKozjBGHMIgbiFfH6HnZ28/5LOCloj8IOiUg
huSpRLSx4fKB45B6IEnVuvBri536+pYAQp14PR4CilNFkvF1DujCbn//w/Os3Ys5LhqXWtWoscwg
7XaJ/NXCXl2ONoQJr4R6r8EhpE+L69yU2XcE8Rd8/zkLIv4+AfWPDodh5EpfMC07SI12DltH+kaQ
+G3wkqPqPVK2WpeZJPgjvk02ozbeX7Jbqf9b1lwN4zhuXZiJrPSi+BA+XRxg2CqmDW6i0T2FT3cQ
QrI96zBsJPTugP2EDAf7oxy/v01IwiRkyQmlA9Evv1MBn7DTit9nohiIVdiNhrvZb4xvK80Eb20z
LYTssi0joSBTaif7QJn9xYp5Pw831lp+8H0O2A40h81oPIGs/7MOVdn0BysPm/Ri4cnYmLH6Ox7H
NMIJKkollGnudXaHhkzxk/vEpKITnQn3w3+KaAU34spIIsjcAOdeO738iBAi8Z4mlt0i5ZqRfW58
e++EQ4fMDY6ekOfC74CVh+jM6b0lrSO3NsTX9baFiBRRhSnSkjt36CGzlQTu+TspWHki6jRdc0CY
OOw70QNPZK6OUukGZ1bXWr9MDY7TuV469bGA8CexVkJTnPOsY+cLVaYSxgt7DCqm5yOia6DOuAH9
jZlTT89BTzFW/hmYDgxCHGCmbdV1/URIQUlbh26XZ29HG5x8M5LCae/ikidgvh3Tbiiv0MGy5ag0
iZvaTvEFLL4zXYwEIkC0lrdRBAIR2gVjW20nGv63peQKYMSJhSrCqF3ec/bYR7tgTDCpuKMqWslg
q7rkl9GYefQFgyLY42doKLjE6uuEbAvL1A/oC7CC5pMjXqeZVmufYwmCt+6t/zBTsfS0qRO/IcFl
vvDmVmjw3h1QfbNJjSFILY+DF/cTJLFE59McPjoZTxNlmTtoTidJSPh8Addk0aHFG4MhZE1KWtgF
Tz1Nas7FfYl4MR03E3oV+ohY0YZ8qDiknTTqeoycGByCkZfeKikOP+VaqsGSZLxNkWXLfaYsCd8F
qBNyz43cqJkbr/wwAwtTGIfanAMzGdjSAo1/rZi9WZepkVZ/ev3EPhn8OyOiqlQ6CSgpRvwXQNNa
Bw6T2rRx4K6GxJY+B/UnV99kwAixnginqd6X7IcOMJsveWV+IlJkIv/7rp1LwiN8A86GzxIisvGB
cN7nrKNNTxqsx203Lh+ooSHl+2Ks4uxCIhovw9UdTRTbMUZfH20EZoJ8Ener2Ub9y1+D5AfmwdFo
mh9r1Dho/u7HzWuFNJ7KYaWS4OaedVaXBzBZlh/kW0N3R4TUwJ8zwpAC2EAgbFHJStwkHMb4KNsO
sxBCF8rMdeXA01DEPkPsiY+4AE624qyIntRuIjQBK70DHZckEpbFSHxLrWHcjKPOlW0cB+POoU+Y
pL5ceoUzKAsWA9HP21sOUCykXlnHPRClr82kbXvo/CTvcSgDTJ6QKxNKSMYZchYITXqRFyREZooG
YJvjqCJ3LBOf6tODNHt5MxyusSOf8gcBb2MtKzUI2GbfiF+OK4983NOfn15xXDxEpoAxSIhjLWer
7Qw8G749Wf6RMMo3xPg7jE79mYUQh1w+nCsEDjrcMDDQacADZx9O38GCXm2w27AGf4yrDMIlJElN
cwK+/YpVp1zNQkZheX6s/hfPYAQZXoj1dHENL74ITw31F1pkeZmfSd4tm/iSV0qjzHBJokpZaOZX
49ZoS454TNmLwnsmVOBobm0mkdSYv6HFnFLQ+bgJ1vp4IZhz8RVGGJw//F29BdXYYuHHDAF9PV67
Z39n513rkUnbM94mXJtY5oH4LcfqesIayWxte74jwyQC6Slerb8Z/nmHuFVs/UgDewzwiOhFW60b
sS8bBDbe6ovQjNqDAfxPyne9tNI4gTMOGLPzNMMIxVdqi/h6TSGpsCCkE0K8ZwhYywwCmDvs9SuO
KMA6aM4i2wtbnoEPXn/y4uASAd62t9Wx1QV43QuQKPg9MwfLhxB+Y1KgWX2WSgmj2ubJXBIoi0DM
86OSy7CDTt9HY3QqxQqXuhaiVy9uYsUR5WVxURMkH1ksTsDzn/E9GUDTTjzoHHCPqPYQ14Q8wjIe
CC6zS7ueKtvn6pDK6WLFEux8sgzw0mInNWv2O99Ugg1fGqEYZwdxxWDSE7XJiCh2zRw3Pxmej5iA
fOctAwlxXPsxmgbGrOyWFrB0h6F8GLFVcvhZFnsf5fa2tuBciBHj0bdFSP+qyR+eWe/l7qfmpmUN
gBkA0Qb4fbAHb7gXszBcHktfUwbbElKi/iMa4VPaDolfKDIcl/Cdfq9pV75du0HfJFxMJ63Iclkd
RWnsNFsqma4fbbGHmW/e9vluEIfnpqk5B05qngMy+6iUoVogLGrApqbAiqWt1gFS7fZulPhXxpa3
DN36q6yExyjXz4KSB83HiS6nrqj+stzVMIazbDiiNR33/acrxKP6WGmhM6vB1S6wHKlPpD+g9tek
0fX5FNVyxATpbGUo3vOSttrMiFHv3KirD5JBmUBtKRZUkDI2ktB8aJ1XFv7tUqaDgVUr1yY7kGyj
7hHefwAJ00wo5E1TKGJgSgE+Q+Cmi78++twjlPlRZ/ejo2ZCoVsUoCcISrWw4TP2t6li95/H3A9p
/cOLk8sxRuLTaZ1gaWD4TB5HwgiwBj9QF7paqP3CUQqf2RBSb9hoUo7Ot1ns0YmnPkestc3UPaoQ
eRgCelUf7vIqXg2cJWi0XcCuS9jg7EpvS09v0ICgL8x/MF+NUoKyqHrFO1YIUFNhjQAc+FdfxBz6
ARzct9F5q61qraP5FHgU+g3hXe+ikVXwtdE3JcfJJef1iTHp83j895MK8l6+AFjkTjI2SoDOCaIb
xSRV3NZxlNu8qgfpk8OT/LNSdbljqCycl8kgTgYr9Cq6Qg0Oh1u2CrExcQDIwn/v1RJ/chlObrWL
cC9n4tuuMn/4qPbZFCv3W/rhXg6MPkKSf54cCfBj8nhztrsxG2HDmMSWYEABthEKqE2XbIAaRCUe
Z0dA3io/fOssuNN4t6fzX8s4lhi7sHzgdsu09GLiBztYEid/XKCke0a9Mi5S0hWUTz6+7eHrxMD1
/sv1kYU2DQbvYrl9tUwdspfs6txkgHO96YiuZDoLVYW7TmHTcjWAZXCELVVnntRyOwf63zgtoUr3
FhONqtyCQv9Z8BxGQ/sCJ7bkcKaJxunfZyNwzpUQbBom+ncKv26eCwe18SY7ZVc4cxIHl8md3egq
a44gAo5iIqPbswZ+wB+GrIAobbKV/7cV66wswe0eDynesaqfMwTYXNQLvJpWl2dL0XOW5bLeCuu6
4FsKYRONbPCdh9ArXThHdKZqAEeOrVk+myikw2G8jeezGC5PIwBWfG1DgXe8spc9SiIiebNp78oY
OwMEz8WVEksysUwVn1eP0o4qM9rdJlWw5ZPHLjedPy/0bcS+5xhShs+z3QRCzMVSCfywVJbikze1
uasSPPOcJ/HtSyLYswS01UeVjEFNUqP3ogZBg1Hh/1zUxHfAf8XFwxOW9FgmVEjsZfuIyRSFuTvP
olY96ADZGd6Z9I64OLM4H+XmuTgGd02Uk5u+KH0c/KbWIk1MgCHh5xFVlZhURx2fLK0tdp1mCbQI
Jp8vzpV/bo30WMlm2UtW/FzsPcdQjr4gEC6nnSzz7/LTQbZ66ug3MKJWJyP0vkaDahW/PQVHRcSE
MCxJKKIeO1a8balSQL10CH9rmoMGFkZDMMxryfG7PTjBnipzi6u5jOOj8X3VrO9/FDlQr+67ZqWZ
G/ycHlGzY10Y15PlVWAZ/JCjnfaTC6Enm1uSlnN7eodZ5TJadRvDXH64218Mq3SP2wL+DLpsxB3U
LhI8yWlBXk0XCTP8gFHziCRtM4YGZ3w6UsgDD1+EFhE4RsO8XznQBM5Wsf/h8G4ecWM/dfOG0T4H
JgY8mSalmVzgheRNWtBe8n9DfKfx6K2QcrK/bgDG/e58FyGaFey1vKHOkkuuOt9ZZe/gztZo5TCY
NKO22pPoItbV2Viwu+5N38yf6Pyh2qh6xq62b+liJzL7xJVRUxAnvi9DlAWddaet1MyszDLBL38q
njZl89mDt/KzjlEZQi1vQuw9wto/3aekNj6FTtCuB7uweyoR5pkdgRC410lDlsj6pcGdIHpfKdIA
qjwG6lObxow7nS75mlhvwfap61X0RCrGKhnnYwjTDnL6/4L/WB4tzM00bV8ZAR2PpNajWt7b380n
nj2FOxfKyMvnyGO2jFLYeYH72pKpxcsF7f542xLGag8L0sIFvTBh96oGiPR8ScS08igwX4mlmHrH
OlZSvHFD2G00Xa+7KM13PTvsFXVB0B2SmXPNGzQyNE/iGTaxo6LCPSzn75K0ABPDUuRduxGF5MQp
7lKT4w8frLPWiUbgI7sdnzpmhLWco5RvHjCa1/p5tc0pN48Q4LX35gDm4+ms/wrtB3MbWT7nKq10
vOW/7YBPj1Odds3mz9vBveWO2egdhPmZIkwbFnFkixsbW9TDYEFy1JD3JpVdpPJsMlhXP11gRT5n
CYpUWZyXf4esi0x8xl4k6LhAoyQLrlJ59dVUkPBdhZH5dhpgnsspd75xy0yzsIy1uZMQXWioMzZE
3JVKIVK0nKtM/ELmQG09nm+iXIYoieODZAsDGq61Gh4R31/wdkaOVNAhzRmHn/PiJR5mXm5tGgDJ
JsI4GJ/GGoKRBaHgMKEOopKxHE0yQnuLg9aXgtMiNQcSRB88FjqbbrAtfCCoaRsbQ2i3cMtVAaOP
tmKn4Z4IXiUdkvawDzc0NNpJdIEdFgnzS9C2QnCwlWcKlbQyxfG/Ziq/I5Vx4WoTU48Ov1hTV8lT
GEEfC3Id+Obje638NfcQihc8uw0W1L8PCwla4IHN/fhkVtzjA1N0ScPbOh+lidUGWpLKZPdYEsjk
s3zSoExPKryoRdgenL7YEdAR7wHvxVDogLSzLwUTuF/6qRUTytcYCokYyXKfuXGpr4KD3LZS+d3C
vdL9Hxz7icxQtL4X+2FWgYgWonjvdYijY6F51HcIZaYLst+QKRR2mkvLCTLGlCRCp1itg/Ha8CHB
y1r4qiAc9jMtEg9kDykoK2KcK1I0SeF2TbBINrDH2yjBTfb0PmZqFcfbYhCriErrpHMTlETcyx4q
/M5pB8P+UITMTl3earAMlvgdZ4ZZAK46xW43BKfbCgZQgc4g8SlAh2U6JYTiTMjs5hjn3BJyJVaZ
LF+tVz5zS6+zKTonWFK2kaGEs6pb1GDRqMHq3V+do6bbEgtKUgBL94rA5s6JIqKgCI3W47xxzEvl
skFdQ/+kcmRrFsSVVfiqG+SvgJ2ueSoXPetVggE4vLMtnI2qy4i3E0RUk+v5BkgPCLNE3oPWbdIi
2oMfMt5BqZSkWsbcIeRp8f52IP6zICvO773H5rSrnNtHwi7E9WHlRgBrWWwwBp7w2PZcwUvroO2b
fp6jdQKOjs5nZ63AG36PRQMdQW/EK2BMBnmIYFpBWWm9fh4FL5oL6pzoLDoo1eBpcDr0pFaJvM1L
CpjNmAk8MY88A01Y3NXi/QtLLjiIJ4lNbTYXFVEe4N32r+yHLMUyM2Mx37+U6bZYPbJ2ZvhZM4hW
GuGOjOl7SNQbNEFTlyQUHKPNwCarhb41tLsfzwaDNrGNwJa5/+5i6q4F+5unZpZyPE34iLqcn8mL
WT8ZV6mXMP9Q0mI2EyI0XNvefBDBOGZv7nv2+ezCEYLep8/plxa5u5hEkd+cyEo7jyseHls6wgfA
6P/oCFHejOAl25O9WLSxr7y0TXd43VnxNr0GVqQFT2fckISzrYXxubrWbsH84wz7UsinYelfjI8E
/IDxjWk2eAEmO4tLTMtGnV1yExNWVluBldFCq0WtWK9SlyWKvQaatH8UQE+Q4oWLQBdTAtzdO/wp
5W7mPta9XxcB08zlds9FHUGuzYs/q2O8oUfDp67dz7VXKw7nQr3+5QASI3VgVjhaTDxxXrWPCl55
7jOeeIdJGgohaE8cHpp27U048qSPp2LgCpd881q2gAspkHw7Tks/P190OJPi7Gg1WiT1OwNzihVX
n/pCmKPleDUj/gzuZ5xXtyPMpzHNbnUKyJC4sS0sV75T1/1Rc2nML8neBKppTWt4qBM+iaaGVfVy
eH0EcLNqhN6i4jpDEyEsgmfRSkLsBqm9uFJ/KLKhfQiYxyP6HFUbF+AcGyGUhOmXUdUCwalxeVuY
nfOGfALwO8IlpnLOd3o8HiaeT1AQxN/GntUQiV2GoLtE884uqVkVb4B3EuXU5G0zZiO+PTy73bmD
xZ+PsWSy1tmDJydvfiPVcBc0bBH4xCJN79gU0yR1UZaMskYpi6oMW76zvj7YTmrLHPQHYnskZoIP
BtPqj1PdYI+5963CXQ96Rn39D7nQJIO1/KQvARzf6mzb39j5asAm9Z6N01aFp1becDAup4wmSoIE
emhBkNCkl4MZGgrUQjHuX96/bvvRzr1HPfUTJbzTOkjSCjbclM1opnw/GtNdSKe0qOg+484Y53Nh
Mq0IGWRnBtGS7eIXjjJO0R3uzSEBq3o8/kXllFr/heH28GC3Eum7wQ6V5bM+3zqaEWbICtqUXAOr
GIxOYZtLol1SgbPOFHhAM8qsC85NInZgcQs+bZT+1/uznjt4n9nQXTboUH7lzwx+hV60knA2K3g5
IkbDM30A02k0OP42iLRJw4EjUjQlbX6fbRktQP+DUUQ/O4Cb43+4EZU1dFt8xgJQdkzBwzwm1LKF
nI2+leNpbqKvPFf0bdpQdOkcTmVzv6CayFYQTw12ilioiLyi5qRisHaQJNssqPdxYQvOkNjeTRwv
2S6pmtn0BVNa4j3RvDe2meMO+PQNDq1T3i/WDQeiL/OYwMIXO7GT/WI4dSBIPcX3N/2WprZ/CFGU
NJu1mEWaC9hJYso0rLZi7tsLN9MAlb4YtgCP0XOw+XKc5pShs9sgdxctEexeIVQLq8aA/7jm7+WL
TY/r0my1mxLWnR49A7IBUYJAh8o9l4MQJRNAZVq2Tu761DWdJPOeYEl/jSwSnT8k1MhgfYXO4F10
ClK4DHHoUrkBklKQG1EoS2E/5NHsay9fBM/OnYUIwuMYkVSnZ1NtlIOv9l9KxIevVoOxpx4UNvXi
OY3NVQHAdbVxl7N0jXGP9sQCZ4opIyAXvcr28OPuMIhSTLPiTC3GpaPE8aYo1W5rJDwMJCrbPNYn
8oI0QQGge2XRVnngcybgxwvu0Km/LKaYk+APk9YciFyJ7HOJRaBkfOTmCPLOQ67heFz4443zDPdo
wy5Trfthm2ewv0YcyudMa9/FM+fPBjFBHlNUJrXa49Z4YXXGEDYx9yrgNCoq/ONVOginfpDmaJwp
lqAkF5pSVEUhR3pE5Hnl6xTYQU7ZiAMEL2w2ir7ugGcZ/HCvUgMljCwsBtV40UDqUPxf6/eALywD
vUAUZPy9sHjo4LIQ9ERc1GQXy7ClXfi8ipnSgmPdO6Pd121Rj/ndRP+uZMwuuSYoVkNLNXtCLa+a
y6+OYYZkc89GQOoSpBMOwJh+5LMlbi4uXOnYrvugg9ZUfRa1lLuI44Sn9Qhyi4LslaWnGnQW8/M2
bz028XHRDnGowLdCyaUUc+9NDsMMlk/aKRucZiIwB28sQcp3LyACLqsf/e8FVhsiP6QJzu1H2ZDK
5NL5N3FmUW+jxo21LiOeE7hwuhXeLj3QbxywF58uwm7HgoRl4X/dcpTsXm+OzEDgJzWacH1YhgFJ
ssnfFEVTt/g3vjmPjhSZCS4roh3fkPc9d0tH9w6xdP0AajAbkV7A3X2xDMcrn0Lcr97P+GJts6OI
PwM5dQ2MLP4thV3JhImujxff+LNZrcIx4p2iNsxyKY6Hx66sYVgiVpa57pdZvpGqrrWkg6zDvH6a
SF/x6+lYN7LbqZKwWOgb81L8ENF9UwgZ6HksPikRxoEoPMPnXOT00mD+Sh0N5BfKemCCCr0wpvAE
80mgxsLcXHDRfrVi5KmVPHQXYRbc68CxhZeWSEWY52sv0xqGMLzfaoky7/wsDCuAVa8+MYTgKd2n
D7d82PnKeDeZnvhCPM7rwxE4JPt95tviQNoP24cwY3wSNXL6t17UdfLjmk18yY85Hs0Ji6ZrNA7g
5GiprOzXWUqUwucIeWaJH+g3VxvWXR6gYbtzvy8RDsryfUQfl/TRwyvsdJtoIv7i7VE+F2rvjybg
FrydxLLv6GsyqnHzrgFnDAcrsm2mO1M3xmRVz9e8Kzy7QhojfCqJL/eePNIoZqpTgYl6ZOwhnRmQ
5Aqk7cw9Wb16qH0CpAzJbw8jcos/R/AS8px66mlLicIqGsE7dVwK7LHaQ3j23gGltRhFZB4C9l52
2lf+/bwsLbZfpi75BkM0lp/CiMl7JmxTMM+W8hqdt/Hfw2JPd7HfJ5d8A45bn08X1cG/R9hz/AL2
Zom+IaeB6HAMwL5bDUCADKhlIE+LohSrfhhY16r8Mm/xQtUi0xQKiexLyXAtJ5xQFzBajP+Ipyr2
QA42F+9mxorHzGa7F5zcu/4S8iiMkDTk2MacY8sPe5iAg0CqQPEzPz5jU0tUADgM1LWSyuuJsz/Z
iwiYtn5cEIb/BFS6niqheA3ablvjmAand9niC2lRFLEQqgFoP0BxkLxCJ4HnT60/3HxbaOvDGjkl
05l2TdmOcV3d8VFocr/xCj8LJEAQDZLL6wCupSppWXMGTtCcZXFL1Q8SIVY9mjv6J8s+Kzhd4Kmh
NEkBNNZe4GKTDWYeBsQAIwDJR7OXiHUYEa4WddLZfjbYDN7/FVC/VYV1rzVDVE1uLcnED+p6oh23
phzadszegBOXK1bn/IjtilvKLOY9gTWdB68t/iTMD3RkpU8hlB64XlW+e+rxynyMPUjKNg3hVhVp
kO5jao8j/wRvBPJkHf8+eEpLwTjjiKree+DW9T1Xrte0oIYhjawT91GNUdoGTnPvhuB5+PE+YGB4
kgzJcCMIrG+WbI0W07jO5qBNPzs2PH6Tvxoy3BkRz1k5EZptBtO6TkygfO/czKKxPVWPhJAPCCh9
j3u8wSfPG3WzeMaVodn3PHHyIhM7ZyNxFiQ8h59JbardjiDepQLgfD5jTd7m4RV/w7qjvKADyo2E
6eKj+9U7sGc2gsZI+2yaF+diGPTLpMcXM0P2BOVdIiH6tZuWlhir5TLQpgufNMdqKksTMsx3zrOd
wBqhiokXbey3OaMGjv5+7qi0ai3YNwvQOLdfaTflqMK8q/lOPRsd7e0zHl6H3GS6AwqIHTbsKqjN
2NIlF7psn7AiPjDJRof9R+uq0OT6ElmYicFeVyv9iqX7i+LXeV/3SyU73dJLzv0IyUMnQ0vRWTpv
7d5KJADOO0L6wDd2c+v2Mcyxb1w/7/5N+vQ2y6+7TT8VDUJo+qjv4BpH5WhnoCRw/LhUPPTut1Kb
/GPqkETpyIzrf5/+G6RbFsyUkY59zQE5R6qi39M3LXGh7GJleYRFesEy+3RekvDb3Nly3oetkPw6
u/mhHiuaXdyyixEfka0kD3VhufcUfcLvMNLjir0SuEhWkbmqoU77mTiIC7FWjtgSNWk6j8R5AjAy
+e52x2DN3VS3P422rEa7GaILPa0lTLIJYsogsOyScy4TrmIsIAfIMEd4P/n0bTTMVZ30C0lFX+7S
kBustEMIvcs19/OEzh9UsFE++V8DaP67c0AXirdwKHxxsYLXQw9UKLFqrbSqSoS5gIImDeesa5Wc
wlFzghgK2DyQTE1k0pYbwBUYh2+qIIDFeQ9cbn1fstS5ZUjWbamWF/IPR7zSImRFFaNDnuqXhxeO
7yb/50JdbCOdCMIXHciBLAoiOydercK2bSPmFv4V55tnvIXq4Q112ZrGWBQlSaOV+UbqoGL5K/0O
O8m8L76XIZXDhf9LIqzWPdT/sDzU59lIXOc8U6bIjckr7lPbvMECOS8KUK9OEeclEFtA9H24b9gO
5G4ocW2HDE89ePqqjqjRdbnQCtizR729wjF9FQbCefJnhZ4pM2OH/mwJTSgMASl2rkN5Ck0d7ujZ
J+NUra/xxiPI/X3OzhxQ6He8mgTm11G9czDHAH9StrdfxyttYF/BEECGLXELJ/nm4FyE4ZNsRnNA
taYGzPvxUJrKmyXmhym+ZhOdlkbp+zUAzmjw6jCJDfTbVFAvEF5ueGsT7qWvV8CLyEat0atF81lP
pLSmA0u8XKpPto9d9LqjvkRrgOwBaa7er0NDk6xxHwF/zPGhrK3JGIHHCtMCVQoG+Ei6echK51iI
XCg9XXbtFbri7MOD9nHh4FlSQXDJkrqVwusTZL521QFFVsU0prD02tn8TGDOrvYZgEQk9aTxrcxN
N2Xk923J3DZBQhgDYrqXoL0rr+kNxCI75q10RJryjk9gZbxypcrx46ycqg250ZrawcLBf9QhNwhi
Rk7yyiwBVNZyXi840BueUHkhe2Ibx6P2T60ZjYlX1PlFl0VSX2qJdAR43lWmnW1PSxt+A6M0kh1V
Enue48BaUTnw+k39MfyNoax3SR5A2PMR4oXuG0DfQS1xsLzd/wqsgWGvmRSg3oG3xA1Agpw+ykn/
1lA0aW1GVnGHz3dn2gHllRTlxwmzY3TzPZznhd3A75fzo5fKiAS8hg4U+CQrM3/9I3lIJsN5nSAY
94Yg5saex5WOrR3MPZ1pn4rxOpyzzsCCM/O1hwWXNnhqGM3sDoEOUwWQv4mCbX0vZGjy6TWypYht
HLIqqvwOG4IfQwnitpUbSKfp3FTeUf/GUNcjqSCltHWWFvQukM2wq2lbm3D9R7g5VyUA7Gc+96tP
L6u1dVTULaKdmj77zCxpUYru5X77B25MMM3rtNXC/68whdwYuxZpx8ugDn463AjyQhYZ9XNLI+Xx
selypkVP8tTQhefWZ9WTsAHyuHb+nsGfVlTy8QnLVrnksB7WTbK2nU/bejFgVLVzV1ucdiWP2O3C
YFUVKwvgLYijfL8CGBReZwraTdAEzbeeJx+dkSue/Su8aXVt8sAATEVZTz9nC4Ilwg+8y1344oqh
hX3c8GNJfB+kQHWKJvAlzCiNW9U7guZy0N1T6asf5dCqHAHqUWUW++uDYe+7MwTaTiBW5JtvNF6k
WYsUBMzQJ8wDkQC05aNpYofkyJv8fo7vDq+pCyD13cce2MpjPE26eZo9VyB74gqC/ggOR88HmBbK
xkx42tB067xmyyUYoBP+fVB93iFJP/fSrEciWSHC4CekbbAuclg5ooZOxGUpZCbdys6bU0RUIQm0
aQljtt/paSaSRx7fPjvqYuFA47d3p9XVoUYoAUesNyeXF8Gdv/nNbHK3bryA8bC99phDHTNxM35M
EuEqFwkzTtWXWVtLf5XbERCUdlhpcUJTtrY4728kUdHvx8dOmXUxmGrfPkg8IIYWJ/57LmYxKRsm
NIjYANp/e08CRB1XVtIhyHANZ9XKd4WZSP/Lc2mARVaUKEc3DihBIShUDj/ZFDcZbIVG5SyHDn4X
MeOBzbDrP+XS/ie3VF9zgRVDjIqnYnxqIFNNEMq0hkJEYTkp0PqyHvcHLkY69USClIEI8Xyj9DZz
kCf4IFQovN+y77FE9+Yq/x7xOwgouaCxpLIBBwYbAf8+yiYyXSy68uCfAUvyHPcWi4IWbbefTKzt
84zsEmtHtF8wojSk+KTzt0c4zULretBNmOXNAHeO6dKdoN6XE0Dt/WEfE0ty4jjWXmnjucZbJ+zl
YEJLofZWBeQud/tr7MBXqJwRrZiUuWNM7scLkZdGWOP8FDGZ9G/K7k9P9o9c0153WrjgaKnw82VY
S+F8Md+sc6sJvTlT4Rs6dTSkuqtg5fMMRzINPLnZiCc0jnNxienONADOsS5jmIXpWxoPl9OvhbAH
McAwKzaLCZf3X3vk9cjm49QfZahLZv3hM50Poih+Ct7a4Iomgm/nxBe6ZuVxW2AYgWpXFVkTaS+4
0PDCQ64Kx4c7XkAX0Zq4kTN8VD+pqtyORsl8JM03KarPlpzswIDdkXlR28UGviCmeX61E1zuGv/D
n4Sdontrk3DgX3tJyxpblkdfApkbaoNDzI0eNeV5lT43e3Dl6iy+82+Vi13Hq3ZZyIeT/BGPnWXc
fXCceAc89EHNeCtOW1wfo2RzA9p9XGkJpcNSFM9LvCu91hhHMzyOJtl8ZIIdNqeA5MFfa1bSESF2
2l0Y663k0b7m1eoXWWx4Pr+K7KRV9H260b5mFPE8y3ssq+XkixDa9zROOZGqs/3IoOHlhNz/TpCP
ko5D7zY7VGWUegcDa/FEZsTW79Y8LirFfsAFPcbVr5fsJCfPYtoyRf+Bb4ecEd/LFRgjcEvqQEnU
MOEsxRO9WcoK6cK0V1+d4bWrCTBcLTRlcjVJSH895zYyiSvsvbEpvjGE1Vd9o94o7IiFrizvUiB3
HjYvP7GPl/uD4GH2+qNZ8kmINNmf60hK7Ge5GquqyphwFeNPvBGbZMXxyS2MrjvjKxeE0hfIqkOn
dzty7yjKPjyhHoeTxAAjGCeQ/nMs3P1Q0QYRlwTDzkodcsnm/MiDTTGgiWflHhShboGGWDkj5uIe
/c7pA4QrFApjskMnyki+cBt3u9686rvaWevYBqkqZBQLPpqTr3GpCB/MsA35NYCjCZ/UD63Twt+B
z2QL8M3RBM8bUeBQ7EGhW/7N44Mxq1nK+rNt/Sj89rCOHpxgJQS3bww3vWhNJqcUDTyzNRjFvIdy
zXc9LK1pCVLL2+waNmirsZNaqwIJ7Uy9sDPCYDla3gdujBGdmoHPOiZc589zv7IdDDpaDyFSDKbv
NQv0V+DZixd9wsnQyJsklSd30ap8xZOX9V+H58OaUSN6gmrxff3rCCPljP8d5wvLiyv4jaikaYe1
37POPCKwzJF8WbAWicziUurTzvqoGf3NfKwD8ydO7eAuFqN994DZ0d2SCq1wZUVisuhTg77g4rpY
x5WjVte6LKxfDeLy1SgaCzOv1aB2YVQ4E006wJr4s8FQ9MdXzZfkIE3sZ6c5Kw+TreYINR/jNgC5
y35YspjLZisCD8nBRjxKe1CH6HPjDyNW6i5+GndU1SMWQasM3Eb87JUbzxTz5YIsq+W8ArjbVArq
JvJDFee2PbaJ8GOvi5X4ba/To0gm1Xdty/x3G5tk3ChYFr99LRN9pVywTcJV/eOgnoHNttxIMtV2
uNBE8ofaEfg4l4F3rxVps6jDcU3cWtBmTvIJFejVTvchVNyutwtZcioyBVvxoYjRaDfLsVN//c/V
jXNUNgAVbKTJnPZcBLeGScSLHsZHGY8caf5y7sBc4ll1IT+H2hOmak5YeJEteTi5j4BlFGguHdKQ
7CXM95wu0/nv2j4uauJJjdBP03dA+lRyzweA8KzOULjgHtcrwhaPUdMZqo5jGse12ZMjVA/y3p9v
9qtrGX5xu8PxiOufh8Tw3/q1ZgjAdGD4ITdBgvT0h7a0opY2vMQLv8trr6zYLnsyYqIf4CJOvvHh
OxffzXE+ERfnZWo58aXqZYcoEjgMK6AbDqAqy9jHNk4htLRWD9WCk53kyDz8Vk9RtKtoVjIgQ2fw
EQiBZCUw8wqmQFSGzeAfoIqs3ozP0QpazbTbRkm3kCeOnE/UBYP27u/qtDKNKG65CwLHgdJ7qQ64
d2kKAR9QKrSEpaVDq4/8Qr6R0+d74dzyHVKIp3t8wXBQZnyF+GCjTfb5fvMflI5TWHulBng01L6D
SeH/vSp15lbmbsqUSvOqIG/OHI3yOjLjx1IwiOI3u4DH5VjfS8kvmGasXntaTUGDfDkArigSsKpF
ZmBSLDMU/Ln475Z38yvQ+DhcTpNEF5vNjBdVrsm0l6JINdpRQyYHrhm12HKK30Qf5D09jjmBjWwv
VrC/5rez7lT31Zmeg1LVKYLFH4ron6cH5jbH4NfQLunXmrBQZSPc5SvbZvHXGY4kouqKfgmDCo+I
27ShfMrqmtm+XwqDhKHGGBnbBsWGavGN4a2abbXzAuDsbFhOHQCBRoYgkqbBaoiYjnCzXEpjEj7u
Szr1Swo6q0KPN+eSpNdUxQt5qrWqcekF072HqUH29wiaYw8M80Cx1qrasIV3z275iqVbHRzbQo8O
GHbRE+YZw5qEF/fs0Rj1CURi3IqqRcuK4eNxTq76OSV9pJ/eihzHZ3CCmL8elowHh5Lp569WvmXH
JucoYIT4GD3cc45JrBIG41GHsA/HmP+W+jl6ezl9o9c0dNzKHqNZSgE0jQtFqKb3x4SfJOhaXjFZ
Ls/Tk5CdXGstHn533CoMhzUAB3qRI1b4ljQ3pR1kb7FJ8APIkU3NC1ONIkLdKEXrDMnRHx/t+fD3
vQIdRTqwQr2W/lvf2GvE6TkJ1nvO4+mx/aUnnjIW6oiyIp8iiS5x0UNKrfhCq/7vmcuml/rZvdpC
EVndO+Lh/OVg34P6SGvzEn1SOnlmylkhtD1ZO0jiVykTmRrSFT3/2J6rvcf1kjMAJ3UKt6/WGUWW
+82r7p1x42yL/AsT+Hl6KDNJMU6ZCEgmfPiUD9HHb1K97VurlxPL3AK6sVdenb5jGGpXsY/u2Zj3
hhXoXOJBQjoS8KuLpYik3tJXXlCz7r9nCwBiTcNeV3/WMzt5SC0LSz27zjLFOusdHFKMKV2X+LRS
+ziVOpxJ/TjwkJxZjMtZoP5IrB1SfOZ4HfxQ9DDeo63sJDAih92nIwc2T979xiEqrsZL/j0dx6xR
QU75EqbpDVdP6iYkws1FItF3oNfo6VvDLnUC52qVhxZNqik8TMTq2t/dnYVw5GCLJJyfZ8OA3YZZ
N6sWXXNJ82KPk+KhejH5d7EXucTDShZ2GFtoHvV8auyTbMJhIBJIiuusvHoSLq2yavUKLYWgVs3o
2rAcaCcvbNDOK14Sz/qAHX+SKI08e5pVS6Pf+tgSRg8AUPR6qy+lZWINbGtQzLkTKTG4+QErpqiW
JTEcFUBvuA2WMuTUpmkcK44fkeobpk8YM9iObEuFPq9Ppwx/8L/f1QdjXnDZA0E5touyrBEmoKWv
Nn10Es0L21nC/E4+1iZTIq8+h5poIfJhfJCIr8CHoKkDIzyZ/2Dkaq+c903vy4AsrP1HFJz93Ubh
LAnDJMY8RKkE4amJ0+T9WWWTVax4jNLCxqOarcDPKbRobueNcKapDf4Xs8o4UZ+ZALjiHVnjTFJM
8ZTp8TlmaR5Cdmc9P5VoO197ZCPsajkfwtNWHjvjZF5PFvrXRLxh5kYSIoNvUwl6wrw8ZG2zYaeS
wnJ4CTpkNi8KavbNUd5HeNwZzcJEiK3uDPqGRKZxFQi4eJ+o7xIAIDq6B6RDe3CD/Fpk3xQDP8uO
yL04eNwPiIzxE8vPFMw1FNoRDlhAAmxorcBSVYj/qO1CnQBG8Mgce406ghGBbzmxixXMqSnPvS2L
2HD5bRyIa00LBqy4iTnY/a76U5JL5C3n1QOqywft7HUiMWkoW21tTQ1+9uoasb65IXI1Qoh/NOG2
dE+Ljo1N4cIBqfGonlKBkKbAb7qEhzUs+uZGHORqTz4XbuJ7rOQpJDAw1RyeY+PYYRMC2AP87C4p
ISya9lYOpnFHYE5p6hBMX5Hi7YXk/gQSt6zPr2Lkrzzv//7+6Cax5qaZ99vs+B1QvhAncIS9PpIu
K1eqvU07G/acNz9ILsoW/5+RhO5eHzGAtQ2hOu3gICbAngv5NEVCdU/kJEpaD9EEkXDrcEfBXPTE
Uz49gb6RqATFOsXrPEBktE6lzMsQpBo3somRZ4vtlxAJ9TJ0YHeG4bcfaL+aao3hND7hwfqNoC4P
0LNyKY4SWN2RaMi3R+FSX1nwxh2JEUeegg4qKiLEkhQc8mxaOQUAuT8SkL1NLtgw9pnhbIBK7aoX
FF3RuzjR5YRhK8BGFqAaSXPmfcnSrgKJvZ/Hw/SD6dSCaopLdrVH8XrrV8dboKgHJ0dRn8bevgP1
oM2/zY2BdV/bhuwvqkq4fbLfCt9j3huIhYK7j+z3xA788MIKaA67ajUPjoYJGUC1cb7hVyypZiKd
Ju8nNMHPw/cyr1Iklc+Do60Ow3KHShxtyignXoY006Gmjbk/FLNkNkqcuAj2XyxgfYObXnIDx+Ya
GfcrKTWKeD2c4JjPX4WI5AqViYjgbjoZfm74Jdwip+9zF+BJ3deV/ueNMSNs8Jj8CR9yg6WwIdNZ
LOqlZULIvrZoqcv1M3UnwbpzN3inc2pKMWjd5lq+JfI/7sk+See2lqw6HXNvC+nOD6U5E5hyIAAg
RbloknMC7DBC81v2FFSxd7VG0w0hOGTY7O+C0H66ckDt9iRgi1TA97o9xmMbhTUqvKZzHX8oihWP
hdIlnP25NW5HvUXRQpvtAlj6D+kTMf8yum86l90kL0zIod6NUINlDviw4hYC9UUgvYi+oW0/6eCo
HVKbiKn4MhSo1fO26BozVSF4+ScqICxKCQHn4JXqsFYzOl+0LFDj5SVcbDx3hZVerxfucx6AFTm0
YN16WN8F+vMC/NEP7H5eIU8q83aDjxWFFu1Oe0/Dgrkvn5TIY/NQmiob0W3EbgUYSWSTqp+uo2xi
8cQW/JNnS45v8Lc/UJl+bKTP3bmXhFb+g9I0NWnqD6mBhAMzmW1o94f2YsImN6RSLMfCawwfU0h7
BBzGARG7AFS23+wtuZCzBqlF4zdmNOI/tf6kinWe033dBeBlKUTXXFcEmVYgNsQhQv3FxuqBedvU
UBncVu3WV3toj3tIOtG9WImJrRNiN17tkHazDuec95XHImAjQXWvv/GjNdPsyHI+RwLHy3CKm0+W
N3LtinVs0Z+Wk+kIx3QxKG7qJ7cz9K1Snoij7CvsSPUSHupWL4qQ1EzL1cFqwo9q9Gq2WhADfZSK
bldiWigXxi7xk2AJ89Jr05EeyVf44SRRGLVWDv6I6qd0VE9sPT0JPB/kE4g7Dgzs/qPJcJYlmXDB
tQhGi0LwmEJiDBfP8yE9sgetNKQVjvcBnqzivS3TWz0D5/xjlnmzUiycKvCSSc7T6GogHZybCfXN
57islbSnR07yof29lvHfuT1TEWErTwRY9pYnVVj+K0VOABY6iJmYD+C88kv4RoRS2v9+HOzBaZD6
Afo8e4oOEhFJfAFzloGTGgz8WKtv2MpGuWrmX0uNA1lwYwyAmM5FBG+LiXHJU/i8UjUTas2uWK2P
ti7E5M8Xxq3BzqyoEQMuZDzT2p4kQ7wW4JTEKSP6aIburRvtg4WIZJuBkw+6GJEo24xGH5Bm1QpU
YCQjL7mBQb4cS9m7c4XS4W9SpibjyT0T4HZdi7BBLCoJHlj0KGpY1eP47RuPSUn8ZvxmITC79taO
Wf1ZFQsvz8ZtULSYOmxPCSt9mfkZC2XgWDjtRmKbTpsIKgHFIvaU2Qdn2ZvbMoKgqYo16pkAHi3d
2hj31/jf/JlCrL/IsAkEc/ZY0MPlJgKjetFtD3LSHaWtYmUS8atmQ8h8BwgueCs23PvV4B/FM0Ge
N1Gxy9RTvz4usq9nV6mWRRiOiQJ3b3EH8FnyCzMPQzEUnjSIk8OsTxfsKp319uEfWvDZmrXCo0FG
vT2fbmyyiyc0ZIWhdpAtsd+I08kPQhmQMPeZA397w+XQywQGVBqK5V3iLMnaoP3zTsGvPzdKstX7
sxArSQR9We+k6vnFXvTt1a5452c8fBoMxhPN/JuqgUehD6yezdz3AudK930Ea4NYRneNUGr5e32s
hD2o7iTzXdpnN1boTik2lLpX04myeljabTaDw5ZoMjQ0e4IFOoJBlh2320iakoclPHBUotN05a5S
Sst9Rk3otNfJ+xRmMje8ZnxGZLAwJeuiNrPPBKPlEmH6T5SXr729bo8E95mWS30Bdt8ocn1w/fvs
oYq0SngTTfdrpIO8aCcCYv65AgN/O8Gpc3jJHQ4TV6vvy0shYgx0WI/J4qKwGkzORrGlrYa2osQs
j+LvyHGVrYBUpEXjcaho8HQZJtFpE8N4rs/CEaqC7Xzlzj2n1KoD5I7XS5hWN/g985h+Y9nTbziF
NwJGUbpl5tDsnfxtIsgpNmjfaaBh3XQ9sQiTkdtwbOl/Vig/bJD1BJB9+BCfIUgxrY5hdlJ1As+Z
IXMzxafUuk9H3ukMrjLtBRpPcZrm4uuaFaeHGLOccEzUymLHl3IdxFTqclmZyPxxfMoSBUn3rxyr
OR35AWr6DVv9Kq22wVfRHIDQ/1Ei5uTO2QSoFLzbUYl5wMA4N8p9Isw0xZ/nhPlimUYgTwyIcCZx
9P82iH7nXyerjr46BM7KhJ6efrKdVaKxyG54KkD53grMBDx8SaIifmnXXxKEuooCIQK/SQ7bU9Kd
exedUd/jUiFxMTzwc2SieOizSHvPW4RAAscDEEg2p0r4SXVjGHc49WjdhRSnmKO6fCjGhrDE6+0A
+qa4cQ5hsuMTyX4+pNNqdshWZRTYi/K99f/9qMPL2mcf8ZC+C+WNHKj3NGOfufuVjs1hLsfAQ7VM
y4n6r0dIVVUl6OwJGjXdOdldUUvmPgKVjM8u81zF3MLWvFyPDN/rubFYeivuwIMRBvKgrLr9TMvs
ilVW8lsYRYbZNXJoy0zsORhA9EuGiTQb0OJxsEhkyUmhwcE/1T+m0ejpCZEnfU+QEGw4F56J8F+y
IBg2YdByRtplBBK9WJlSpmElCcH2je2pLJ2EZsfDNl7oLsrBW51CXbepX3bHAkIZy7ZbOVajVED5
N7MX7RYLf+FPDj+KdZU3/KrIXd6Dbra9+77vJ/gccyCcU9KbybZWuk1gS4kAlg4akuHRW3aCu1cD
BFfxiIwHAuutvV7gAKqWHcKggL8Iz1zW4kGT34moyN5J7VtVQNJ8jRDrBCGHYOR9BCsrTUxnzH4/
mwNauAUMKbfkvYWfHsP0WvHlMD1toyQh3DODwqWTvYqRCA2umRkDc5zPeWofP+U5Th2XmpkVAOrR
yyw/4Zm02a8IEltr4OkwCv9cWhLq2QjK+ZX9BO8GxzkB3ZouHJhbCajznUX9tZnwEm61YP8uD8Z8
KJQHILqK/KIpt3c+zGVWvyXWvrhLNN834Qesa+zxsnssR11atRyOSdlANKXBe5bgFbmXhgLUpAmJ
NaXF0lxe54cqLaNgK3FDk7CW1OI41qLLo6DLpnNMmxT4hQupOvVXDL/Fe/kn5xz7e4Fdp1ZiO+A3
DFv9aqZDSRfEZqR8ASUc528Y9RmnIY6TmyPtm9+WdNMiYOS+wy01Marf7KzOruvNSyaMejg/1DPS
kIyZ1TBpxktIQTadMh6JVnAmJeiW3FT4ajyoU8fyZmg0vcG6p9QLcmiRXEpvj+TGDFzSVa2LkEmZ
UlK/cnvgvaz5DxEbGqylsQ+VdP8fcjLURSo3fj3SW6NsI7yulKbs0Wc6HTAoAsacUeufYIowJKX9
ygxKUhgMhXi8Yv/XjBMI9UW0SNdIHYnd7bz2vjg7oPEpMeR0Klvv1pJj4ql09TuRc7RbvFbAEbgQ
SPYqYXOqrfLXx5aicWHQpzEm1BOo1cIYU6Dd2srrEv9/7y+3/WzeMGcPsq7QZ5uqyo/bF7AIeMVO
ei8mkvS+/tNlNx4ESEz/V28RXUwcvejfqVAv97t+hjnXmZQtmfoTHpCn6XJY8wJsZMqn0gqkATe/
F1ia43/EGwvD4JlPE1Z1DRgXUf77kmXkYBxtwc9aH0CxviUxUgq9DVwi0hLuDQdxIn9/mYZCzmoZ
SuHrTrk9hxygzUAHZrKANiHWNI5U/UX3NqY/HUKtXDff8VIQLIrz6z2U2C3fflY7R2r68mc2mqLH
6DafEvzSMB+sUy6k7U3D5uGwokz7ILlIRSu0ud02z4YWcH1s4gODWNjgq8noJt2alk8fdkagRA6I
AnD9ybjQs7nYdyMXlIsrNNZ/mplQhwXGqTCrqNdWTCsz9Wtn6fJ0zC1eDWsuUaf5UvDjALF4Sa6J
J8TlbjjoHS7teZu25qZIeAvcjamA+Qa2d/MjCxlisNCiIP1/FAUkRg0HlMY6IhjzcBNbVQ02ev5p
I+VvdsnCx5yBJKtEbV8CTZkSgB+M8mF4U3HPeJ61D8S0pcIo5W+n9/JDlSyT7x12ovWmjqHtplL4
mSgGybz6ihJhzTtNuk4dxXT7Gbo9BaKX3EEGxRhTXqoH/KwaY86zEBrXsK4NlC6SlGcbaYVQX3+5
1T5cnoaL5U6SZqkHTnZq1XNemHn7BXrZab8YrZxh1Fsa/XPaGO6menYcyr2U718yFES21tD2+IM+
Eguygn8szVfwAfDFc9fnJUA3rdZtSBT5/HVLGf8wfmrfp25WUZHJwUaXIw3+DLYIu4GvgQvGXYzt
PiPlKuvLUcoBVsuQSLqfc04lly2jADhLB9nyTPh0utoIpguB+NbU1oP5XiE0OCECrHxBEx0YOsug
k3zjUdIlrLva3UIdHxQblCp5BPe4XSZTnv5HRPkQGUZeLwneyOLSvHbkEHUjV5rZg00ITWL4Yd2b
jBRtQFkvsShqhIi6YoRDhHp4+S2h/yDZ7gkJK0vjRwalgfP8prHQ/du3U7Khx9yHcZ+r9PKCi+bg
77E7nS5P2++OCbRlj4D6yqdQrh1F4L3fzevRKWfPQeeXSVhFLAIoIwmz9e7jqPIwM0JZEFFuPtrO
SvMrCjVNV3CeVPF9pn9MWNxn4dsUzmU9RHf80nLhW9dFz2pLilwToB5OLTBLjMeHkOOsaOzQCo8w
M5Z4jLFHztgVozKybMZSxwG8mohJqOb5u2OUhCOOyJXlXWlEDRjRSfshBJ4D6/CxmIuaRfyMWahb
Y48CiHNCTaJtf0FxdjIo4IhULkSfeCdbyyqP+t8Kf/yn3qlD1C9LAYkGCU6LdRt+G31YqPsZWh1d
xVKN0SqPs79w8cP7W1b/XOHfxv1qHtwWcgM1Emy11Og0OuOucoKRrEi5iMKFuv6QEdnkWxjYmoRO
O1AAE0D2jTlit/ZKiejDhfU+fiLArIXMt3pRa1El9wH/gUAl9TKEtFVU2O1n1aKdJEVEa/cRmKzJ
PdLhYmwFpmKR6LnSaF+pGVrmwvwMKZPxZxcAEfCQFZmVPdYCuVFVWmZEGV436ZIXpOKCogBDkfnb
ZP8n/f6tA1aCylvI0vrQxjGPJ0mMndFYubdqXJHa45HVHZ46bBbApQuo2Ab9gZj5IETePKMRCIX8
DCdr/0QihSLNL2iWnKBXua8CF5sPc2mRZ1iia+4LtjWXe8CO9JT/uGsPy7NzxOa8MVovvfF9FlWC
Xbf24oCKoCHvvsWCzXsqr6aWmFyl8ySMgqeWNDvLLPL1QrP+2LrC1rcMn679Avm8ufSWh9bjvsLU
D5ikEjDkRW1B3Dd2y9nwBiIc8WYHe0StCknDbCE+yhJ46Cq7BGShr6Zm/+IQbUHmqdnaMwc3ou1E
A27jT8vdUr+/5KD2xDQckgaIeEZ/6z1njXNECugZF2WynG8wUgMtZ680Iq24yCBnIjb7w9oeEpyZ
IkEGn+niIG3xgORgC3rU108G3r6gOJSh8l7TVkodJpE+Vl4mDR5AI2LZwLvJdoYx/TJNJk4JdMdv
2kKwGBGXNUlZscnuD8aFKVY/GfzAZvRfcmQC6SQ9TN+aL9gBiQLMKyafu+Yw8+uY6WpyRM2h9731
uWbQWtB3rY9DHuTsXepacT101gRNTcW1F59tRji++O0p6PYnDh3EKaDr8ccs/khe1IPCPYIZUF1j
MFK/9wIasE9/JJzFxhFlXjMEMKctfESSWMFoqVVC5DwTyRT3wYkMHFNPQRoJpARX07xi0ICv7wrD
WU/8HKrOBnYeYKqK9joSOZJAccOj9ggK3GmC1Usy965EZ734vBwkDKJav9p2DZfdyd277QHwAyQ2
AEwCy1zos6Zc9Ar+tTXIma1ve/Kyb2/9lsvpbHJAwuvChAAvjxdmruG/oxLWf1XDssjw701jNIaC
n5S2go/tyLo+LZaGVX2MpB9q1O38d4GohO6t+b73vVdGEqcUYWn/6Rh/JJRfC1CejAiuJJir1Ndr
kXMpBz2dRsXWiTWlIuIcTnWb3ogYmksG4Pa3LV+J7PQeW0Q0zbLqwwMu6vzCBQsoCcgT5JL0zJdC
Fv/O4+Nss/mF00qkhBFTY7tMIYx22mkIOJlRMy4amHscVJJLTZ8E2fB0dqCshbxhJt6Qp0gV2E7D
X1pnRyBQAoX/0ElPwOgQ94Emyh3715GSKT1X9VUHIXrWMnX5rQquhsWZhc7LO7LxjunQPFzf9B03
iiyz9aAXVVIvstgsSWi6xsAfm0B5erGNHVsnNuQnWl04f5o4wFImt2mN3OPhwP3eIt3/cTKbd5Hp
DbO84yKewpoxDcEg4HMHIGOiaMh5EAoxv4afSg+vUOg4TTYLUL91BJduhPKcc7Hbe16oGbgWZ0QV
gmdNO/I4kyZYlNK6bDXPRKiwnECSikxQgtLkGjWl5I6+LfeRcNZ/f+W/lF60dUk7aGgsRvm6yv7v
yiypXv89D5RWCaWdSQ1ZLMGx/vNULRWgK1By96RvReZz+O5VTY70u60wz163PbnFFuzYT2G0KccK
KYNBf6K1/gWadC1CVOXjSl0DK4ZsfzhaaSGgFMkZ1o4o9VDs7eIDJpyFh8x6DKURjbHyQVdyfTcn
2CgXcMuOtm/Z/WrRDPiWh/eXaxsN6ltfkXGuTSy+ZfYIfupTNVSU8o2TwklzMiCja41C6yvPCK/u
8odAvaYljLhRBFRaxbqiQ5OzFyna0JoJL/s7skp0UuAIDliu8FTAfSI5s3KPbD0Yv2UNyyR6sG/8
XC+5VmjsttKqSdY8Lijaa16Auk8AJSH+uxixgIjyLWXJMi2mlh4QDRmzxrH505OM6hkg8TDM5Tv+
J1TBQwkdTBdOZqOqTGPFgXpeO5ngPlyogptDHYl/mJbLkzeCe3ZmsK0TENZC9ybESf0zoTha5azi
TjWgTslsUp09whJr3nZv3ILeR6eiqYIaTxey9nvishCzM0RJompZSZDzav1lp7Kx9V8wus7lEe8Q
Uo2p6Iq0g03JDVnLlayX2g9duUBvOsKuYBztdSFnSUdw2AzBCgl3NMB0xspp1PSD9XWVKc2mvtdC
NbQ24l4C57yHVk0/H5E4gWv9LF3T6xb8T3h85EYyoa/ZTc/4RITSh223HiCRIfyOvPb0WwFoLuyM
ldGT8fEbFXNnoJDZ+0E23kJ1eKx1rvDd30NljCd2or0QhuqAjs/3hmhxM5m23ISXtixUDJw1xEjq
PgvWr4dwuZA6Ybiha+yklX6nLafGjita8urTDxBhb1gft6M9lnSrq4RXkAllNb8FEOS3Sxzktlol
MQnd5B7RjDfBf2NpcMfNTWmrj1OqzZ2WnYjYbvzeAdHxY5dnCk0mJpm9jhjnf5NfV8ozz33Y5fY2
qs765QaslyHaakZrMLdghZEYY6sEqI6bZCdAUhdgJZTlyiGnZUDlcAKcoliD/PXEslj/eo1npY1s
jkwcJMm/17qvlRP98RLGgshO/hujO5InTRYm9g90vQaYMdZcCTeki0ad5aR0iLj6dhShJZmxPAND
zi+zwEqEg42O1rqsLyB9ZlZNL0JT5CKu7xK6U2DYfZFw7eKGAQ/4ZMEY51KyzNG0DkojSetENrGo
oakWT9U0txawiX0QEp2PJJ1nFTKMPC9E+I97pnjeIZ+4UPgQmjCvtc6KzMkd6aD8obpOzNQEymM5
vneb2WyYWxwyL5FrXY/gBYqlVCWi8cpP/hELj35XwQi0yrlLzzOzHWLuVueSZ0lk+SOGlrLaGctt
jTnI/UtK0crIKGjtUXtW8bNmZ7NNga+nxzbhX5lYeHhsHhTxhONWjEqkvbPHcJikkaDOL3zkhskM
e+yP+ZDAvl2N0R7gnS0wSlqVK68JJbsdZPsfo+Wn6t5v7ops5G3+Yldr9XRdmxsbk6DbFnHM49S4
gCia6dcvrauc6BDZpDsAsdf5RXcYgtDg+qd+5vzer65Q2t9ilJ4SoUWuDWCxnvRuL22e/4+hwqQm
UT1Yni9T7B40G33yoCUKS11ndHe++h2BejplU+4k7lTQUvYODApQo3MbZ0T7cROa3iIACj5OoSfq
s40KQ86xXqlJ9f9NCJriqkUzTDnFtgX6x+MCHl5wZp4jeq9ePOCDgvuH2FcYUzs7RCvUKQiEwGa1
c3+EmHbtNEbnEPZeCWAKP2NysVYddoU2k7hN3kZg66PeHHZdYfpkFZsh1ORqRJWp+Mcgzdbnf+4H
nMPU5SuA4LtqCKFMnEQwJ6GxPr0h6jlpT6ed4P9MO4vx8e0RzkLjJiXoVk6gp7n0+rxhwwP9KIYG
QGaUx1DHTt9pE0ZltR/4hXBLkUEdsa/HAAYgHgpap7nDN2DLh+gQnSs/tRPvH60WsbE67SqN0NBp
3oK4EEwH6ITq/TOyNqPhGJRugeApij7WaOEe1QjiUzvWUEAQWoo0Eu/xtHTFGNUAoFldwNxFVWx2
7Yn2WNG6vQ0EyUJc1UC0/PfrHeQ10XBfY3+FVRZqX2o/zF7TFRMy1hHwhXXPqQtjIgvJaWXvUGjw
Lchyeob66hp1WYGylDwGQZkziVds6Fz847eFw9ucK4MuhueIytZKvY2Bo56y78AtIH8okqpmmABu
2P37NSLpNNXpDXnc+gMQ7sBaJ9LzVGIpgS22mQ+n37iqPYhLufkcrVLzhKLCjP8Tl9Zh/BiFwzJi
j57dYsARFmbjfYE/a7AVezTPNSjJqbjeitQAU+CzaUepyaPzAbF8v4aY70IsOOS2G8NN1cufu7Nc
VWZC+U9pd/bKw6LygvCZV2kGxG0jMH8/7TqdlIIPzgDHLHbs5wuidQNJT8sgEoT2gx4BkBEcMR2Q
AaxjZYnPmICkLmdxfQ9UBFs8WKuJ7w4BzpDtUNqV9Wb8BU5mKTEP+KI5HZS6MkSlbtk+/NpAwhnT
ozfUyYitBW41HkZfq7BccGlLenN/S9985CcmicF5tUiBxw3yNuC+s2eMBmHpzi/Z7f3cisqIq3hU
0r2u1m5I7YDZGGf7+nPDG3pgI+sXuwNF3o5vg6BpJ7BGmI5mPkEQIIEbbJxqhW9PrjuSb2km+lj1
oYiQ+jcOAnIfosmNZ/Ir/Q+WCXDiINttxqfL+WO2qu9fOJQ3kLLFPsUQDcINdZFPSVM0Q0aBjbDJ
+GZWrulmoMA+F5hwrheqMFQ6ygMeT7AIMh7xDRQCw3VIRbDsXK243g2YTJAIJLoxon/MYD3I8uZn
olDAPIuez5CQ6KHxQ2719msuubhJAJekApQOTGxIdAVXdTHkTpNzPkn6CsVeb9hZckEjVwziM+sd
8Fr8LYfYL4vmtLhBTlP751Y/7MurgySltARSQvm0GiGJtdd9MD3Q2ugU6dNZRS1qi4n+g71ObZto
Xm2iPb2jbK+IZfObNRutS9ndPZGZKMwOVZYonJIo5wxvQXYB+OG7cOuToKmIJqr5dpW0HL+Ke/8J
/IMaXXG6C+QHH1oP++ElSYRxeYn5AILt9kJ+WDyWbTLhkboeJAErOSvGsxZwo/y0B50TNgMDA38G
W0TDBPkJARhyspb3mYOQjc3rzaEMK816Mq/PbMw3m7R0nDGMY2cz7VH2OpIamHkWIwh/mvsLYnkY
1vq1EvPwi3VBxssVQeQQsOffx6W2Kc1+LTdXJ0HKv3GsZ6Tw5+a214K2r+OjOh3eLGBUun1LLxRQ
dZcVI/9wbIAfaXeqS2dxNS4j4u656XRT89YiIqhNsVlxhoCMq9zbnVMv7Hnui9KnNSO4njPmSfy9
YrghlUglw9K19yYwvXJvLwhbSAlrtuNM6eEaBisK37ueEgYsR3yK1CYV/WU6n846FEqXcTqCuHX2
7+7cuD8wEfZMZTd5wYtyuH5w0hNZ50iNl4LRMTfGQuqSNFdLa3pdc38XakGSZXD2sraBO9CmaNtM
nc9al0ioc4+KQKYAT5E3ohUe4TwJAA+/k/bhU/cCTb/MfC2FmyqIEtqTatWKOhmqGPqC91bQpuPw
IYzK6WQqnA5GCVaofquddKetAgqHR+cwK7rQSNiTRv+A58djMUhgf6sdLMFv2CMWAH+/cyPXfXQV
T9DraYXXGzByxDrfhiKasJUKCH7EM4Q4tB3He7pLCZDMlS59QrAoeSV5yZAYV2ev6iqKyS0tZutd
/H5m5AQw1a5FZS1jglrqIfI9VZ3a/r0QhA9McdwSgElNEVSTW+Q8TRWZLf/eZzcXVwgqdUrq2cVl
dFE5pJPhYPsW2uCr0hUiH4HaQjeet+QjwbAUlPzvNThj8EeN+Lne9j1eblOpw4FLiVExQkqDIP3x
JJ6r6RlOOXP/u3iv5QIpuuRrnhja6aqG7SL4xFkwe0xcuQqTdyJs5vUICysT/W8VpMyhOWHtWnxB
NiOF2DTDl/fzG2ecVi1GILpIlp32uM0eCGh1TblOY0lD/PMIj733iD8HomoFlkIF/Fupw3HutwLc
rm+TkshJR8YlQk6UET9W1vjQUk82r1r/UcJItnzY0kRoGnh3tTgmJHk8zjTVE0TbhFUpijpTm7nD
syKwwDXVXhdRX3Y+cZibc+8xnd6bbaGeNdZfNZfcGy+Pnjh6bI7CcC9e0O+LEa+ClejAfSoC7slw
kBqzU+GLIX646Gshs4bFY/xkfyXhgJ2xsNdmbq1/AXgNeDi7Kuy2nKMH7gPVQ+O8lki9is3iGZAy
G9Vzj2IuOvR1ACns8G7PIhx+OdjG6N8qxQ3wqGbT4chYWTEFPwLjLjwGW/f4vWjat7jB3ulBSO4K
AqgCJ5SJJM1wue+a6H0ndbX8m6J5f3NBHCEL0T/kf8qfMgiLn7dOerX6hcx+CYCuE3F5pUMg/Eqt
hJGiBGa364n6kCoKX+jSdmxpVfhqFEdyZV6TXCAmRlp2FWWtaU3LsBLj29gSmzxZayDCnzpN3NQF
vEvFVl16+MhaGUuvkblbGk+TcgKSPwuSLC2+G/LGq9riL83/9+c7NIYD4omOuuRt8LiYHy3UjGn7
39vQRtcWDI7O7oHWK3jUltLDGJVWkZwZ6q6sZSOBe7j0Vuw6B0CuV4VLxI73bEg/86GEQaC++ymV
KdzAU6dn+K8ZTgp5I3Ld05V8ER0LkKW6Aepil+uNd9C9aNYul2m88DzJRciD1uVYJBLbS6/rCDvy
TIC/lAWIpVFQKUCgLV2Xl3bv9qnE5GamJhQWeLjN/x1TZFbLjw8NSPdN2wBi5pUDSElgCHPhoTKb
Q2oU14wDwm1G++qmSddfegoIO/3D71lIhwXWRX8hISEesGdsXsVykz9cvd+OtAtaYUl9C7Oa4EgJ
N/q+rRP1S3dnneKt6dD0TuACLtsk8Ae3r2lRXCDizetexlfmaYPl6mxOvzLifdMS5upKo8CRUqV3
bWQ6b/0uLl9F6GXrMbmYxngf8ZJ6IBZC5lMI8nTaj+Xi6uTl6SvtjfvipUXpL0ZLzrfutGTN41oq
JUnZ5cRcJtzE/noYbHCap1qI9UnId9jZAXPkAPt7B2SQ2NRn0DCbli8WboJy+lIDfC3vVbwClr30
kx+NYTGVR5eMOW4wSxnVhOl/YfZL24138YCHaCX21yYWjR1U+WBmzpIUoNILp9mmvcc/kaHOAwqG
a46saU4oyNbpp4xnMUhNcHMhf+hvV8GBl04AHUWWBv3JKsQMQ4kE5XNv6G5esT0CYav2eSGvmw11
lqHNDAT/fok/Hqg1UAUHqBaumd7OJYqIP92q9Y4FFIa2vGetscrjwsocwuGfeig76JjHxIe0Voz5
SWELO/8fTlbnWE/G4snF9UAP4VjVSM3Z5V05lCdoMrmZJSXAXJm1mxL0en7mvbGkEFcU/G33P65k
+7orIjY6xjsy4vgh1rtLiiaDKXV7W0oOuezCvydDyLX33FXvB3YY2ZeV554FkkRa0taAucAqIdSN
Y4B5rV8oly6MCa4KdBuNse+fKvmxAP2ROIhqD2Oo5+HVdwjWZKoa2kiNUvnBNxfb+9cJ/5/Mvd2S
y1xQeRyBzFGw2Q0FXpcGH2AKcw6UAKh5OYjxLqVOyB0vKy3aOI2k/4b4pR88a1OKj1BCuIIVFuZw
R8oS5UloVk+EEMl9LOzvY81V8lxq0qh0bamSXu+LwGnNGMTgU2H+ILr5xmLCmNDHANmkDOGAESTw
3qmKHGQi3B+NRYce0HGVM10AwSBG+XFPD1SVJtV+jiHI8PMDPtxFd6LBr30Q+ULHpiPp60wGQU0i
lwZsCnIEbFO4RP3tVvWdL6ydkPcG+I95sM4+HhFsW3LJ5JTczlpnGwIrSb8gEeHOdiOSPsxwf/Em
mKjlLyP43JA9jYTL9o91vS8IRxbv6klLV1kANqCA8Up/YuPnYY1Y9hb09FWsiL+A/lxvu0EgzNSn
8pAPY7MGc0M97CPBS7YF5Jq0R9R/Vn53gklX495N3A9y+FfppuKslbNOHgMydvrxFI9v/wadjBrF
YZw86M/YQlCA8Pywc0ufZIzpq5QDv0bWuVh7TLJz21gtZZONoV9FX6VaovSfiQmH8xeyQPgiSGCb
JgddH2v8fYJY1bwkE6NAvu5ofKCAf482ggwHMZI/KsebocfJ/YYgC0brTSUJhuGqVH6RUWQAVwVG
Afxht6xyu8kvFXaZeZAqOO1c0gozgPVJPT5eFNRMZk2BcbD37LC7WIL5qVOBVKm0uxO8cRdvQys2
a/UOUggchXWIZGRjOL4v4ARLdRo8y5y0qR+OePYgxCAcmg31o7qBrScf608us3nKFClulV3ethQm
tZGtOlTafxiqGSufEBXvsKQEOgEJTCZiUtHne//laxJO9g4zARNbjszZIiVURjwQxl21F0qsA2MZ
nFlfMZY557n0fW/oyB+6/Mj00MjTewLHfssqnCCHuwZri5fVJ7qzH+91nDz628Yy3HLrNSpP1uqT
oV6XH3hMt/Jbc8YbWI/q1jiHRM9zCIheu/Aj8Wok7JPlbnFOxWa4QsEXa0liDkfjbHPzwuhaDXiU
UK8zNRUSnYp/sNjSPwE01hB4WbaTnk4mRzwXAXy6gsT1HObTxR7buBR3C1Exwhc57cwn6MYIv2QW
kf0Yi/cwfK95fxlMLQcwbLU7RIB8vZOD+BLvhAmhP2F4aDEbomZS/SW1nwkeyzLmoGf3ZbXPsCT9
Uw4b70a91jOk1mYtZoDahsH/r2xXDexVnqmo3u/bUC01pZUJWolfLSPvdzBF0upm8N3VLGvW/soc
Av6FXBFqYDKDwEwtpzS4ysPMdrDQVrheAL3CtCLzrfIyxnb3GLlJ3lE55+qPW89uY2XGngX18UE/
mSmbkTcsEvICtwa5OPSalNuxi82O0qOFBF82HSfpM2xi3vtxMLqFDL2/5rTt3mBcxyFDI4nBhrKP
sx7u/3Rxe9/aOmdto51dPhksDyHACupv772Cf2tCHqjJ2ODuSExZYgAzvBz80jBLVau/gvksxtXY
PXl0aqMk0RtC0QnYf9BhAntIqbY2Hu9aikxfKV2862D+WCuBuOMrNvYJgu5qiC6dPGZ92VpdBKi+
K7lUr+o9IK/7wfp1HJLsQQYkp6LvfGmC9wBchmSdYF+u22ws0jW2HXyrszR3SDfVxaSdm0Oh2sch
owM54cuTzLUH7AaXPmYIbWQ1JjkdBtDQTo4V+1BNfF4qywN3EW2hl37x4/EUJMskADS+d+nS4htz
GQEI4z+2YMWHY0iIfQYpVpgxW2FYCrmhCk8GVdHD6YD4RHHiMpuwmBMfiIWqMtsJci0rH+yj6Us/
eE5csjR741apu649lgrHxp4Beb0zLcQpCUwIxvOV/WG4Fq1AejVPyi+g8U3EzSXEqK7kCxiI8TZc
lX8LoOofooHzWBvoVKb0GQ/6xDk6d14OrB7egSmQm+X6E47j8O4LN+EbJbMTQ4hGthmhVxBplXQv
RP4gg6hWW4woxYvJx2yEQ6kJBPGQ1bThMLH1zOSlq/4iKxtudp+K6t/w2xVGOMkLxKUSih3GK5WU
Nz+ii0M973Res25yDT3FohiqiNOnb8wTSnzahDdZ4FZLpZynd3Tatxzda+0lSEwh6lf9DP00yc1V
JTVKXNiuU08rR6HgRY3QLNCMAm9th1DHCy9MLi0BR2fxgmaUqYQIQgqjnikTcL/LgwnQIo6EGRS1
HYBpd4apIAgr8cwJ3jfXxBBy9Fl+nN5N4jryB+lorFXVPGx3+IIMtlnhW4KfNCDbucoo7Jg4gp6l
UHkmqx3wgadRGd5OEuonAm6LyrGZPR1G1Enwhz9mhS8tz/Tib8C7aFoNzPQaKUd3OKoOSiaPC7WI
P9Q6P/6h2VNk9Pf8zCRNpxhzMs7MeERsmFAz0OBw8tpgGVT239ZcrcVAhMvTykB46WAELfBt4caL
MU0LyoMoM4pzqqsavgUN1G3J5zEshlkLfCw2uYRG3qyLhLRLmkISWCpTAQ3bbeLiNnJHRMSLta1t
6VMUYtNlMVUILcTEQzwY2/eas/dmyM/5xOZ2UXsrtNjECoALf24j4kj5WT8VR2RKkokUMGLn0hP/
dtsq71YjdHvK1LiFQ6pXtzGa5jUMMtKBIrXBKGdGb16wefkC2ryOIDIbkupKpyY8ZhIp9oLZT8jF
fG/bEODvnpyr7hiPuYdnPnd19OkwB6Ikmj3EsqumL9MJ4uVTEBEgWDUL6fMotwF3iakqEgtEU2Yh
UA0qGNIURKdvtDCNn6F1jQMv/2y0IOtVbQxiHn0qSp2fU9zdw21hwhWwBCLjCh+LrT5F7+bCDk+j
dF7n/wIQ732HdaVb/Azz91UKu+PS8Hc68aUNqMQYo9SHN/Afd3ygrB4Y4NToZjqB13NYE9qRsJGH
E1fsxpZI7vEXme5yeb0JWa0YrBj7teifyje8V30Pp42mRSwi/WvZLiIUvfAyDV/vOaAnhlk3/57Y
zS5Rn3uq4KBeAFqR1NGYp+RH9fup5ZACCS8AZOubD6gk4UGslbt705h+YX6l2tVGfGeaT4v74e1G
b5BXh0b4IfV2kLZwj+9jZSfGri/EYEGXz8s5miTwbvwNLlEO77AbZCOhxKP8GhmQP2EA4Bnar/Xw
JAG2tFZrKsVbxTHRX1mNk2TxQ/fg3/meq/uKzja5DmVm/Gn/W2j59FBeA0MOv2KhoNTLU2JzX41/
CfPnourPRUOCF9PsNne+0K4F6d7xcDXgCnyvBHb/I120hzD4OmRK5YrtFjELX/FZihcIWYgu3zNo
CZxcHH+jCOePxaggWqg7XbXlqoogxCfmCnITbWJ1is7E462rOOdmQeKzaTUulLaGaNM4zTJTmqF5
2md34VjOm7NEqY8MSR66NKZUExpTCjGXn+AfgFd6WwKCKIeqbL8LxluIAaFa0CpMiqr1XGAM+w4l
YAiiwxy9eDJN0WtqLluTAyaJ6NIsuVkJ4ZmvWUDjcow+0aap4uCH9uMpZ3rGw54DcYXnAwYBKB2d
lrxJH1vIRaIQTyMuyn198v9Tv9EcYvbOGA2/vBdNyxS0vY4kiwRVBtHyBo44mpdDfezw4LYUT/Ie
EZEYXVA+/NEPOzjzd1wSpFCthfBF+OBLUUmKTvGimQR1gWdRPiWZV9Kqd7Td+g+tsrbxYXIirtrh
5wANRSjX9Gf7AzkMQgN8ms+gMJx0wWId2HfO4CE1jC6CU03+vPKDITwjAHs/nHSpSuZ4peTz2sEr
dO4mv0BQK2/ofHnjcfhst0AXUxhRmf0wMchbUHxGpIUMvCfUdjYsjnvI3a685DML074jX4SdVnlN
8Q2wUa7BrEkYD30WfV+sF/74yeRnxfytukv5hXj5fm+9m6Mq7o1LNuVLmschdeIt+RqKkYsu9/Qb
k96Ao1WGB7oNjyBZ71IQoSeP0aJ30nVWwDQ9Fv134+bH0Y/MuOp6x5knDr0yn87uIsSKg3l2wF5H
Rq2YARLKIihYTvlj0iElD9g1rOb6vrSjiH3+KpUu+mv75+mPy3+kV1xIeG8Qz6hMszmilnJIL7Ur
G8ZHLvFs9WaIJVXEZ6dUTkcqsI8Xqr+itHjnZwZ6kMx+zY9eT2DwBAOkVcI8S8+pkv55qwxT86Tc
f3VrJXr4V+FU0BzlvKOi/tHunbUSOMpC1dAHDt7uhCz0CtQiNweLSj2c8tgHBqrGDUIiFZocoTQh
vFeduetkP46WOHkY7oggD67hSDyMDESqmyKPwkcrqBpUCFHjSfOr4mnO7cQXS7Da8F0Xjk/b7fiY
r18OQwyFR5QA58E0j5gfEbh5vwcD9zZt6O+Gu3O8jRsKk31RxuUzCsxh6ywolKNQn/1m5WtYVfLF
g9VkQLWCyKE0JMxNlXE3cdhNEZ2p7MdFNmRD+TwsDcIavWIVeK2brqA2YhAFHqaeJvSbqi0patFR
pUMNDbCPrCWuqxFBmtpW2ygHIPS+KKsqU7y0IOYpguNr9Q+d67l3eBG8ZGRN8pSXIyPUbYC+eXjJ
xZmdgysOdJ8UyJGwhur6giHFzLC946C0rR6HcN8W13f02qHjmzuZSgYst4cS+SBnry7CnI3+YZhT
/ZOeyHZWZT649ltcwDsn6hnqUPCloviDpYoa0QlOa1fREqRsPUmG0On0MR/vQw8Jl5kdhMLYDjEr
lftjg29FlIpon/hLLKb4CiDFmEGuaput9q6HRl6axImmQezmfOtLXk1Kdi5z6ozi+uliuiTTZcyz
97JFBTgdMiyVfbsv7mmOibHSFXSKZA3ktjdjlEA+h9uZlh690x3ZtMFUCZ/VQYV0iy+RyF7R4fG8
zRDdLkxu26uctRPSGdZ1g2o+pbTnLwqSAFFgebwi27fOL0EeuiZH4keihbHEF1tfWzA2u1/MhjMC
1acIx/w6MEai+8B7fJJ/Xi2v17tyBPabkDRKRURf0fi2ZwKtc8mVLzbQqVZYOUbEJskoL6qqnsVb
SqTGc91CfwlFuhmA1cbgV3dF+beCRZd0QsFW6BT9ckjiHrim9SgpU7DwQLe855xbfH7TdhvzWaX2
S55k+UI8hEEy/CemhS+I8P6GDHPEk7ehWzqNJ7YNMI+FWr2z7sBTM9J1YHBLhLXrcUdNjndzFX0x
wd5UXnFVByCt3cEsxfMQZCr9NuH8Wth6LZZIezUbLolS4nwZewVgNEXWGF1WtejjUNXfCKYq7cAa
xfGFVehF+Mns/0HibxtUsmtDdLqSicnzw5NJcRbZZVqewfk8kd/SOdxTC4taJ4zDfZPC/bym9yRU
E82f34wh/SUbkdKpsbs1ZvW073vmEt4mT0uiMp2Jmym7NMUDCklrwN+TxpGCBJMGsF/6H7Nbb6sj
e1DpZagQzNcnQpZcOxefXhEkmkY/cN+iNXNs9WDpkMEEMcdlHOAk1RGBwR9nPt9V9FtWsPAUDm2m
/1Q2i03LeNs6zB5WrAB+OEZFAse9w9OV63LoYAOXlbakOwS820H8burJA5rdotK9rEQde9VwcOlx
V9UHHcz4ZohV6P48yjr2fcxvWN2WLF2BKPWiuKjloX37e75NtIbR/Mc9fE3muwGOOay0rZHzzKMB
1ez49gNbZKzqBQr1H6+vWf3PjATIoPxhQvLBDk6JFnffKLGBhXjh0GjGA+OpjUOXARip+AmFXY6a
sFWdXBuAkem6t1pklGNIpo8/xEtRB86AZeUMGidYn1DCWtQlkgKbgTG5miQzFpzXVBf32wqAXYij
k7TuOkGGgi1VWwgQmPISSwK6Ead83ek8X+2msDfJ4nccALPILgVtOWtdLND9smjyqtjI67jyKsqz
pG0yXj+8KYY664/LTiIS8k1HXgzYZMJqCg4j716sFAfd213iCY9ca1cqtRKiuHlO45Ub/YS+3MNK
nlcPzUn2jqpiYwZ5tJZjjZU7D40rrvUjzlN4KlVJfQfGtWWKRd9bWlQWJ0l7sBMjATAeXo+nMFRq
/o9izmBBAaqatvst72d4pwWEu0wXI8BGkmYf5fB+vQhLmNGZvsws6M1K/mxU+dDrxK0KwBA2bP+N
XXI4Wja5Qs+iimHvcucm9mGi6Spr2GxyqChNrDokwkBj/Fdppvsw4LKGPDeaITi1Y5RGf4xSVGyM
vG9oHgaIFKa4xITAyv/oTHlwGVrLFV6W9kEDKS6zRq8k6kM+RoHuYR1DbFWGPZ4iK/N4yL0HW+WK
hufXDOwXWwSS01vaBFM0XJRj5TrM3Pam6M/saby1Fe71mH03hSFIQPKCLO75sUNsyUy4FRai+egb
Ir+ltpTB4PRfnZUdD3qW4MuF+vliChKWh2NFJ5MZzywHy+AV27neaTF6FjkgBkpWVbejayiyWOab
CYGgcGGqOmYTaP/o870pcgS0bMvwqANt2e3KMaT5nCAtQtGIpTgWIpUYHz/TvtkIb25/4bFUn2oM
l3Cqt4s1xUQo2FsZ30XZmn5q+8EuKn4F0O+Fe1H5qrEv4E57lWyTPROochmf4U+NRYR82ngKO7ID
P5aP/R5lOEMWe1fhqUbehSpNFwa3bvsnf4Cx0wEptP68JDY7bNqmmMPVb1eWvf7A3RVzdkcgXJ+F
7ZNvbJhfWywHct8UWlLQT+fb5gh3vNKXAnC5h94Z3QHNRmYWO7d/crd34uefVN+4gDYlc1SyP+5H
NzEL5QiwX1XZRWL8GI7564X0MjIGJPhC7GfrIPq9FnkAABGU4e1G6ok7wjwSjq4+euhpd2CLyAcO
oSYLjvsu80xfpYBgZL7+3nKHRGxx5Nh4WZgsdEq/yEgdRZwf48MgTag6BhhMMA4LHO8CP564H+/7
tx7MHKp1iY9x1RHFBTW/iRlfsQD0ar6NllTgnw3hAHyJmt2foz0vqOrFGDZ5OPxeif7GSz6z/+yR
M3oIwWMda6LxAdlaeoiye0dPqhQPsDJa6XOOOdN0IVinOXnFNi36MbzNlPzjfotU39lQFvCIz2Wn
OwVUb+N7LLd2E/xgmMgg/WYi1WU/dt6AphzqZUNe97AYEA1FATL5n/V3XrYts3vLsL98fqtmnnLR
f9Qw/pYNY9Ht/Uh0/FUy72QqNhkS5NsQP9D11g2EY4haAtxZo4IgQnZAunj78KBM9o5828fv9Okn
I9Pl8XUEHXZZAm/qnqqpLIuKYZTLQTZYzZUvv7gpkJxH3VR7qQv1Y+m4a+AESyBiYOm9/QojFvaU
6vKXl/EpTqQ/bCgD69TTYZ516ublK0pUFOj19iHttYA7gN1A8lIRh51ggAuSx7tJpgtioERQHmid
G//RS1pDhxQ6KfbqN0zPqrTMULZ+Be7c+vpTA6EtJvuJ2eb/SGQU7rWwh5pZ4DIJI8oiOyltw7II
mnOIsw6xTsETH1ByHgNRrgD0RqwH5uaCgObA2OG7z6l2A9zzUszlLXQVsiXkzJln762CDPsMnaI1
zqNNaOf1SdIOD4R5ZPQWkunr0ApRMawXPHffKK+SN1J2vhWku8IJBYcda9tZtTG6NlcCNqVaUdHW
oKmdYlgGcQyuwQKaXteddMYC9m6URnLlNfPCH193U1ESCjU8SMLk9vPUPfC6wzGhAl/uyazkDZEY
0n7zr4MiSFz29w2bMfox5rvLZEIPIXataoGJpyuncal98R4CVzEKHokAzl7uVPX0fjION/bAVFq9
II+29oeWpkX9MrOBZv/hmUJ7Fpnx5wkFMOc/S9g/xdWaL3z+ag7rng0g5puQcCWvQZp0uNvLkV8r
9IMtrOg3sKVF3sr4JQsD3631hNS3/zu2pUNkeb3RRM+OpkrdHHFqCvlRpHgATTCbVTCoqKGzYBXC
nH5lWIBLQU+fW0e3Pbe4/9ZkzAzSg/8Y1I0VM6YkVoNZ4ks6klDMS2jXSuHazqKFtTZc7ymSrz3a
Lv+JQQZrwCI8uajixAqMv2X83BiYBFcogUtB4vDJktdt3thxEog1H0dHbVDdbO17yC64Dumet6lW
4bkWN88v7HFHDdgTp2aYjW0o5/B2no5BRdx/zDpdryC8+vsfU8cJDvV7Rj3qx6zMOE0EXq2rRmWo
xY17sO4webC7g24qAmCp/fycjOkAQgPnPBmJYFL6VLioHhvrOgrT1Eu+qxTjyBLmcfyx3HtGfee5
RLZfM1nDCtJGPtLyBCY2f/w19Trs6lF8qRKwWqAnbTop6IH1mAx7JCoUuXTu3tgDte22qQrTmNjb
C/tkqER6lSEaWOuPupl+PmltZ1t7p8MQiVhzwL7uGVo1zdgSbxpBa+MwknQA+fOz5W6T9r3Hc5cd
jT5SILSvGhGoDI/bjwIh5duhlYo+bwiyD+GzxTP3amYX9Dyt6ZplaZvVaxB21S2NG6OZe5a6EQ6P
ld3/1/f2kg40bV8tWJfMT0qaft3POqlC6iOJuQ9Nw+2qfLKDKkbMvL/15X5Vm+xNna2aehg8NV2p
4Z/Zjbg27TNiErab5raSnkjpM9Xdepz9QSiCm5Nb+TsEX3bBru0CzRdHugPRNRcqzwFqrfVXtjjX
8kjrMJnUIMp5mcXoHC/dSAtWXjqLL0YwX+vbQYZUFss8zIrbsSEBJMtAm7UCYjwH0puVnF8g2Me0
k7Db/DAl+up27JqlIKKUutIz85ancYPTUQzs7oo/WxQKNHxYOZrXGH0TKaudGcDFLRAIy7gh56Qr
lgseNzF/If0G9YFGoaJ6BnXZR3G4ug9YoGM47UUUg4x3H5hYqupdwOW142PVedbILU6A1uboOMBL
Fjj8AEQhOfXvqUj6vtSNxl0tMn7lrkeQCW+OcwcfPI6a+/n4XGcWem0ANVFTtNI+wC4ekqGIqcei
QhrtKshtMWenMzDYln2B7i3Y0tlLPmX+K3GzVQRtSAkPKqSzJ3gtosWXgsv0mTjGrfeEe356DK2h
BpUyTgrp5Pl2Jt7jlyxQl5xro6FEcMZIOOnnlaOgeP6WdJBHpFSBpL1WbYEFes1j3W9J2QfBYQnT
G7SlwzxMDQ6G6KeQ85Ts5OwBWrfQHUM2cuAZvramuam6ppLVWU/WfuZxQZaYO+KnF+5M3MF6n2yO
lyn1rnqP6XLjVyiGc5ixB0OqvAWlViB/3s5M5c+RbWbuffD7smq2v6I95QmiFbV065FwS5FtcRqX
Ang/iAgAx+95p/QDrak2l9xRweBgyzkKlkQ0jSREcU4tGTlQEMId8FH7ApCMnGaJr8rfxO4yyRs7
LP16Th0QfWUjz8sgcYM//s0e43AWyYg8X0vB43FGK6GtedlHa214nZyFV8b5oJm6/p87mKJvtfEn
Mpr0KrHbfzdvNIcslxEsKsk6T65MFh5F2VKzuUTqn2vHuD6x4gasmPPHwobILi26cLu3DVqCqntb
JJrIpAYfWGoCpvmmyHEJhV9dPb3bBjo04fE9p5lfwggv2619I7yctPhSjwZVQmHru/l+2Xoj60Hp
J2ebYzlKZ8/I9UorSaVXvZfXTZBkpDerbDjM7lfh5b5i6GjuumMLlwYQH46rQ8kWsPnuLxFSYu21
6qkfUlcYEKmJNtXQZtManarU2bLXtGcbb0T8pX2cgLDv15u6W9zNPyFt46zuiHS3tX3T92UyGVNV
5dHAujAnZqnuNwUllFhFMTQkyEM8RfhXxZf3sHVMeg3KfTYsVX43FoboCxoo4x7FS9Zm62Qo+cob
Uxd2a/JDt9k3+bHzFjUVyK90y7oqul/hso8nygaaUwsQx7cNfFAi94nr/N0KZDt3dDloLfHXshrq
tUwvVcHHk2xdcwOQeOcIiZlkgYL7QvqxVqbq22M+GFOm41Cv6zux6Dxrax+uMRB21aTkZ0ehm63M
ds3ktf6QYx4WUmppv3QBFJn5OrCZCGKs19D8N3cRipwL2771lB6qsGCZSRXXYWk0UrvoANFv/JiY
rdW4MadDQ6Ov6L21Iul8SfirxBVdPVfTZZTmM5kYtcyX7QiDrty9jYvOhdSsYEBFZCPf82hgr/Fi
LnTbLccWMx7gv9vSmiUiFXBVOkIU02oi1/2uadbsU1iphxhPCsW9g1D1DmQlRReGyQAV0YuUihlv
AoFVcuu7nnrhdF5Ub5dmIrPzWyDvtpb07iJhpXIxRQj29A9NVfeQDcXt45PcOg4qZY1UlUsw7MTH
Oz7kdH/HD//a6M75LE98M33G0BFQ7g8/9EdVUIV9/rGdEHJ92WcuT8YO7PyPMRe/DIBbuH4bh5a9
6xfgv0BfTw997+Pan1+3ClXv2JCPNAkAiqIQK3fQLrS/XOXnhd1Fq1thN3vez/zCr9GiX52QHc9K
WONL0kE8kI8xax1EdAXUsKgjYEQpI4jqbgcq9PSx7XgbmUOfC6pZHG62LS2Syw5evdRBMTdqtJSN
9qQeof8qY3J9a60VMeCAA8EBWLTwKFJWnMwzI2kmrT2nIfqhCTAhOWQ+qgvFUZ2ThqBc30gYW0ZF
5pTX0aMXgBPgezRVxIMWhB1tiF2Ibpsv5uYUx6XCcOuimWSImGWAKNXlaWSChUbtq7licxVyV7jR
tIyEdYhGhxfvaCI+PEEOb78DzbUKAfNFX5DMcGGCfcNsb2JjUN3y7LcnUDPW+23bRLv/PfV/X/Bl
yYoX4dVFmkJYIpYX3iqkBCiv4mc8KUWeyrwd0pjup5tpaS8v3Ty9P//sD05nUzEtrF8nrpU4J+8y
gk9LX91T+x7+4BJlh3fDeRh8Jb8dIzQa+16eMPY+UGa9lWdGdzTxi/8ekjfmIX36cf42HQOxtjtJ
sVY5GmBvG7at0lDUMvdDJC5i1wgrEx4EQKQx2jhEhGa9Nmk46z78IT1/uMRc8SLmqeR4DGJIBGBK
L77dMALpwydGeH9c1jzYxhtm2XB45k830tONxDENMiSTJUFK+9eHGM2qCX0hc+qBVv9/ifqkTF0E
KhGbJo8QEwQ9QyB+yryhPh5Ek9qqJU6IpwyNqjcUmqp+XQ0Ug3Tjc4CpS/1M78sc6OcxNvyb9b7+
9t6ADHjIKWKdQh508XolBnllrEVCLigdSO9KRZnGCB6tqnFlGJcOcUqJj0O3UeFDsz8vcLxPMM3c
vTgcnEBW3eDFzTOwaX6KLYYDRHolRfFzBZ1vIwhfF6FRsjXngTpRckHLIaDKW1/vjZLA7gcDb8KC
tkqYEEr3cyRIHD9kfnBXexSFODWtXv2litkOH1yRlrrOTKC/COWd4Bw2FoS1G+qXb/AnY/5g9sTV
r642zYAeEMmBe+c0ecQps1jD9cdRkzsrMwIqPtajM3kVaM8hkLOS1sbhEhoIz1TkXn9jswjXfb1L
EOx0ccbgLJkIka7OdGMkRtzvzr3/4v8JWfjGMrfBBvMtdxnRhKJEDGcwT90eWTUU0IJ5obR/A/S+
KF4pa5v7Yod6PCDwZw2kXPvKM83NBMt9K4rhoQ+PGoVh66sRz4F1XNQSp0ifewMMmzlaYGh18fYp
wXmyA1wYbgVT1Wexd8ZUBTf7IrWWTGLECDq1F2KHAAdeJJmVx98Li2dI0HVI5DtoTSEnE5LL8Gsa
EgXhQPTo2mmK1OG1JhUnPuKlTpOKnE4+xcm09gzKXHDJXrE+IOx5N26NzKhxHFS48Mv+Fgbf1Xsk
KaSPMckoki0M8ZEWpuBI1b1KaMg5pel0zK0nUJShf7QznMzVfaYzdPmhysc58wD3zR6BAymaXAfI
bBrU3MriryesjAPZFLDTztmb9nGlSERTfGWXtFNBV8UFyGVv3PYxhTLC4cKUpz33bChky0hRz8Od
dsRL2gHTRPYnexPddjQd+qAjy0Fn3/Mk+JZf+9QNqzPG7R8Iod6eQ7rKYoWa/iQw/S0HhK2tTBNO
l+r+jE8gIKvWFHfRaddL/bjdpfmzq1/2pCwAbVXH4kNdwg+rDIUi6gsBwoSgYlQb/4G9oQmoLzI5
SuY6YqGNBTJHqlICmZkoSTQJV1/1naSigyz9qaqEFDMMESUgba6mtin2VlRYD/cgNIQ1KcdflLuR
GB3392Vsehb/8YcYQ4jJUI5oddMG1yDXnGZHr32r6JEb6hQO4efTzV3YeLhdZ3oguVcZriPDISDJ
WIXDHbNnntYaPGyfiV8h1+vijd9frvGiZqVZpEswtsk2nOayM750+2X9w3HZUWemoZsZaHFUTLtD
TTKwKNahVM7XQ8sessFdzGyKZS0+8jCg08w5wIk7uA/BwLRFGbc9k1DsF/X0GO5UTi5NcyDxUsED
5EDIAxI13tRr5HCGCp3h+DYq6NK7Bdhj5VOjEgMF8qn8blooWPewBGi1f2PNvDqWyXzna7BAJQb+
pSkEGUrhCYScvzSdxCzKVFJWBHme9xUsKMxlOX84bL5gAQeoqUdp3wrfsh5R7bfa0I+v8Iz3A2Qm
MjwjwCP4KewIADZUeM7S2kKZxrMdmyHSA5OAdd7CxRWNiwIanWQ3EbdmxDGlYy+CSVsm5hUaQHa4
I/2Gvhdtkw2/j81GlmOEdJorpDNz9UF/sH+3WHE8iLXOHqrnC+HrkQIDFPmmHowcBTfpoRkL3xNr
AMTNqVTIyWdC2jamsCEkNRjpq1YAI7a9AG4/ntntqIxA9qkwv4xGqpHSSK41LjRzEhzlhd28E9aG
2z1Na64RPCdngUp1nRtxapMrNfHSZaV2T4D+cFsyG4VRmze9SzUJlq07807KFs4auQGLrEQuqma3
F/x1G7Nq7YtNxzsJVXEypqApcfRTJIJ2Tvr+edW76xmL0F5C6jGdec9WmxIjN5kowiDk8DmbpAq9
PgHPyr9YTCbwDb2Y7+FNflNTSOkHYyKTGYonxtviladV9noB3xYZpWdHRFzcb9TGcnq+MJ4ho8Hx
Zq37Z44z+/nIVfZB0u4vmzHOV9gGv6dvT4t4zgpNlSdUlvuc7EONT2jIk72jWfziaG/2ivwAdRjB
5fTXBF6kpAZaEwATVPdmbW7QDuOiAo0dkpSEFtkgWFdCK1XGmsjdT6d9WNBP4icvdq+uu2NQgBTi
9AreJHcjx6wEP1eYDVRicjxbRNqi0FLt80LH+3T7ZT1hGzvI1Iqi1h49bfNb4x4KkD/ZaVZUQ3rC
TMsDC5IXhze1U+PyGppvYOwEDGCJxhkBGISYx8lZHrbjVXV1UF8VPngHQZuhulSh3RM3pXbjvZZE
FTGAOf5jmzoMscUgfdxFk11DACUifbn3Bra5+tMcmY9SBvnTLb/2WgBvu4MObjdP7HujtYhIF0N5
QV7dGjGScm/uC/fIoHAsSyB5PNOqOzk178MZ168dOicBp6ho3f5GuThvyUuUI+zwdnBeKv6q2O8/
Ryt1SGaXagYVnIA15LOG6eCcLaJG63xleGjuYNigncosTe9vxAXeqE5dRqg44LJS8nkNyaxg/ODa
Ho1S5xrLp7z2rf5H8C99PGvzh6tu5t7u8tRGAv7vUBXaHLcNfNLoTCyNvN3oOAxlHhaE6Dk2X020
2Fv7hCbbHrsR7LT3lRTI5dBW9iy14U/xiRp/m+ZvUY8mU+YPHdUll6HVfVmeyYXp6N8+4fbrWSvj
Dh+CfLn5IN5CbNMdqi/iY3VU5sT5V0eGICx0OGZGnEJWMzCzj4tleMy8HSso6x4L4aMpjGMt0PE5
xbM53FkMOPGHw2KaeTYxbpCvF4okuQpjglcLEZuU1sGtAnpIuYna30HBObbVrzOXUkwRWle7hfpF
DbQgf/KCm8YKEV8Bcxyxc7xFkLjVdxZk0q6BnuuvDpXZppN/M30oNG57eX6XoOOfam8ei9XIfwdh
Ifqv4yVnuW1baw5xEjiyVxjNAeF4LGM4epR3Ej+GU/ki8idcDYgFFms5x4vittKtPOxpQ9zGNrE6
8A/YtfXgI2oc0hGx25tO4TUdXF52DZHXe8fIX8zwkRnJom/A0jQ/CiN4tyt/X0wPF8/uHEgJL21+
y83jP5HZnd5alaALcV4SQI5cbbdUqP51nFSSJsceYHtJJI9Eyn4MpeEeznW7ehKbf0TZ0GOuLk5H
ebiDlNIcpH4/y70sSt/9o3ZBkzUw+aBmTzOo7Uf70xuEpD5h7+GyX6L5baSWx4h0mn/ZtmOeq/5B
neiCGozVVCBbRnW7z3L0YzAGAiPzZ3q2XU09/GZq7DMyNQ9mqbup5x6vnjOXHkzh3f922ZsPbOpA
APR7BmadPNoHpFnRNvANOJ5RZ7Kmon6V03tsy8wP9iGCJnmM4GYjlvCqox1g9gteGEScOWXbjZaZ
iun4WbO+WDWhzzRIVt8lC2Lt+YHTcNShWtFUlEAYrwBLLC6zSGcA+b216chvejbyxpGder6b12gH
wCfisDJBRMOvjhElnymySp19qrrzpbrh3rA65mDUBhk/yXPt9My5u1W8NQDSRqX7+gx/lai1u3L1
N67fFWYoydTK83uyZ2cKjuiny6prgQoOKlQ/xtz/QFIn7yRWHBETRWZPLYt/FaR4M4BPxhXU2k4O
dlEENdfZCwSWYJdehqMjhR2H9M/VB6WEiiStTnZ9eH11fgcrgSzNlIm7+TE75G6exS5/ood17I20
Bc2y81dyfUarnk4ZDTDNGnrNYf28MhMCW6ZBNxEOvB5JlSKEzOuy+stoPIvOAaVldw3ygaEEjIT2
0efg5nr9hZsJZOw1V4VOO6GXckq08R3ivU3ykgyep5bVDinEqZr/TVYuXObdHoFo2/HlFhc1mKEt
Y32kJibH/49iiLg1pOMs1AzfQrCfbzrcW9lY7ZWZH23cZ8NTDNMY3CwQEiUYC00w+6B2AcrE2dDh
G1/xWcOaS4lbS/CgXWNJU0zcHVUNzhTdKPF2henqMFNXdTp3Bt2e8nGEcsZprFqcCK0Fpq02tzge
rJJeAW3Y6QNcGPUftiSZgQjzha7O+P1cu7iPYCx0MOeUUWYDWArJvr9rFNM3O6GPcLzX/g+G2E0M
jxlGgPuZGY1OsxpkHjLAgh223Ae8YB8rMMfeJiYd3z8xAI6kkrxJHfF4Lk4o8dLQ/VQxlqzDmcFT
fFhcO7PUpH/+tG9lnaqpKoDU1utBtSDzppDh8w64ZCyCWndr6mvonQrkf3MCxlsPZD3h7k80VezJ
V20vxdSGLCmyeEFbPxWJGQyDwIAJcsr4WP7cXx41nLebIMX8bI/KsHwgi3e38WumyqiHsup2UNxO
6p673QHF0xF2pM44t9Ll6AD93hzukHz/zjkuu+WUpB1IOqBEiNQpZnUn0CO8ctScsh3xNqQgFj2L
TEsl84YLhW6OZIcoFEYYKEYVMwJ+mDnzej+hfJBqgAZFPRxysndgtnkSnFHslyaQkfffOGSsegGE
x5X6PhMWddCrit0JjX0qt89EANReVMsvxob9dvXvxjAgOZIFcNNJQPkalMjKMMPSxUItfepzaKHI
Vqm3j1TVR4d8dv31fNAB50zeaz5H3069lXoNUZDaFQl8TviVcZHs6t7b3SmwceDlZwsek7cioZzU
sYwNhrIFV9LbQunO/Z+fLvHedzWtlkRauAJDW4L3DNqTa44PQfPTirEALR+VReLjQCxzZ+CGaQXe
aTYmBXv4xl/Suhv/ya7YXyW63M4++XVxUJQmVhjLptkkTYk10tVJ7UWnPG90qebiXPv/NIQqkOMu
QSvoTxqO4iL5DMPeaPoWb6I/uQleFcmcPFsUJ3nuQkYAVaLXpS1JOBIdAOLmRwYl6/k9b9Hh04nn
kJTbhkk1hDA70pYN6E5CYSaslEq85OQE/ifkjWz+ZS03Uc4Xu4YbPnOGSFWCEB/ZRbLCoiD+pZSG
Yb+sxSoo7D/bMX9TDGvt1yLQSqfHUMz8TgRpfD4TzkpjjXoZbJ00cebnCMeALlXgUEQeFOIau14M
IOAE0BQ52EUCcA1hDkSSEWNo3pHYGFR9ktT4sAwnZjuoLwxzKPq3aSiOn3DwZZM50GUTMSQcQu8g
IjiUncxPuI0FmjVm5PRyWI5SqIw94Fa5BCv55MLnkuNGhQmnnCn3a1wTaFbw7ztBpd4tPxDv2U2s
dVu2ddSS4CWl8JD7vzNDnbpqeSpRNLJ2xRTS6X0EiAsTSV85mshvPT8n/ZXGrsVomrOcUscd5x60
qNMXYuvuK9KA6c6nrirVjf0n5UY0e499tggyElgCr7zZsUQhbhNMkRKP01JsVJU2HoqTgxA1XV/5
T1O/gaIQPSSva5MtTybN22i6aVlyxfrK2b6uq5LBPUkx6Hj/sxpy/fl2O1dPRqLSvbhEKhmQkJl7
XjQL0ZK7jllSkEpRiyex5m0BIzp54uGzJSTdziz1Mf61QvoiYMRAshCw5nRwVJdx+G+ebS2AGuKc
9ewU3WOdkyaAF5jYVy8AZ1OLdmSaKWMVUD4BsiCyLAxF2zuH94u0jY2MzmqojYg2/BCXc4z0B+v8
lmM2/7evNycb5yvn701AS96o76buaDGLYYF0FIouAr6l6zVngKPE5vaGHgy7n5Mm20tnY5xL9n3w
/ZmM+35507C5vs1VZq3qcj7kd7J9Ky1V1x/r+asCDBVU1c7l8P70/dDfAjbyn3M9izxgeX+QIcUH
54h/+7CEkm6zlaaGB8ClM4wij07HbMwohyZawNOLrjclSMhP2phosaYtjqEsgK7VfGkUTksQblrP
SOtawY4RmLbE0BJcv33gERnD8t/IwaGP2rLFQhZU8x4VsXFC7YI/H9lrVJwPDpfL1/x59H59kHxs
3BzdGbvi0bL8YcvHJ6VwH5iKP+kvwSctbxkE7CINzJzH9HGopWWV46juZBuBezfCohQQ70jZMxs1
0fLdwJm0AIDNNWvasB9bwOz3kTwCd5jw3gp9ZRQD/xyyEER99LPaB0bu9NYXxPwwSqH+QOzlFLs1
yy1wTyyzftxmo+cI5HpqYADIYGqx7IDMOGZvcjM1EAF7F1d7eXJM9OiBKrJIgoypdGVj8hrLLUcJ
StsTRv7wzhiSBapR969a0qj+r/WHFbBX62Vke7DGkV/MrUMoEua2c/Z9o0UYKJK2cTWA05elpz3N
gr2xT6co0sdXOl9nA2W5u0Bx4IfxjIipbDbMg2Y6UeC4iP9HNy/6KALc5+sZcl8n56xxpQnmpo0h
LS16tgWrLQMM0wmjJRTfnWd9iPPT+6vFdDoAAvgxPbYJIJ57xugAUr7+JofdgAjKh7cFFxJi9ZgK
vhgW5pY1an4dxnXROKPKZRHkhf/PvpJh9UAq6z2pp9j4G3nAYK++HPlfQURCr1PqZ28iXcC7MdSH
qd4SFFAgvQWuceqt73AsKm8m+jdDzUyBX98rWVwp8Y4n14yuVn5GjUd97rLfZmfBC4+pTgrSGOnG
3xpfa4I1lqbWqSYNLb5b8V0g4Llxq7Ov5priI6fuGp9nxWJ5dFW9g0ZHwiFewX1koW7M+0pDnPm+
N7n1xwg6aAmWX+7qGD01/55T0mTPz8G6lpem6ImT+eugwH8fspSgWY+QQFO+wnSfLiWoS1SOY8z2
5jrsjL76ATfRJkiJ0PAHkzZVh4eAAvbGIbA2QGeEdT5PiomZX4dFI66dszTtQJ/6IiSTD8nRq6vE
JPIT8EelE7SvjbTR0BYVK3rYlRI+9++dhzGyL4xvRXXNxJBERL/qe1ib5HBJw0aGi2jIg6skO6ZE
kYayH3VQiYY3AKdETgkd09rq05LuHtGuLVytmiKWIYC5FqYt+JvjNbRLKAmlzGND1whlQm07UkTw
/nfHx4CqIIzef4byVIeL1e23h7PdHeA6Gxy68YU5kastw88nFakGDZy36fj6JoyE37t9xrKO8lSE
b8hYQWB7kssKZAQYRUPyW/X1f2X6yVbhtuexCiiPjApIF00spT9QsGQJoywuEEoyCjPaHvwUeIFo
oSXtaylbTWNjAEI6vQHXfCTlS90VALLDHWYnRviCznWAGvpGlrQMZw3yBAg+kWtH1vdeVn6ywx0v
eCxmX+ESpCEVP28m0TrcDsnXqYYNbSVySlBzOVQxR9L33Uq4ZISQlNmgPoHKZPVfQl/aOJEAMTII
FHJlkb33KiTDagzghfdteATCa8H4LcZt+m/WXplg9rVrObEd8mbu2N3HAXW2z5aI4U85RZywqaGR
Uz42WaPBXGF62u8gNfmCAHe5nxN4zRb+gS/+5U6aUpRJXRtTVFK61+kVu5aFXu5+kimO/OLJ7Wh3
nsAnAcChBhx5DARWITmh+7V5CL5sVIb8XU6ZavaESI6YwYm7lHAwBE6zjrrJksT4Hj8B7v6HaOzc
n2Udal3BWKELi3TInlpQ5izA9RauXdCkfB8PVDyllO/kApc0fIZas8mcMb+/bfa5C7fJHA1MsAX4
j7RAeOchtSA3ucnbtXF5JDyJsh+S3oQhmFaIOvREMsF0Qiewb8GKoylIKMFoj7SOEDFuppcEvaIp
cCG2UDjJQa3b4IIDDyJkdg2T7bf6FkIFBiPmm+sK7v3FiB8NSQhAOGc4rJH/x0FDzcI1UO6+acIb
AkMA/NL/QaVpqQucNfL2Av4AI1EFJSdwJO83yZlQPshVMd3gN2IncOR+/Ty7ifD5qW/bEp5ZxUZf
Pte+O04YRuSbMF0LCI0ktQoDMfs1gfLo8nXy0BqgNz4tM1026gPJTsUuHJgY2ApwANGyMx0a4Soq
J8frQS3ZcJ46ZJMKVmVhHuIc5efvr/7Sy38fx4jTvaFB5cAX0W/yRsUIQikOCOs/NZhpmTg6+kiZ
m5QwwPhq7frVFZ3qVp4EI7xwZjrsJfHe7MIgDuK58pYlRyJpK+71ilu7PIqOUeb4EFxKra/Pvrfk
LsGduTTqZn2IL4IJjfawqVzJK5OtwVbJALZt2A5cJIRfn1MKhp6DqIlKM6Ydhqtm70eCZhUEEy63
1rkufcYPlE7SIlljywkXhXPqLUy4gQ9fweY2d9JtHWkpW2Z4Fc0InNaxZAogc+P1wVDkbbBq9GgI
LLLpLAYiBgrfvJfchzS7YHJVwBleRBed49SLimFKSQMxN+tZ9Wmt8Ry1LNU50JRMiaTsFxjVOsfc
YV47QJpStyuPHfhRPcvfRFEOuOoh9BxvGdtXmAZRT7AOcH/JP2TFYiGu45T+2qdtKtnWOKAvhEwJ
irHnJ1jGVNJjOdsKUqKmeP/7gG7vt7I6n9y6MNI9aqjHb2nLrmCaWxid5GFHFPJszrEIHVuSjJUn
KlaKgJ1ekRGXwZS8lo7UVHfziQED1aVxd3ijNZI7Y0UnebU2Pw9qHU59YG0gj6WijNQN/CTXBJPr
/UnpCEL2y54r+UVUrO2dRDuHlonIpioeRNKWVL1ntc8rF1zhuerqBVKsMXw/9xKmFGxrJakiF2xn
oZ58mW3ssxQqzTWiArAvz8msrjsW4kB0XYveLQPDoJwcIU/1U4m/GHrHPvYvgxNxGS5aZiNzsnow
DCNGyeS9Q+RmeGoN8JbYEqK749210EosqD3t1OVLiNHrXQUkqCoL9wioQ+5EiUA1eM+F+wwp/0wR
4INMaPRP/7rBXWYXOGyZwBD9d+FViCs4CQVEINO6MJFEAn84FunBnh0TQWp10FLVtYhBUXRV29RD
77vw7J4krEhKqZVegCMDYGCCcnoKfIVPnRrcxaSY1aCH27dRy/EOkM5nDdve8KqkwN8XaV5jcD2d
XND9jEhXzwlFPEy6StbVJCF05bsIedKTFXuYWy6I6zWXT4XcAw6e2O3U6pcmN9x/eKDi2WfMKW4E
zzxTAhcTgk1xHcokorSsKCjycv5uYH6ZRYRqvJ6LNf/CxtkB87TbcLXFHvs8OM506lEN31X/3sFu
UJckFfu8WOiZqUdbrVmALt4r9zTzMRw2szIHx/D+mglO8xM5l9XUCgNjYRRe9HiulV5Qxc/LKnpO
p46TEUEM9pXHq5OmUzOH7ZypGtuWguGaDhM8+X0gZaeHC8lVTAACrYFRbwi8Bvc5XRtyhbeEyVfg
k4rLboKjAGE9OuTqjgXYjyzccrHFPMaZMSM9q1rw2cKUCKQTaovP9p5DTSy//KCDBmSKlp+Y3pG/
vtleFxvlTH+PSlLZKxQSghoCkMuS+S5Gys7EJ4z5cx8bRH+f0inMp8h27VFZngUE0SG1nVWJRdlo
x3khaKR3Qj1YzvFghM+lh/NBkOtjzewMDYxQgGhSMiGexCu8zZArHkHjxnHYtmQ32u2akrxwH2xW
+qFYq1lYTPN23DqAPKsW6OZACvCj2/S0j2E2kIkKzBQQxzr5GZnUQseVDO+47LGZBcSp4BOn+8U9
rGXv4RTbpbR+FpynYlsgWlBN76txDoJU1cBnBUYKZ8R+lm821v8JBeNYWwasPvc7ugcNw0ttewAI
d0nvleGIH+qF57ROOxZl49bxfskF0ceeYA3uD+u6DAZJ8usR+EsByC8Gaa+uxXaIO4sHQMHH8KXX
jVWOil1rX+9eiAVl4tR2bh+q31dwhCvD/X/+4GLMiqhmWXQZbBRB2udVDgRFEJPC5FBc8Pqcdvog
I/v8/2i/WNF7jZDGWIn/vJrDNxcHV3/ncDbcEiGN6h6APLBr0NwKoEOiEA2SUYPRim7of6nAHJs3
/AY4fgRwRKC3UnnKj39cXsVH2M1LpTqtj5kMeQgytcDOT8yG7V63+XKRKi0YUS8j9jlLxyWbkyvh
Wiq1B9jPhz0FnmJiL76HkulzuYbUf4hMy4dFa+p7+LaEf7h0DW+vrzb+GysrCMBmLPxC/BQb253F
MgC9R+H6pg/iCsaHG7oyIuyV74napFA33Kn0pzjAOZiSehN635H1tzwuzO+LAzdU5AN3LriUOzFE
HN9m3ym0mTOPBEvGBUkzbOuTTDyxYyVO+nSha/c6htLIdQMasnV7//SxqbOoCeiWKKEbIJFU0a7V
1Bq7Mxq310cLiB22isW7bLhHUnaC+hKm+KMva7sLIrdTMCHRljdSQrKEAQ2sKMGAJv00AWJbNszG
fyl6eUEbXWq0OeJzfNR4Qvr8ADeT5ngiwQhM/OyBZlztYGd76pycVV+D1JkcwSpyfBcnsWT4lFT4
RFZV3zoa5A4SNMxB6C23r++540dZTAiCWvcvGqvznaM+RwN5TD0EKerg6K27KJOx17Ws0POsWd0P
UYZUbgMMtxIvainCB/Sp1xLF1TWzfkBnSJ4NidIAYqhvE7KkaCJXYkiMqQ1iJwjnw4KJoYlp2CC4
c+aaTZmie98HaYrsCU5rbKMDD7Gz+Ba50khTDEPFPBe6lPVccCz/XsMEhj19hmnFRP44p8JlHytF
t7vBqpOO+nVYnNs1Cq7/2yliSTDwTYwiuM44to5nLWjAjrqXwv11wARscd5xyIQD4QZTfU9YYWIh
sCZQt1VaBCxy2SPlOEQ/NFOqj5SqZvtnBUvP60snIinlzXh4eQJzmeKyfVguDdD0E3V0Kqrbv01T
S9v+ykW0aH0GThC8tqXoMRs0QJhCXYGQQW07kebNCUDDbP1arBacXRctSYsCNbn+cjlkRW247EZz
PsZrNFSxq9pxoq3kG+aVHeV6NZMUyTshzcntE4uKyAOoPkoJUlGGIjiF+0y0fo66foiyi5oJmcb6
CFcj+FNHoyRKNNZVBuuxSmWAI7c1PyPn6qvsyLUbP8fUWunOqLJXdrOrC1/+ijj24BUsSbySghNY
czXkf7Y0dGRAzihS5Jsr+YK8Tyvk/91rBsUjU1VaOY5AA9XwTBiSgqjlt9eHCni3BI7OWIJfkmBs
JG6vteQGnevz4R0OrxTDtg6Onmd24zkOPIvbRUjhAMH/VV3RaN0N7DGz63YfcIxeVGqQstwKjIUy
LOipuVkGu+VTZeJiAZoTngyKvUy3nzBG5/NuzI47yBT0GBcdHf7apF1HdAoYzAfF8xd3stxe+POM
I2W7k+izt/LtMAwGiAwUsOTzAntLs4aYR5Z0xgoXFDP+z+DzxJsSCVP/bPqMx+7eJSHxsRjwBg3L
7sRWJHeg4h57Hjb2J/JFxrtFfe4XTzYDN726Ab20XRcFT/i27U6M4ykZWgAOizzphFhfsmix3EQq
lRTyL+1Nbhwjx82wcXy7ZfjziV4MwuBOMKlKxH+uU+9Zy3zQl7nMu6eYovOlscV8ONNMimKtbqyG
vbghOy5Or6izGqziykw6lga7WLfhd/yKawh5uLhX4Yx6gvXODfFlfY+gfC55t8fOznZTOXeHUevE
bgPTskAJM7JZSw1fhhgGn9tQ/p1TcNqPdfzRHqaqWQqhjftd+3e6Kcz8anBYRuk7jevAiq1oz/Mg
7yz0xuzsMKdRUhsVRKfr56gPPcBGvlbWe7j8/yS2VD+R+juiUDi4wcwHuQD9hwYpfL8W9R2Nh81f
1GtdgszWVQGjVgAaRrfvEYuW18IMms3nT5iiCu52fZmH5e2m2ygFhrvC26LEdAwGuGcTIqzAEXGz
Tft1OClF/M6FJ/2bt7tuFj1QJP6lNhasmVicce1NtKExu7b4lqNw5PB87rl8hTV/OMpSH0+THhOP
RJsoRGrWp3xG5gpnFc20NPdKF6lt03ZVZry98jMACic5/HIj3xCSNSsbqTQIIzQyBXicJSLiKkNi
xngkhSOUKqvea85mMYjp5XVCZ+rPf3cz07MUGdKyPBrbZzj1Z8EZtyNdHbUdHtWG5fVwa+okze8i
GPXWxWGGjuUWiXxQhWuxKHYjRFHwdWe4g/n598rjJtpa5AqKvP+JjtAHbbpRxDeuja+M8KUSJYYW
NPYxVckXnLKSEkjBOeVmKc2zM0b2rxG0sFj1j6ptFyF7jvJDAQl293qc42L2iejBf4qO/uZKuBYu
wkqH0ZAbb+cG7tmv5Aj8eLP04wvyJdbI2U4MLO2YhINPqUAcOnNkSpPY5OoK0NW3f/GuIr3RZ2lg
HN25QbsgHGFrra3U0aXMkDFJt5BL1aI1/5dJROlhAw3T2OKpCGOziclB4JtdPIyWHWMyW49TGeMG
Azu59ghRWZW/wvtKa1UC92ZAeYcZgYoRzEPoyndHQVXaApAwYrpS+0DSb7nWVkxDDsE9mMw9Mpsk
s4385eAINUnY0RwL5noWtQm6kJGpOOq7R+j39BbPfCioEvl2tznIM4DJEx1jrUg/aMsw2wim5KpD
aj0Y4w9Yhc5BKUKbN5NPHB0Mf1jgzHA8/+Tz1wmw+Cv0McoDn+dRydDbwZIsBpf1H/HRPXWK6W4F
33gIJAMbdYUPxQu+saaSXhKf/oD7jsvwj3m8yBa4Sew+nlf3gvIhGAtSvBmCTrMvGmMkJFcQ/PUh
N3kWWc8CbcPY02WT1hQm50AKzkvohYAVFbVorG7vwdSkvxW/l5ODwQbdLbLjJDh2GHQ8lnV/HtWN
jJSxMGDtKQwAdDO5UPFeabtsTJEuI+4mZNoHIOuAGG2djyFdcVItVRT3DtMRdeIzJ6BEdRZnvHNE
coCHhPcKZavQpdVtiDdtk8s8zjcVghQOEE9WC//7vEtcoRWyLQcI9Q9ylwu9XVd00FjybCQpFNEI
T+aS5ayg0zc2qlKmZI9RGG5qJdV+/4RVrtY07jiJVjASolyqcGJ1SRs2F/1s24SUlHXd5D3TS5wO
nUSJQzCaELnLLJJIk+R0GiTN+dyRZXD5QHfmV+ysx21v7a2GR4+/dDRYREgtR/e4ffcW8OdOGWBu
Hm+t/4LEAxHnvF9sd9eLlzAXPbLQ71m2aa9IwdEonUxTeETlKFf2h3APjv7RvvITaQBBMk8P4V1r
OPSk3/IucilhCJSeqr6aWWUDmZnr2n47vkuflEsoLMc+GPXOSTj2hoPH3qghvkVXzGMCFdBEfvRx
MqCojosRsOsNcTSPVLKUlVmEkPwqtrcOiHPvSniR1yIJSdcspW3iZ9sZ0im/4OMIAf6ywQ6ggiVs
mAUeiQsLI+rbcNyDkZF5vz10Fi0d0vlFJYUgt+sIJWmDkyTl3H4h0D8Vgr9Z7B1lM1Z1BgIT5nPw
T1leqK3Owuc3NOVFV9h3xdfksJy0gNUqhpqOgryRb+Sxo8Womgkh5GMQfuKX3ra6zs3oBs/NE8nW
l9QJ2IApBezDBzs/0fj6avnRZxaqQNdl82CfaaiifI/MPeW66D44tJRZxrHja8ZvsYPqfS1FYVGS
5L9fteFqHKVxkjB0LBft+GURyUuIpPo4IesT+SpubtA9HOb5Lxxx1hk+UGchh7bItPfhfU4ehQ8G
jHbYjMFp03TzcGC93Oxp3T6C+4zac/jVdm00G7dHdr93FYQPQuaktsJQOR/BxQi3BDWr4j7D7Lbj
Wxf8kz3TtTnW9iAjAAcZa7uIAN9DDD+HrMnYjjrWnau2Cf+1uMPabkj1fGTqQljrLsQ01FVNb+pI
ZyCq9CZznll+kbs7A2jiC2feDJaPqTB1YsWRFn+tMxSDSjf6Is8Cc3Ogf6Sel0W0WlZNWsm9MJIL
Djhcsft3D3Q4oirv8K6TRy1YLmsvThwgKtrUf5aaUJl74q7AqkZsbc5DyuJjaltkEC0k7Ef+54fX
b23iT8pNpR+Mqk5zkjkNRhOzaKNFt4TXGHahiwkUHHXcgEYhkt0ZZ8jtsczUEh9n/b8xACxf3az/
DnXAx4INbPS8MpwqYaVoav7la1IM5eMJ1dhTbHhZqeqRFYsF2hmvmUD9PCz0IdTnmqj5C3ZgF5yg
4hGfeW/1c9UafrWg/Bhr9g2pBe2UOAR1hJJtdbYFMuw1UJ7h38DS5NvbrNhrv/IAhKacyUheOEzp
jQNrr0LmVc6E5xkcdsxUDqobq4VwVDm2Wbz1W2ebLqhUFt0PGJGEGaDBhVvVJKR3KiIa8wXBCxPD
LFRkXVbiAW0wOXH0bV3Jken60Pboku7HF3WLkGAFKlzc8kOTKPGbv8uVWStAptz68GhJS8x5Y52Z
PATUaISTlEeQQpyZN2nGKF5Zr+Nwbb7C3L8gK+bas4qmYZzEAcCiIhlVjT54y4oxd3nornChaEs9
60o0XhZKf4VCh1dXLkXpVkIXODe095CPW0LFS0hDBK1d8fVzXqM6GFw2u26J/j87AgktsXXQvJNl
kh8NZgd62YhxzV/K4hXHplTw8m1nQvcbBCQB3T04BGIkNgmKxToFBewwT7jcX2AUpBKEvVZvevis
tRyFORnCzZIeF+VIbOmNODoR81f3aKdHR3b1zDYxZ9MKE5p75ESaTywsdhPGIIJ9LsFzRqsp9oSg
HG1ujZjal7ssslW2hLqDyzbyBKvjuh2SCXeakjd9kmb5RMhf3eJFe9WZqS3p+RK4lTyRHFqNdS5D
GtfKAAcN46pGkbzRFpnFi5FP7xh3laWFN2/lFqvaYOqi0y4ynx3wRpMRbTppzxRgn5vA5XiX5xlr
ZiV9js2AnKqn32EuGMifTro+7ODdCihigg2xFXUH2nHexvnoiCceZUFGFiPbIoI5hslEUz+AtiU+
eHYZIAOeClzxVF23P2gBidOIHZYf2K/cHgH2lo8EAHDgK5ZWMxkDj66UIom3Jtny99ytHKpZ5jZo
u2U6VZoy3N4XhNOack84wQPV8zEoKBOpUE57GyUredgOksclko7cqFLyNXMuSmGaUi8g82dtNjwU
RJju/QjLXY6z9vE/iBPNVqmwpDTRrOvYnUk2hHm2GyN/h/ZTj6JyGgLq6cmp/66detBCVHjr7gff
ng4sbnlHxUhQ+4RytFYTXp4I8zCv7oCCXEW/JNwThKgQO1YZbe1J9sp9dKM1VU594dIGDFgk4lTD
8mssx3Nk3FXM2uKSZD/JV+ngc1eQpggnIojf35MAdD9vLHde2A4Bid0707uq0Y9OjR9XdeQrqLi8
0A21Lj71ZpE0+e+9BmSzKKrivnQ7gpP/yRDt7d7hhu5w/1nPfClJdJx6g5Qs4X5Nd6eQ5GgSDLWr
NmzF4lA0L6InHCscExCU5E60TYXnmXKHqpSiVI4eOnttBheqXZ66GmLka78XF5HXDOt6XD4szB/5
IEelFzNghIj/W9ThYfh8JXm6W1Vs3bx7x5Gjt+m9HYXFkPl4mpbAKkLzr7JR1n+lEG3jsjJUHStH
zNPKsoGPQaQLZEOMYpGJDT55ayNX4WrZ22fojddjxm3uoPP1iasqbAzyI+nUf8L61YP8/kGWkdZn
vL9PQ6X9Jz2cVYMDtm/L7EHX2RSIZSpRlv/b6MbCH7LyHCuiUIlMsDyE3o1vGMhUp28sGhu2Qr1P
yFZnK1HkgZbv7YneSgNQd5w+0bKpXuUdoSjbAVxhgMTJFZa7GaTPJyhGu56kPyx3tVHx+mVmbUv/
F/elyHEz72dITYDPk3Hofp1YJNQ1dq02zU8bVQji3ifqC3hqUFDZmdYJznV+D/UAQ/m/JRSFhkaD
/4VHT03KrSUx5mqsBLJJGvQhWltxlvmySmqZo+aqQuRB9UaJ/1/QplzEH7zWE2XR9sq2kC2XunlX
rQKEIyqwSwvy9EgOpTQQOUapAjNuN+rece/jb72sc318Lr5bgIbooVd/BRbQu+D5j3XBGicSFCSy
AkTYqelgXaTa7QSpEcASOYkx1nroQml+VZoAuambmTR7QA7pRZotKnc0qrfFuIK126GyuIVjr7ys
r1HpOv+BFwDONAT5LT754oyk/7RxrF5OUxpK4ODCiwSjXtcwoCJa6sOOiabVuM9533glMqCWCaAL
esSLiC29eSZLfr6MvAqxRgnUZYbGmKrexpHwLkp/efs9XvGmfYIld2ZlOUMjy8LbTHhiGczS9zDV
uN8O7O8tChpcwyCQ/o75j8wnJ3BaO0SyoOLphPMDJ6PlBRyrwJwAuUean6X04jOUeA7s38NwPLF+
TEDbxRKJpqPlb147N71YvMTiZbl5+Bs/lJ4Evfl/VtRtOfPHTk4OhR5T34GBB/CFb9BN+lmrlaw/
77d5BwLQq8BAIiA6Ob9RrLe964sgmG9YXwdac/xXaoD62T1gO5aHSIJVKdB6TPXMcRtDN/n5N5BW
B8i5iQH2Rh4blMndZ1E2WyCf4HHVZShqLrlxpGRSVuBvkuBRZr8sQqQ+qkyGI9XOyXsYzMDtv/jK
Q6biMSra5kLY9TzKI/ze4eMYMH6RmOD3a2vnoB61bN/98HArMSPU/cGGa55WkMkW4Ah9jVXmjmJ3
u9pblthra8Cxf0TeBS6tER4o3P8QTFacFN2dSJx5HcPpIGfRwQFsh4r/o2vKVlSWRJTYDvgTJy99
Co4sQ/tiTMzi8XWpyo6t5qo050EHI1RoXsFyOTXkRM+MGEfPT9/56YpZ/TUgiivkTMPxAT7JmYol
JVasxo73aJuRNkXogNxJP2qyRsuZjqOr1muAZ5nboWSE/rXxQmigyeh68oXp6ONzd1jhrIAO48zs
cnq3PJCB113FfogT1aZL8s/py3wwMG7nnkMgk2Xjssy4SbUJr0t7/113vU7UQcfXfcMxKNWxLM9+
+XsDN+PMCj/0Z4a79fDh+k0xoC/TWtH+ry0EZsPna34aUHP26GYab26Mkb/V1AXU3Rp/fjJjr+x7
PugJAWVhae8IVuUiDr0T+UIYFzE0hDgAPw0WtEAO7cjZsNupQCrw08yvGjIjZhGqjZZq1s/cg2Yz
rn0iL7y5gwRyOFa4HSH4xt+/esG3aXgpJFVgEWQTtfbvE+LzVABOF3wiPughR8ED8+pG6qIO6EdL
WULXjWMS4ze8b9OCFA8+PJj5r3kg++tZMfvDiJS5rctjzjqA73HF9OyYycNDC5aA5bBlnW495qo2
iH7lWeqVn/M54ZfIrI+yaruEUSmqSf8h49HjTtI1MIgC/8vCMpKROGliMimmba4VFETPp052gDdf
Bc+VMhUD9GWm6IEputUVT3XYM00E8WDQUmCAoHtAm8Bbq8cxLmuvXWQnjmZimriaME+FRU+LyYqP
NZygjFjN9qLJZy3Ao2eVd180N80UP4XzL5vwI07ZAxvDXDQwcFBe11PHO81swl+AYGB//3E/bik/
2wGW8smUqi9QAecEvi02WXr0r1mIyHPQ8u7clmNQFKKD0GloVlzYP9IsYaKid1vYi4fnXZ9w0KQh
Sa5h7jPlu5JuXY6pYyXjF0PT1GfFqQyqaGGecXmI1mF/DnRHKKLsaWqJ3/XI8A9P2fnLoZ6L++sF
Rlozrmru3QBdheJdaTyJJho4gLoxt4o5iiGwKlGoJiyf7d+lV+z/S/KbviR3nEuySE6R1IgatixX
9iLhuJfd4TM8W9zJICOB7n3xbOouFK/vVGoUz9ea7l3zXmU+iBT/xhF7662+WyWNjfs58cQNIeUY
L2Ozm8UVeIOPlrvdpXopEs7Iv9oNyQkZ8LWH1hvIPOcJWj0F9nUE5tpQo4e+Wsa4Wpisbq8yYSKf
69OFUVei9hO6E65yi71HUQCN+JgDKwgwIEvv2N7LxT6DMEKKTmh9wAwDxrx9BWFtDLYF5MnscPBm
t/nqDNyxJKSuGmLHUWajdLUtkTHhJr4iCwapAt1VD6EyZ5xEh/PN7oVd52qhjvC3FGXxSk1FqNSI
S3nvUzuC3NQxsdPClfM09ul/2vIYXMSYxss4ECH9GRIaYYw3gqFcBDGEBMN8mQKyqp6wuPX2A0dI
Dc/rJnZCcpaKbOtcjZd92IuVhTdnnb1X5gRAFuOqoQJ8XHtmHc/cPy3YzjJkVFQCBWXT35YyatZa
2umBj5PU/kITh4Jva2kpPsuLGaRYIcxxcRLnGU31D6+SlHKpbDcrLQ0Du4qVvxqZkb47dBHmrRPN
9GhoKUYSAKiNCJ8K0Y0aTlrg/1oY7JmUunQ14mYYLcwPUCclwM9lmU+UXXt7r5wFIYxHM2Je+LJT
BDWKXcvlWTMzxd+rSgfmy8NL7NcNKXqq1xddw4U5nIv18VkH7r2YefSx8hmaGlFgemTQ9ikaqvet
J0DqgJFnLnyyUvz4LCqI3ZSkaBKsyirSdBaU9E63QOTmpVYDyyjYNbJoVtW/NBq38kPS0DxZJdpb
O49HnIySO0b6zVKcBOc1kRI85tIBRaaNgYxQSc46Vx6x/3O9iKEb5w/rlINoI96uUr6cm/+Jp7H0
oMwvsbSbmwAtZ23deO7x1WJ4aIu52nsjQTciU35GkgwoyMjVcI63kWFtpl4dwGUjfzSwAT7UWhqg
qZezVE4ImijMEvvnpNVA3yxZIhRONDHVOxhIk1XP7YDjsnNtSUgz1HNLdyI7UNqGl4aB2I18j4fw
eTV6oN01irWlVeI7VROswjXkc0ekrzSUtexVibMkqOIJYTwb0AThJPg/sEPIOCwmL+ZK77K+cSPv
iSW7cqUR8AyVwaK5Z/OEYf/Nub00gP462PYIMvjkfapjItb/j4+cupyngd7FTerUoIbiFYgV1LYu
Ieg/1PR2ZOUliUmnx/qAeZ+Kwu8vrcVy7CkhURLfyBxsy/fZWT5JA+Jhc/LQh7IrYn16XidB4jWD
xKSkbQb1PqutMhMFkgkGmcPgTM5k5YJYqW17aNYeAOiTBvy3yhRaAVdHxk+9/3RC9pPb66jtQzYI
KJHI13pU4VcKgCK0tLfiTSx+t6JhZwPmxntlM18W22cR+fK4VGt433ngThmC+PUe4TQSFA3AiJu4
nyc+n/skmyQg7tfXMQidkmvUToQPe5r8ExeZA05FRCzXCPvkC+6PYgh6MXvqY4raTKcHpAnk6gt7
9xzSOohcTNpTvZTdsC4zTMCLy4ki5D0e59t69aQ7sK3ZRDkP7XPCjYFUkLDXGk4H6XXulNkeiHMZ
61dppGrYazShxrBdVQrNOaoqfTbZ1/BYkJRFix5dkDC2ui2Rqs1bOFZq55UyNQrmA0tC60gNkgv5
jBFVhG3RUKbL35PqwcGOTGfWhx3aMcLc9vXZAiGnAgSOIPVH7IBLKnQ/0FwI4jv6qYNn2zQmNzqZ
RYX58M1b00Vgx/cX2HNVuBS1c+zaeonZh1U7bBw1GrST72U/MaVsqRA9PATJoDnvmnFB+A08YCmh
rB7ym6SkLqqssK+x6YmSE2G5b52xORlpVBqKCZOFMAqLYo7XJW7vpvvdBfaLtMKbVPf1HwblwAIX
tN2IvlKUMFDxRnJeyvFI8rX63mE/Ftqfxl0bM93thM7jT2HOZGRfpjrPMn6V/P6wBQ3ht5lGpSwS
YWkqEG2S+Rh97js3vKxhc2x+YAyoX+nw9XU1FnRHO/ms4gXshNnvM3kQ15Pd82uPX8OnNDHG5Jrz
xh1P1aztITCwY1WX51DPJlwvKF9RwIexaXoEyaX2PZg7kSy9Kwpe3aUhZOQGY+bnZpZeIT47UsSU
cOgbNIHddg29lTBIUGSX9cgemklP/FtOxd9ItWPMBu/gUHzDwMvUmE/vIbBHZ2wxWPjVrBvYfzX8
0B/634SIGcfTQu78EroaQKyxDJ6IO3429bAhyIYxqahwfDkXCL9XUsNnzr4bnkE9QXdcwDYo5tip
uA3Y6HkiDupM+DasLR6eTROmRPz1OcUyi0XhHUaFlxQGAhC/T4YiuSPUSjX9c3OeHvuJ+OuzfTPK
m/UidsHnfh9iCL59M+N7dTePTknbSFRCGYeqwr5QvnU3OYqrTn8qDW8+dJKXuTAJTtUA0cn6sZ5S
U0LgmOcG282dY4vj+jPqu41WO7OJMlEQgmr06wAko3Un91azZchBguMb9zypI4rkCfOBvaISjomR
W+mTdEgCEf1/MSGEEcMWzvCXqPSkZTUzhsSHT/hQadCeoiX0TLmPgk/4OjRrtl4R5gMeXT+StJ9Y
dxgx/KqnNJghhPzUJnDYHYeBVhjLw/KwaJXUqly3fJK3Ulg/4qsQf721Enr0KCn4S0P90jdcUBmD
gFcRSiEmPp0yn1CFXQQHELY16z/UA81K5zZ2D9FKs2O00SuQzjefeHKW2k3tOZaU2KX6iGaPBLLw
SLvwTJ+so5O2Ahe6nx5JZd7nZ8eGD8hUsi6hu04L1TyC/VPLRjJ4oB3PP38K42zHOExlMBg+twdR
jV8hFEdBb+uHvvUuCjdY3NIh0a7TEEwA1tM9Ile9iyfsZbW/HR3uEKzeWWhUUybvNj+tiPK9RGiP
VDlG75U/soQ1OKR8tYsnoSpkbcvYTouQA6dVIc7EygEN0Gbys7bShONCAt5TnZ0nOBq/xeAD18x/
uzm619ToOf1QaygTAgoZWWEWI21VUEm28s7LxUuuKet5AvBfMGZjzCAwVbLZrJEQ7FCy8iPIpxq9
iU+JvGBT8swpwaOghCdRRNw5JQZZnnWctTIza0LV6KFu0Is9owBX5aA35p+tez9uVroIXgd+fVOj
puPAGOBKJdXYqOU2Yx9hA/poA/nJgcvsCWaKvzNz9FcjcQjKshy4yMD8K8lwUTqu9adSgMN2CPnk
7ugxhjHfjyEF85Ai3V6SctRodsRIMq7urLlqJGXDBDnogER8kLXRbkBkTSzHFxfGp/LImQJiPHjs
bo5cjRDDYb70UdVswzfB31Pj5NC35iYRq6c/DRg1ItxB5a6zgf/zusOttV30zr9YTskzyGCmvZ8Y
LnR2poldcqgvzoVF7V4BKq9olyvin8dUizxzgpSVFvjAqLXurXNvsgve4thNniAjYbnq/zIIW9lw
10MKE9ZgEQPMyIZdGw/0s/LcTssLLa1IF1wTSWj4FJDE5K27fWXh9B6fyRe0CUpIDcIY8AFkkFcO
PAq5EZn6xxyiwjSz2goN+553WvixJdFRLbnGHQcCb0Rin043dsB4RFsYDtRVUCKOC0/ifunpntYV
JgbKgIdXPc1sISdH2ngvRzh29GPFJA7a7gSF6BwV7xB+Ux/SBz9NJR+DDJrIpujEBGkGJ2MJZhZV
8amxAMIWrKiUVICNvRTTNv3cg07UimcASoWhusGIsFNJZrKORSB9fmd3x/UCLvla6WOG8TLavJMT
l1Frkhm7cClAdsLGQ+qv5AWPqOx1EXMFfuU3WINAUbILlBUN5v+YbkkbD9FdQjqAouqbvfLnijku
lJtUsHsmsnXdrgCBHmLC0yg+lDyiULh2MWC+GGvXD7p1Zb3LjYVHeeljHFFeU1FQqeD97+EqddlG
823VymiuArM3DuJHgG0XHcAav3AG+4vFv3Ve8NFaZqVZGYFjqCEwZV7zNE4beViQ08HBs5QZa7FH
qSRzXcb9JTDq47ZAplqbRCb8Qfq8qAN8W3fncTex6RW3Nwj3gg2ZswVbdTt5vOOB5djKjQFCm/Bz
Nh7/DJrbmTJyKfphfdEf4LkPSog/wcyZRHlleaPUtfkuIj2BuEFVWiCZJgv+Yk727GxU18pINUJ8
7KdfZH24aHv4QN1N+I4M0dAjNAp6/ipOH8nqxKternz+kHurxwLHBBjLA66H04o8YZ0SMbOyzGln
c/qIi6de6k+wMH6BHMBT4tbvXNtzpPSIsJUvP+pcoteV5LmWEaQVdPLDrMD1N5LmRr0Ch0I28ao3
wB96OR7MTvp5fuARMSAtj3D2Cita+EG8BY+GqwvlDh8Xf3PzSpPyavSdKwnIQcSOq7y8cVyfoYZX
SzKI6gyCMocqJ69FnHPIXOhMKpyuSKTvMGlrhOyRGzBML3ueOUOwqv+sGXENCX8Lfa6z93BNtjDe
skSdAt+jiju9eXG2HOmOva2VlkRKikC3KeaqyX8O34JFtP57idsmaKsGCbqgiYKyBahmWpd6Ekk3
evUNG2GLf5DRZozxoNHE+kDk76DmUDr/q4cGfi6T/Bc53CunUBqE35Yfs6jX+7TZz++kKFjM9Bm9
omqWYdlqWZ+Z1IEkUJPrIZirgcoAVh8zIK+JEYtww27JOKGMjTgybR6337nqqoN3o+7efIx501h9
G8sz4q5lZCm5DW82WZafmWnPodvtUdyX9C4BgFXDAIwJCehBNIraTbAyTH7RUSznIAINymNMbrXW
owhPzHRLUWSWGkFxBwlQVhQLzDqmrQUBtmc8GTiWoLKuP/SGlMvhD41tn+Q+BXdHjfef0GXcOeOK
FDR00OHwciRhVGPtFljpG0CKICB01a4tuVyPFReSKrnGspRlU32CahQJ3qkohnBH1i7o2Vq/VKVZ
tE4H2Z1IVMUlLXlJAlIt8CHrq1blXeDKBqgIL0TkD1wAaIIgqwInf83DvFLRrGnl82OXbCxXfaRv
bIEs9PFI8APN0hEdOlsF5VJt+7iwt0l6eu7pzF1n/3Nu6RDjIDhJEAgJUnHck7RX6b8ICLUg8s34
yyh/2rBtiurFUOjmsxcLqsSa81GeEEMPHtJDGewLGWDTTCJYoR0gKRQB57B7eRSRJ2/EbUkVoxLL
bkx7ocy3h9xzSMHIdZLf08JintJZUsF9KK3ulpeUgfAnN9uv7lMa22b7s6y3+Mle8L7U2fFOCokM
JchHpAcD/sUuUpzgCnPHbEJr3vy/ysuCNsuK24FEfkOtzamt47GbUtt1/ei9w20AmEUmNhT3Kuwy
LOtrRy2g+95rMcOHfo4hJyXxgt24LcU4n95sCc5dNMa7XwFmhe9FTHClSUIMEXx+FiDufhn/6VmX
yVNUPcl5KK61lRIHhcQ+BO0e3etPKOMV87mXo2XDunUJ8DQoSZDAkNEx5XiadvGGZ5KCEZPUpOs7
OAwB6Io4jCtIvdQvy+ur9efJjVXHEhM6Xc4LmZva8kbfarBzE30h2scHX3RlwDaDkMd+UR1kvYnC
bxbidt/DlAn0DcgIQSw7i/yOPJc46zbAV6A4qA/lxiCupabEr5UTWB/hm+wMxr0ratCFyQsQJ3SJ
zt+5MeUMrSGlfu+1rJA69iMKSO5UrMgs9TKBZ+w06Nt4txgZ58yfSn36i+G7lrWx3bM1ggVpy5Bq
/ysa2G8GpJYQJMNS+SYucYXQ6YFaE2xF9OiE0x/kgwccx9FXEI1GvKN9JNa9s373nn5ExSJLukbi
TmT8hXICupNoz7oj8HdT8RS8UVuBuDdUmm4qRvrKNAMTTAknmMp6yNRtjC8u+jn+739tpZqQ7avt
L+QKChLF+qF2sYNB4wu0WSEvWWNlCm9/lYA3qTxNKlYuLNZKaWdsHryzPZE/j53dbz5kvHisD7c8
TOtazUnD/lYGO2PHKnIQwwNnJWqXn7lvYHI9/3XeCMxJDplIEgaOHR9G+fyBaJG5tRyrTSn0AquX
qi+9GArZJy6uu0x0w6vRE1zUxwKH8ORq+u5vEpB8emLqQB6yDATdw0QVMFfy+cv63Mdkf/jWxpTA
kBtxoQv/Np4rQ8P+nV/MF8wonnecjnc3tIg00cq7ygL6Qwo+046+Ja774QWDB/Ccpk8IpmoQ8/G2
n8qJ4B+mh3zgpEF096jO7OLLrnSGigxo+SrdO0GdywAMmxkrt779Xu8bd3w0Qx4ZLaU89JEQIyAz
ZPnBKGPgve18/KU2GCaKzHFhz332wVD/Vie0lJalNV8Kau9DFLQd9sKgnoN2H+A4buTNgZ49ejl3
J0b9iIyKLXY/0FROe+/fLhtVmM1cjpGVRuB+lduYZCbLvq9X9ylJIaqavp0Eva79pzAZRpXWEWje
XAQY31joliQVYa6d45cvbYcz32C1lkKrzUS5bf5oxKPvVod3+4mATymvBDieXGguLcGHBB8NSou3
VYSoYvEP20pYr/gOHN+075oPH1by1rGfGe7K50w4zT4iTCx1AeW6wp7sR+4d2NjBoNAAS12GK+Zi
EPUOXLPgQH4pwHiWfFOPVuokzcK/7V+WMLAMGKNOGlmF1pDBoSc4A5Y6OXSCokJ8cN2KRJvZDZy6
CPx9V7L+sb+is9FhRuVFqxfkWgzF1/Rno3O/nH4msLYZZV+QFWuVlivwW+FyV5JL4MRFQO+5oRa/
1fPS1WBqbi30XP1tVyAa91dgJ2Zb/+M9QMt90mGRgyNNcelaijTQz9aJJ4qElH/s7bDFRFfcRhLp
kkRFPGhsEB6eLBCcdC+cEj1mtXTjQ6flsLCO6s4OFIEoaVuqVmUFEiv8SanEcDqtr4gTMvQWp+1V
ZgyuiYKs2SoL8fyTg5NbkacnZxcYcji+cokFFNBL1b3U9Jg8gBPLIgwpO+gyk68GjCNOllyWRRPM
Kinqchco5cxuyHX6rgRPuqtysJpUdWWGClw43M9xOpaTrQvx+/QKk/MXCPD6zsTXgYeHdpc7zjjM
im0iGi0v95LxRU+1xHU4vLxdwzCoCnSS0hmNuls8jzyf88hRnW7RdvLiZF3H9ppQhVfj6oNYODHY
3lEnWQyfrWi6om8jfTufoNxHpWU6sBIRtDX8o7Kg7ZCrRXo0VGlo2c4Sqj3WvLEz8isCCuzDLbsH
S2HJfqvvz1qROcHBOrwGp9UhrufSU3/0oiYhxeiOGyIIMrZ5fFNxLbh+a7F5ZCNQ8gQVCrwHQrlz
R5DAE+dd6YnZF9Mg4yaFwaqaDFF+Vs+CD+dPl6OiAW3E1A9j8CGodejG8YQpObFSyww7hnVA6vve
wv6QU/hAGoRiPFh94682pcqeNACPhFS4TuMNPDzEwB2x7UVG1Ff4E8UKx/XdmaA+uHEC+m171+J2
qvS0eriU3khygApgIQYAVxkPvjYHRgCkRGN++ccSeOwXrnaeHd8ltPcCC1Yu0PiWNCY9JuwpEpi4
js0dVaDxjBZnbL1uCmfpPZW5V1m6TA7+UqNInjJa567GTX86fPtO9kIO0f0THZOjK3TkTHp7Sa7g
72H1o24lXOUTPDqo2NFsIXAAdSphUBPuX0hsVsTxsTmhcIPTS+8HH4ilhwKzKySHvVcNQVfVaCDc
IRVtyXmEs3LektunFye4kEC0/G1ONENjodZwfqmR7ka445MabxZliA6Iho7scWts6ZZ5wveyWcNZ
aU7k3p5WbCnEooa606n08CQVsrBewadt/o6KDzr5dASLEoz5+rcPELfAdZotxkSLtwkQU/PFy3vA
1VtLpbL0cRHmy9CKti7JXJqchfbPbn1dW6u0Ih3+JOWaTOm/6n+TtRZbrsDac4jehfcWRQPxdEpS
aEQWLos9Q+1gUrmB3TbZ0t66LgN27Yav8IGcBHhnbUZBdyIsZOgxGHhbF//wfk0qYB6V/GDbc+Ac
9V3jGDLuiwsyraly0eI+exjWMwaWgDVmUw7oqdpB8CjYqfBCnQgB7+fqDQ+Xho4nZuHPlqcCHEV3
sEeiNtgptwZH4OWWezR8U7fOLinaUh7r+tBe2F6gTtRg0JPDhcye1jwh+XOx/0SQTOSkQICYCBWA
7fx65TGKjYoH3xXBkSoupyX/9/9vBU2+5IF/zctBThArCr+Gx1EtFVjCJxMnw7AZppdsFFpCRk2G
u+2h7Ivs2XyGTafeyJQx/FY5yiewCqKKWE2j26UMFnxnDR3wO3eC4MjKE3TxYrgtYKhgVVydbNNB
OSSkRB0MUyp8lu88wOObMmdHfnTss5WY73ZM77qLh4NrVIzNjZV4y6aXUZJ9m67Vulh/LwV55QtF
5EXDX1TGC8gfYkWfOlDJmlsmTL/E1GIWheauwZAkRPKx6T0O3+WKXxqnjqiSM8Q6WBmv1viLAyzH
g4UjvPoo1+8C9oR+N3ElCxrvwRJp6nHVouvXmOtNfOorZ78/F3uK7F6yxVsGrdNOTFgDZBgvznwh
cRalYdLjqxzttdG0KKgqPb6JNKlnntJS9ggKEYKRz8X4JppZ0GFIMGq79yjknsmAYxrKdJAcJlUv
NGCnjTIPnhNIKT32/UJ10pxcfHIr3iJ/g/I3vE/nDBO+ozYpdSjpqemCydJHjqWmEs9LBziVXJMF
etxLQyfBeVdx3xIEo4H7vYpv4iIlV0bQtA/DTY+D0Ky7cWeyMLk+KbFYxdYQLjZfNFWzgbfebDJg
8StYuUMn58AQeUPPqUrpbdmf3i1pEZ199vmnrENqLx5Psx3dPOqD9d2NC3xutapMH+B7B1nNcE4a
O6IQF5ZEE5sve9ACNI7FypadWfuyjN+EAIXufz6wMbDHlPZ6WQmQYNwdzEA6UNd/25keaIVYQtKD
pVl8UxivwHUTyT5utKiCXuDTrLibr9IUqbIuYthdWxPMyrmdmAjz570XMApag7iRfUkbYQfpNAQy
YPPYEidtV4/0D5z+smKZ8tWI7G0PqlQ+G+xNiH0ljOg4tFu/+pUqUV/o8kmLCbgwYfzJSkiwHj7a
F9BttseFhsQ2MpuY71dP99BmBhaOi67eJwsDY1qKFUDY3mkOZXeFs7b3Efc0p1swWPL9M10NLc9D
mJXet83Yzz3QywZYMoxxEvXmYgxd3mrUrd/cekpQQv0Y3DFuXokmz1Dx5gkUD0yLp6RdfPoLE2ks
lDZ5OGDBGaAIBZno7mGtOCxOgTOJePByRhLOn+8V3ar8ORRFt2Th2t3GTRx5omlF9mRSZNXugdeh
+KUvq6Dhj+tolchS/x7vDncSfqb5l/xhcevpb28NJZd5TKpbpJmZulZ8XJjpUlNjYSHMavydHAmH
W93N0HQf/V1NEzZDCoUX2Bex8dCvIv83CajjZ+fnfwA3OW0WRtYpLdKS7+X/3HnCRsOr9Qkkr5Qp
EmaLqmRrZj5dhZBZT3suKaX2Hjf+D9dHpvmpgsd6/lCOLBiVl/kks6lMWY3JfFK/DiaKcE0CyZDr
FLBaGeOjsIpDmCiPc9tlJaTr9gZbetWf1P9yvDBPi5310/frr1X40/bM0i8QmkmRb3OlO/arlCdS
q+1AG0B7LAmm6eU9eElqUFHACDpYsPo3jHFYdftrbTlEdA5ln374BPnJ6drjprz6U0TLBzoT27/v
zDrK1qjRHNsE93roWCCsr3VV01Jl/cP+3ddzQ5Q344pJR3VTiOJWWvmvjUY3uUfN9PRESDD0sUt1
pmHAjZpWHpbPfpDkWyrj48J7oztPaqCdjzwDtxAEmG0RjjHVrE1ZHPiGbLx9qUDiLyWvDUxy2oUj
RAvCu1ro/5+NM0SW84cZV4sNwYg53b8IV0+m9hYemDS9rxK0Titcgt+dTqeXPlpaNPXG70J7gVhv
nqOFNlTbFxFFCBcAOm5cs+hSzaYGEIOuCyfU1pIRrvb07xEPD4NRILgeoOnuz5rah6aVEtDgQsQ7
W944F84RJ8FEz92lMDZtuZ9s4xTwqf7q4qVrNHh2GzB8IH1UbybyROAkbr1CkP0iUshkjxXDqqmS
cbr6KgVc08ioFkCZ2orVsIKXP4IU8Pi2pJsfU06v0b4sNt503Z9MEAG4WePgn31JNtuFzt9nV2PR
wZfsIW69UnCdZPEu4b4bWKYG7e7VFbyJ3BMRzITemPV64Dk8EGs3JuLlTbmWrjTdYKjskbVc4EgF
N908tgWirf+comdg+V5Rk3JpELrhiAnWHM6pM+UBrxHUtnvo1EmcAwBQBOOTFFxFMCjTG1oQLWdW
zM+I6DFPCAvs9zTq2QTBczHrTZZofI7H8ng5gviJI1BGyj6iaVXnVpY6hVRPx8mD3M45bEw1fLHM
I2S5eJ9484x38QPfkBDR6tyXJLne18LGReLlKFw+bJ5KKMgrtIAKuM+KQ/yogqow1tcepvH5YAhb
S6ECkpv2zA4bSFYAy/fkxuvbSGxeWj97KDoI6iI8WrudastfejfqmpEKEHEDvhJOpYTMfmVzhlso
rhy9DIyYgpLnpYBkZ0R2dnVPZQvS1JM8GvTeHB9YzrqrFyHNPXu71MhcLPl4fFfWAMX4abr7AeBs
QonpdaZ4zjbukITfdE7EVCpmCL/61m90qM547+9LOVImtu0eUUE+7kqUYCadxiQgZm1w47Pq78Dy
o1xWqf8g10K4FU/scDuRua8R6mBAM2qMAwgjVFJbbj6vkwGqoN8XmNfvTDcDqR93IuBKfjg18xiX
VWUOd1NiWj0DsxGCuwUAlsJRLSbSYMrJ0EqT2keJhsZxeXW6WUShb+6ufmKdV9QZpssP7OztB9PO
ZV60BHoWzyJsFB0QlHTtpkFGviPHqOw1DkPeGWkIk+zrmg7pZ/OuLpVTr/n68Qj0MB2DtLGD2nSR
FG4XhcVDBYseBnAAjUr8J0GMKx1hpz+gZWuwyD8s/36GD3p/ACzZQPyMQ/sYfI9LZrndg4qnAHdL
XIGk8QT0O0tHWV9+he+2XURYU8l2+Dx1DsE6CKYfsRyzrBqbpt/dmS/L9Gg9wsLscb+Tljgsu+eX
1E9u9+MujQ+JY1jS+AW4aK0mAGVzA5pmUQvTv9DAUVkvVJrLSGYLwi53YcJ3imZz9QY2foH8CjXM
521RQH1GwWW1aJWSyU1dCQFcPMD9feWrpbLGQXQV+m3ioTG3QL3q2fS5sEMnNI0z3HJrDLN/L/lP
aUUvV4Ay2q4Mn8JlNbyNsIxBethPXIDvlOMhT8ZCvK3qk6nVVPAW6+Hnfzo0TSA9KCA9eJsQhMEI
uPS9YJR1SSTKoOHnAlsCqfhH9YlN/tPB6oUUU3IIGZFzB7avZqKYjvIBsOdezs4rA5dtflcJn7c/
5dKpM+pvumk4Wzs3OpNBjWo8OY2ty1Xy1ffBxrHt20A0ExKTP4NZTrgQK8oahucK0urUXnqGamnH
rZB2iBeoJPfyzePqKYliSRmG8hioP1iiG9zBYKepGj6jRxAAcj3OoFUHRQa4+0XDKCQ0Q3jZRfyZ
UODGroKVl+HNzgFO9vfa0wRD2Dc6QinDZ+/TQNRufSZMPZb6i/lRFUsn/k68Op9bM2kAjrpy7Tkn
Afg05PyzyFy9d+pGEyPQSX/mqnU/sffYybEL6Xh9kEZwXM2jeEvMcrC9tbNZ7ndD7wTVHzX2dZpe
YWRBLtvukD3MJHaYzDZgJ47hhI+hNUaQPbE1wSc3O6t2RAfL6Z+CfYy8POOvSiBx+ZgAayd6C7Ub
EL0mr0OxAbtoYT9s/+uez5qdUIS2ZVOr/D6V18ZApb3DItS0O4OL4XM9C76MY11PGsZWsmnQJ6E2
Nw2i7Io7QTFOpssfTQra+cWFH6RqD6WIDr8MMf8gBhxQ1IjxZSful50QIHiaLPk3z1aIriRXr9S9
4J9blHej+otH/Smoh8MBMBSJglwG46ih+eFovkAvoDAxQYaneChVOf9L1p/QGW8Z1GTCa5e8CisV
nnGgSXMMtN2EwtzPWtqaT1SfnE5CJMXCKQYJ1Ro2v5wjQaVEq9VW5fhHvZNQpxLyhsw7oizw61aA
zdAo2Fk19KFVhycWzzHGeTE5MynTKfdn+0HBtGbgts6DNGSDNlzuORkidmszYFi+Dy7EAOW51y+f
FZrkWa6LheBZHDtsrzI3GLFB4uqC4ezgq6tsHiLOUNCUlFqC8DMqFGKoXiuQIhZC0bWNwyfz9B3n
4/e7HWUUXW+wP80hQ+0JquAFH80DFD+v4mUTUe20mg4//OGsfj7BxG0GMcjyEX18og/1WAbb4ALr
cYWoSlzxZOIxYp/aOjp3FWlF47S7/ows7IftEIlF6ijXMzvkI8uhDyxVekwuOb5NddDh1XQeztLx
iF6qJOxL+6R04i+Vg5GhrbChGusuS8TjVSwha0vVrkh7b7siZITfSEjmna4a8+5pUHcYw9ZWu4J4
I9+bQY+STGd+gBZVK5cUME+8+M1MZUPofPJUZCHk9ZELJXqqKGcrssEl3vw06seuUqXpLQDB1fOo
AmauGpBerlLBQeESDYHAVgosdck/jBZ6goaL/iZNIIRWzlbRHFn/xtxBRgpuXgFvRoVFoRsU5jya
egpXxlcFll9RN5lQtJunXsVi7DVQS1HqJPNzDFXtmL8kZLvrtwXXXlj6mq+DcVIjfU0lPGHe6RLb
iFU0AFLhZ5r3amt20RcgtO1Oa8sdjw87WNBSXMRUDvJ6ngS3slvLqnc8v/nBxvRjl/2N4FQ0oJpX
/tmOVAkSYDRLUVcHL9WLhrJVke9qAPVTuk6rJKz8+aE7ihohkdTawTnxBfMs91T/E8kOM4kXvGmd
abavehzuvE9L0jnuEtHJ6hPAFv7onSmUy7xHrsJvZkZOTTokNCMK3aAM/+aEIyFvrKvghd24t8gD
LNt9+vNDx5HlJ7ej0BMF8A3n5wbeIh+vJtdRb7tkJ3pmoxFRczqtvjcMIDk6DsU4qCQBEK/O7p+T
OwSfB3273OeUhm+FmqHyIsIoAB8YWac/zMIVBbUSeIy+3gAhEILmKCw78eyF9uHvaoM4oZqnjwJ+
4SAR+5/Jg+asV4nsDvyNiFHAUYUwI3iFsj1QFjahoViRwTNo7p/wTMQdiuX9/Jnhk6lP4/LTdjGW
I3SUs9pbdFXfbwTZBSh5b8CSBD1X/wwGMQQFxfnDf+pMngmx10EzSP65ViOJBuwtY7WE+3/w+0si
NZHpfsmVYuH0s36059tXC/9vLJXJJiJdqrjo41j28QAcGTtCQVUQdIBcieZohPfOEhZBjRYAF5kT
4bIxG8WsbiJdR60Ni+fkeiiiGCJhNS7JcXVN5dQh3yM47PgEGGrI8OOYvQWO+GRtGcPowB5Qtk0Z
p1pp/SYy1TRxlOMVnkc7y96clcOiIrcPfS51DdNObguLjaiQoQsDIJ4OJFY03TCBxqnDQv/4E+Ga
X5h0zGbVYqHMnbkQxf9mO/kf0DDTa7cJM16t1R/DWx7QOO6j3SoBc6c+/jFOrJiP7nSkngKesYQj
xb3VERmDtEB9i3o2pVgrD80yp7mdb9z38DjEW087xxll0lW2UqZykP8FhGvoPITvXDMXYjEFDyfu
S2s1cY1cIkzAxuAuP0VkyImBBDIgeY26EHfqRpqZFSJrvIPXT1T8PNJke40kFX2AUzGO4p41jEKt
ZNjSGXRmasigh8pSYpEfFSRA1qHeDAwhdZjMRRwmo6iXeJ3NDwYW2OKAtoDCQCvcJUTJxCYPvlY2
RRbg508iormazHnA1+GnSIu8fnmv4KxDkjPIJbaFEBW2CIsDWspzHYUEBj/pY0Fe2crUDbWj/Smm
4mFKilSzcgu600Izbbs8xmxgaY/bIQsZysqWkZQVqbsUI4C0lITnb9bfq9jZ5BdiwGPWGYD1yk1a
OS2DW3e2Z/TPM4BBqjlMj8K8L5HsbmOH2zrxrfd7BB7rEeGmZXvmfsbIweB869FKTzM/HZqZdGLP
jaYo34HPsomJpK/BoQ7K5iztCnLzzEsg7I1FqogQ0VmAqZ2NMogFGEe9Jw0PVM8XlbZUqRcTKiGo
FU+0f4SO5A3v2WYd7UxF4yN0VPQXH+TfAun4tpHt/w/dbFyIkItEBUaOVIr7uq6d1X3X+rr15YF+
6sjTabnOGH/FFKL91PGO4QkEpjBleM8f7upRzRYXKs5wnCp012K9iilIdiaXg5qJpNw86rv+btbp
Drpm2BaUew/S9se7mlcdyUWWiN+fMXM1MBfWzgv6C9dm6B1kzHX6BJbbV9eaDTf+tXoAENuzF9/T
hQs1xRoRf01/w1EILWgKtO1g7teEQAVhiR/jaRyjMJSTePdi6t2Ea3wdYWSd+tijkOvjow7/pNlD
PcPAG8WlhzJ4CD1lwQ4QrDBDSzr4JRvF0BxMxemJr+T1BhLnvx35Uzhnsxa+tLQ9U4qDCLBbtkaX
9rDwfJuL+CA1qmpdrj8+Ltm1TPL+PjHpQmQgJe22IToYF2T5zj6R63xEbwKSmn9FoWE/iQvmJHdM
cc2z4sQDxyrMe7hrcya10mh4rZxouQS5bpcbOaioN3bV55br9Q7iyn21dGVv0u9BcR5VM9azWomv
93QcCI+HVq7xKJxxzPoZdU2zSqaA9UTZyDSrHutvXHP5+QWbJF+pJCJ3u3i/QItelRzSzYyKP0Qv
dyrRQiJDIXYopCmY8yncx5rE7IiuOmpAepQQPvY92+R9fv/EyRyjN/UaH7teDs1okRmw61H2+JBZ
7bldYJZfAl7xORaRKPtRttlzkLiDd+smy5v4jbqnUoarL1P+HndC3exvOAe591YmwR+zorzl7YgA
oAok0ek0oHeS6udKU0zCQPc4k23RROyQcH47cbDBUUblDfGgKmNGaCp6L0zbuz364//u4Jj3GU1h
KUeTQx3OiV02MqPH/FESkhwWKQTigMKcUvjZ8Cqcsl+7TR7gUV9ly4g4EoNP1Oalk40MjQRqRsDd
WjucG8/uM+LJ2ZKFHjj//+FnZh0SVswihNoq0uvHJRZeojMs0TfXX24y5FJ+fMf3cK8FuOHPMwTu
f5gsDzXwlxIt1J08yLdLdhPZ6iRtOteUslhANLJfQ+lPqJXwKdbUU4Apqq11WyuMCrHGFsczhUke
QCgw4lAiAOY/YwOr/7FOuh6Gv5rKrhSDI4cXjlCLJ6+KN1kKnNR7kfTq0rOa6h8DawL7R0H+ECc0
ZYfYFpFsF+Jc3hrBYqPFAbMVNJvnLkpJqXApf0SS3mC1CJJ5hMD0t2MiBYme4x9/ZrErJCQAeC63
PINPUPgZskx5um3IIkfGwgN1ibDrjCYU+p3fMXX6v2qVB5djdw01VY/P1XxRAT/E+S7k16aO5+cn
lj/sixqyFsOABANGDKKFksKQW5d6Ra+6CLKIGDUlLeoHyIOx7Nv12KcOds/9O3N4JClJjG7Fsd5x
eJnhrGIaxAFgJ8eKA4A79ECczpI5FZrwt8CM5pQTZ7OM4sD7x8MskTChe8iD/AVRqTwE/e/KvO6K
fPj+SQRB5V0pCPV+KJKUv/Wa7lpovcxAXnxvnySaOgIbDsMIpWSF5DTm+YqRpofe6DTYx+JubjuC
xxrK+4CF0NNXQmX820z6rGv9+h7d4tm1xbye5iEcMwM6RHxu9m7zJTn3PvLJydDDl62HlbJI58hj
1kzyMJQqaoepR2YTmvc7h2mF0kJ0uCW5KSqa2l76ZLh3Az7JNy1oWz2xcZy3iHjhNc+zgsAIEKA0
9cBSCwPF2DjOs9h9C+ZSHXPdoBfx4j/WSHZVUUk57+Qv7fdl4HtNrbSj0AeV4OxlXUh0wa/y5DJW
wG9mXIAb/UOoDXW8GZUT+sXAi/1LL8apfcA1xjxgCGlt3+KqKsQq8XPQVo3O5f4gmzZnOS1di4Vk
d4iM0fRJoicT5iBqZ+cfuYOl5H7x4/UQw9JBdUqtghjf6QaoDbXFMR2nbL5vgOx8wa5bCT0dhFAQ
Y8uTWbiZyQHop0HyMnizmhzw6Lnqq+v1Szabv4sHN6HGUyiV8UpMdbG7YqlzmAePbI1SYJ2UxCtz
e5frUUGmDMxKVSlMiJVi53rHuOglY2bpx+/llq/h3p8ecB3/sUHIl2NaJuT2ncKEKR4WiqzOogVg
neQ/9j71WL95yDnoVdT3OVc/8NjYTJJI5Y5cQ3xwUeIsPs8JhR9UejeseYhns6Kn2LPA28XrQU6Q
XbhJVfznYtriQOljn5BSiyJjXbBPuQOTnYW9WWe7RD1v0ZCJmHHo+HE9tNfcKP6se3vgGO6Q6ZAn
Sm6jIjXNlRBZjPEUsaB53SvU/LZVsPLg3Xe8LX9pstF5eLe0P8jPoZTDN7VTFEiplkY7q2RXtpDA
T5jMOvR350Bn/ER2bbz9RImJFx9Ct8pvzMvgzGymMIyVey+r4niSelN5U/d/+k7RVxDhupEaeF6T
FzO85f1SGHHAnolk8AWz/Kmz8H0LWHs5eUHLO5+YiPs6GBUHgyRVYqfAe3jn6eA+CbALLVIB4vnu
Qe9ookBzTgcRfP4iTnMLes7Gli2a+I4CmYihJ8+4b4PeUM9mOSJJuNkmvAIL83bJSxn/XfggcaKQ
v8TDWvQ6iUO9QsReWsnGs+7PdtPPAYJKpfmfqnOw3XQ3d5YL7I2WoT+kSd5oYojqGzzoMUvA05Sl
rSeNSCQmGc9SkiQY0GKzLX6kD2kYVWWiRwYrJPE1MmKvnKLiwIk8243wD27Vm12juX+fRGq4SUZL
PcCky+Wse1iZzznOxonAg+QGqA4pv+XXzUB21mmHGE43Sig6pudrnnc0LJbj2c0AHMlulxYsFZmV
bUDQuDunz8qsWnyMbQrKZiP6pmzCeLtzH2JD5mObNJ0xFi95RBsjL21mxdPCYgAbfpdInxVG7dMV
HH0LgwaKz+yxMZJvQS0z9C3pyjwK8qatsBs/c/1w3Y9VBluTPuDffK+FLXmZn3hm4BOrfJH5XLdB
qnbo0Jc8INylIiLp7Jq6VRUnbBdEYMNlTD89dONimt9Av534rcgMYyvs68ccXCLqXBTE7Gd7qLJQ
kFV8hVzoPQViUN3DCFQlfDyJOI3NH/m5N0zRVu/qK7cWNhXaIRPltmDKkmoWbCasTUhk3+hzDznW
PfTwToLj3S0/IXJxYKfeeuGpkfxyr2VfDWusRYeDFwWncNpBlShdP8yC2wEUqCRuUzpXN40YxYoX
LCqwf/DkxmY21KE1/F/59Dns2uZ9U/a0a9KVgTB0IIwekwe61Zv9JxDzT+59jNz+w1KEgBDNa41b
QBLgZcftWbtHc+KbHnJpJeT5hKGmz9X9DPar8x4NkRn6tLDaZF30TACm/a4vlCVl1QhSiD6SiaSk
R6qH//SuRwD/HlUa4dvfMplqw66AFAY9yWtVZQ18KQTOUbkXW9jU5rgLpvBZ2nmZzdyDpXn+swdi
uVyt7jXIyeh8+0RrwogEjURaGHmsq/N43QxIKOwA+yGI3hqZ3+D2xv+Mlv2j+c2xTp63DI1P/1E/
7SnGm3OjzzmM7T/pKe7WF4WNXO5jifm6GS1etPWut0+poyeJdwuHxKyfVNtvLeRGrkwjOTKTNdTc
UVw11XO8ADDzF7PXf+/QqsQn8uE/H91RoI2DzNvbpYMywU6hApsrS4Hob/s5t8OiHu1qy7t5AyvU
a6BVkaLvYOqaMK8bXNTD5jZzbg5V3+ChhwBgBm5MUOH47ojn7zL7MOVKvsAlf2OmXxwC9Shgknf0
vTlEP3Uv8nE4BX8+PyxVgpcLrix4Pu8SmzQZhPkxtogfnpoMCDcfu1rrmKujwpTycMxStbEqpFHw
WQC7WQusn0X1AdrHurAxdNJ2vRYFdZb9uKeD5onUDKF05FTmW1xQPRtVYVlznG1ePlyW8Qt7LySI
1rCNkknQ0E1ZFHaAHFSw++WBQrGwW77LCjdpO1hZbVLroK1D3gYhDAolO12iIZzmri7an715vn4F
rJDs14AveVzKyFZbrnV6qMmmF83mc5oopUdr+Z5VpXzgTbpjhYpbsF0mf6Lj798jewhjAOUsSB9s
U4uxFIhHFH9ldmyUGumPYHshXCmkmYCSS8wSERP4hNpQcLqnpCtlGObxReAw0k90nj9T2I9bjEXU
oDNaOqK1Z7kfKNNx6je9HPXe0LagsDx4VaH0jQ7m8qzV7OJA9E02Xa6Gr3rHlLrGPYBdD3OcmBl+
rozHd5cGhT0+jgFW9ZFx6tWhhJOGfdlAeuN9tS/paWOk1X/khjEVdX3WOIPpvn4RdITuqeXRSlws
cwm0mEabkV8oD/k7P5HulpVRcMluvLGIe+XWKYp5Bqpu1h5BOM7WW7P9GUo5ggj3eEa5LAEw0lRy
pbnX3K43D5Na8cwNSNUYXm9YlO8/87IMAQpYSCF2EPuvuMtopfMTHnqMpyy1d/NhBf6F9PAwSGBJ
uVyfiqt0xC3eKrM6VYEw8bP+9h+PG4zsD7X+RJUpSXfbnxVIXacLosSrj9NiFYIpiU54mIPNI7EX
T8/46f24tM2CjE07SvxIZsN5ZCv1UfTIUBQbpaDlDIt05NEgSS4D81OqsVWBrltn5JI5XUHvmZ5v
o54Z7Jozjt90q1T64EUBnC4MJty96DQ7LySasv6IHLc0iZ+aL0UQqOcbXmyP9aX2gyaPWQAa2kuV
+TnM7NCDdFUYLxbKw8ZDz0fg5PRFnQf5QDvJ49vqcAJEVWrCNJUl6zW+4+vtDAuUFtFAl760bzhK
LBVljWGPnbGZraZXoY2jStyU5RADzMQ+b9l2bwgYk9EC4CsDz80Y4k5OHiF6oGAyRDLOWb6nw5Hm
c6Eqj6UiBhA0yCDQrB83Q9it8bbGT+AtLepqOunj9l70eV3GmqFtuiHb+oVOqjlXY4Vq1sc7eRZi
Dv3T9qhGzUASMkpTvG8vh59cj/rQJ/669SYsxiS3ZWngjyICYlJieN893wRD/SCPYPgleF2fWaWL
G/Cph8vT0a9x9IwyIjniyiMWLLbKjxuYezv6C3TR1H8VPyKzANeZv00wwNCkLcVeMPa85YTSU+1G
sPUypQG/WYzOjaVWm3S+LKX0nFGHRCJVQPGrrmuiQ+6lwCttQulmzZ74XWuLkrIy+h5Q9MKpWZf9
im/b08mF31kjGr2KzWshQ4EGuBL40xUecHkmEUcKhjpu+yrmYVlTzgDbRKHYcBszstDm9jAQei6E
xoWejZFqnoS56V4wcC2V94UWHQSGMjnVcs+A0U7FBe23iZSRfJoQMc4D1RanqiRSEXDzEBBjXDIQ
wEJrhI+foZgN0spEIMkT4Mu/BaQm4jbERpY8KBCGkkP/xp5AUhcGZuSuvVflRZzoqy5XHJRCM8Ct
+IpBKQYP5xlmGqCsH/FLb/FiIKQb5Q05curCI9qpOHKB47jzjG8/hK7p36gXCST+It5KCdINCVRQ
CaSYSTxOCq44pu35ndMAyDzO5+No97UBV+LsrsdAQJykVMneEP6EDu6dkKN1hxsF7few5ERIPntz
zkujhplzfz3JWw++ZfTPsnAfBwRMKxUq29LP7JaYdWN2UeXql5f4mXpUK7Cdvo4kyyixRRh6lKB9
LnnuVthXLY8cqRnKmWSJ2IXXloEyAE1xDi89nBZ1n7YUoyFeGUjRanQeFqz3KAcC0yuSYpRmfdGp
QPr4muvhoYoPuX4YJLS3j/1sJG50yCPyMKGr9/NmxNmHUlhrYyxv2jHEQ9EJ+gUbTxghB2PIecsL
vrdVALXyq5lhIlB1s8csJx729b2skzLMyG9g95cQ2tLHOCjnp8Yo3C3aevmjR+Cf2VAl/i2/RO8p
z59G/BixzN4qlncGEv6WOV3jHcrfCzVldk9j0eCQ7wPHwKLljcJBOWHnIsAhOM1qgW30ILwZL6ho
BKXaAkCcsrXecteNQRughGWhznLJv3fdz+MNKilerDCACcZEvfvAHhBjSytlSmn1bs2CuVzd7Ti7
rIfBOrm5JYWPZ6kWeeKZV6iO03IMHJ4URYOIizclSUDiUWOq333bS5H+cHt0NLH9WqgkxuhKZ9TL
pz/Mse0uat2fh8veOsv32j6mbqLVfhfGHm0ECIySRJwVW32c2w3X6UdOrrNAeIJ4Ez1WVuy3kup+
vXWZGKGjstZnytYUgG3lPcKU32nOlaC+YKqSHhr2u1iOPL9MAIkC0auwm9nkdu3/cRsCkSiSpI7e
dONYq1sLpwObmiAk2M7Lob8rBNY/Zopz6ERKRXF5LYR1mFsTmWCKoDSICCmNOHgsIk0nfytDdvOx
i3ebsCj2dB6K+3wsM71sPgNXF1X31SiJny5W37pPIf9LdgjnP2ARqYDhck+I2uaw8n1ceWkhVpPM
0pGBnv9MzCEneHB1qdUWDjLEz7J9b8eaMAT7rd90z7yMIzFNhjMnn2NFTr6IXDntNb5mguAc/jqc
6mbV+xhxl72rEbTP1IE02sSJuZNkO1dJ9aXoepmLh0f/+VHaAw17bapvQkWlyhGvBcon/96IOR3s
iGJooqH/wlKk71MXYghuPaym49jHvdBlcp9+KV3b7ru4VJTQ1DZSMBOm1eRMpOnPy+vhOJabgtjt
dJYRI6O47DU83eP2jBB18boaUa+4pT6Buf/rtAy/iSCxo7zzlEMxQd+JPYTZuAex7PlYjcBGw8uJ
oP8MDu0EdFYIXCqvsSVjn7HkmrkU5ql20rK7NLuxeaqUJSbPeqnFurjxNMhG3bDmC8j1i1Bye48+
3bWeACFWIhVIb0kWzVzyryuDZqC+ZwrfgoW/vegWrJv25nUmVFbqgarmTUo34zZrotWFIT/oC8bI
Ne/DCJKyWGzMjukzuoRZ2lpz7guL7l+83wT8QRA4o+nSZUcBzdASuQXsPGWZQX6XESVhU4S/yy02
Z/+hPmtVnun+mtKfxcySdQlBSFOMhIlk9FoiMj7G/srZyKZYjpxF32euZhypT/HsDbm4i8LawJR2
jYkm+paB8SVYu8hyEQqk8JyxLYUBQVnsniJCoWRnQ2ACTlvRBdh0znGe/NHdnmVo4bhA/qZYlyCt
VmSD66fitsfDfHH6TZ6uVD1j3jpXSe1IfTen21s8xNIEOZCnfNl5EDW4UguchFFRZ7Z3nGCDqZfx
NOSYqZVE3KRVN6uvWMR/DMiO4JoJcx/VEwuvDQ2AJd/q4ij46ZuuwLQ5SyoTqnOy3BdunsWOtoZ1
FPqjKAb2KKCLNqQqWTHIuZWsHILDCjue/svC0J8rOs8fXeuCsV4VSgVvGfs5MK70/2rPq4tQf6B7
j5/PWpz4qlBKqfcICypVw4TRaiUXcxD76A5TStH4MVOGyRFldDkcTycXOOTZqljNc/XmzV7CLNpV
yY5cj4jUe+G9EaIUI2+hwxptJZ61KJJ5U0BFyiH+LKTfXsIDoMkg2wPAkJ1cY1Y8RYSTVXRTOebM
sRJp/rIvrRXzkA6//KNmYDeUZkei/cEnDrQ7EpmQEHvCodskqTiJc2oFpVzBzq4hMWAP3L0Jam2x
S3sB8Sc7ioQYbqssIAfz3c6RoUyyUvQofI/lLCKHio2ipCYGuaTpVqxMkXojVNw5m3korZq3tF0Q
rk8RYI3CWfPTkUxLIXin6bOtyp1U6IXcg2w0QbHzHKIo775PbVVh+rmllpbMIDrAebGGIaQY2lMt
BWcQHhtnWM9oZCquztFoOpnBvqX3HfAtl+9YP/7jqnbYU0xgPRhtWYoc3tSPCp63CtlSc8JljC3O
dSfmQf3umf8T9gEE0gmRgZE0nIWwwRmLakEGmGX6HLvMsPlKLwscnKDwlERaX4GXrTGrKY15fsLx
o/VYsUIsDcVVx+L/e/VpxtNX+d+Khut0n5j/VvEz5o0kx9jynhis4c1gc2MSp8NAezRKZlfCQFZi
BenIyzaUD86ex5OEsiWWrMsMWi45bxmz9/4NG/powEKt4KiNM0fK98yXqV+zdDw1Xn6MajV3ZVEI
RHLV1IycGjJRflADcZFdKhyXJ2CtuN4QCpv56N02hLrKf6GJIWh+RNcIwzaUIZrO4QJY0kTatWuX
X7akwoQG4AdK8kIbvPoGbmSJi86DewI8UGf8xLxlFpf3zo9wPs78Wlfkk7j3GATrKiYXklNreQq9
KHEQ5LQnF2xux1ayU7b1Ba4Sil2bt+TmWsZpS1RX+P1tirVTYi2kCpahSeUcdLEhZhf/hDduDLOG
4GMqTyDtlOjFnxN3ecJdz4XvDnuwn1c/kBMcsUxSZIsLoVo/W4aPyaHlo0XXUrgZ5BSpagprwZ4E
zZq+yw100DHK56rAB9vzRIhQEkMyLKBVmjykasTR4ZzlcwhMWtmFaqtUW2ds7dv2iNoxvOA8yczV
3YehOAFZGllrwO0WLcJu1x2yj87N2NBRwlmhDE9CSx+JFkm5vQpJM92ZcRBiKphRLEmivrpqpdIl
ZNFnLcbF0PKYM6SK90fRsXTrkOjS1ofxuL3xRLu1ungHMaLmsFyEPJiAsTwc+9EwWV2TQKf8yrzs
oz9Db6UU5aPh44CIUgYMKc8CpzGwtUBz+4wJ5om3gkKzNI+6xPdOvG+6FDBMb9iwGB8FTHCOZ+83
VrKPvO5kYQKOOb2uezK0jvIw7F9whI7aHpOgR53eIiezx6jINCOAstw7ecBcKwGz3fabe/TG+fv5
R9Munl2r2cIQzqa+1qs5DqUFmO6/U4R9XkFi+UplpIsoyW4EtHVA8oWtESiMeR88JFHWFSGbaS7J
deIYA0HC8Kzhs8bziT0CA8rFKNpruexoLDNJ2kDgQ8hjhANMRi3DyuZ9fvkmmxCiJ/RIZfO0/5hd
4q7phX2A5S5N6X9Nr7s5VqPfV5h6E04yrJRo92Av1vava/rYSNflHndopolYMVMgRGjsyMVt4igv
8DvzZDVqHw7TGNGlQeV6xArBy3RQ9YQi+XzAXJBFaW7kJmtsrwxRG3xocgqahVjX0+w7rxG5LPZt
QtQgzB6XFVzVk+RsmosRXF31RCSnWfhnJD1s8JJ1uuRnpEgosapRyEU8UvrHfPLyXqlo626LUOsE
suKB/dSaEDQ37XGMEmuTUE/5LHdLEmRkA9Ai/SMxYKPnv4x4JDKv6i4mpjt4Ndn0yvl4hXFrzKqV
yesYx7atFpEjkpUWVmUebH5l99xS73H3F+pYvRtJ8bBLktZwDIgnot47zQhMJlXzNF94JC8ivKqi
6FBOK9x3dRlpR6r/tY0FQZ/DcwVoExqWxmjy/PgmNz7CdTutkrv4Om3XlPz4ObRYTdTJEuOTlXS+
FLHNck7CjeWDWnSGqQXm0MjBZ/pf6k3VHjGbrw/ZZIryMWzfbgaYu72JOGcEzzBLHhuGdGiEWTFx
8pRkx1lYeK1GWr2KaQKNhRL6njPz93IPb2ZfcFORHTfQGHcQY2R6ltZY0BWL+HcAnzmtXTZoVevA
YYG73tx1y3ikPTXxTghTR1PPeLFwJ/6DymSU7M+Rp+uEJ/yCC9uOSn3zWdNAjWL9kcIVF79+hlqU
n1DAHjdOsYLAZhOdhVya9JdcJxdLemBUxye5Ypy9xX2KcZPO+vsdFqWo03XzS999WUTPFkzzVRMF
4Aib2epDial/bwd94DtK6vljclp5v55cgSVuYGDgLwUlYQaIdGNijqhApYazcvF9r8S5xGvslsXl
qGd1qNKMU0eJd4VdNRvpnAIsgB+ucfYCtu5dOtrDApz3LY8h1uXFkVbObs/gHIn4jhnV2CoIzO+S
uuv1uybuyG8NgPTdqCCHm6yJfbp4hUSIyFSo4Ot57Lz5Otl5zSsseSKx3dCPG50nNqaKI4i2f1m0
IDu80TpXURUUp1UeXs82QRjaaBV8cE0/4KA2YWbXHCX8nKjjVZE6OkxWUqqg3hBzIksxII1AGLH1
UfllGiL/7huASyUcvUAt66GQQGLyzV34jwfNBE0V/ipI1Ls/LtdWHwOUjqVKfu3DWAQmVhWZqi14
tJEWGXnmqQ/iWFEaUo7OraQpWgA5wugPnxxbDcrIJUTorGXACjeYbr6jg8VwgOC4gJBvQbZYsg1P
JXWJtT/svLvXbdRufWKxRF3QJNIkvO10v2Hp2vK5KAXIwXEgb2C8lUTMn6JtqV5V+s5QrnhyXrJj
WMuJt+8cpV1aYmzOF+ZHQqX2Jp07zjT660t/4WoRAmfv+gUrppzlpDoOSRktfdHGHc55GdCFK4nY
fVUG6kTZtrbV3lfIE6fUxwdoA2HGJaiExVFjs568it6avaaTVHsdnmMIZ6pNnxwfOn+buUJeEqTZ
pUCIJtuObW+3TB15H93Gljr4z6GmmPsb9VIRqxeGVyeN6AHHs+q1YrtExb/VEpG2PL+tsnpDQDvY
Nu5QWVsoc4ijFFJotv7EdXNTSPCCJ2kg5LtgHAGkieX/HUPANZd4Nw+YfnhzdoWcrRu0ANzCyEaM
eVhC4j+el2KeA6/1itTf/i/GnNsyk+fMFZYOEZkdAW2Cj9nZLB+Ujhx1nuuCBTZOHI073Bd8IZ1L
v0g11dFJulF/7nOISZTK2MEAszBNm/+IbHrqfNUlrPmGj56JWIKT/9hPpD7BnDJ2NrKkxTK2I7bq
wnU3ZsRM/G0JBd3CgJZYFomDbq1EN/RRGHDqiUAF+d7RAcW4vTCr0HfF8K3NPIdGIBHJdol/ChLg
vwWzTXA3ifMsuMXLwUeUWfnBmzs3w0Ips1KouT6caFxTaOxcKd9cnMV7NdvDKQQKVwDAiculjGJV
+K7LQ9zH7Mvoi5Fu0xxEmghNO0Q7se9EuIytlm8kOlVCat3+XUvoQMIg/GPNTaAIoezXZXYGMPzy
ym9u+Ws+yNHu+nW+OSBPY/ZirDUNaiP4GtGnH7vpAxf5IrBAhomtWXVGlycfU6pSdxcQ7fYt7Kux
c+vs0eyudSDR3kaBO1/lOSJTi+tb3WZeNaunfGRfwcfW7K+Z9ypwFKJFooEly8NfyzS4YthI+OWL
MEvljeWUO57PckazZXL2ykGrqWKOPw3ih8EMSXLYBfOqLL3U9EAOg4PcEBQQ9YZFJc/0HNh5D++6
JMxvaDXT50TgSpVxRMRsEaauD7IH5RizYDNAwOVPN5xKmn7Cl1L7HAH/gbvj4bYMp7goK+iYl8j7
uxTlSWPR2WC5i39eTUGo9vIN30RRDZSbfh86eBeiUMJVTlEaQWg3g7iO88W26RTuftYC3KpDF146
17qEf2aA2dVcQlv8QeDli6hiElh1OlU3Ao2icCB0zivC00bUZdWJaQZusIL+Q9Bz1Ht8LX+CI9lL
tiHQ8yt1MgaZ55QQjlcCvLMfnoIIcDEqAegrNNrdgaCB1Ea2+1zY/EQcEy2unEq+nYWoF14EtI8l
inHgLZDFkxM1gbLOQN5NFfT8h0CvGw9YimMqa1x9yZonWGJvMBlZOFkkRFLBLXJztSFv7t3n6Z3S
NXYWJw46ytoRt/g12/l0EUyAq8Um9GH2voL/HWOvhtGlzf6Pms8uT1T5yQWWoe/oSkzFoh+OOnuD
cHxnzmkyBs86+h09m69ZAICkhXj6P482VmEIatEsuRZHU4N+AsFmKNzTWrJfa0jXMulqIAGeYHZL
kxPorLu75/HuGM7sqPUCmB1Yfus36WpAn40bDT4Pq3oYG9+Nar5o3xDGoVEqVSgnMLRlVxwoejLE
dysHeFKppzyR1MmWAycgmJuq/uhQU7Jr/HZNPTbt7d/QT71w3FKgy4sjdonDnRLkaN7mhTMHy2WT
HhVioIzoJRtOTyxCn/tvytSkd0mndANLBzUIJWxY4D3t4WCXn5wRdOdBwCIYYh7vbd7z+Cjk80Uc
9NO3qlc2RTUY2TQ7SFZuy8aq5k6TAKOYkKBoaR9MzsMxHEMY6mPaISP3AAMTTPv246g/74588QYt
5mISqO3uBvzbIQ3SxBqWZHva5Cy6tkGxBnVT8BaEtzr2gjynAfXD5rM69gZcz5uSY50dSXKWZhiT
3i9f0XxQHS+QQBkofGG8Ffj3itoTFG9kXlOdiNQjYGx+Rv+yhqEt3k/15PbT7qceWkzffh5tAtgl
RSdlRskVDaDFaD+AtAhHveZ0BbhXVgJ+2r35PptKi3ME4E7kOrKUTRYmFw0EscLi9qz7Koiqpmtv
LhBSdAQt+UrmLAHIo59+3L/Yh+bIKTTcb9bQwoB/bGPiZL6BZTwBIgiNdD/6Lz9+g72P5X+Vzu13
ylS3jQPJNAOpCTUOu2AxaCWCm3/1/XJC32kdzK06lJmeintYzgHbLL5ItLiy0FdVc9hd/BEb96U7
Wjgr9eg6czo88JgEYPX+FpUqEy+AQJ/aWdlw0MpigwySaZJUImWdIngJQRlLb1K/AZm4gZsQ7oxu
hODFczTWSqxvrrUa+dz9fPoyi5cSM8hYc2yuxaL2p5mP9mymh7Br3inZpvYqF50CXFxd2v7NSJ/f
9/j5clFBsNUg7qBA6NukFXako+J4z+UruikJFOVVImUDsMVKxGRe0dj/XDsZfK7UFAeOztUBiGZ6
wTnRNcvNHR5vazT3CO9zknLwbcZILQUv0Kdw1I14A75ztZm+3d6Cq8QqU/1MhwR1gdDgOtahZhPi
kLDkLDI/aveilK76ORF+FqEGf+Ll+eGic2ig5XBEAoyzeYvYkO/htCWI1j/pbNl1p7gyZRW+318w
NEZnsnuxMW5qRgHqvbH/6xoTPR+MgggVSPL81Xfs4oObozrA5m0g+2fFrFyTpFFL1rxcOoEyvEWU
kDI4Jr9Io6WNM6MmqZl9m27QAkD5cNCEYgt2TKb50dkCr7SNjZEO8TjxdWQPRBz3pZXBO+aX1lZ5
cPyHEhGR1EmBce8tBvnRDSmwq6Pr0f0+BDW4ZjQOisdwhE+mMnYTjYyfJ9OYWPiciizSwIUa22W4
RFBmnvjRvgNocm/qWdccQAqC5SRdumIk0ROm6pBM1E8L0h3CcI4wjBLQvYkz9RnaOC6JT8pK+aX8
73uegt+fCSaRd6QIM3/ITuQtt4eyF20rRi65Jg2jPZHHOa66+lyvJwwIyjayp/IYhsjrgy5GNLU/
x6+VoPwpginoErvkjD0E9NpO0SSYzk8t0W/B3ood+3jnl4t1Dwq0m+XiM2l49Hqd1YCQR9SJv9Da
FTM305Zi3Bla9DMMKY+c/lJsCH+JhAwLKIER2v69HMxykaRv63eqq4s+tCYGtKMKVxZ3sGKfJYtm
69pb0y59h0kvwxsKdo4/MhR1ZbcK7wYiZe9FfRsf7GILQbwi4QAl7kzXaDdRJPFgWQDq3O2tn2sJ
RYp8INsNgjIJJmfUIP3HvB/aTAG1GZHuyn+DUuz0h8nQPl6HJVbHEXDLC/+OjaB0WGu9vIHyLA3e
rsO7J37t2z5LfvOcVYFXOtHIARfHZAXv+BkqefTltzYbxRcwnvU/l9/jCb0z78AcmGXaN34GuBIo
T8+rMHJjUphrWzy0byuFMzyYRASIWbzV2UGOG3G8Xu4cGpz3kTA5ISZlBDyvkYkYRffvXmtP8nrv
Di51z0xLO13mcJ9Pw7p9XMZ9MlzX5lF78k5M2qSEg2wqGdM6l8fTwXPCu+B7p0eeLOgO6ecv+4T+
C9JtFXSOvW/VzKec/C0Fz7zijSS8jvTRr9Nk9mJNScriSZ8MW/9bDTrQhiLHMFESZDdHnUuEFJnv
AyCVZDtjpXSYF8WN2Vo0ux9/Y4+6UYwnxIWcmy1vlVx/P6LHdcV2NeO9OMOtGRf4lc2vBhvKJ7db
DFB2/267drK0KzcriJ6EMon1y0CLobx2YTnP0s7ehgxUzJ15YHnoNyXqIpQNi+x+v3Xg4fxmB738
nlGfppGjhvjBrkLHfi6wzXANUFBT7Q/lCn1zay3SJCVqhgkQyrrFwFVP4hbL6NwHM9m4eB/wmL7J
G+tqm6u93aK7iDglUScdBguFAiJJM2q+SLeDLStbZjlsf2XVh8tqmG8T9yK2VX0hnuPKl/z1uqF8
sOnWjHZNUnQ0vwKysrmIzvSFWvAk4gf24niaxJytFDBec4aG1YuYKfKi2OnLDwNyVJM3QJTTns0E
N83s62KBfyL0E6FR6uRIxVS/qEtA7ojteg5btUqLFj4BkJxYm2n9JRigojg0HHd0zbwMI7rMDwwt
JWj4QgDlrSHlLoygQ06vu80aI5tGHIMg6DdweL0xM7UurwozxCXSZ2zYSY6jrgCkpsZw6P683Ul/
gOjezonthHozGacgmmeATml4xHj8Q/ACrxE+5U/QdApyH78k/tDB8AJMb32wKYHi3kslzNNrSy10
bLuwBDLfl6YQdbAjhg3aFJPg4QkVdw8tvBrGpLv4Jn8swz+rmII5pdu8PBxprgTjGfj5rG8OI6cm
p1DoPVUrsyIBBbsWboGwfbv0uMh1MLh7oOU8ubArp5g66YoqN5cWaLMkSOtBuqSpYedoepZP5mIe
fCM0m3pdgUEjBGboA0pELgNM8+ICPa7B5t5Cktk+2mw91Rt8nkDXhMyB3owesXysLialKOJ+GNBY
Ic98xuI9eJblaxzwxudr9JT2NDSlGcGVthhNpLURXE+QCvaCFgZk118PWPaOVZ6z6XPYe/Yuhh3r
NhRLFlJdLQABympNU/Bp1BfB4HnqvUrYsv75yNo2o/EiPmwfJQ5GAob4MfPGOWigQ3pYKC6Ic/LU
9hWAk38O1qD7ghnFVqymf1ABcpbCN8tr8xXOH50uA3eYOyRu6w0G/8y5IY/KX7UEd8Y4y/54IH+I
1g6IF+yKiSY4DH8qK+SrQA5ujHlne3WSheFyDCIx7seRnPoyMMYpan3kWCgr/wgSurI9io0Fci51
PyZBcvHAeqewhW+btgu6He1KC/2vZ7zsZp/iK1NdWikJtvKrBi95CwmPK5vXmn0bBcpIu9BgN3c5
I/ODlSoTF3feX/2S0IRGrYhqFJwv6Ri8TA7vihUssjnfj9UIxwE=
`protect end_protected

