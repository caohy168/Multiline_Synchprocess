

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XIV6+/PXm8FRNU72sonnILYjpxjtmIZbbVLNSWrsf17Y2ws1SDZw37iDqiHVxC1cBgNo/dObQumt
yWJq0muisw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZXPA9HFe7cAtyRoNz+yMSPw2Pyn+0pRPvi5XjdJyTktT81Si/ij5SgLi6R0lagxdDco2VlsuCFt4
OL0Tj4wvHy1Dp1ZlmyT/YK+4naDchHt6lXN2dYFjXydimftHAQxst9Mhv6lRib5QRDOa20ZQpskn
yks2LbBSk7XEzudIYJY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bg8I4RzLDMU1lDDWoHaHEhOZTFPFr4IVYc8PI75p6rwLWa+GCWy1qa8WABJB734VvQ5wpTCQEDJd
rxf1ecFNcNhvHhCyE2wu/BzY21WCLI1aRAqFQXE1qi1Z2wDjSCFHJSnGjrE1LDefRxcxG6Tq9XbG
It/MsawBNQzhK43GHNj1+k8zbaJGp860b374HkhV1ZfNQJjcX3XJZ1QrIoPuFXx4Jhi/vjSlVFXp
pw6iybj5y8cMBzzatmsSoxyLcoJGfbq6C8apYs6F5VefEZxehY+hYk0iaREI+yUEx1YOnm0lzVM9
0NDqetgtQD4GK5VbO0+mw0/9k6lrl7kHG88ctA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uEnR/Mi+1UEzM6gOG0vkJoA+Jn3kxV9bb8otdkKTuCLYdJMYTfeNAGMqrDN6fOncHFTG1XMkSv7C
TzB09OOLPZWwUC5RHySY8jhavl3U2T+KX683mdCktfKMasAgiszkXyARiIK48HqFwHJ6chQHZVFP
PHgr0ToY3Xkuv4qeSGPvpnKroN4SGD/mdjKnjoQHGMZuZK8qyq5742CAWbQu7VMown6q0X0UZPcu
1EmiqSozGNEg6NBdiKBwGO1I36DQN4XENNdX9KsMUX56OEaXF2SCnvpLoCayaA9H2EsYpnARgVrs
/vwfUY42CXp95G0sE/mbV+1ahx6recWmvPJSDg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NoPXYyMJfSM1kcGd9d2E0y9DsmmxrbygZhs9LH++zh9P1OAn6hS0Bk8t4Ndb86rV4ZNvh1uF6+XE
APAfkag1Joec7lZ031DktS+E+U7heIbtHrj0Z8txcCoU4pcni4l4NRM4qg2jau2rUeq4Ee2HKgWS
atNnstf4UDlnanJjkbw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EsC7yizglwjm/VQRLhk4w7OZ3mJkXIBqwvXZeGGoI2t8w43A9I+u12UGUeBgq/MHOJNvVYJy+E2x
CC0Muz6vedVRM+FhA7lG1BhtLDfdhf5tyuZ51k/7eDcVeO3IHHvF7XSPJrUQ3MWUinYFQ3+Gsygi
Y5R+qlsaaGcS2CMkG3/Eih5tpkgSHmLV0ktNrQA5e7TmEG0rhv9Zq1LfKnAJYbEHIFNcOJuSLtA5
plx+LBg8QKQ+k9ZVnTJfrTN8PCfGwKgQ5n3P4POrh1PP11JPRcM+bn8OQexcyQJqzY2NV7fLOQVq
cI+aLpHw8NbqgXQRENmxsQ2ZAaG1oapGd13YQw==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qGiQK3HCCFErao7nb8j52G5u1V/rXhGG+ecU5rXKOUf+5W7QurCsJoepMeRrQbXCDAHalCi6YEjP
SXPVc1914DtWdpuOJR9bEDnAtPisBxcDbhjyAaA5GzCo09H3cDy5rQzcsoGiGTT2ezg6Nk1pmUz2
fP/pXAS5iVEWqPpMvSBiURlCFQ87/ni9/RtdB0Uj6TCoM5tkOiWtvD+IVC6HJ7yXfevf56YqU0CE
qkKXwNZZsQ2OGwuT9rL7/cvtRSms1VFzrIDIdrlv4cDuAG5rFj/CLH97nZfGWwZ7B2Q4iiKHlcJt
wt4vxAZVcrklHBSJLO8VzMXOGbZnbCZmugsMLQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VSFFGi5I+8eqPTjkRlMIk7PN+dnGGbWsm1buYkudsXq7lN301VzY6tMFyneWG0aA/kEh6PynLm/2
wd6EFwFZ/CX6b8btvoZd5x51dtWrAg1xEwmnB+ttvr1gRv17BaIzDKRP3nrVwAbeIrguXrfzGUUK
s3UDXw/ik3avc7EUEHARenGpG1MkKjjnV5jUzueDFEIdC1NuYD802BHFg1YFB+51wqGLpBMwLm7h
CC/EmDTGGZYUJAHMTXNrXI7Ji4rxad7i1Rz+hGhk3whN8mhDdU762+MaCF90usEeFK/PE4C7MhI0
3sjbqKNFCjO3MEcV8pp7cgyujSgEWcYVd+eWmw==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lkdsksTGPshZmOBDJc4avUeYc7TNjcff/db8BrH3sr7m5ZC4Y1oBlYsbaqVkMalTZKY9Z63UDWXZ
AfhEkvl4BS7BTXTkLmETGWV28hDtA9OrBk+Eim8hy5x/OQ3KnP3YUrkChGse4nMdIrbWLmb2d33O
1kr2UzGclw+nqYyjAYWpbpYRPzVjkUMp+TTxy9b73hnEPvTwoisEEXB3ubzMq1CGEsUcoQ9+5GmB
VaRWjX4pdAVuuCXQceCKOsWQW+4iI9n62RvZjTfnS8VkElcmAbPOhCFrpH0kt5KaEJodOswVExOa
cdByl8ewewezhdqPRoC8BU6bxXhdis0m1VS7qw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99648)
`protect data_block
HzyGtEGpDzsH05QN7y6aeN4Nh8LFwnqkwYOOTm0BBvhlq6Zto67fCxwP8fEtlqT326yd2EjLbbjh
84gKNH37X+B8ghoYuV1SH+pAN08F/Miv5+9orapqe7+6rZmhL4u8rMrbCN6xQgDaIN4VRsXGdu5+
rQfnshQ3FfReAKVOxkSaJjMoEG5Neny/+jxl4kC8ZeWaRq52DurARHFXjJafO0ld8Amk709ilnLE
xTYuuOs47ihY+MK5Gxh7HaXAaKDss6nrF8ujDQ4Y8e0AeYwb2ONKVW1ieWFzWcSI85DIpsVsxjAP
f4PXWiwq8SWBN4ROmIcNU6q5q2oPzACYltkKHi01VznuHj3sHMWE9XMNVorGjLByggNel9amq0vv
V7nR1ZYoEGWGui7NH2fGFvbV1U6Kaoyh7y+kBMw76sqnDlKtjV1ezpz9hcKbYSyMlWNEuIXQ8Nd0
6Jgw/toMTXrvGkWnNYcxlCv8N6d1xb7/ggXeloc6yqOiCT7YRiJP5S9Jt+254vO+ZN5YTp/BUhhR
BV5y7EYiwh3x7bASV57IC6GMUWB8CDYQ6y00AEMcA0ISWqB9RH6VUtLVaCxMAQ0bt7DLnRZSmuJ0
MWBmu9urSA0zIkGjbpLSBKCpGkCZW2POtomVK21kLVpDQgtlCX5RBA2D82Ork9zM3l2BMHYDcsrf
OW8z6jkB3bzyT3VbRRtO6ksrbt/sC76CpxwS56o5faiBj3p9NGHHLHZ68Jvc2WH8umnr5cNNu3lJ
yDriX6090mqih/ZVVjTNp/jlR3Cso+bar7u91BNhHGtYQp5+S4m5HuTEs1SpcSyNFBr5eOYVaxiB
weI8OzCZNqhBOIe8dRN+Z+MydzsGNeqYtB7IznuJas+4jA8ZjB9L7oVszM1MK5+zhYsFLNHH36xB
SZzb95iwYSiceEtqH/Cpb1YZ9p+5atMNcHOxtjv0gdahBKBGtuk44j3SzDisUVWEyGuFu5BVKkQ2
ZJ/C+EMw/CwDENUhy8mhlYc3wcNMji35Px2WabXQ4SLKsocgfs3/GVACU+nHmbQ7sJ3MsARPrVFI
Ou9RDgEdGPp+PdT4T1f7hUZn2sK8HSiHLGqUenvc5pO2iqODJIJ3sjnvKhYVnfqErje7jtSCRWDj
7W/cdlxE74ru73jzJWiuO935B/9XADmxgdfsbPR5Se5tFEaql1v3a7kZ6z1JaqHsqZ355IFJuXqg
BpOj6ZCOlchYR4zhFAZUlTNy7mZoMqTx424Wrf1zYq8AOytvd6SZKAldUiPtUkLZLauvTurFbabo
k094im9fXrwXPMfHsP7Pvo/GWcaaDi4r/rU6n93Q8NvwAlJkkFLTjjImtxuI0eYc5H4ak93G0roI
PknX+FvFnMbbiqaRK4vbSquRRm1YeRvWk1ufYzKFBWNeDuWnGFAvM2qAQqZ56UnLvijVUroHKoy2
xzJ7gvRKWLxZRCVzfn45p2LUnPHGuucKGtdwgStvtaRfJtVKL8nIYzZtt8P8PILd8tT/3qIVTUff
+aIJxuly/AC3tb0VvHQi8WmoFPhrAD+VKZWZAZRRxpySxdjlsn2siQ4a/WBQ69FN/DMyxLSWyFME
9hFKcM66D/RhA+njsKa6F3uGHnZO6kSnrvUSP0Xq6RIy26BJeRCetvX2Ocb/sThGhXkblcXbM7ny
cEygrjUBn+CkPo7U63+HnyGYYQGw3+bfh3MnQRpe0j5ftqzFC6iNhnxaN45MqH3IoZ66N4ejRFMb
4RzUqDZfmxfKxCGa1mTAJcmZeNHW99R2fZNidRaVC6ryCzrdDT1tzPw6AoddIkT4pLT5LHLyoSvk
0ZwHS4x3A1WOsv2b476YEX3waGaIihtnFoMr/vh/sEhSjofmphtNSoSQBx2A4pK5fHT1xdxVSzwb
nAboR5Udk9oSaWkyNhbKC4Ajw3hWNK5SH75BBggVFZkndeFcBdxwf6hgcDA2hdDCHnb/Afhax9BY
G/z6bgjAKmQxgk4ta+7cx5Rs5OfSg1yVvVLKJlv/DF+r1Jm8FOjyO38cqEwAZM8Gyj6l5pBPuPmd
qDwtZlRplaFPU9TRzkPYdDc+o8LNEUxMzRzszma+G68aIz1wzHIEQPiGeqegeuxuvpUfR1qa2r+A
O0glhTI0bM0BpQriIQSt3d2vU7f00lzK6WOa0y1OF3JMqNaeOSwKdjb9xPoJGIxtHelPEBn8tusH
D4Mq6yQozxdNHQjN94liOyWmAWAg/DieQz3Jqj9hIA11VdCi0LWtt0tEx2rykB1U7p7hB9e8yKKE
rvPOSc/oao2x86s+XR4PsCYx4HadTlvHy/6AAPE4psxmdjIE2r2s8qiowjUPXBAQt+QjPvsSl9gp
jfueKkhZ8+YtuVnlupW8PZlQJIUxMDOhe/ZnO/pquBBcRTDFN79Wm7LvyYxoVqyWl8FrrIIFxXyY
hHlsALahvj3DfgxXYhUVc/uCQhTQoZdWV58JAzDaZI48oC+VVJX3JaSqiURcf+dHZkDZcwy/bCvI
fTi5dH5E0HPoDb16GQX8r42MOb0AeXncFsVVCJDXPdy/n3TkrY7DEuLeVZwarKBNTOdR153QpIvo
jGkuwDgozDdD4xRyNG7wG/K+9X8WNKoGeRWmuu+9gspWgnSC3+x07LhSIugWdlu/skQURHNMzeeL
ReHkp2fE9RA8WkRPAXl2Lnv78ToyjsE3rl2HK1uGn7wlMTEHUAEr6PzYOSHLVdhLFBevyn7EJ2rf
eEi1KEPdBDk9CrTVqkiuyQbFXUxXiGeJ4deoMJKZ81RTF8xSSx2fXUyE9cvwsIIrsnloTjwFonJO
porpgwPhuOrrhaPDqLKKBaNDHWNZirkujRkghvT3pFDGVygnvJXpueNB0M3toPY7dIfOXsvp1fjK
FOU6FnV32PpqsjP5fmjr2oNht96iMQYrwqrK0Oau7DwzTt0CnKdZYUpOrA6SL9iv8feAsGdzZhmu
c8dTRSoL/ObgOyVRSOZV3hFbRJGJI+05SRCYJsrLaED6qJm7QqKdFW0mJ2Zw7WaoPTgZYVbJ4er1
U1vjh6Bu5a14gk3gGIX1LG8nyAXdy8PTpld06aPQRGspPuJz0a9J/aNKN6YoCIDNR7wiP7rCiIBh
eWFIUiERG24Pcrm5qZDdUBRKHNT8gO9TDzU7jNHI/BaT+hjPcvcid1piyJ+CNrExTvpegej2+sR/
SvVFVElrAKj86Ytmgn3FlBebPL0p7TuqR2h5fDtKnlty8iBVHZcaWM1og7velzs3XkIccJV7ba4A
2vidx1kKsXVOIneSEX2RVvDaX3Tcblyr0xp509Hit39FNOvUW13mxJmZE+B4LwljQBLQz8jigr20
n5xRQtiLbmF9le4rM9MUICCPvLD6olSLBesxfpi6z8uFHo1/rwNGEzpu63lxQ4PCiFhwvTg5rXTj
pcMVruKDAQJr3WJNa4LMmDpH2WJOQnMy3X3siVCt/fsKHue+Z11ZrUjjZdkaPVA3ms8GdK/NNt2L
+4AfRRYkfWCIJlzbMay83i1w/crxADBBJzMFpSE9MiF4XFVBa49ftb/WE1dSpsrdvKJp59Jbq+vW
xqMQVcPTX2H3H79q3VMPjK3K9nKr3wWPOry0QQFUx8bnpOk4kyK5I1ruaLnxR9hA6Rw3nQ3rHDGH
Txg3Ce+rvsizSR780nPrzPpkAB4VSudjB7AcEshQczkcoOtGxIiwmQhWwhC0wPtsjrNd6zSLhSuR
ZS0+HKq8zhNrf9DqsKsP6+atS7Qubh9zUsnnwKSkLW5ySz5sY6bdPpGn/WfEdNqJhXTqqyvCEFCA
GX3fwKKIWFVq5HbpejfV63buHoRl5Uiw6BHP2bejWpCyqo8//Qf+MOnMPWDaFSAxovrJFz9WGp5X
z5BGEbQ2l5EsGtM5mPu+yfyNM+DDmyWloLQPyB9NelHoLyoHd/P5pyvCZVuXVs+xMyH7qO22MzfL
XVd6QsogBZKxuNolQIk5IxDCQ809DCegLug2cFxJcozWGW1PSFh3xKubAGfJ+hJC+ocaOwuovjDK
HOeI5crUkpdbw4gDtaxlOXdIbBra7d8/sivlSQECdlQgP4eYW/umEA8aU5hkhEw0LsTmjoBfChOA
A706SRlTebokqoePeSoZzjiDXqWRJNZpD7UjmYew1vQ2Yet8qD/72SwdUz5Iz9qeK5GvoyYzWr1b
SA8Xy2ed3zGRFQQut9Ak4w50PicKo7eJkY6bUtgF03l3Y4k0eg9CfJtUwjVuTpt5EPzubAQh3FP/
J6pLi3h3rXQ4LZtufGM0nxVucH1EubRNXBZdzymdxEQefx6+vUkxk4iZMyDU8VAGga5OwKxeIIrD
qyrnCl7BGNxKKOSgsn1kdJUByGUaIqylJjnHDYg2tzRjYd9Tzng5z4yL9GIOBs1/Trw0wVZDqLPc
WaiMLZ0NcY3kXTzLNZ3avM9MKZjMlmRUUOEjeQlAOLLscd8+zpzo8TOe+GewQFuWSlwF1VdgPU9d
6mXskFgzmB6pOF3jwdZT7MeMTZBmWbK1JFPEwRH/PJs3P7CPY26ZdxAQrVR7BbYUcYVy//6i9jDq
EV1O9ZxyUgdHcIMaZq7k77Xk5y6xWZOZlahT1y5r6tf8CjrmVE65yOq5SsZfvlQYI2IXs1DzBQUD
Iy5JxTVNA5VlOPUk2UGBm1p3y/XUkrLfProN2T2pyUydJjWJtQ3bLTLXPVUoGSdQpEkhqpD9DWLZ
UoJpbbAH2hjX3HGNDSdG3tyRVAYdcvMJdttnJ5EKL5BTfIxf4l5u8fu5kwyHsdwCGC4XXwq7RQuh
wsQsgsO0oH/FEr4ud/azMxsiuhi3hZn8jfcnWkywgVYS6mrgymKNQ0c0GdnZrE6MdLhNr+hM7bZy
PfNWoOkGvpmXi1JbBf/ilcsjugo9vidDaah+lq6ayNw5vNAutSQ0w7nP87CqPYDBqbuew/+rEAkB
ZB6dYiZdoBoIPiL4ZnHKbVAm53Pm2LdmXgQ6Yoryb9tiLaLNHQf8hGZDJD+xx6El57srnbFd49AV
56k8nGQe+4nfm0YQiAhLWgRKPV8EvID47PM4EWm1kx2XDibIFlfltAdSuHSKk1djIYJ/qONt9z3S
M81rry/NRuCHM1XnyEawhUrJKUk7x7KAiYGlv3rGeog0iXwGnGC8SaBX4Rq5ZaD+w52JFxymPL6S
XVP7Xr2xYEg+KuI3941alRcdyseUqv0NWwUenmfli4lLU1mlmC+7yZBwI7kVOutVcJYqSDKz3NBc
sW1av4XRPTHEL8SYtOyRDBSsYNqZoZrmFUfrlN5qTbGhYG6MByHv+VvfnvKqTUY48EhjDuIwHAnB
Uywdfad+YGozBRjK3Zx7wwG1ooYqP1JbB/j7AG7p9cIdL3f8KI3gW5AJCJX86/3/gETGski7jK2d
H/1WTmBRABuZXxxCkbMGBYmUpybWSYX0JXPTHeXzi6+CoGFaDj/4cIK6i2mpm/u1PrE6d4MPrVMn
NngC5QqLx4VgftST/d5Iovu8FAY2pZr+3SD/53arrwJkmCWXHDIl+r0J0UJ14PmgGAvR4agL9vz1
WIEjhw8MKODlcEPUTKV1jyyoKTx5yOM7IflJUHwkGch90cnu7M0IlCIkG+znRg9UVNvIulinf94u
zjq//JMQvd3dwVj+u2SzsJfsEDKQ0l6Utq0GiK0LlrzJ0gLJcXQB0eEsD5M36lGJtXd5W+4RJw99
08Roag7XIo/fJPIiA0rzNZ9IFm2P0/bB5cZNnJWqoXvO8VNOpkW5DisedyAnCVdCec7VHLgBufWo
vKN0gVhgy4xFXhbF9Vdy/ko0MJuXU23TcYgvIV3Hrw7oYhuk2yOoBUSmogCfHDATFuTMsJc/BlLk
rn0h7csgBSqkTzylU7unffuVp8ExCMZHVAkdSgd2/hTzDTCv4ToSVBWTcQLcuc08QDN6rLhYTlwD
+sWe/PxGzv9T0EnqNIM1z9VZ81+mAV8jfls9f5hKbZs9U+nWrYZirJ08uZyhBxgIwhOvkQW+Gjg9
ewiFZ0xiy58S+jaDKq7l6cA0o1zZNRwqv4ZqpTf+ll88NV6UzwcndRCTRSrxSzCbH90fTCcnvo9B
/hX0aSH2mU3e3KVyMS+0rG1WDooSKrLytYD7Z0uJHIy6yYf7cqF0yT8hY2KW7KWT7T1Fhzi970NC
2EaFj2WqvuIEIT5r+14la1iQLfichp6BcKuOi3gzPRsHqG068nO6O7zkVA3zbnoGoH9MmJCEPD8k
GUh4NWEaI6tca957a7oPoUQnlvepBJdJrq6T0hOWkzqZpD2XvLJPhS/3uRz8RF7ITKeQw4ES/Keu
zMCDltH4Y1WLA06iVYEJff2XfTqVjObWiLM4BOjiC9tpNOXIhBeE4KrzxxxmfpsPo/3TXAdeLPR1
/Ah6HNq/7ET03IYqZZTEDyQczF8WSTtZgosHOTvJKHAiJGNz+U87n9ES1+7eqXd/Q7XwDJVgizJx
PP3DDBVBji/gu+bqtaW0mNetv/gcc+kayTo+03ZTnXuAVZPG6RCnSW4ri2Hhm6/qECuo+6m2Wy9e
QyxnncdhAH7Z9z4iuCV3p2i4StG2ww4+FnKz/dYixYZgwmbEb5bgHgVdk7AbY3mKh6UnDoeTekm8
YzggLgy5B4EBKqNvDwkaRDZAzy02YphEpUVRRlgPTHXTyaXXo51GH55UsTDkhMbqdrEQX4DyUsYP
oLOVPOqDBacanROWXsd6NOohPsF8aVuihv/jmNU17qoTGz/Gs1h24xmDKKPdZKwI4Gxs/kdtWlsn
1UMqbnxyQOCLxNB5hBxJlZ5wzf7/lXqIT7zqj7+IhQ1ehQkMLLaWExPfXCAHZGqDk1qkRXQPJlXW
+auROOwTKeFIHUjyyDooga3lQFcaaeJ5aT1kHsy79Wqt1ngRRYYaQMlPeWup8lFRpLktkSCkgPZS
fvH2N7L3W9Kk0KIXfKEadUWE5m8cf1kqt0AzDjBGzDGUV5Km/l2QEwJ3s+s0oxTpucYt/V30A6Ud
CcnuAVDVJZt4jts4PqDtifScDhOler8mKINwlnvTHesWPOWw5Gv74o+PoSHn+4foqA5q9ZYyfa7T
+IANbX4AgQbWI0ePdTwIZ0hMw0DQ/aLtMWqS2dFXDFfcGEoelZzgRWEpkV4UUB/VvMtxKTgaJh4d
e719J6wsg2zN0h7+eYyMtvf4gYJCurJpzQf1URL6skK73dAI+bi1WBoyR41Mkf+miU/3JzBENEH/
EpdjqOslfij2EqpYuA/BI+lcuNMXPdt5v9b4S/RHhvR9h4FMSEq5vnsthmM2EPk/0WKrXX3Cveml
Vn4pf01cV+BFYWCT8kZO0SP1RS2HYsbhu7ah4zq7l+bdkWJm2oEEDnaPUGzGkEBTDrsoDX4C7ICX
JmO9m0ZcFPZvX95jkAx9qi5dlKsEjNT8SC3DA1wh3/fbUiETc3BPT0FpkA18l1/ANvXoC46FZSTF
fCVPFxaOYbWy0bTxW7RHXjORRFSYDWJCGFu1MP8/POfaMdPEdOCLW86L7b8xmyIlqnzFMmhQ38+W
4XJufLLDqpyAKH2PE7e/5kdQI2hnNv563a+5fFAFjPcWaiPDNDFbZpBytKqyA+9pKpI8s8gQYxbI
KZXKHWuJ/8g/RUY8KD5iVAWVIeOQL+T8YWAQ6WjvWSlg9KPapinXN0M5eTGJtiY4HQNXQ2F2xotF
+sxTgZ5J7LJDtqSOeown+wafoTgCcMoKqeTZR6hBxPw/HHfahbt2ejzMB+bL3jLFlLMT2rVEXtld
/rEqJX7n045UzISjx/OXf/trgEUsicR5X82xHxpYuoXkIGlr3axExl1uBsX48Y2aDlTImaKJ1dJV
hvUf5OX8N/qrM5OcA53Cl8lYAAoiugxIQsO1xR4hIRusNnd9qyEmkrMhO8YGSnnoOsdWgHQLgjnc
6B+MoJQZKShdAcPlAmTeLrmtH1UuVG2vNlFCBlDVaWuWJKAYX+z2HcXEAPdoKZgfydk2ErJYaKL3
X9WzCh/sJYMkID/y6ndCG1jbnnX7L6BBpkwBiLIexoJQn/VXKNSxvQaXKpvfrlK745wHdnc1brgj
n2DLRx1vrDsqWuKjMVagj8zAky+QF2h7ElGHURDAS9LLuDqDTEqyQugUBi0CMoihpPRT0QR/kqWt
/CxD9jQFR0hurC0ZSNgRLrKSY+wVve9LDvoG17GRf777pONdOwwSRRANTdazjk7iNUum9ojzYOsd
2RI7C5B0MXamvgCCcNpVSsZGgdRIjC+Pge2WUMr/StGQSwhZgmQuF8LBaqtyo3vUVSO61Cb/AWcY
2+tAK7pw1OCIiy75MslnCLVvHuFLyS33BmUQ6xgtPamh0ln8WE8C99RRmeH6hPdKqhtYiJf7wZVR
LeDq5LshghbQiYBqJcJRphF9rM3WlfF1PvnTHCVhzsr2ubaZ7C0yT6YNy870VLz79zOoqr6/eeG+
vKl0CdddO/SExGaDBsVtmYUZrSIE3ewfMygnPeLhA1T6aWlhd7kvYsNOxnpT2XUDYUQ7Azv+LnPg
nBakMVIBO0weg91FyFPs86TqV5+1/ukijxvcxZBv2M+M1cG226s7BqoA0pIyWav12DP3m5TuMZhR
PYPhHLcdAj4/oVh2xE0qj/djvDWPNpVx1VLxWY/M/w8vDGKQq0sDN5sKNCYxcyV4NKJlvXi2Fk0/
L1HRq4wTUyVaa/w98vSx6OKuixluebyyBf0ENCyPG+EFwrdwP34sgnkZhDstl/BBaOyZbOBLlq05
Ms+p2+bS0ylDm/l6gWavvPr9z0GijPiqiYfr/182SKk7ul85F5k0AiyYTWc56sfeLrbBgQ5/vF51
7lS63GBAaWHCmjd0wuIrks5Ye/aoicr1r+wmVQGkLJbL47oRb+rCB3rm1fi+p9w6yl8gmsoKuxsv
skcbkuNaZGi9Q9w0mcTAkjKVFg7/h2/uqduwea48j36I/1yUdzsiRIH/u3TnXwdIlF3/hRUls7Tw
5WzBSXSMhbKOYu6HpBXPeAvgKeG/jKE6E+rh61dzbMHMAfb1W4YNIRNWm8UE9PUOZBBt3G6Q+P+n
Xgy15YzzlhSZh+3AP9CTj0GPVJo6Bfjp3okkzzLcvXDmFTN1vwTB4pJ8QlStPrI7GwRJwZkCAAfV
wKz1h2GoE4rRHWBBiCmuZG/ewFmvQ6zzjZQKbCJxOjKE54bjZPpQeow9pJCMEkXfXjTD3p1T84Rq
NnNmcURb3s4hHLe+pAYPh4aGWkhlGSA+VfNL1RW1/sePFGq3TJJ9cA0RBqpY357zIbY6j434MTyn
8YEY8mRjYJdK3a9C6jxYWsemILGWWMMQ36SO5OOAN27MrXLZxIMwOiWGrI4ENfQAKlhCfMHx3+wn
j5TNhvjQCmq+aPkIjksrK3jUaVPnC3AZ6dVBMiqYNPtDqv8GEN9r0MDbb/Q5InJmKE5XyX9agr+s
sVhhiHbf3nO6e7XkG3Y3Z8RnJK4VeS48GPLZZe7Fq824HBB6w99BoDG4vyoWQZFrnrhJUOP0wLIF
Sba3jWeAPurLQGzDBFt8FKp+FZSudeW0hQQsQjrrY8BJHZun7xlgcJuffAzMEnBEukQ47NDKxO75
fp82p8aC20SI8NuPbbSQlDI8KMro/7wdARbVfRa1v2QJUHEszzwShaCN+l55SmsYyEelrjuzDxfR
w+8faFTQdJFiTj1fOGiTjaxC8zFZOlMoTZAaBjFZbDlpg5PabxtkTGlUFitWnQyJ4w1B38kwV4dg
2Q8x1yCbnd7TcxYDwGIzqGfh+7A6Ot1cj4cf2yDJKM+7jwONGOELt4B0ZCbR6aG64WgEnlEZO/iJ
qMJdDaVPSHQ7F/WME7Bc+y6g5O776jHjqSlNbApvgiUJ7/MPFod5g38jPnbZ1W8LdwLnS1U5D+s9
/keqCwjlVaZeRCZ7MmrV0ep0M0nz91k5ntWC3ljbi/1lTnVoyTbGxD35vHK6yWkbFeYOk9YGLvpZ
3JTZVyy9exZ2mG07Nr415qdJfj51pqWj+O5z0giLysCu3GvGydFgJPpMUuw9YYlLW87m+rHW/AFA
kIQY5DSNN7i/Agm0yFvD+LXbiy5c6kSQh2B2O8Oon/p2m7/0PEkmeFuZuIdEHW43uk1NNROlHi8X
1TSliBLY+rU7J6DZDIIHT+hHE1tGKL3NAbCVnUf24lqErtR27r3rAOUf11TtfkiHlUL7kBTnDyEc
L/AoJw+w2O0wGc+fGW/CM9Akg5ZAETN2eFjeoNCSlTZ6Co2nF3U/WqukuTKuYTZH8RQsKwBipz8T
GKrtV5Vrkb/Moo766jjHzesU0tZzyOmFTKCY6FbeLJNzJcoDlQYqhcN4BpR9rMKpCztiFvz0labS
WcwYCVkTRGrkqvbOcdagc91dJd/poGm6b/7VUsvlR+C9Vyaf4lu4rNp6kwfTYN4zSb3T2hWQ1BDH
n1+VVsZLx9Sgj/3js3qzuWP152184kSzw8EtqC1Qi1z/XWglMgY3VfvzbipebTSYQulHNnDHwT/0
3Y88eilw/gin5nWiSUwECVOiinCZkclDF3j2q3Dth5L5TGjNXrC2/4+qkhc32bwDCxQQ3Lg4akgz
KKwr0wDbYjgTbAT/HrtShCNx2VRSjtH1F7P7ClZ+T7kQp2QB8ai16W/32hbcNyWaQ9/mcmvvhg1/
CiOFQU0ZcKghzfzm+Fu+KQSl83uviWTVBUZMQ8/Mda7V+db9Xr5B6ITW7I3YxiyPg8nxYFw+ioT+
LnNSvEuX+S8EK3Ww1hsqYVJ++Lh7tDg1XI4uf78X1+d+HnBsW/JNhkJTtIF5P4sNHssM7TSgRBVX
hBt+SYxcEX8B6v02U8tcdlqioR0gDfLPKRKiFRQTU/FqoMyIpbXERDac5sysBn7DYgCfOa+CO1z8
XdTt9+xIX7WOEsUd0dcEjVEHE7lmBqXh3V9JHamuT86lzLSINraM43Jz2hLZmCbfdM1IUkZUjiKw
haKl8yB3XJ/Bi3ktYX3+MZcEPkPo8mJwBEnEMQcoGTbo9sMal2PnBgtFZcfk0LoHmVxmml7yJiVn
zZIZdmm8Uu0eOVFpoe8/tE/HXb+VmqNATe3mkZLXx/VBEO1rfju21NvQemSEbktGSVe9+nLrOIqR
W2nnacL+d/L1eCs0U0EBE96w1OtK64tAAlHQNkTaAfUDJ6FzTSivkO2YeKMtNdQ9DsUQYg7ipYxC
i1I6pHV7Bw0JWWcWv3bMEExuEa7/Tjdl4Z4ukVuKEMy5R4PTjiTHQ9AAqA1XzK+xJyjUHCt73+Xl
e0mZzubL9aHwKpgxloMGemtXiPjvo0qcDSBBb6ZckzPzZ4aJplb+OfRWO+pizRM2kXWL+u7VVxNL
RoOo6FJk3C6GGjEIoKPuSYgsWbYaSqAoRplG6znUsXNNABhQc63laU4Cn9q3KmjYmQm4excmbItJ
ue6tSNlMfUwj2NBtHXAuwPWdarOL6r8x45RAowlauEEhNNYmWTuBWZ4k+fAI5pd74U78kEmLr/Qz
xxPkF9LfWypfPKXM3BqbFJbb6i3bJDurwzmCAxxoKw3zYL7hNrQsIZ2BGYl0+s1JMepNZBCSSTPW
RX7pB4tahQZHb3pXH9sznPzYygs3l58rcN1hVC3i+NFFL9v9yxqD25IvAgRUODwC7xWCCssdkHqb
D6TMh1UDBVasa6PT/4F7CAyxvsRvqHyOBopXxUyMTTOnLy18tPHm9GuNh9ZaZDslevqEroBdeMbV
9XyACrk8k3ZvFFH1tHIexA9NcoV27thg0uZ5G8FF2g4xaOByGnGQUbo1D6PRscuCJp5X7BnLzZs1
cxR2fTlRBOHA8DWuZBv5W6VVEWXa3GMd1qyrGAQTEpRw+YyXrhTMvBSgw4bCIzkZTqRjo09uMf0L
Pdy04hAt8tqA4YQ3rYDV8GsXt8sBYgxheQDMth29jD2ROcxhWkpDI2IgRQIIEmo9sF47KIpazT55
c/PeEP3xoEul5rvUNfSCcKwbibt2qMMAGT/Gz6BfrDGhbrH3GkP+S8mJjAuKodvW8Y4JiM/aiEq2
9x0G4xGzUH2niuTG1n6Ld10bX/xT812nZHDo7sA5gnyVtBDM20K7X3ucXzmq9Mw47W8vFYPIi8g1
A5kGA6zVEwl+lzMfH5kLGoW2fdcCkUGt/h7LxRiTAAuErtlP9cHS+wmLtuWG04N9hgxEedHIdD7C
iKJhH76XSFCyC7kUq0RxtKeaN7i4/IO9zLMvGTKYUQ+Dx7oF+i7EgInb28su0fDsdIH1HjWYVO9G
NkptXCrqogx22GImfHROMdC+GVuwQy55dFWKgUdqEciviji49TN8uGciO8Btz183QoVeQita9eq5
+8Mg3kmqadoqq1njs7oI5lV3B2h/Ldmy9Ww9MS7lY4d32ooSQ7sH7V/yLTRnso5OL3zgta3oXOiV
bMyp2cjUQTRWs4UCIwiOVgxx49zsWsh2BKpeL/bFavsf1YcHwup9EjTAYAzkGaZkSm5tgWn2VG1u
Rd1FBL9k8Pdeh99i1Sa0BrVb0ZOmQ20uPVCqSS/BLbWreWdROwjjF2GKQb2bEnZvCPWVvVBRWJTw
qqe2O9SpHwvgOrpSqin2ZPkzBiAmr/TJnL/VRVrgQIwWF1c8Z5RPtaokAAfjoWmUUezDC7HqwRlj
en+y0ZnbYiTbX5cRP5vFPTgBHP7DQ6LDCrQDSKsc68wAjIESot4YCsw805tz8/tDu8cHE9Jp+/9E
/fRbdS8LytPSpCM+hOzE+PrsbAHkKc219QlLJ3ISW+QtaysjiKYoSZTZSTBiV/toSnAkcTk4z2ED
LVf0bXeMZGr4F2c2aHHOTJ8nNpda9G4BQWv5lVTcr8LEyw9Y9eWYwnGBWxwv53cTv8j8LoaszwuO
E4dW6fzf4Bcls1bL0NKxR7NFn4fK0Qujdxf7NE2FYMVwe3fwgdDV/9sUAsfjpv3s1HyBM1pm3mFU
MIYAOEBJoTdMorHUpOwa3FXP0b+qRHtORW3uv0bzuWuyvQI7TiHxOayecAMYFC4zBeLC/9bkb3J7
pX+rctmkQw6hRP854qE1z0GDeRRDNOORWe04r9rGqBXN8OygNZxDpstTWixnPPqCTiytYQ2CCS6I
QroQZLx8gz/yFlS+ANIxI68Jd5mW4kgw3LMIYlmhpR67hF0jKpJxv2iQww79WKKYGN5u+kA7ndM4
TrOq2VEgs0sr/asBxpgiYO/p2seMlXJIVKKM618HdXRGG4F0JkyM9lDSKYvA2cAwGJ+IOsh7agEn
YqLliD/UBpcFtCFCLQZ5FW/+2badTyFNLxow9oYGi3qHHTgA1Nyd3uQNKpVa1DcIuKqyOGTCoZ7M
TNrcazCDc8VfMqcx3pdF8BK+40QkPW4PDsy3iA0Ex5y7wo3ukbC2MkSIpbFFDYgDeBbrpYHcZLIo
a+M8Nu9F3cvo1ki7q6OVZzBDj4TH2iSThwLFzwphAMK7E84uCVfj3ukYTVdggRJ43BwaoGwH3ffx
EmC3Hbn61IK2W2NdYaHLEHs1Vp7XOg2tutx/RIqVSfL4YJMSOgXlZOkrCdDpyRqZ9xIZ+7LxqgK+
wTXtp42ER6/zJxZUz17yRF12bsjOKRu9vkGVfQKRPSwofU8OU64W32HdE6jSR2ADz44rkrH4DGnH
HPQnSV8J48JFQwX4Kp+Vi6UYDD0FocRjPlFoK9+/NsTLEEl98ykDu4XESBxAyPl5my3rubU4SaA/
nB8dHUMjZo8kl+H4m3k6erD3+Jpzes8Pv10SuSBawYrM+JTsIuOy6mKqV3mX/nQKM8YitC2ilraC
C+HB0VbORiZsjNXBXmwXIcktQDIhV1JFdonabjq+PIRgERUkOp+HawxT/0eJPLDF4fZY98XcIAQj
CpNiuLz8usCkXUgOHdczJZx9dn/6zwvFfeL+5IgO5vAlpP+0aCfEH8uKtuB11E05gqTaW05/Az5v
EK4aOYlAT+5qq38uDm/T+/dffKUUtPtYa8lReQ3U3bHWItvmaPwLjYzRIYcoaIFihuaXj9LEN3kD
JYhewKskwHfFx2bcAV1lYPVUV3yc3IcUrgmKpnPisuZV7NcbHlfhFQ2Q2Mh1ehpbgt2ix+jPu6K7
xoZzN7lsBDYK8v6tVBS6zhe4SkfBdXlofGecD43jiJVHpqD/KLRWXq6YzAkbwD2wFY45CmRdxMs8
MjJFmyc8QUKosXKTFiuI+o81BXjQegnUKW07CW3Vu+VXfiNab3AYiLcqbKVtEY5gzeYXm9NpVfFU
bR/xqC7TrvxgJKJErWxcdTnYrXDAmesQBrb7yzHNPXjmsikIq2apGtg+TJf767PNp51Lilw9U+s+
j+1IdGWCkqQiph4A/71cag6Z3QBU0WiqBHMfK3jH+OdUTzcGXnUUDmuelxZnbQRN4RdvL9bgPg01
bp0mn319Figg0E4aZs0p0LMXMYVWs79a93sN7tDfS+sBKBeOxCmTr36Tl6WJAQpYTehO5lFh7pkR
Xs13IJyu7bBqENs0bcpDd/429HKXGtXUKGCnAFDXWJua4l1/LbzrJ1KNnDhzYFSSOVMmlAQmgCor
CiqBaYc04BZZ0soPSaTvMIxxT0dmN0nTK69PqATNphJC79icKgHmOet09FqHqvvpEuCr9MPkr1nz
PbiWeyDuo6JSLZ2wxYYpnAYpekchsiG25u8bE4NupV8JWjjzxVVYcMs6BEr0NahczOU0pnZ79P/8
DousWlmkVS+yAO+VfJTnjbAPQI11hPQzlWG6VUqsWUHfmJ/PYWIrD/GlPXMfD9Xe5fZwdVw1dynX
kW9anr+/r+wlD4iTyAkdw6n/ixkiaLDRDHnUeHk755CKJfS5Q7StXEGVUSaONNpH1aoXKi/qNzdj
7ZmPjG6ZHrTapflF6ZN2bbw3doFQIiMFpk2US+agLszTh6WH830gEYLe2g3RAY/GIgfiBqBhNXgR
b2nepzd3qCgHuh+od2SVXTPzXAs604c5DtEvS1retBeD/OKEd0nR1L33doUDFg8ZprLMMxgU+wNm
zEczfM03T4lEA3bzAyihE1Pdpi3nVPr3iUARkwZYbqmvuRPVc0bz2yku/aJGvZyNpqT7buJxTbKW
xqLS4amp2EBbQ7oc89HzB0b+33BGdf52CvkcQ6rueCQc9xIl7bgJmbB1FKPttOG2r08BEnE6+Xcj
W5QIXRxChfqPBbwVzhYDcAt8rCgEPxtQbA1Wc2zkGFGJEaCBDf1ExTEFPJzB2T6cKmDZjlR9UQtO
uPqsBQcGCssRdJyQC5DGhwozKBMOpNeXa5M9izm4zSN2OBFO/F5H/wclK7zcLAJhj4thTffseqKB
2OXPTLDH5z4oLV0i+WQWQQNIlO7UaDoGfQzyYLTE8LDRQXMtvkmGSZz4ujaDlx0FEEQWeBb+8whH
Jr+JiDCoKID3Q61CCxsEjwakDBXMGN2orcy7gZ2k9XyZArNFqExt4atGLmzF3QtamX2Pazj6FeXu
li6PoLwKlDa/lsJi2Gd2Y+qEDTeHmYjf3MX/qYJC+n1rpyQECIyKPx8Dvhv6zn2AcCjd0wu5Awdz
I7Mv86QSK18tO9hZ/7QjCGoRlb2qwP4dXRVVSPFQ9deY+7qrUjRroebjH1fyKiaBDZJ6SA/jF+qL
iDSUGFnwrG3U2yy69ESQxWzsA22zPGwUeSQVgW0JZUvcO2CKP+MLjwRQ4omaYt0MwT3kMM5DKM5f
VJAdwVvkCZIYng3oJztJkBU+HEmvkx92toeFwRRWyiZExGTMoZBuEvF3xzzWX5RxwEzXGFsDqQIO
ZVm8gjdVkcv1HX0HZvPeqhtx8FBTME5xxKwMpxSDS0qITxxromvBH3VAJEPUtiji2NXoTnf/fuBu
DC0OEzyYOy9mwEMQxA2clUED/2SE8QkWKLUup6M05MMTc7rgYSkWRZVdmlqmg6pFMSHVxMSUYD0o
6+7H9cdtxAjYbTpEcfczc0gkEgwAaqHGuOfJUoVCTsnDPwbS1G6AshivSYf4Em0msCUGnak7zm3k
yI2L81ENQlnfdu5j3yd/5SeW+zqiNokjIZU/sQ3NZO3cJRh4HazHHYfGrzUA90U2FYW2dYRHFyiB
z9fHSm9h0lG63W15XwJFnsIIv0869NEvU05kMRHmGy9J0ucQYfd/x7m3m7PPxAbjAmZy7+XgRw6+
Pbw0znuA9BN4Pia4PEhbI9IVpvabFU0eB4EX7f7v4D+LliLAd4EPHD0iVHZualR0VTUWZWHVibdn
x8473vlqX5WUsSSYfSTjmJLok72GIkUbSnGRD+4PZnRQ6TjChroUC+bBsA5JBbE1RK4b+nixahKC
PA1wUJeAAatFVSN1ICBlDYeiPJE7XUyj+0VMLWqgXvpQxS9MwCF4I6OG0CxASK/ApBrggnmuaEio
3KkRpFmmjT4Th4vACcZLKChc9zYWZaXEj8FcUDmNW0fDtaM5rsEehiX+mR26DyWjAbqi8ZlzQqUz
3Lo+qiiRCRooiUazg4xQrLRvaccdQnQYrinPWOUnHIi4ItNpjI4INF4MAVDUWiH4NPZT1eqBIecZ
S02V2P/hSua7K5gNw6NUlAbmAPgijkzux5vE4dNNgTgargCyPWeOWt4G2SKkzQxYppT1eZOgD5Fc
2ilZ1Wft+7OTUe4KnYORn4oMvYE1+q/0nprJ0Qc4Ovs34dseU5WzHn6o7S7KREZKZErEMX90qhBq
sVWGTYBLE56T++RstthFAVURatJ8CMjEUXZGnsLzLWxlCylMHwetsTe5XVEYC1AilJJoS8Hf0oV7
yqwOezYuNTAQ5FQOPee68HJmsCbgQfNzZ1V2EP1NOTvRoxwG5FhFJf2nx4VelbNTVUjqaCCgJVbY
WRbmGq9+4sxJ+pw+dkVufk46RrP+hKsykztnEV6JCXTUHlFS5OBN9jFl5JhoUi4yOwS4ZfyC1/VV
Cbk37eihzW96AhT5L1WuFSIlKekiB8oJINbfl1AdfPmUu6zZc39saCAG1M19ocFVGkzEjm7xVoCW
Qr3K2Eka0H3pejiPzRyfWAJwY0nKaKVw8JqwV1cgGjaFmuA4/twLq7uLO7P5dAXqjHH/iSD+Z74Y
yvfw6Fp/dT1oqMzB3GbDtcjcprBCO5Hq7PpxZeosAodP1Nhd0WzG6VFyLec+EaJ30oUijc9bL3Jv
rDTMahUqhZkZivJbvkRh51oH+n2NWSDKHVvT/5emt14JJN1lV8EH2lyr+vwMCS7SlDjtEFWF3jx9
M9a3HfpIOu0HRnLIORurT9WltH/l8Qg0vuhdMZZtL7w8Vsrq1iKoS5JwIXsbBhQOPNLfLTKm6mJk
g+MAbLR4yv/o4neHXgM0JRfBCv+sxa6TsLcbsPHkXxhm7DmT7Dj3rohVbzNLIHmzwYJerBFd8S1m
dN/H2AZ7fvqudGC9zHcHdCQ++UJuE1v3rDtT0qQaiInwjNmSbJfjwEffzoqFn3LkyN5JfdyugHin
4Tm0PcbFkQ+gO6xBhr+em/T9iDSiH8U6KAJ9o/Hm40ItBPSMF1MiT8EZnfsO9oznmT9yfGIzBQJw
DNTaVAfgw5pZIW12jVeLgA33ooLrjzKAG4/1LDbHAVOZOlr3BEByROhT/cvh0ea4Zv8Iecl9hfRx
Apt+qnUSY4GIer62EGY9waiDYqUYBrdZNN2tcyvWCEqiAmEGKz3QNB+MkWsmBFRBHB5Vc2+h9Pl/
ySmIsB3UJufgLPDTzBf1fOjCM0XJbUTAa9l4tg9knhQJL8w/gbV8GV1PomvdXhjkMK57/jKCMolz
ZQ/JNxazGaknukFerDRb5vbBlsU434UeR4sVMqIy+/EBYe2GBFXh9m03zS8GRLj7RaXSVZOS2JFl
CpcLuovAhMx7L2/D3q2CrguXKkfEwagx1vFefGo9diNYihIxbijeS1XYYGYTdzl1G0OKVEZVMTql
s9bmXR8ddxfhVTeUHB/LvUAE3hK0KDyMIC4M+tlq35Hgu/XdRst/3e081AqSK5WSXy2O6CCKk/6F
VVz0bjp5CHQYd76S8i9/34h9Wcvanrzw4eB9td1ehMzVxAI4p/Byvlcwlm7ERw/Zt/QDaEr1GMjl
h98ib3Q0DO/tM68nt9nido1mJ3XHBNshzNQ0mPQhYJYLuCisXLj838X3bFjFDEh3XIrRwx5+5lRP
ij6NCY2GIKuMAn8K7wtIIJ2d7ID0UaM8eJyLJ6E4XVkkhZP6oEdQWuga/lP3yV4EVdTdOwPwg0dI
tA8aqt+m8Rmxv3QfwZ8EGEQBm4/dQmbvf77p8Rq2i82ZRCg/ccDi9Y9vCtNZhTie84Jh4iIGM9YZ
gP0zTRFPI8Tnz84ZQr8iYsPNBnwX4rN9tFFG0R/OhvF19NfOLifXQ9EdK2yJN9vICtuS1ta8meSN
qFf/5Lr1kDPxO5fw2cCPfrtza/A3vNfzW+M7rxJVHUQNAzeqtBG4fuxcwMBvfasDFCbHCTKfWgk4
FbUdrDU/zUJDO5bTG1ZMeYZT1qHk/t85Oof4SPmWcnQ3Q65UAt7ay8hFTR8xrV/QlFVeOzEakucx
luLO0lbdLv6aZkzYKKoS/lxLR9k5dd9UG1YI2PamYDpVs+wyGhzXwdpp/cjfM4/OBpnBG4mQOSY0
qboA4seo/nnSngjrNbhHadZuA3sr2aY85N88XhWw3C7eLbYnif+G8ifk+w9GXjwAq4LCEHWvwl93
o/ScOf/9lxb15M9RdY4HBicQfp9EtE2cGWk/vvoenIANJmLNokkrIRv6ThKBkbzx6/7U9+4+LsVF
XrjQpKEU8U1f0Gn1+BYkezTbxB+vRGZ8mm6drPUBhRT7DWO0Pttpzk0yhZjDA1rv4Z0CfbrhJAdt
Aqwl1Pb7AogLSP5cMcTF11CoRXkRmTVLPFLXctDZE0AMwJrH1vT8HQlAFK5F+oFIo3Eby+8rxfRl
rwAXfoeQqWKu3ZK4CBNSjdqFB9MDT/h968+4GoYCFNB87+PDKsyvt5MF/U5GoiyibVI5IXelobUw
GY0TMUspQITjB+oMSI/Ww7TnR0SgxyT+WdFIEIJZ3vcURTSTFzXe5I86R9xeHDukOegKGLgib0vh
j5/JxF7IncW14eLrizjcjSWDHU37e0y4yZT8aY568Ir2dt8E6buhhjj9N2yCXInNCbiWLzsQLbmv
TmTpsp8El6RjckJlQdn6CE5IC/GkPDBJpqvBlKvcYfIR9NQSsWq7FM3Th+pGtDYNhfUTc8sF/G7a
Ht/mvKqe5PqK5WNtoJiewNYULVP8BICy18Zp7wL9Y5S0CblRY4I9htImSbko280X+bvs1PzUxWre
kI7QL8rHSZDB8UzlvVn5hhW2M/nfSfm2pCUmbmWn9OvgB47zwr9wqlTflm40kon4RC1/lmkVe06t
6GnhRO2fvgvfDEMOhldxgoUM4E9s2ZESztFqnjDNTvydyNIfIiDGyHYtNLrZHF5zncwmKbNVy4ja
zcTxG72nOErlnNH36OaSRoBpOGceLXQJksHymbOb+dnXlsTEVWj8t5cRwGxgawhMseSGVDlBUG4x
ckEg6ozB9azr7J9t2eGcpHUhz1up1kmmMW5ILsfgEthl2MAKKIDNYMdNVniXYf3btszXJGC/+S6k
8bzEMgP0GawGISV6pWhuc+TJgbIDg1mDcFfgttkiPVjvPeIG5YZetR0thNWQb8nnNo8J/ogDDWwl
5sd0XKWegORJg3s+cjASWb56qPWiKhdKVEgaPPUzhSRumpMRTZCJh+VrQNb3TICoBvZdNSVyfeXB
hiVBdzO8vfuA4yDrmlr6cWaxHn+2kYleBADCC9TjChKORNj6IU02hWiqcOq6z3UA2JDaRa9W8iF7
bgcCnO561XCjY1RjpcEpvKRljrOlwmvcP0D/syKfAIgm11qdTevaiBU8KcFoSAezeml3VUGQ4Kd8
3p5GnvwIuUB0I9A5ZeU4JuVJtiYRlg/1eSbP5ZNVA2/JsaRteM+VehyobBYaYHzkuNCobJ2gWY77
61gIox25L8vkl8qTaTxP8bKWkoU9wrBJGcuSsJa4R7BVT+0tpPX3IkdZFvwhq7smWDmXBmzJ7Oai
cahC6iU2ru0ETxhKDkU4gy3qUDHn85BFWHhr5sa1TJvMGlmcXsowt+ASploVA1lfZhNLJ4v4d1AC
C5eTa44mDOZ5Hsaq3FlqWgzfhhodrOWZ0TLjZ8+OJFZpRodDndoyLfSm8nrNbdmf0DiId1weERaH
/4f14FI2uLhcnSVReQhZoL3EP1vNd1noQwOwjerxm5+pW3OxpGSiovgppMVs5hTR2TZ9D7KR1cyi
UOZpD9oD7EHOMp0e3rOyxWR2ZXlyrLfa/eTcUBVXZQibVfgZRqT/G8/wJ7bcZbzPsquezXDBwO8l
5Sps6XbppNKvLTs2FR8o8gAbHgBy3HEOiDpRORpgTT7jAPQCGEwh8/otmvRTD2LLZvW1owxgKXGn
rAlb5AXv2dA0CQHeSwc3RH4t9s6lIUSrI57UCO3VxqEzePsbKMN5OFxTtdOpOoq34c8msqUS83cX
xLMZR/T5vtLoqrNxW0/DvoS3wdlQS3yjYqIooPEgccuyNyycnr/dDP7R/XROHPRulugO0pkY5JOy
4yWu31EV5vEcI6LIrIJxd3x/Ab+uBLbf0Z4tpR8fBXYhf78r830Dw5BLTFN4RtNww8DqjQw6eiPF
Ym/BUh0we7thwdfhBHZ8UXS9qo35mIvNOJoF8KfIyhb3l7rkBr8EnQTdIpR+m0uM3p3RTEEqrPkf
wLTpCw1q0wc+1txpDuJYBcHIDD8QBvcy/sdMeH9WztU6bakIWoCsFuxOpJBwBMuvMY1+6t+R4a6W
eOgeGVauwxJ2kyMryG8zbcg+jacH4CAS9tryrgRaMhbmaC9G5HuY36kmw1atxKG4bv/nNKcHz/Jh
yW/bNMawT7m17R8Ezdv8N8SUA3g6fs8oMCofFarHHPb5qeprWurhMpO8fvhfEBtFpycOrhQlA1K/
iukWFx9yRY+ZNBquXJ2s+2WPbsyXZC/P5gmO6OVBfMStzgU6hQZbZvRuPkE8pNaqMjM2C6GeeWMw
kd0mmnsiMx49VMQLTyUJvN0hHrhG1kYBT/rDLmZ6owRn7j6muutG0XB8lkjZ46xmIhb7zrOSNZLC
a3pCprsnd4gKe/1Vqcfqz+MuxlqlwNpngYzYggSvug7ZQlDsKmvS5TX9nLJsrLCIwkzl2sdjVxNR
jQU5Igs+JIGOKpHIPa3QsrdqqelBW744nJ3j4sc73TPogHp7Om8VrKjeVwyr6XNC3BauCEOXtO4M
ZcKDGY7L1sjE6nrVcLykiuvrqa5q7xgx/IMOqZ2+hKe57Nj4yH2adIJZwjpczPfDFZSQG207Yfkx
PfMEmlAhih4H1/ObRIEdwoknUZz/OJ6jHq6KEls8Ag9CwhhivXXJMBClUzfhkk6TrEILQ2WZs3Qx
bD0Jd+cifHRy/YxGuqyv8AmmsuHjIjXhRhWAHdtG3HsgOzrpx022QUoIDhR0vQy7QhUunZmVPqnZ
WTY3IpeBuZike6PY+agWQCBJfnVWSrHlQXC6HjLiSzoeUtpZGTWvKRxHoezvkz7ELCDeZm22U19O
PK1Ub8zvJSsyrLTaqG98d05f/C+P3L9msZjvgQa4owzOvUEcLh+UyKCD7RJENPf9m5kIbdXIdikb
UjCdrSCtQUNT79IutWhV7ceFS2zFfMesAvhPWZ0/0dNmYVTZ4Kk8GUn7YtCud279955/l37e7qMj
an/eJLvuhlQnbYiSLZWKI3dCdpPaRbkNQ5lhz5JxDgY4SiJckgSYLOao+SV93UJEIb8/87JcbJVO
bdrdCoxB70LuecobCFZZJP6tPpVTybNCZF5MrQgBJrtCfFXrq8gjAJvEVE7vwHTAVUkPLR4LxqrZ
TkJGh80+zsG4NTfUMI+/8JJXrcqWWvEPV6YoKuJUAVQNxU1WHORZqsXXfG86z31aEbq8yyK3Vlwt
te3I9mOZXjvO3xqyUxIW6Gi/WMiCnjVzp7oB7jg/MpWC6azHgVLt/J3pyPkxB7gE12as61ogOa9U
1wIBM8FmKCSUPiUd0ATUivjI6ovqoUuyHPEK7wHe90jNcuCeUjQTalc0FLmpMsCa1xLQwF0bLyWV
dMc4MqB2KCAl7ZRjBUXYvcghcOq7s18cZldvVQk81po3upXuSjM+Pqa/DFNpdAmqT5GLiokhR0bA
DGn+wMwoBO7k2WyHvYSCPCiJf/cbR2fd7UaKqdvquVvKbA3NiTjK97Ak8c7S2UUAPJ9K5sH27PIk
6dZ7hZT5iIUkTvIAciv/xw83OdPBWtJYeA4hra/MfwKIlbIs/ujwCnK8ZwX+GGl5UeKxdtktfqor
vXETX0/xPLFSzIxHr3tUkNOT31lgHvMZFlYf61roHmNOuDu/Ws5IEDoJ6F30rOCdD8ObNClCHaWM
01MOhJFhNyPkW4wYRLLbi9sFLNGoGXcMA5qtO6C/2ZUAd7f/gBj4TEDx9IUImc9Bo73z6GZeoN/H
Ny/XgEWDiXmZwS/cC0y4c233e9ctFT8zjpK9chQViY3/tbGlHl3spI5LUMJGceldIIZS9RhkF8TT
URXsWH35kRHnfZfj2lxH0+QW4y4sgjcIsBCRujmm69J4rSrlfvWaaP5wvGmdAXQU13Rb+ALQTJu7
m5QsrwnWvGjEDZXCQLgl9SaAImBzcqp4b3yE04dW5Q3k3Iq9PHCIsRZ8r3Y9oA+dleAFRHlKCFHq
mbVOuR/K70VQ9YUkcaGdhT7RD3zTjzPA412vY3/jpWJifpXWHcWVvG2gJpMw2a4yw+vNvVPBZdvi
FpPBzseFEtXkB9V8e/MwFgyQiEi/4TjnPcGN6ZBHpYdev5asWeETpzLtnGfwttAOx5UmyXVB48SO
nTQL/rvp4WZkY8vORbo/oSMSflMWgYz0CGTy3IuSUATbVMu5ZD06AnQLAo8+ouT8HguXy9DFrx9h
0yjNXEUCxer4+WxwQfXW8zYsOg5bSk+rc3NCLyK2Ypb5vai/3wY5oHWGetg235cjfokleQFRLSS3
F++7zbMdidzTrEUv6DdfolupQSjWntyNLgBLCIQD0+WgyN7KnPJLwADRAVVmHkRs7Tg/JaJzYh6q
6aySfYu33uSBe1cwDbBfkxdqlFo71/UxOGIhpsPoqzRHGEnDQ1u3XN4S/RU+QbdcpvRwF0EgGhQO
mb4kJLl+MIOIZ3Lzp1X1dLnUGi+QITNRTjPXqSEd90u61Nhnq96UNhp8SK7BDa8Q/Hdr+FJDhFuf
QS/ro1nIbJ739XyabzJbfwqPMixWW+RV9ZPFfb3tmmNUtaPZBGpEvur43MFniKjGxYZ87OhszTCo
sKKrumZuflV8IvH9j7l4Pi5xmqeZWdVh1xZxcX13DWdgybJ8WnHaYVF6YsabzQWlZoKPRv18bEBn
uiQEKT7H7F54nk+iurkn/m3krT8jU1Gi0bGodDJKNRS2xPsz6eeLYLoWrMVz8W/HMwD9Y9YQuLyr
xmsZ4LAwgmblsD3tXdw7weJa2GSQKxEkqb1lqxAc1HIBK1gntKO1ZMmItPQq2gTg2gQu3rn8lu2O
1Ya+mPU3geggAz5u8JlI5JU9QHYaLQIpLd3JgahHo6TDU+tCsdYAblqfHXAjhr/Xj1ss5mE7SXX/
icPHnVtXnepJvGWJrRCiPAt1oeB6YCBrVWLv4euBFSXR5G8hWRdG6jHKTkTUZkcFmmqttBvZuvpT
cIN2oWfKS4npW0KsVEVLUQ1emuskDO0Wo3ZM2q3hNiJgOCpFZI2tKt3Y981N8bYEWk09P5X2vHQi
i6zULialiSkHtD66AXEYf5WbOUSWDQ05oRt2undiG+shfGErSNgfmlxw3p36T05RWPXOe07Q3B/Z
LV07m6H1oDomYAhtEuxRUpk9kwgR8MBpJ8eiaE18nk72Ia1CpHG9aCCYK1DsAbf4zZPld5kTmsct
JPsRy6+haiHzykMditYm1AGOVh39Q+vX8My+nrmZoGFEV3A8CSJwgPcX4fA2ed6PS3KKASfQo76G
RGH1o0vZSsHNFrU1LgMf6UhkuD4rjhAbyXqTlVHoqOKTrpW89lB/Bp3babACnXSC+ipsyVC71z2U
+LNLLBsdhs2gGwmjTtJ9TVGW9VVtPfh7ziB5Jqv2PogJSx+fYAFoYIkJ42GDYYdILBARLUaXPK2D
O8q/UNNE+3Dr6I50Zxj4zIHBa/U1hl4jxvHXkPHMlUgYTqck2sAs9VtvczTRrKZhT11LK3VzsViA
Aws3wTlaETy5pEVZOblhNIraf3Zbw36XsCy+VjqVx4mUPjACj/Ci0Wz2bpOXCS6pxy+WMiarRo9o
djaQC/kq4o2cCG2PHh3unL4DD52LgapygCZ+jBnYmpPz91qsfppdB2V42mpu2iJEGSHi3popkAtC
qR5V6mvrmVI8SMJzoACRqOA6lDcM9y/fUM5j3zCrrCU1W970Y1Nw4eIwE0g09wt3EGaI87M1agK+
97qKdjOT8jxKC3Ztct8puAnsJBbzYVduwP9CPNj6WA67fYgjMSb1blGd0hMSCLN45FT9Wa8jNgWt
WTMKr+28Aoe+Nu1tc68Vq3LqkvDKnIaj0euYLXifneONCGbVEGiObxfA1SBHRT0BSEGyjXPSeZH7
JHR1qfc6vJYOFtXCZa33n71699jkZCIaiJaj6SjbWd+zHylrXS+CU5pEDaR8+DXB2mGwWO70nLiw
FIekpVh0TL/m2rR1z84xLW1e7eiksq2dFuuSkUgcXn6CBeRC1eCZVijoNfQMCYQ+VTVAZa919ZUq
UgfoGGUqvpGv/hGF1o3NQgUgKANvObnOMquij7mcB3opIyaS6Y6++X6gkPg7y7IpEZS4BH0neHQv
ce/7TOj+6ceZHu+jtf3XP9WhAkvMm0dKrvyIbvplEEYx3ic66tP0UFfbXeIRLNk0cpvOaQ1C2sGB
kQmRmL/OMoJpbAGmfuw+GhLVUy9dhUYLmgT3kNBtisfU24quRdps4VSVmVmc8NJ4pi1/at0Wi1gJ
Afb/6v20OCPesEJRBm8bomTeDtsVJliRjlL9YpEvHqPdvrtH6QkZBV8dRjFLDSF90Ex0A/0FmhOd
1iEqRHbgb3aERRkAVtp2KOcMqxmDfYmPOc8ZH4hWuSh5kN9aHsPLd4RU0fPvoUOG/f481gZ/ZeQQ
3Ni9uVSjAxm7UNQNlgBsqLjOwk68Hme/9xtk/EKdzntjEBece45uT7NVyguiTxziCFD2SO9cpJ4P
JZBbn/fkDkE/842IbLZRY9qDVzKRzwiKPEf2R0CGW161E8xdDKfS+pselLDTu4pFj6oW6mBCLZFS
uZtEfIGM31geP0MPOGMPeZ+qUtTghaWEUckjBFQopG1RNxLUeKht+rP3y7HmnbtVBWa5hiKDk6uo
CdxeGlirR83GkltbBH8ZGDw9nshUgfxr+Z46eA6EVX5mhGuHvkDNGhybRlw67e2JfOtDEvpuXLQ2
ehEoOZfLlk4r8FT3+q7aKRGiB87IkiVwqy5DU/P8kMKBY2CV+WrTT9Hjfml7hMl03NUXXti5eLm/
mr02Jmmr+wnr4IgYw5beYzHKBY2atbM5Y6Tk2WptVsB/8xE/3V13y/8ZeQVp51hx8ZFZT99w8+b4
UTKzEj940FXM0/tlkxwk1TM4EitIcf8Quh3FM+HpaCAxpyaQA7F6viQW9/stBrwvFZ+RWu+f1w7n
KtBRS0LWm9HSnyXCLqkmeJsvjeEkXfhi9UDWtlCci0U0ULY3MQDLIZqdXExzuPRPDXoAXTlUioFW
CTfKVl17f/fL+jgNTihnQpYP0PgxEKscPtLwT/bKFTzsrls9I21MfSZLCKXiEsDNvKBYeGC8AtjQ
mW1OypJeczjQPGldvGahJp1/pnU2e7x4Yf61ZuNCxLFmysbgJJVPX5g01/DvWVkioK3zk5z6UXpW
Wm9LnKhESqsWd0V0ofI7IE9gHffAi9xTq31hI2Zfe7psYIIpCBO9uTLOrWqyW1Byo7VuaRsLee+7
0IdbiOHLUMchWA7Y3nyqgRl9z2tDqryvRit0AXCDcmNYMsnsDmKOvnK/6ooQMsnVXUNwGJ6Wl5DC
p6J1Vw/dve+O/a6L6+U8gbOf8Ko1IXbbfQEPCY92Ot0EMxJ3Ww4piQ8llSdS/61SdOStJz6AzJ1V
H13q6t5sEqnikB/zts9Hq+vwjEetgAW7lI/ccY3CWpeJbDyBVwuGpF7ifc4KaOPbflRMXDhcfAiT
p9P6BsTytEN1P7Sdl9cB9yr5CgcMFpLKnQofaG/vLyjzPCv8hI+c4I88OsxR6k84WlGw8iz3jQ2n
6vXLhmGay1Zh8beojADW+T4dcwuzVRmYFBLvYX+0WoUi/qGGJlHRxDl9WpH5cMSC6Z+CGZnjbx7k
3v/HnsFomQZqX20mtqXj9V8FY5qcCqLeHRYhArKdAeVHwVq1J2LV4sluNyOEBz/oRFIQIsZOYvj1
pBiWieJLP4gXUfG9/4b+RCckS55CAwt0g0nYiyxOMHeoGvieCGa8skHTXuaEOJg/aEv2lwmYNinH
dJfUWK705X1TeYgS70PHyvb0ZHoTBJHYKMxH3w/+gtdb3OorHYljdd3NzpKudK4TT32iFq0LOcbT
WfKjBOZQAeK6uPeAS3rmiCeBiy1eqtd6jgxXwRmTyVtLbEYyDq/sSOpsghiEyHlhTpEnWAEKf49t
z82W170nAMbeESNcG0nXai0dakey0v2uJYHosWdblvZHd/nz7vWNqhmdA3fA8URhFcPwKkcig+Ku
YqYTqH0QL8ChtMGh5MIb8jfdCxOeh5aOczC2rLiQ/jdls2zOs2R6Vz91XgA1lVuEI5LGRff6J21Q
PFSBCvmHs7/ynx2sYNFVF0OhKeOVB9OFWFQTX5WRbLtASLivR2HLi/lu5+g4D8rA7it5FysluKOi
7s/CQmHOpqI5ZR0hrdb1swAnnVwhXdm1T5pqMht1QjC+aQvg4ihXeyW8qAjy5owCxunmWYI7LrpL
6WXP+tE3IRjwMlLXfYpE2HMQtg4SmqWI1AVPoEfmTB8yKTYSOMovzoiSFKjFFgY60kV+cSAelX48
j6QdJsqwUxswEFctAZtzgyIjIJ3Rifvy/+gXBD8PrgL6tphayfJ/5IYsziOZoQ8OCYkw8DWe2fL1
SQFnlrCq/USUKRVXnrics2i0Fp1SwQr242QBMmqxUJakFJTM2bcdtReyzAo1H6VuHwR+DnPzW9OL
owccGJ4XzvfAaW/ufDOg+UJ/eEMqPIsINH02i9AG15u36fTOE3wPvtmI8UdQ4O+0+O7g1/3oU3o4
4mlE1X59Ri6ZuD2mp3YcNasdiVUbdSK0P3TJW+cM4y77PSEC7eQphqOFpP7r/Fv6zWJB3J1/pRGP
QEVFN7X6uUl8IQGyi3ZqnXhRs9NawUBruP2y5cPmX08Yv3N7VrW6pQFSyQ07RqhkqomLz7UxcIat
6fY2eg9AaJyn1KE4HxWnbh4PDzcMIBaU31uVLKU7obT31v+N3ahXZ84bK787hVnj+ha9X9+uR7Ix
SEzegnETigDTkJKNp4bIXerNhIRJiMYmB0URCmUsiRmkyTPYzJ6TfTGkd4ykq5plE+KfGFiv5vG1
yXtoG935b+TeTKpWaWFN1dui8wgLpIDm5kWUgmouawNZAxx2mJgPO9+LxvseHxyWmgWai2iERUWz
oiQrwXrkOB2wgk3YUa9CGb6QhD6B0SH82TiycG0+4MmY6X4rUT7AcpZEz1dnDCU5gb6JxrN4sD30
hkEroAtBIRg+7m2WpTsHIGekhTFiLicSwRzb3bLNSMHRuEek1rFX7XimIFfb1T5cCdhXF2gVliDE
XmwCSKNM2b01mkfPGvsgeMrbxT5qTxPWqxYtyM9rpc/1IAofdF/e3kX2uEI5U+FS33SbgN9V6gwh
iGKCJq9yTqpAPz1ENqYRd3UjOJWKq58wQ6zGlluxIz3O3zS87PC5JjyEUF2lTmiUB0xKs8ymvp2n
qYr8twz5+IbTYkBjFfpvrsZXSgTi13yA/u6STcc3FU4Qu9U9fW8/NWqOkqP8P++mn6U8xQZKhPeL
i6+BtuWYp+xFJtqPtznnA+cnkeukZ4c24IX2pAllh26OmFiHbvTzUAlGPNMVSXZSla+ZgVi8XYu9
tYPhRxQJLgAag5WBbxOABbEnMHLDWY4atPpFl0J/Qew+ZXYHtJMf7DiVEulJvXdE9f/GvRqaLkZX
A+YufyBjShTdNL4nHvvcZ2nB23IGRKBcLQsmilG/6WoinqHecmQTR5uA14qdQ4oTsXJQ+Dx2Q/Ne
eNOrQCSnGb0KR8HQLGYDXZ9j1xhZOBMzDj8056GjZbTr/UyvFGCGr2jj+suf6QaCyeHhmJ5xW4eY
esisQqBpZI79HpwNDs/QgA3t94adA7ch0fKHbemn/NJNWu1B5HLsS5V44691MCwytn9yOR513X/J
CThDgD3/dT6r29CeqeY9ksA0mdCKFCuH/rYom2a8uzYe1SQano13znqwc4J7ZBv7q4+UrIkymblt
pwmLE6RJv2FOHinz5fVHqi7sr9LnB9fo/xJXCoHqaeAEEDE6WD4JoZa45PnigBGBuqCb3EKGvdEf
TTR3Pz3vrEkfZRUt9vYC4VqkK1dKVq9+ST9VAKkEl89M+73cwNTWVZ6iddG2lNZCQ0JWlKOyEkW4
Ym/p/naTjKnQym2S6o3ueD56HE2/t/OdehHYX8hEPHe6zPkQhdeQSON50tWt13l1GzjaSEuL0uts
goVCDsG5VSE0zxwNk5TFFA6pxjgwTK8ZsG/r8Z3/8PCcRprROySE31hBKPaGm1Zdv8sDrlcnE3LI
HJAiV+G3LGeXLQjkPoy/d0R7CjVBL4tjz4vGohxnUwV5vZizvUmm2Vn5R9nUiyjXwxW/ard5GO2f
d1BWIHKvUFyb6+cYWc4QFAKEkp1ngzo2EUTk57nbEqAgi7//kfmTAiQBl1VRJD5iF3om7ECx6HSo
pHbcj5ebNwvnc116czDIjwACCc30ZAio0aqZiCaPD1iRoFSf1ZAIMZtTSHZTc66I6dP0B8IiYaS4
54KMbO8ZORF7ZxfzYsMWD3que87ZKkhoEGRWFke/AGycNptwFBfRcGIl6Gecm0I48Uu7Uv1f0oPc
q3y/OA/H/F0VyVczgeMRxZuDqp6YUnxj9XF3fCqLfIof32Umbo5RCol/mr1BmAmpXaTpADP9oHOB
c/VDpbAnlCiWfgWYEr27vjO7hD9p091h5qssstIMdYov4+WhlmiOz4mlmOpSwpGm5LkqbTyol5j/
9M8v1yBTTKi2E/Vnqir5p4oFKbxZUIaNer4+NKDR6IrhqNMDcyfdi8MKLn4QXAcXehKv3jDch5xd
TMCwYAdIUjGtYGl/ydsYt/SQ9BpW3oOFLbxEkWzL5UUvWJVgg/4R41I92vnJrbivtRwHY8VNALEi
qWJGpNfz7Pqye1gZHipSwLef4MRi1FTJaEqJ2I62OSCtaD0FPYenHdKXSdyrQg3MihjsnVcjpiQ2
nsA14ongXvb2YoPy2YkSm900tSy76NgPy0YZCBLfAjAfHzcZmPUad2xdb1RWg3YSbsdFPYdcXL+K
tAmTaEcFulgvbwRqg+D1Vc9vQA6cqOODzGbhz26vUkplEnAb/eOhCjygb+lDKb/OEK1him3fCJ3F
fgn2HS70G7k3FOYoTAsW/hdnT7aV6HhZ2sqaZUM3SVKjzfSYghpxoxK/Fc5V3peL9l4VZLH1vrXY
DgkTGfSSC+zrSoNyBbzHmVDgjzEnYfxkpWRmfwQTFjjBvsizHkOfgW0Hw1olYuBvIvBaVWEsCovd
AMJTI0Z3k3FQe4Gn7/IpmthXQ/UNPpAWIjPTl6+VBgRww+fHizYwfOGBck1tEpPhW6lSsWrz5N79
mX9NZfkbQ+jLMfU2KTNxMgsi2SLNfpPAh7qp3Qzfoyl6IE0ddJPTldNozD0RGtZlETyfNwsYVybv
36LmOwI501FKWGaG/qUT2Vow5NTD6Bj0ewTvqhW/nwQ1VQ47FPbeyXUyvtd8gF9yr8ao2N4CBVrG
lWi1xLRyo5j+uJxHG4P1esJCNQgAn69E2qLMmc9nux1rbd34zIn2Sev+75/lZlW0xT1eeMKgOy/f
8YWRVdHvZ04qOFWRFo+tSkM5NzQVRJaHaWLH9xjKmz7guk6lBe8SipAHYpmko+PVeLFlPgUfDoTw
RI4zs9UAnFMKkowPwcq4ovOwHZz94PxeOUNziW/gOmhRp+t0Asqm2HJ0NYN6XYF1t+hx91ttqu9Y
9a1z1YXDu0CGGT8N8Ig8e9p2J8EQjZAsbPsIggwLsk6QbgUI18jJajzWTH2jUkmKGSO/3lQiRupJ
JlZceQlYGQXls0k2xsZblpPx/n13sEKynW10xztuPNjT7hgqevCctlHcyYVF7pqk9BGjLnLvD6ct
XRbcZVnDUgX1xQH3B0Dpv8cLKAmiP9wlgaPVglost6aodKpbzak20KoRZadQ3LYvzDQBwLS5cG/9
vsE1bnsqu+FYXmcWt3dlKrm++cwrzrK60XwcF/livvgyx+0Nj4oAfFP8ETncwxqhHzps/Ml1BtnE
SkmLzFVbuuoAOsFeI3V747H88tet7gyLFBYDRZitVQjfFrDSMeMwzJcX9J+KzWM1zc4rFFxmPSEd
mzh7Ay1di8O10MDPRHEbmoQIhVN2to//nMnY5I903MRVGWv+w5E4+Zpji/IP/FbHWgPsdrkO/zWA
SWiRNFyGGOzscVwUJsKC4hy6KLaaQ8Q2SAJX97zgeQJok5/A5wXrrBWQyGilpCSUypPkpaCUesXG
DjMP9DWClXtjLTtXnYCIv7o6dPvGxfDi0fcjKfZDRpbbLgHqFZE9punp3bZeGnnvxAdv3sBqft2D
H0qJcxpMsLW3JyGnAVugqWxnRoPk/Y+FNyVvSP6VDTqOjvjNwLROJ5k/SYDvPKVdAStIVdCxjaKP
KeitMvzg22/fLD0EZCcTECPdXcE15l2AIArSN1QOFK5Dgz3yEDRnqLxGQf0p8V4RGfrkqcs6dWM3
Bb/3stbR7wn7G7oy4mNK5d/roRsCyeayfKCQzEC1pi9ZSdYRRqDBd3Kv+FsvogqXup1q+Nhr2Sn0
cGuvmKwPRNkv0yaGKYknMcdLup8JFvpFYiyxsI1OUTgiTSHSZeHIO8SAB8gaUs2/8sLcivvxRpQx
VMQxM43IVWMumQPU+HqomS8c901P+EBlMo58EdhgW0+hUpTTLxfjWRab3rYIB5W81hOYXkc+zeyQ
JDTE0hsYABvQ8niNr1/0+kelRHT1e5hRPXsCCwXj/yMLb9AU/R+K9/AaBvpfkOrXUdYubSvqe67z
OfRc0ctL5a5NY8rq1pMYq2hJI5+yziG0MORMAuaXLLV5kluH5i5+z6QpNCEp5z3xMKLQI07ex7hv
7/NYK9ev4rgc6dWbsN1wq0rGKe3tMBx0++UzETJGUUzbojxiDA46kgmKtzE9L6wiaX313noeQ8h9
GRSCO250aQkt6MfRizsjaYK944Z465qTYa/yDauLn/m2XeoU/Pp2BIDqXsU1KqE3F2xUhVI/htCz
3eLeBgL3dzs9jC7NxZUqr4mPGKgsOIOSnRThmrRK/L4veSQqIK9/qb5ELovjxx6AcAcABYUMG7QJ
s3qOhuvQioI570vK6Jq9TpTMp/uGE4UxxJDQfapLkEu8piHnf11J/q0sH5aiNXnZo/ZHnyoQ7GaC
N5VeNvRpRUm0mXMrBQypg7s/F6ISzcr/Wkji7yf8t57bOUZ4lupi3CdPWvpxq7SSjrxCkZtSn7te
7/ly+ah2kTBTAUUt2dxJb1ebBtdm4FNw9Miw0Or5zz7xqUyrmIfmSZBuZRbAJ1xDEKAkGKqa6pi2
yOsrPmclW7UC0OPK2mQm7dqGSannsPZCsKFibkJpygDHaUtQ51Qro+LhDKDkb+O197anAeAXLKRW
MWiMT9OP0hA/QcPJ+JMQwQoajymm15peweRIgEyfZNB/LqFIBzMymPEQ+lWokCzoVqYvNVN1STN3
sbGdyzLyqGXAwWjvjQ9AJOmkuPNhcUnvyThZO7p5wuafDJ833Psd5rT6RkA9MmMYKeMZnvw+3CUs
n1nu+mbxbCQvcRNT2QAW8ANGP8axNBe7FyJ/9zfoOSjNcfPNptTDkQshKsNgXUt1Gr4YM1dgc0cW
cSNXRWHVDILWA1oR/BsaNAqOnqyjtEwN/nrerlzw+/wDIo/dXH5vixsueEq+8afYNSXlkyGUEhu/
ErHEaxBvIlXU09vRFjeHbGe40kjLpAvYaZADFYF7E+tmyG6Al6aU20vwGcMvbCFVPPldd3WBfVg9
JBg2vEdgLeP2hnp8WrJ5CHJ0ZJyOokDTlaV/4L3M6h0SqyXlYUHVaEe5lzcJC75aDPGathlBv/xQ
8NCSBalzE9CvO/AIqueIOJ6RFmWq4OFSHNz/bSdMgRDvsrT0KGHqywrsAjic5GnGYFcthJl9+hwC
c5+VHz/vSFz+GLcKM/TaAYTj9alR98deGcPq5Myl4AmPBAEK4fT10KecUu1UpR9MYZNXNlwy1AuL
7bD9a1Obudw6Uy2dFiLB3j7QzagH7/BBzCH4zAlHg58l1+xsLjghaSDJ9JYlmOn8r+UpbqUlOzv9
uwpL5gEmvSyTiWo61VQdliUPR3VbK3ezew4lTfR+hLkGbyPZMGWm6cvv9ZKV6XJMktEsEcm1t8TR
e0oKLxZC+P/zEN7SAevvDSIwmVDc5agw/4IE3zSmoCg+Ak+/+FiHhNfCs41R3uhjQKW11+pG/GRR
VcnRUTdTu2cTdhtj0ZjMfKvrSVgx2hGgRnO8R4K92zQgUffjsNwwppWmLzue056LNBb74yJHXEYI
m1S6XpdwmdyBqukXD9mZJzqOfGWB/K89bOgt06u1mlt9hWZhieck914rZSFpMBLbMLeRgBLTapS/
W4QKZBAW83xluXfJz34Pkue4ByikPs2Q1vzsPP7UegN9QwqsUai61vCrKkFP8RpPXroU16lTsfN1
6K/F5fTcwLEkB72q3fgAE+YSSmrQUfYjVY1ISAiVZQ7HyYRcz+0AOOlROF0fELxS9Jbl8IJZoJQK
bppkL8oRNsMmTh27byAdOMb/CcT51NVZmlm8lvPnCgNIJYepJW/uAWRLezWXmJHlqBtu6NZ6fMV+
30OOCJ3jNyLQ4Hf14aB3eAT8f01a3hgD09nl0osATO4JQemFeHkLwxyIlDhFK+BBTdd0SjmwROXY
dOwfh4UuKBoLca4JC0JcWJ9qds3jaRu4y257bRDI0psWcfna7pSJoddUnnaApI2J9WOBnIZo+YrD
/eC/PT8iZO4fDxy+74KJsgEkS7qCYWb7UXyVzg32wzz5TRB/ttl8f+VRrwgFpu0CTxHr330lDm2R
tl4j6z2fQJEMQAaPlStSaYCl/yyjihtgs6gtrjVzy1wIZHnVlgShfM4EnZDtqXV621W0cM8P1daj
CyI4ep7n/ky9rDL1v1PkeLFVwGw17nTnVux41tCBZYorROUmwwqh6ugYIzk6XaK8SRNfJ04ng8ux
Oy1QhWpggWFvXme+WMLgI+U+X2M/Mu0icazsRZFp02mn//6o4Kp3/6s557mE+bvCCEeACBIRLUW1
KSLRqcdF/nRzcD9oBRzpkzjslmtszfhgLwXh8v4ZeTLJN8q/NAId0FIUjLSmVH30czeZSjsBBgI5
gaO1qcpwxVWuWmsoec3UlaFP8BxN8SfJ/PGmE/qmVgfGRhXZp8D+8p0yUghn1mq2EMeHkEWSCKwZ
CQlIa6NtWLUhTYmCIsDFYDSMzvTWOBS8ammSkrVceS1f40GYPDCG23lqSk1QpwsQ3YRNToc4/i8v
kD/vrxintJ5Y5mSHX/78ehPLq1TzYofjJjrQ/bypX/xSyJgGt/BPhF9bRDfG1hVCZNEegoOh3caM
LkanPbf8A12owt5wUmT8xPCwjKgyA+ZVKx1BqPV98CaeD/8DlUJevp4Vbxld/j5OpXgBuSffsSC1
YdHnRNU+HhFxdUxjEDBK4TjbKX+jZXMdPCAWmeGjjqdkaWuSzOX363IS8tYEOza1cSfBQKDhIZ7Z
PDYtnZfRmEEcZ8euGnG6jMMtYDN9bWuE8gnFtfjD/81QOUaHJMis5NJfIBwaoPMMoaPK9BPgkd3E
6kuE7KUzRWD+jkF+ylhW7kiOqvDj/76pITUPOjUYWinJp7og9uws3+YPvj9Rq9Kqr+qzGLpoZxC7
2xys+QunBh+sfcZkzHppRuoytf1DnRwKg9zU+BUmZx06aqzcyFZk8zjFVxeuZdFA8wVTQDWm1QHU
7dAd/jrADD0GKPbQBUO6jfkPdc/uONbo9yxne7yYu/nDbCclWeKRIZpnCZ4ltRWzXRAAR03LDqtv
KB/uo/LrYjUy7PybNOYB9x3LAYMmopp9clWj34EfCXe1n0C7DvelLDp8/zBT4wAKjuDd8xRd5VKB
EGKqBicMRE66iMuiEOsqIrPVMCrvHaDibaoWIuPjOIbnbkI4GAnHCB871UDaW/XdKEJzVn1bTALD
YXUzdxuNh9wmYEV/gEaBlsc0l3Cm4gDJR+wnXPgCc89m9lR03ZAX/rRgzoYi1a8I/WimyRTUxnNK
tXYRD3MLuAAeLqOab8gzl/okICt7Uuvl948IdDnkvm6xLgNWXfs9p9qKU2oBKd8ieX7wWqZ6kxGH
n+ydSpHh2xFHnSFot6HtQANG0kWDLyjJW9GJIHfgLrEHgI3s6wOURS7gdMTN2iXaf0wBeIn+gZsB
sPriMhCtKxCquHQO+uQ37VIezNV5n0q29pNwPIlLEbQyxZp+Jxj2BXycWfVVm1oQM8FWNH13eMIJ
vGMuoakRIHaXDMlxrkeixVZDhYVuZau0V4wKG0niFKW4wGmeP4SosQV4yU4xEjCKszeZkcxofkCP
uU7vhoBzHg3ydEme5sXEec7DJ7SBP2YmdgyJukHji//+dTxSHhcjAcmQ8G2nHcXIikLfEuLZqgua
aDSIl5BcWW+vAkh4QK8u+k/EMgYJ+S8XEtHFbngMq3AF1am0oQT9v8k5CGT/CqVyAb+r5C+nQMGh
tPblkGZm3w4TztomX/mUgsTKB72jyUAFxdz+8Gh4laE/RnSJT05O2nJVJZmjQJX9LVU24Nse/YrX
2dd+9fNMB3PDGbMZE4wkluIlzOsjBpKU677amYl9/+/QZjvGi7Ucj1LybQKtSxNDmHoaJ9+TPHS4
rnuAfegAUBqFieIcaGASM2/Qoq47Zgr0WpjzAOS37JwdT7oJpEzMuG74X22PdFQGinTLgXaNwh8f
ohWCpOq+rNKTvlem4gwnSAhT0RpV+Kvw9yJ++TtOqfG1jTYo4nJAAhE1b6yTEE2rySHuYV51zJCt
+hQbJTIMFAd1VHNabnDzsoyR6HKMLLbLWC4q/Y9tk28VV8GZPmttbXzquzyJxaXL1gBnSePbdN3h
hngCWMX8sWysV7XLiLekGV6dGZ1pBaQTjRxZVQ9jUqtCRNTfdhNP7t3I9hxnsXJM1w5Z7vmSrGlu
uZ6kcMMZ6S4ybF/Zh8Tsi56H/iVKPK2GhIDQZWQZ3dwn++yj+aGy0goDJvK5rbJl1zv8b98yn1L/
4YLyrVJErvsmDv2ssNnaufwZ6nY0a8XN0XvX16VfHRSEgRvo9HgE4cvA/A81zvRPNvop8DAlVopL
5G5hhaAO5BbYA2ZDuPV+22s3Ukk7Ue6WJynr8CK4/pTd7r043rYrE0kxNMPIDOspaAaEC5HNXfnQ
xEI2f0ExvgIq0h33tWUjIOuVPnyfD/RAnpUh6j9H4iS5ylSBXGap+ujY8v7dPbF7IzFrbhpj/npm
j9MY6q+Tw5WCkrKRzn9U0uXIjjIfxKb+la/04SCEdgZFy/J/qnFTfH0nTzzPdF2RmqbIjel9cVKX
MpMqSKGIAf/oqivakkIJvTMxTuoQmbiv5DskTecr0mmB0DAvE33FFaBYdoGha7Y9zk9jc/fJAg2S
NJ4ZCWr+CIGgVFxaSyd6NaoGJBXh29W2CoMpLCrEBBf7aIhKUb/qLOZfpYtEi1caxukBCRA6+bmF
EPyrnJ5CsdqyGWTxbT5blEsnbildPhlRAvAE/zHWy9r2LpK+T9ILKuv6zvidKr+y9qY/HRzeWHyZ
+/b22t8H+vCrHzNyDxyOXdnWWINaHgog4pcdo8ySgoWWZQNaUZ4jg6LK9VixxOxGI1YW49whfXtl
nifRiwYWcg42pOmNW4lq4o/zEz/7BgtCvHb6QWg6JPcKZRuDm5b8kP0iXqS6mti+9Kca43c7bQUF
YBTOTfFSqkefXXBUw15pPoCk+Yh6mJf2xCiyrI9998cgiiqjJ2aDTDFTEEa8VCXEAlXiq3Do+nwL
VQjcBgNtvhP/bCOvBvS3CxiwukqHqmV3M1R4H2YsUl3WbF2obTZR+6zdegwUij9lUwDWPkcCdnp5
8EmHAdXtIcSWKl2XExllg1yFKaU0BjEfzTP/XPEIrAg0lni5ZUsXZ1DfPJfsSoHF5Iun3MFN0cEm
JoYgMyIbhjdkKJumzggP02TFEbNovUOpUugw6Er6UUg7kB7Ge1p6JGgbfEI9FDsHVFJHhN57Qwa6
rPsRUMpmnIxT3TR0unhYASDQFWuS3rHbIaUMYcVg3HvKW4FsH4kdri7eleyPazqC5b3Y3+xyxADH
uIccvezPWGkdUwUHqv3skhWlL0e7vg/fXbD6OGusvQXsrC319vdbKKveOi4DA40sQ3ExqX8zhcDK
tskeX/fKm93yopg4bAxmRpdLmdGZjzNVwhxtuiNrMth+6H0AQP4QYqzOrGnnf7d1GTl9I3T5ivrK
jxch13nhr4NiH89ojECVBfVw/M3gx1qOHBx9g5Bb4ikn6Mp/343pXSVnoo9WLOmjPrRb7EuckTZD
i49CnSzraKqX5tFiRk1MlOqWJnlx6Bq4oaktF6GJSiJKj85HFZCwFOrKBLqG7dpJ+AlQKBYZaB+u
/6+P388tzSFcieWPX5PB2n1wMZYd6+c4HqyhPpRYt4uOUOzHxJ8fEWV/8v8Zeym8uRQwioLCAxa5
PiLI3ibpu4yPMWfRSoy3oJ/YAu8ShlG0CvFJsY4aJRMAN9JZdPQD16W5UPbi0Ut+6e4GwGGM5usM
askE9Cjo9e8OF8+E04ePowaGXnFM0FDDC9u46zSycMLZ3/zO1Wd8Ci6FhumV/WakT4xa6AnVzX6K
ZLjxlh2FefCW2GJe8lsRGhbOLqfrl5DT2Bb21rOrh2RGg7EwucXzNbXDi9Ds2RZXvVAo4MTZtJEQ
a7AOe9FsDWZmi7b/8F+sDzzr2nXrWNfYgiOu2gnuLGRz5kmG/vS6nZE0vfMBZdudRZsKBp43fEcq
bbfP6X21M6mg+F8Ri1+3yea1V1Ux8hzCKt4DqlgaCQOZr3jrIWSnCYpV+mmc8Exc2JYGMzalxFuS
hE05yEo2MyY2v74695ZByKHY2iGOehZA3q/Hajgf48mhI3QP3oG3w5O5wtU/pGuf3i4HjvDuLsRG
o07oSO2W1r7dbSOxGgr8QTBOvTJg2shpqCZ+5VzEDzryZ85Qz/BAYhK9uJAxQuNYgNTXG0Lq+myk
O38GJ3Fa0xvVVM48t66d3UyuR4NQm/iyDnIM55yXe6INEeEiWMoBGFMi7yJZ2UUNWGK6f/z8UNNP
+3eRksXdLXwRgtFa6n5pe4n8+3pXGMCOnnZBcmLRzMmqtmGRKymEIotHrB0jLohBskswXGb5ALtQ
7FLoGc2DEfFsxJnttSKMGyLscEeJnutZhNNjO534E5FezToPfxsKI2urNyEcIIf8imZsohdOKyZx
p+rW70PnItvNFvjum+OZzcT8N0z+0hLerTQSasyvjnPKN5xSVpl0R99Zki2hJ6Xw4DV3T6Gl+T7+
mejzHhhv24GstbjgxEVIK2OU41ioGFGH2F18SV0Jtx0nPyEXCMmJefwP58ub75kX0c/7egtN5ED0
hAGpsF82Uf0pjAF3hlKf/17Qw2MwKFOyFNmjlGfVRNbKlRfMHYmDNpwlW8rWcOep+bhLQTW4fS5+
fzbi/hOh9UX4d1GYwL/OKdgvSSIqgunStMJRhUz18risf6mAGPEimuqq1JqSRBVPjdBZvHFF1iEq
nmYBC5TScQd7Y8+wC/QRe3uDJV9EPXmDwT93K01Q5UFbjjS2kuaERib3V81zLITvHr+e91wvC5sy
2e1oKqGD9p8ns5VNlM814Y9Jxn/RjbZeiWl8WTRNCZXpb7sRh9P6WEc3NSilBRA1o5sQOMWxNmj0
GwM7FNXOqijVAKW0FHNpiHybIDgdm+vQWFBBIoSGiCPw/l771A20s0m8hUkywtCeWXrj1h2ZER89
1MP7qC8ebKPYrJv6Fk+HL4PZ8bUup6E0klMtEITqCIavFO3sOMy+GWXsH9ITSDCNbYIY9bprdIEw
me119Lql7b+Q2XVZ3EDC+GP66fuoxu8HbrJ8NV6uY+CU3nK6K7xr4s8A7QNcsB59qyD0Y2Y6B54X
vvYYF/1kxkpn/oC0PA0E+b9bNN60IQN8wrr9+tdVQlgkCsMwCZrOW6UzDD4uZt1j/Fmc4fiOtheA
1jxlvUUNaShKWrYe39KSbjORxvP2sIf709OvPbPL7yih1lKLLvpwvVN7E7WlMTFPDtHEd7JwhXvj
qF9lUZ40dwC7+V568cOJ+chXnHZGhQJM0lB+8Iz6NLmh13e+Jih1jI3l9b+Fzu2IpcvOT9oG6idm
gc742VgOSiBRuwENJhWzquA/jHUUm8IFJeJX4pkLkgYTEq7YAGX7VR6+LAmYc2KPYI2s8CxM6+At
4crtn54rlbEroVROmVsIRFSI/ui8B1zxnI0z+kYzfKw0EEBbWWw6N3NbzxsVHVbPPIqhzOPHm0Sb
VkOktNF/EZ1tfd2qYPcTuMuyle5eYM8QaAjpVky6ACk9Mzqhi5qPD2GXDEqaDH3vK0HucQpuko53
AyZuDy5Tvg7iPPKb8iVg16Mmjsp8+UzUhNux3oz3WTbXtDNxBISYMgvsTi+8vtB7YLy7V98WmSch
CKlyEf6ZC/2LVrzKoWCxk8EtH16uX12P9fDjI+1yhWoqSSGXhduEOQtQJLb4UAWCkx76HCsg3Vli
NogkRzD9hARpG4ZFw0aTDxv+8Fc60e4aP5eotNf6kgkBVXTwfJaoPvABNwUaJ73cL/wkXCku+nhZ
4JXuqsTp20GF8ueZXtmasUE7mREWtuSX/iise+0/uQrjixFz0oJzUkA8Q+0gbB7GrrN2ZU+8Xsmz
3KixZa09Xwi/XOxH/jcXfRq/cpUgVoKJqs8Yo1RHaDvagvhjefEW/TIgpyFAdDKiTkwvCs0nUa+2
leK/Gy4cVi23ueTj8OVAlYQvvRKQVJtC+BgL4bje/zH9w/dZoe/c5xFZ0Eh+/+8dsH9fYXhNT78D
enRMonF0uOyWIlpjy48oJhG2J+0Yfs6+NIaX2kO1DsBRjSOuuhMAuQt/KipIImiqUoz6QrXBBUiR
xE5IzWmKmt7aipadgdI9+VKjCYqB3SC78wOAM/82LeR8o/6mobVIAqB0rK66jVxcAxkRGR8LuwTj
Cnq9S1KDn7MMEXmtHtwzmcUCqXqE02KVqUEIPiFoDIwRvayv/2PF5QDeBZGXA1X9M1jaGp/s9f4H
Lu4n3wYpY1rFgmZaWtl1MAq3i/mv1lFc+JH1PeLDvzRML35CC7i4QU88ZwRZS/wgFlXPt4wHJcYp
aodQLuFn7y8LFaDzyvwLHuAxdO0svj2n0pEU8C9HM8AkBq0y9JyRhFJJFUAtWn38uJHpxk0rQyO7
pFFzHituwLjsWdH4y4qnStLpHE/rvllNLEL+cu1KSHlK5GteiYh6zbPni3iPOHCWcc6TzUkT4A2C
zPVSUVW6eRTgzKcmAH0E4eTS2qCfCT7QQV0sWXoci6idaJjCiGiqU5D8SKD447R1f+INQ1heokN+
z589wR3l1XRifxwBbQxkUnCLqNYxIzoVABAr1mwv4g8+ZJIUifCnpVTOOxIqSJMmYrvOjs8ftLV+
DwsmCA4aIlWlupGuQ13USBQbydARDH9kjcwPmc4rJqQ7S8QtROfzgAq4p4ipfup2rKVeZtr0mv4/
gbMhZ99a/7kvwjGK2YgL+fZqXlRDZmwmswq39gPPLsm05ywcz3dmXmPnJe6DeXnefWmzphmIsm0k
UujUQ5mNF1hdv/BErgMah47DH0hm/mvr/i6SJfKrDi+5pO+LrOBp8HDNGwz0KDqczQZZk/CQBa3M
SaJAFr6q1cZS5vcH00ljO7S2TpI29yZrFfretJlDdJdlJj/8wf85Rs6Ce8Vv80vQ1v61TC1/MInF
0Kqu2cIfOXbeBWTlmov6fU7Qkh8qFObStHqq0gIAe8/ulk1pJlz27m7shoakhK31LsHuvZ2inCo0
yFDWfoGAxHaJWKcwrT6r9TvECpr7NjrRityKqvZuu5H6HPA4N/3E8YMQi/RBatjm/x0Q+fajWLWz
IcVb4GKLgeosOdUDK6nWaxJaA1S2hsUnGYsfySF3aAfhX//eyI//errBisk8p0KBalTCL5bvM8LE
5dz79d8qV8tvkSSqy8BmzUDsP2fDxJRbqvK71dqUJY+xRWJhxYT/uZY46pinuO1VzHjEdsLwMnoP
Cg1FdKdEhIj9oP1mzeF/f+EEseL8SwR4lt+MrBwMmuHXY2GzNyM2xntAZV83V7hJGmx2VL7qvNbQ
Eh2vqezs/4G9bwuTXbDI43Y5yo24SW7adXWfVAOPR9Ks/eXUEJlGo/FeDQKmGAexi+xpSyU8nud8
JvNM7MO30zLz8WNDcJwfA6ORHAug6apoh0e4YNp2hklb6DQHGwVPoKmU+/ZNqwibPTVh6rZlTEHU
oGc5Vz+LXyRN3gU39Z7pzOjGld/98o0ciEjE68rThBAD6Rzw93xdxvZxZ4Eg7vQUMDasENaofFDd
TuQk8a5D1ypGtyjupbFTgrm17Kjk431Xin9CWTOCloNDDp9qAHuNYmbSQ9rXCSBtkFrH/KZRI93O
wljBkC/EVYOgUP0h3Vxte+pLZM+MTuQSREUYMoAj6T1IPyYcQtrF8nggkGt8YYjRU8k6LB7k2xj+
nI+lFfbC5JkfEcBe5t2ZYHSnPllJKErcsGyRJbKEj/ag327TW1Iszw/pn2YEtC1jZD7BVC2lpLuB
+WWFY+6v9ekTEAwvIn4Ll9NEEIF9bR5UZ28A4nL1bZiyN2FuohbF5RIqbUcm6Jiufd+TREsXCvLM
BZDpF9Z7i/eGIb6YH3XAXNEGMspYv5QLi0+sE058a2mO3UPKqec24iV+EQnQCuCnl8WqDnrCfJbI
Kuihre/OAl52uTosfuioSt00AHAF7nFmzV4b1bnxbUTU8az0BIyF1ixovP+GcjlUV/CkKg87bV5H
ukcualdjd54c5vr2VjtyPXbtq1UCqg8Hf8muCzaAPNAXDSkHDcrR8IKo3dlhQd2hrDyaUHQpfFIs
2jbPEGiVNDCCjH6Hb+hPqAuPjFngvwqITy6DBQfMDQMsc1iyhNd48LCOBKv6VXpMQjDTg2BtkuiE
+gAeaK8u0ufooaJhZZ7OhNmLDDnHD/xZ6okaVwL5YlW4PoMykghtUW5TiytpTGCSx/pVu9OvkwGb
9RFjukQEK5IIpQd/MgOokvVPLCOgO2BcCrAFlqska3VKSQd6WR8Hkuz2LkEMBTKIWYrsqAT9KTSh
TLBh1f7Ph7r7+rkzTxoyIVVgzqupDKwK62jyqBFPJ56x3+TV3tzFqiXjTO6eoB5FkRrJ2yWfW6o0
1wfb4OHVDny7CJ7HtaMc6Te2wuUJ14B68YQtgu3QlFMp5XKVQyUluwIhSmSidzJX4Ur2VZm+lV3a
c1dDUGuQYklNxX/hhvJznRIRL51AtOnodngvAgRRl+6pK+D8dQ78ofo6d0mXIRYYMye5zT3DI2+n
atuTIm9d22hyU54DQUM2zYs/G861AgUpIWMK/EER2RZTj0EitG39dn7uegMepVYqaNhmLfNdiH0s
Yab0nCCnJk5TwFw9qEUVPs17P+EyM28gMD7F0FHsBXjYwmCIHdFK9wvmgdKghnUNWd4+U0LbCcWe
eIG/PDnpbvZ3QYcez2PCXuFIUSGXtJ//t37cNOmiYTrJ1KD6xEFN3jYyMZoZlQ8z99V/WF52Aaku
JbPqgN+JDaYKaW3Ooydf6C6nO3TEyu3nZjBS45w/fC+KyXMR2fHUQJcOBukds+70i2oMZibzpJmp
uEU0abJ8Yf28G37nQLXvE1t7O8kt8pomLxg5rul+87mmYynQuDjZf/R2rmgYX2FPND2n6qVY7ytP
fVVWdAmwgUhBEudN/NJBk8mun0lJJXn/HAamv5elitccaOp5Ss8AtGC9GVYOdovGhgytbBVBunXa
iBK23wGS+x/u6ReTv0552GJBEVzsAn7ZhV5IdBp5yiOK5U05fSHgbqGpb5Aya+LSFNNLL2NzhFPb
045vtuEfJuh5Luxe+/ZENiQ0eiqty8diUrAopegfRDpdtYlAdaFlIrmhCW4mmBA7NESfn2/rz0g7
ixzzbfzfmNId4PP9W6rzH5dZwVezgI+94U+lnZCNcxC+OfqD7fNg3AojPbTVg5xHhzXV4Wwp6lDl
k0qB+VWTaidIfmLaMsrGlSHN28lNmzjJWQoYucx/rdi4WW7xFtWrlN0n0bPXfaLs43OoXUWVLGbO
4buAH4Y9ik0NsNYxpwVMNx8kZuFrcCgSVFECdS/COrS6nRWwVLuN3m12/tg1H4Xy8dNsdcPbOtZG
tsRE1S4P8oToety2ZqYMSbKqK9hHxrBg0nQjIEDz7zZy0n/e7PW7081evUSuhCbCm5tZBwR0QIgI
f6iEeWc3ASjxClNkjwbNu3+ERMCBVDOKEkiMhND6zPgdrGIxzrJotFD/b09J1bSqLjfN6QpAMUZj
D/HyBOywmu8vPt4KKlW8Ai1SqvBHxyIxU4P0I4BH79JmtPH0fYphsPj+B+L4QaeqVq3s9KW2vycn
IiwzMgu4gYkReKzWcunQzjNQUJztMGhYswx6MCpuaqFSx8g6zFJaBjLsz9n0l2OEWxPY5XKkMs1s
muIuUK53PwEn8CJDDv1FU9N/23v2CkVQjmHk2VehbKK4bmVJTZsJ7Ypr5wZ654MzTVW45cagGuQi
yNirqbsSsiPhLT5N5wXlO+ca6yS6kS3g8zTXJu4sD8vNkf2mR/Uk6QK6GSJFoKTecJpOiQHZbfVe
zY9ct6G6kK6oM0YoLfpjp5QIeQA+wol9PcqS521avQ6JXuPFcrEMQ5icZfKvTPUWfQhJHylzDqL/
IKSOv8yf+uyy0KbzKoKqQWHVezeBCWeTmK4N+/jf+iGvCGyZEfsBasXqLdGgNCCcA9lICfrYRmsZ
s9WE4lG1GB2pRI9hQ44CoDQZ3RwQtJeDSMdFFE5PJchXZIn1gCR4mMozYpfUFO4IU12xre/k0hFv
Wi6PegHRx7Ivn58ffHcIySJORiqG6WwhSiSLj41L+LuaC2o5Gab3O+PRwy7Qp8hvZKRWB9IHyU0Q
FTs+RrRt8LFFMDLR1LcPxA1roVZgACE9EoqMx8maKsN0binhzM/NMrWaUXf0UFmA998z273d4NdZ
r660aR4eoJ72yQfr1+2r+1+EC5KheqvNEQ77OIqBsTYfYOxWIPHdgXpIRD4wLWXcyWOcHeqSZ7rk
e2Oa531wFRB49vK6QTJ2VMV+omIuDUZjJybYvLOb4RpakRxaMGwSDy5pZqfnqpwQ8FGoU2LdC6k4
8j5+cM/lthK1G45W1fAqSjxwVLoAkkFBf/I823Ta2g6Kf36LWiivW2ZN85PFpuin4DsAni5cpo+S
PxXF6DJqLfld31OmynfbT3XdSZdaUs54u+xNn+UddRfWO0IYf1f5mE/JN9FSjfl3LLRyAg534ZvO
V6XFikiAZpX7IlONGWUMsscxwM5qhGNE1Kbu7JmcI3rmP3C4l4Oj4t9AfSrR03UG1snASo6GrpKU
Dq5snXB2wRuMIs/B5eAYREGAIdU3sF7TcWd7KF9YmE8F/c9k49uI2pzZsNALeBGZzrftHpBh9CIg
Qc83bZHoZth0KQPAqjMlmkI1wdMwxudeRAEvWWABJB/FFSL2Jvzt1VB8mtDftvnN0eZGnoaCAOTB
C9wsDy+lZAVGYcLcZpDu/AIz3H/PPF64bdntY3eLXlYuGCN3/2UFF0+HI/NAy8prb5PjPjPrDtMT
vnUnXYK3QWAszOqPIuDdz8eeCZzzmnyDW5/3Xe5hS/3YgjKutBqv/YxMTun1aEig5TEXzB4q0eaF
2HoE7TwsQzoi+WT8CKFFKYrkMOm0XI3q1SlGU+8pGTDE/eoRP4AHDK6eBjwFjEbYq0r6mrOHG+z0
ffRD7BMukHKsuIaeWmjnlMjGIHSuUUo0pFKDUZNaCbwvPjtuIo4WlW91G0o3T3SkSZCEmCwmjrt4
IiOCowywvFgPpV5vAbebfKlyQSYjxopgkBtOpLkrA3M04Rlg/1GO2onJjFngwfN57f3qK8XBI0UW
KrOG3Og2XuOIxIKk00dJdPscX7MpnoVTBiR6Af1dXR/W2i3f8BU6kLTmeL0/SbGPjn4XNxH2W3Uj
gBiygHXVmMC/iLT8+Ogeh3DXfVcGqa3KK3Lf4RQmR2c82PLiQv+/dt8GWUBeRC8zVW+dePQ4uoVy
RXDk1HowamGMP5zqMA8NSYQWzPEugze/1Tmc8I2eDP8qTFMQzC6no51Wu1L1Wn1JPp+k1jijozBw
ZFFxLcgxidYAN7yT0btVBPhs+vwKEEFpMxwt5Ehxy8zMgN0xfjGNgm9m3QAOOAG0YMTNvih8rqsb
JYTDuIAMaJUV46kQVds+57/L4/k4DMYeiIMniTaVbzIbAE5C6BpY3Ig/RtYhQOKkuA2mpdGJH6Ka
Tj+OY0gRne8gPMpxho4XK4iKGPWgwHk2iVXxAf9LEAq7a4CdvFBJTpEA+u36B+HZT5/8RMNZJvLy
csu2xJ0UbvMzaYNKDlHpKdpuTX4dF+fIB4d1bEH1B6XWzKod1aO8xP9Q07UNLjJU/1+8Gw7BQ4+7
1NMWXXY9EcnqhRSKpd2X95swoq6J5UYcta0hz2LPvT1V2ZBNIIHjQd8iNKGX5hncx1YNCgJfHV+/
OF4HSNWUmEv71sRIg5spvMi+wO8F+4DuXBMaQjjKBdaNG1QUhTeMtMqj5o/0OrZ2jZt3Avk/bRRx
X6hvy4g5T5cxcZaTy3Yw/vtBnASAkwt17ivV5t/CQ8m0UAsvDWRQxnAGmLSt1g6fMb5WHdIeEBwv
80tEMwWEJuf3tuQXPhNW+I/HAe0Zy92f2j3abNo+X+qnBJgSB4mPypAIzZ78HsFDNgDmXBROD+lj
6xFInw83pO8dd/G1LfrzzaUN3Vii8PMUSPzKG4OM5ymWGtQQ43+bNe5NadPtMXEXJtt7pelnmg9M
nOkJKm6OvTUvfUrUkuSrlSWyBtr8X5xAuhaTLAYB7n5DirOUTssJnUiYa7UduW9X8DG8PY6fEi9o
M9clEocXAlB0rU6+008h1gAKcLqYdei5WlzSWiSf8+t6PYVyVZQZLbsZY2Cw7v9K5yc+ntYa9Mjx
duipmuTbRhEbNh214tin6wfDxLBujCtk/DM6/bT6+h6S8Znzr13fOMOhV3kIwJe5YhsAeL1nBfK/
0gG27MUUR+LzIIjsiqCSaXn6paq07s4YdUFPdoeub7XXNF2VIj998x3vormq1BzeI8KIR2TOLisx
bHmuRq2scu3raFp33PZNXzIj6befbgIlDag1gnVfX1U8PatQeq3vGFHKrzpCTuX9/XDAdkmWCvN6
1kN1GB25clcJr5wz4Fy73ELPWkQPEieFQ7zv1Yrr1Cizi6ROajRd2ksQQwDKyMgYMS6TjDbuiEGE
NZTh+kgXcRFN8lVfIh2Rv4Zfz/42SJxcspECkm9TN257zed97pKP7WwWQ21nRRIwackGwdorO/ET
AT/hnJ1zcrjEwW4lvK+CToXU1sMzt7fLOu7Rs/ADW6qbj7D0QxT6Fa4JVbAaodfvZW5EbTMsw8lD
tY9iLJzBEDVOVl5qkcnMNw5ysiGx47zeJ2JtapVB5ocUamnlIsBShgBLiCm/uhH+Y1YGdSs6rdoa
PH/8whSHT+vsrJ944cf57TgSiCeHPEGgX4JNQEdM5bU+RXnAjhqvx3wTnvqT6r/OyVtWjdIdrZ8m
aGqIE/kGeVJ77t+CjAyPqeCELPiDky1s3Xq2EqmPO3lMHH7owzDp0pd9H6jbQwk6bNIpzPz+Zjwa
HdEe6Ht/H45ALgUacAYjVQ4KiBhjMraEVGuNSg7fW4T+g/jla59jDSQYyK70Ia7ILKP9Pla+TZfy
FTl1jJIHnR6xLKJfM2c7phFo5cnfH2tdb/ZzxhB0QYDrIZwMnaivcBXVmACKRsdt2Ghdu8Wbg9ig
QnbBudo8tCpiHMXj7HZRSbd/beOh4hvxYuZH7AfvlHEMJihwdNgmDZ/fdgxpo69maOZE4bv0lbct
91AVQAtmQ3IAiOvZMVT3Jdff76+rJCyEnZdiGZy1+389lGA89yMHE6+bOWynGNix+EC6FYKY8HvJ
YCZhWeq+zUT1FJ3vn/XCtLK44HFy8VrKZSc/V4i6OZTSuyYleEZdYvRiKMjpY6m9HMPuEDT4iK72
0GO8mYIq7d4YSGrXOmisOwSimceNHvfbS01cCE/+mzta8mQSgmZWoD889gQfOu0Ku4n0eYThaTt5
mQ8eQW7AC8ndlKwy7xn7EJ3DHF+pTd5tWfom24bQ5sdJ/b3vyHaN9S/w4nQPgHefgtTXe5O827X5
XlOE17xasN2+/RR76tv2BHQeRFHo83rUk+JXKmQns1ZiYLxTgPWM3S8MYhz1sSzdWr/4ooy3Rhs9
2ZxEghg2ThsDdm8imiyut9Rsn6FspKJz1x7dWSqnrUjEjL7bQu1IQ1xTveoya8fAa6MZTKZdLl/N
GXPLRaaSbcTigEM/uujGfmqqR7llDleOXRw0xQmu3T4M9GUExDzKLKXacQsKBzXZx+efgc2TL5Tx
rEVQehfPWMFdjTK2eF1hY08wF3uCZqBjHghG2OluZsuYRR+FBil48xZ7Q6ZMPaJr7ZrDtH5hSdCf
FT7/pjcpBAKlK/2Tgfc2huGblgGBe2DO9DfzfwocUJPz0HrNHq88CIqBnlwxUzrMAZQYjujvMzBQ
pzNbuOsEwLW9me1vzFSR/qXhuj0ZU5NnAKtzBMoC0WRNuz9RaeIPgJZRC7SJxHwW9wuBJoXTfqMr
1xIDIUw1le3qtaS9jN0vOpCbQw/JnV55Z1/syLartyfYqfqVa9JkYgWBSiM5eW9mNgKeCrqLMVqs
L4byFksZw/sKgRZHvqsYdMFyh/0WZvp7w1L9M3OpVts4VeqoAVqq/9E3z/gOiu8wJopKpYGmkf2R
4Jj7XiG0Fci7ZxS2fpfyKKksWULj/qOfjmno4R3L6aHQDuHTZerZIdvasRq3Xk+mcCozYvloRKw6
spCfiptvClpR2s1tvDTv8fVnY0wwn4L17O14qf4YtY120rMtAtvAZX4lLziLSENy16MlR4O/i0/d
KLJsrovs1NAii0YicXABz4Bl/IkbQDGjF5fMf/yxC5nPnosWLgzg9y9zCDS6Cy+77W5erod6bZ/F
Lz5PagWuBT125QjsXxuw9wZ6BCtzOPkP38m0EdhxXgWeqsOh5bNxVdNqQXAC20wOso9QmThohQfp
ykeaZ/t18j9He1xfPdxV1mvjdOgl3j59GqCzioyi4OrfunhItwCo2rjK5kmIMtiqM/uojrytIQqz
HeB9JIkc3aJq34lCrQTm5ddKnOXe4NZcx5eDQ17TzNckgKyL3T5JoXn4VgX/vKiyUBGsYChorTGC
PgO6q1wnGFqVgI/3HvvlKInkiBhvLm51pileokovTz80L4nWliPnngQKAcKkcmo6gTGM4yuFbiy2
uqGmW1l8IrJ15gmsQ63pXoWY25/9OCkL+Bd3QL30e0k79SWBsbyuCV+2KC8Br5T8HXpD3+wK77mu
JZi7Oo3oQS1BQ+6tDPtKuy44YOmHsxwiTHQldnGr61xefg/M5ROKsXyQL3dsZRoVtb8WehlG/q02
uzPodve+MeDVGLyAEnfwPXI7lhZ4VAArbhm6ZCq2xX3wpmpcwJqV8N8Ipx8iXr3fukRcBElNc/Dy
UccEQtvfmXkYKuRYzI9d+v1/InNkwzhxmH5HY4ERsXEgonVvu0vvjXBAtoG7i+6aWpczcC58Tktv
fkWY2L1xeV+Q/KLWmNirb4LvD4BmPxhdlshL68xOZZ05RXMYdAAfUsDy76G7YXttifk/l1u0xWot
pEzWnNjCCvLNcbfYw9BwO5IE2oti/eyqLFZyA6buSUBBeW8xhe5m/EhWLXyIylKbWXi7WA/jIB1u
5xtXVmRyxxVl5P0dhNi5PKinTHdVRKffeCklxvKnPV7QEMQK+AMW40ENkhF11uChApdJh/5+td1f
9r9bAFP6PfE/Ay09VfrUNcXb3GhfU7zYiDI0ZN8yQv9S4G4PgROQs4LSi5DiUU0Ynqp8R7nXnzLh
VzKJfwldOjwZdq4m9JSZ02qqkXbHhCA1W8PoxTNGN7AgsW2RoL1YBIuPNlD2ZJnpavGCkfwwak2U
WJilXZwiVHMPXE3E/8Beo+npsDDnf+S8C47PRqgRyzMq45nbENeFpM5pvqU+k/6Ym3y/P9CTBuq6
TufBAPUDHgL0ncAA0yNRuDlsbp5DYEJBwbmwymTF5C4Pzn/5J47pJDD162ltjMMRxPdY2DDjwdBK
VZs9jOyoQ9KyS+GnQ594MCXU9gGPdU4y11y4gJ/cYE3c2n6/I2I8ZH8CdmupLso6q+Dg2tN65zo7
N6JXvHXnUE0bUiuVIaSJ1JT2TbSMplwF1jrKFs/jFyLKJYJdWnawXPX/BLiDWDlDJkyPRu6f+77a
J6iNjP7StV4d4Ux1Uo/qPfQaC7mEI+2Pwc3z3stw+kEhVy6zODfCT/LGsPgg7Z1d8vZQuB9wSS+g
dUZIIllrJlrnrt3id5uIqO/rr1lgQkEob0yvNvl4NxAXNt3Oq3t9Mt82gRzTYiKnrcoG2GqktWwi
4pE9JCl1skdPh/WDaDB4NZ35eJigd1lxYOybWuA2N4L18stvRsA+G/g6zY7KDMBgVrWjx+lhPN/j
gqXEWO24K5Oi/6DXth75aF0Cm4zRDlKOd7/XAjK0o0gmojBle1K6E4jEYJLRmDfzd3UA9p0CTIfw
LWV00y+ebkNIxCgwOdkcKnA7FzrGECvq5sDQIXIbaXhhkUkdfbsH29xceqXhgBXF8MFlTIYPOrLQ
KMBt+Ahz8NLoICZwxyC0QQ1FGPuYu7FDo+I1DHWlaskxlP+E49Y8aKODjiVzmMFm5u65313Jjy1R
XcpcYbUCCIuGdSSHw9wMpES0mWPBcbHE6yOpdbLcfB6TrKFSp0qYCg11MuUhTGkeHaveLvdzqOdi
5z5NI1YHA+jvU0fKrZsmLs8m8w+WO+ORYJmGEntTFWfIJ/8aG5zN6LLUwIiD/aVP0E48xE7QJLUP
sAE0qUS0v9iUoNVsb3a2i7wXyIFvdu0YfW2YWhODwszXcBbWvWHjWTgtiYIOJ1KInH30bcHaemYt
RJJWg+v+R6zg1XI6fLML/twHtdmuqbbH2K96m32YmtEosE9dqyDcrbdlEVowku6kuIvB1qYx1Bxx
9xGalUycO+VTw1gZsKJ/M3YNOn6VDIsmjWfYH/nd3SQxvggQK9OTiUcfQb2I7GvyexQDEAMhTUy/
O/yv/qOc6Hc4gRLrbIuF3/fiMRglDzGe0IdU12GD3vRdqY9pqoJ5PNGQrP03eKRpgb5CjGaHTafw
mMN3I54/qAmEOl4Iwcpu9SD6hskXJuUsg5cBUpvWmQvfMYLruG0ZgQ76ca5VDju2gjrEDG0WXhK4
xECD1eSFuAGjcvxMz1kyy+3ctO0vOBOhzSPRp0M0GmoP+FPLDSRMe5dz+8fF75bMUawVgoiNZutP
gcLh/eNGbA4aChR0WwwREwn/GTP1Z8KaS355jW7+usp8Fv9GZK1PD00sWNIa0Eq/vHHRzspHDdvo
IUKwA6huz9DC++O7dzDkROOarbXcgoLHGdg4XmURxWjOnKh8+9N5uvrx2ed0NUgnGxOgOonoMiLd
nFwvjxa/Tvr5Euc/rdhKAFs4MIS125NHsQbAl0TM2Hcgei4U0Obdjn67TjsCdGtEi3rwDfneXsVv
Jsl40CA91wxngS2Mgdb8ybdxxiqQHiOs8EsGsBjh7cFwrMfeam3mNN3NGRfpT4mobD76zDsXYWa8
IKUjzFul22odJFYfQOqKZYSQt5hPJejd6b1EIwoIxotLyJplaNQoam3gCXtwJckVrw+lg/rapcd6
kza8j8PEJIxSVZmpygRZud3Tn/URgkED1VdByEXiK2hXGNgz6vMF99mW5nUdwdtaewcKYSwoyUmu
DhRP5doyakTVz7ca01Xa1m4ljp2mFvHV/X48r/3xuORLkOzOXMBgICoxFSU8Rfkgyhn6Wu1EZVHy
OWdhMn5FZhK+mMhyl0u60sUuhMdQWTPKyWFIpU/1ofdL5COzSyH5k2tw5TdD+pWzbbHCpO2+K42N
DZ1e66YsydJPOdb/44pN50QOYDEvA1T3E58RA+b+lRn1ArchW6aHIjvXpfLBXA6hFtWY+Srot8Xc
x4aaP5bPFGiFChPP/3SsEbPSzU8YOza5pH4PIq8fwzKriWaxbo40f8d/v9UhUBMhfJtagsDPstTT
qlI2DE092RsBQq5ifhf9tuvMNmor5DF4JqwOmwIv/cpNiItYnbst6synD9SHCNFkkdb7OcnVbqC2
sPfMJhlixrY5Vf97kGDdadYxEyjM8h6DpSGf0KW0EulKVyq/Z1xyeDdU2ObvF4Go8lvgK9PVFWac
PcxCiwSMoy8Ufqo4Q3TtbOHoScFaNRTjrdxDf7mxQX5WgmAQHJ0hfPeFmcEgZFUhMhgYYs8FkxWm
OsEt/9ikLLkibLYjVwszxCDgYh0ameXlXW/MwMKiu7Efwu8fRtWkLRwAek0gVJcJWkeUwS7+YLZq
y7ZyaOHc8EClPfLPfG1Wc8FCMd8U7tkEteP7Kqi6tU7SNOzhpQJLGTwbgPKG0HaGFGtKlL89/8W4
Sao7FsVZs84aVYdPERH4C8DyVD6nZxlX8rJH/6+JIJ8fPXDSxd8K7+qaTn//L8YDmxRRfAKMPiDV
Iy5yDp19tWG3lCFR0EzSZk2r6NAHTPQHIWVKDZ67YX5YYaldh+/m1xdF9ubn1vg+gcfSuOvfiJiD
3o8MHISwwV8HfTeP+a+WAlKxSMMx8WIPGMA34ULqlk1Wcco2/bBLJ7OXY9mzCwOnlQs7ce/MuZl/
IXZva1OFx4c9TejL8aMfcNMlpPoaI3HiLEPIW8zb6sWIEGYeQU9IM4EV4my25n05znc4tCa/GUbG
eufFePoI+bMLQvh4PBQbbDplzqNfuCZxz36PqyI4puOcTyc7hoYCFcIS812yeZTjlBTlYvVGZ5kX
M4g1HXKKwnvq3OpNFd9x/gFO3k0BclmAUvBUlxcFkvE0an+azwxJ3v5CckIPbUyXLvx+IKkk66Q/
aX/WanE6dst3Jw5eL2UI6n1XU+ajkdrH980ot3qI15d3ZcpqFP6DqDynLYw9hlDJKXUv7pbhutaS
XH/9QcEMWOwLopjMiE29EU6bAIQRaBZwBVyrkhR3MrKHMKq4lF9v15zb9Qo7LjG81YvmuH3/D5U4
qxyoSelnoWJeHfJ2OW+JlQhiBTdDvmfS6Y62/n+XTOifWJlfuYGH0pwU98HijZZLDnp0xQY03Hkk
OFv4KZHPVhkvDcEk2vyuPgW7QDnFplpAFrQVyZMiqYC/n/iZ6eOpmpO+Otn61sizlOhSWXteVyUs
qq2zMLkY6PElNRUEoBouyEUBTrjKP3slvPXuZhey9lwAE1ksMMZMy5H61h1z8H4/imBOXDC1MhZB
NnjG+sfwr0Rm1wQ489ppeLGOMQ77/V254H2DKclZqMGqQnYfEEC/v7wTV1grOt7oPW9TKROygWNB
cNHipWj6bPhwInLnhyzeLZZGBZOw4g0FrZBK1RUc3eUsEJd9Plze/qrSGO8H4S4x54I+hvplHA3W
SF+oZmFS0BaGQc0++pYVpcvpOd0UCu6d7shdliYrtquzacUTmRSxygw1RydgvW10th2HnXYVGzSk
rux+eUYNf2O7fbPGx60rFzuYr7Um98+lXQ8MzT6XyT7Bd/m0omAkA9BGCP8LYmlaeWrzRtImJ+Tk
yhFdzGOZzThT5kb1JkslpH0p2yNt3LsiWwuMoUVMk+WTLWnwL1xbixnnRxNsmuaKlq5CyXaQSpM6
GBcKDe4Am3ftineDTP3LVV4/sjRl/JfGoLj1asM/MODI+RB4mwSJdc8gHueqCCTXKX4st6aftoxe
g4IyPDjn6e90blLr0IFQplP2mAG7Ju6FAp14HD9efXlx1hpOEhCvH03gYjEZZRLN1s7vfGSUi9X4
u6MOHLel4kAPvcI51ZFkCWjEcCLq3S74mXpAlytv7To6cijHiXi7heDnYbet2VdD/kxFYMXTLxfL
YQnQxiBM1PwwCYFq1tb6iPhbTvTz9v/14o6YCkBgUN00xX8kE9lP3caZMlwb8+6Ftnsa5mjgD1YC
0l/E7ClfIaNzJ3sUwrD+kv34nQkJ6XQuADwTOZpxIDrFWzwtn8gMGidpnBH4YQJc0clnY2AP6LAT
CnuHaAV/TGK0tNloDHq3S2xfT6AP5B2OWd6MYyJwYnhtdkwrgc/GSY/xzLbE5Zt9JUdWLtFFwzIB
/1wceZ1H0aN8wvglBchB+UfCy68U+Ewcw12CG9o81h6nw7kSwQW63EpD3H8nMjpivzeLZManbd7E
Qhfht5gP3Mo8QGbo9ACcB5+Z8AKaW1bWBi5cfjAB8tCpTCUPD+u6crJITwEW5LUcRpZJxvbrD328
32SF28CruqAffA8JcLSZUbn34WkmALiL3NgSVWLdszSUtn4VhSVPGOBLQgvfsvgQQ8hs14u9l8Ds
EVnZkIQTInp51cYSsfVXmBbWyGRIY2Iz2EjN4/+RMNxTuTtvPUHD08MPky3QZddb4XqhJrWVtV9X
DvTm2CPbn27RQXEDnYgi4rFhsuliDU20jiRKOdL36XeTNtORRJ0VygEN7yraMJBrpmC+kQu7hkCw
lT7otUp9+1DWb80fz0e9zPk7DOaDZzjfN8fyBMW+2iTfA9mGhh0t4/5IMDp7zToehDQMAlgUWiiq
bElR3F1DiufkxkW7s43x8aihTpM0vpc5QYZEJvqsTSivJVzX+ut4wFYOINL0nAhnnQ9gsvjJ2M7s
S7GaY0lwzHF0ha3mpjDaIH89Tkvz1Mzh41zu3WPE76Dpre143dYOOF2rr2A/OYZVj9437cbNFZqa
MvgVioKru9KohKwzB4mkgoEg4az4HcVxa6GQkueeU7bKKa54lb0qyzCeTEZUsPsRK902bX4acJN3
dBRvfeMDaDDoDv7JAPmO1qFHdS1yEMotzUSc0ov/rMj8PHo8bskOECgTg7zyV7a1XsihJHsJqTyJ
khIiqTomyvUr8zW9gmyK0DKbwJkHOdt6RiubSFXC2oMFPYTw4vlUxSGIUjPO1IvDWo8s6MeCSe0G
CEBxwdkK4VNkZMGx5c5aeIRSomCCxl8s1C5XaJJ8Gzw+vHOuWuiWDAOMAqMEe0LIKvOekQ3dheKT
heg1iCCRVt6zMOA3i2BdpD/rLlqbk6TXB+ZC1AN36kQyrfrj6CPMcFuZxQ2fTqX+UIA4Bn5WtEu4
+yZpTSR0E+aXOyORAKysAYKAPiWawjH2H1npc+sETpX4WQU0UcznI5l56tiHiPwX7jz7hibEnvnk
CRuk4umEBoEFFxdP136GDW/0QhfXFWpDkuFoy5xid+yFGVBl+rb/cxBLVSa8dQ3hMFg5IJ7mjku+
56nlmRHpbjdZTrap6OKBjt/x7sW+WhTs0VZa7iOdW0jf7hvZJpKYL30QvmOCKjChAywbpBOklEUn
MUstKjHwdf/rp56rzfQVdhgN6/+LYeCJy5ImmiGI2yAD2cGpkBcWVDmjnpb3Eg/EnSrJrzdeN6bS
+k4nRZDtsM9yTCd5V1yaMTZ8FiBhZ+XGFQIOW+8AIwGtbXw12lNd7AuPD7SYmyaylK/XIUGlcLaK
1kOmEnP11vlj37/CWjRsztVijQCY6esr0R3xg5sAxdnw4xwdOfRqG00VyjLsvJVJ188yfHThFVWl
fVwGish7qrik+LiNrn238CfXtPo9i4/p7moCEX4h84WuVX9n/guYYh8rmLi3jeMMx2tFrQl4aza2
eoG4hUNlT+2la9+B3UWCsAgVLwbDxJYAS+i2kv+W+DVe286owbiNhdQhEIityDq8qCOdufbiz+wx
KJ0uV1ODMtasVzIK2B/FjLVptCnDd7hU3CKUP/fPYzSo9ktNYz95Sb4riFdoYIWQl26Z7PdiEsOR
hspK8kfmR5MnCEg+4YEP/sur+pmHeREPLOzvvKeg/s8EjRirO7r3RaeUTiIxdMHc2c186xIGgg7X
gpo1SU01p0NAuLbRT55yGcnyl7E1k8sAmJCZh3fQ73VGVoTtqN1uIhvXzWCsURr/MoISBUHQC+Fz
V7NdAI8+UsEAJrdq1fSvVLB0VP4gEWioonBYSDz1Jcpt3c6y17Z9TjTmrtg+77gfZ5jr6mKGUP1n
s+cUatGujtHr4sNAlPXQTZfbbR10lthxma/B9NrGWaWF/2HB4bwaMZy4xsnnxDUbacN8cI6RKTTB
2ruuvIIcjmXhzCeDaRjDoZCbePTbOCJncbIv89+5hFQRhh2HjUFbV88TnOYAoC6/ZlnxSG2chKxg
EVN6gSvFowGGXVOeKwZWkg1qCwtsnUl40v/eCpExR7gzLPWM52BOW0SQaqLAtV1lBsDAdA0SFnno
KHrDneVcYdMwQ3sKTpIbYhujEMkbAft8HbCXErPFeFX00208X0aolyfFPKUXEhQPjorykBDR5eZB
4/CCRrcnhX+CL8d3/Hwy4kXYwCUBDvzV9VgFmtadX7mAbrU1G3Eev54MlqO0zqgvpC6O9io9Scmj
KvmyOkuHAWMvotRBDraYkcvU3l7FtHtabJB1M6KCWu4PaoRQ9S1o8Do4tg9n2C6LkJ6/yYcfqLaA
jJPFy4w7RrjjpXwZxne6i1suspP33+VLcsQN3GiaIlAz+JRG7UszpDCfNbqYKQaTgRc6Irb/A/Xx
9+XW1hOmhHISGalVZu1w2+ANenAA8H6EnZ3RiR3Qfnx4L9hxQXDwYMr1PLlLMZaTHT/NnRYG0C6x
8XKZIzy22F8wHqlpDPTcgn5D6Rf9P2YONxv3RzTiB2IpeskGt0eKs6KcPSTsBEi6d0Nz+EiuOiwN
L6SBkK9LK7ajkqdM+8wL8iZ1pl0Nmp6btoTf92SVNJlYJg1ZFheggFGkTPW0jpgxL91aBTiJ6JUv
o5y+HeakKB9Rspe2ukJtqR3q50orDuzMyPCzGOhEpyF0zMA/t3t60vgkjHx69/5c0+GbQwNjB5OS
3v7uupdtxIqEeLEf/emm+cl5Umltpm2PQVSJ/rWLUHaifh7mec1tjMbWGzDmligj30ZMGKbuiZyg
edN4/hCMB8b29cu9EFLOovteO4wpgXzhZUIS4rblw9w8eS96C+oK1eoEheibEOCmasx3rb9wL2Ce
OaYl275daYAk0AxbHnAxuJ71RpxhDXINVJZzaFWIwwOTG7/vj3BXFmRaf+x8FYY2JmOGVA3rkcE/
ZH76Gth5A/ZsTmWeCajw2bxnlXTdSgOfGKZjJNgb6tgZWtKB85R4nC18nZH7gNkTE57oEpGcOv/X
QVH9xBHyfizos0QGsoCNxTdNzKqM5P7dZVCqEiLq0bqCElUwQ204HLkqLrSl/KyUUavTNmBkZeRX
ySsusSPJLn6qL2PtQMxPc6fHeEZLc0Yx72sR3bGNKekVmpA+0Nw/PckS2V9GUhoYm2tCcq9tlsI+
tcMrg8Ainb4kA5351eqH93IURqZMLttsrfkryY+b8oJ2VmEjODLG3hnbIhaYQBO4FLdOmpqOpY6h
M6XTKnzhhno5YsdnVTkDiOIzSGrQqOd0kaJ+0EEtMbNggEXCx6+aI9lBF6+O90T9yZPlENHNhCPa
gNcZI3AKfpY9wAzF9aB+uKRK/5a4xjGv2r56hWRb2r/II1BF0idEDhs9GC6lv8soyn5pMe195Wr/
Gp57Wv56wZPq9DSUlEr/AoAh4ztcOsQqhdX1AA06gfOANjSmYXswyS2Qa4yYKpTw/GsuwHg+bHtf
R4MopRUPqrrHA2zsWpFeHGjXD9klBP5c4na80b7dktprCRJ+KoxDbYg+ghAQSf4FalIhRC6IEkxV
23y5yzawK785roQVcqv4Ex9Io34eHBrzuHWv0Ik3z9/DslCdTEI/tfS8e67bpgc/yp7f0LPmzRG3
RJp21+8h7cYAIg/yxZEaEJK+AiKRg/5zdSd7kxEjS1aIHlKFRrKp8lbfBegjpSVgqA5h3w6Azgcn
AV5xxU8pbThBgoqON/ug2SvHp9Lmbg+Zrvcz9GuLP8rUgJnpYbHaWcI27b/NOMcf8Y2aW6zolmVo
Ktyfb/Ojq3+8cvLDRiqL/DJ6XQi+LUeVOpbVkXIY0FIjVda1sc+aB03WkVjxt0rJlFcZislMpDgj
31T1/5V5NR0bk1FzCtmvHx6WQFNMt/zZOCir33F4hiKt2Yq0+BasfmV6PFK/yI/0Ih/N0QTmQTFF
QFZCXikgHfd2XXPtPHLa/HC9ak0Dj9WrIaHApXAQF6a2HzfEcx+qT+wMJg73lVcGr4iPRKY8xSP/
N3aRx1ZeGxoWxIn5Fsq2kze6bV6Pk/WsF8rIhZJAYMy9+id9+SATYXIRXaZ1BblemBkAr+/1rUZl
ATGsXb0jnQBL03bcMveGmV3+yKOZiXmHRFPQOzA4SWcQVAHOI4qMNqy9XRzLYLXM8ntGn9J34ym6
+ii9iCGWMxdGuD1+PNR2cTqWc6zqmeQ3Na8yuwhPyqpXHRUcJ1nb7O7Ua9G4L4hXeahRSYaICiFO
j8mo0J7a9GUYhpISe7JTHtzah6EG7aphh0MglPKmRXwJlExO0aZh8Egcpv9seF3OfbSmuOmZCa3r
gAfIW6U5ta1DzNg9esuzssW5sR/QTBLKpy0h8pstWWwuaV4zjZKRn2GKh2CdhqI8ttZymnPOxyn9
sMrY02VN5/OTAfZ7fle+xUTg2zoEsxytzdhYc5xv/KjTIQHAZYwpi2ZS/7sn2pVLpbtef5l3qkJ3
3T6JUGP6EliffZTwnL4MqXQxrYVdy1e9Jf7z97mb34+rpLpWh9Quq7ZoQOC/mkLgag8VS9oFl7z9
9M0Vz7v0a4rt0Sh7BhRv7+ngNLV3vnLDGjBHQEn3/gxG9dCSgOJbCl+oRKb+RtqqRToTn0PFAaJF
zq9t50WQW8gCvsIGUlPgiY3dNs513Dynh1kSATm8two0WI3Be7lI1DCbXQB+c0hQPr5dyhQHqD7U
h2rhdbFXtgCiW+a41FRuKq4hMc77/6zWFaJbEBfd6P5526bStPULcWmFeiHiulOkaQV/TVn8nAX+
DtGUFHuDTB6AyBJ4In5APv/vN3nlGlBtSqjY5G0uTmTSR6kUhdwlJQvYDdZ7XoQbm7pIBu9VGujp
aDP4v35lXF4h5gQf0LNdA2FyGkveJYKFCLPO2UemDjDq1oDL1O712xEy0y3rcUkrQGe287y+eMiw
MTTBnRbZBgAGrY+rklPjIYVM+nORMcRu8u1SkuWk29mu7y3nVwb4U1gNAzGueZ1rD3McmKq2fip3
hXmdWdBt2s59ZLk1AfGi0xn0aY2uD5w6jO+pIm8Gv9WiMa3JXoihOOqGeLyBkJUM98SGneJMzfgU
0/ze6/A4WcBZkwPeVw0ssnwiNbohrhgYXQieewJZTmDIXzYqtSJ13NtjOF9PjW8XP4dfIAzjkKEc
4a+Fd6bTUrr7rEFb0v6aaS2KCWskRaD5H2TdC+szOLIXQqt2aa3vtiP7Paix7QiNLnXckXiLSJjE
lTu1kkFdPRFx6xFNGOSuyTu9TqQlmOs2KaGzneDVPF14hueGGLsZZP0NnPa/bQ1G3yV8zmELMIjO
80UfgjjsRm8RdX6xMf6mOo7PfZ5yWrkBzax+MS/LRq6/i4S6TCigj3t3Q5YEkqTBm1MQrRXZl4V6
TdwEj+psrQjshC4SbwEPoL9J24ViXOT50sepbxOV0g6A0Chjm01pwj1vILDVLPg4Qk8kpvVwbQVR
+huM5DnK6rtSH+bnaKcU78klfKcTbZoiOnlPyqHmNYfCeJOdJ0U4fCVx4LA9+aC5cTSJNb0tZOqo
lo8xEDD8CQf6xBXaLyB99FO6tyHQS1ujcNuY//Np5AIiducf7+BM9GhBto4u7/iMUzQXEuaVxQFz
YzUlfTQoCLYNAVhbFzvB7Ach2pn2ukdrlyL/yc1NrX3IJEo1f0/YWWpKoDExFEulNfdjdXQTfm3A
A2rwzFkTH8rIC0hV26hgCqFJEQOpzx4t69e91ZbvWLx7dRZJDurtZnJmcxulFf2BsFVdHSh3YauU
494jVPtqxqXQ2meF4UN0UBInJxuauEwVCYVlW8u2C5+k0NP5jc0aenXIAneAYCSs+RxAinG414JQ
egBC3qc5kQ4FL7j8fLtRFcbimjtlQLnQ6FsyYVHqt26FrcfwwoJEtmdOe/G2FWKZHHKmZdshkwcn
IuKiGn7awMjZOHKsuhfuIi9cGCw8OFgZToyCln4nv3skEgtE/QV+asGLNK43UuJ+I4F8cRHJ8XFc
3+p09HVYKLNdT4Rj46gSsWmf36txDhlykqNDjQy4nbpxzCh5vD2jupVyyfbT9YGSWm6Y2wt+u6+Z
0CcW6hzcYDihI8H2qKEPoZcPAj8wJlgG10Z2ba2IIxkOF90WIZD8Lg/utQZ8XiSPuM0jHOjuNp4o
h2cI/VEOoMwlSPTPNZ1C7K2YUAeX2LslkT6yTQmGwMv/Dh2zdNI0wzs8zQA68d6S9sAicRA5xXrK
DqdgEIzrViwShZPXujtrfjAhpJupOe+2BlmlmJcR93gn29z/cWReHHkFS4UFxD7r87QpjpkBIrkS
JJBWYfc/cLBRWmjwW0HFNhyCLZs9aRBZqqsFgfbAlQFvCPqTVHebsVMYvHdrFqHwiFf5JqeiS6Gs
owcvx67I2+PZS+ENlrP3Np2WzXUVuQK44Zm+mN+6XXkUoJyfcYEiIiM4LBu+sL9cS8hDug/UogC9
7TL3ZOpQOxvHgvRQ6T9hiHHSgw/vgpt6MOHoe5Sq4VucQ/L5s2tsQfJvKiqDb0jzeehCg7j7wAgo
IWOf6Bi138dMGtAdiYeRgaXA2vto4+K0olArzKMaMA2j9v2Kdashf7RI47CAlLXfkcjrPx8ScGpe
8yyvpGVvEYbpFBZLqkYZNAQFbgD8fxx5YiiNqmMoqPBYPmdKvvRih1cUPd2OGuWFMO3l7ufIzmE7
xb7asakZkFuI/ciLTTFA5V4dLGRKYORJ0d+btRlOecO8QOTZ+jY6kGZwDlL03mPvhex7Su4VTRVc
S7WJ+su+CLDRawnZ4VRmIJjM4g32RGQZZq0+k+CzFyxVEAyElGeMDLsZ8U7Z5rQ5KCemgs6ticOQ
WrqS49yPxxkcBjic0ABh03NbJzzncjdr1igJZ1uagxgqT+Okoq4mgrImetOoLovAmzP8XUqlkINL
XpzKCX81ZOpTwE+apEZEqQB9+iruAoQ0Oz56bkgE+9qyIhQRoFY+oA/Oz1SX1PcXN83JhJsAd86g
VLPzNHqUT2hbvc8tTD2CEEImizXGWFIgRB4wHMjbiKn6OJWWNDvXq9SsJiBBX3grCBxBJZSSsv0d
VoZbf21aeDvvZeX6bJvDE9U430A70XErKGckOD2kyK60EEaUHkYlB3txxV5lQfz8+7N4Z+1wFNoW
pUKl9qTtm9O52Bb2kN2uwm0aHwtdH69lOg8iPfR5PjqVkui/nY1+fBV/upqj/zAg39ZVFCF0vp9l
QKon3KWh9f7hi0V9SsifA8IukrO2ofArGLueAa4bee+qHjnVOicxLOl0C59Dpa6U+i4kxp8GTJnf
rsh+lLkoxoFHZMlsTx9gSKI0PHZKPbid5vHJvpCp4yzUt+VNW/Gd/GU6CvwU4Hxypn6tPfgoVV3N
qskdNQ8BD96bf3DcxQYQ10qZ3mvaxll89vWnS13KOmyDxLw4Kj1An07BSGhPTNBciCHa1gMkdBAB
cLyzylQZSDK+G+iHNcgZ3NmRSudbOM5wN1R77KVVja81lLsbpltnlNzTL5YsNdzxjzw59M9eZ6bG
j1QBo6WOKB0Zou0Jobs4ecl36AJXBBr69tfIMZkr8FzyFFJDqwryKdBNnZNvcVLttZAlTOZQZ895
p/mE66sqxsZO8VRCuXe/GYaJFNivGlMxCAYJ51a2kvWXIvxneCxAoxgSNOGAHX9y5SrQHpxMDMU7
jrLR7PtPNMi50pfu6MCB+qvOJzLu9J4G+XzRh9ycc1W+11XJpjB2LzNQOrVnk800TPTZbyZTYtzA
blp1pStHgH5/7vHrL32tT7h60wbNGQLwrfbbPTWNKqM+I9BexdF0vyynCFDV9WZkt2FItKcGCRoO
87tzcTVpvshYoLdHDfR9LRMqGLhlpoSU2lDhOFav6Vh5vdv6dielbBrFr7zN+S9NRq7xLQOwMqIa
4i/eFka0PPNJpZZApmk3+k8htdxtZeSvSzlEymmK3cce94rq35F1ScJqaEnUqnhr4fLSlqdhR10x
sj1Rvwim3hSz9Yn1+aziGZatFY/v6G1Z4kqTt+czefowKcyGIWhZadPzRV5LdjyGzb8KCEuqStT0
FDopd2Z5xqne2sJaiJrFuuV5aPdgR4Ws8YLxPRc/vM9SLWsT6UedOkP5yUr0cdQvdmre9dHW4oI9
7HYKfS6eGBD0srXotXh9RXOyO8Vn9Iei2O6pCNpTSSA1UdQ/x0NY4mwOlW+crkb6iiRmuAGK6Z2l
byWD73LHaIoWPGgbcmnz5MSO5ikSxZ++Q8OLCMYQWgzUxNp7f4qpC0gVD6J36UKZtQBc3LyETW8X
2oq7aRAvNeeHxYLQF2XWlCN4s3qwGdYscbBgFTsE038HKJ+Dp/osxSokT4tymiYFnPNkOT5dWT/P
BrNIZlIyshlGwI1/gWG8cKgvCm36HPGpmau/kcHu6kSKTUJO1CWLLbJBLe9xdbqs62Si4beJuuwM
tEeb8Q6gSsGHKbMMMtnzKTUGpBlKpl7YikVHCnmBo+7FeHKBy9H3++WGJ6hqJOunIJjN1VeXQvL/
PN8/+MUMqHSwtzrzy27YemVrdaKv0y4baPf0Wo+MCTjoXCR/ENSr0OGe9Y6Xho385/DA0OjA6cdO
nsuEPAF+6T7KELKkCyFeTX0NE20HKrOpyj7giXifcaFLJoKqSXawR7h6nX9kMQHQnfhctdiJOHX8
h8i7bBNwA2xPlk4hQFq2iH4RIjeiCTrruhpLTDZ2RPYgJg+hjsWG1LCCOCQXbFgf5hwqtyQlcney
a6aEtTVDlalM3wwxm20mAaMaJlatB1YouGonYqmmJ2M50jX32y9/KEqHzZF4lvv1LJA0Kgyk34tI
oItYAlEfXaa6OGtbfnxm8DSXEuVl2waHANKnIv6G0I4I/t+kpQDpKouqBUYu8z/97UMO8W3lAElN
74wpXB0gbAeJhp2vk7q5aX5HkSrPMuUUqhqg/S1L0QmEN2XeYIBwy7wmCYEm2Kl3HbvWUDoCcTX3
+T3onekS9/8KMiTtDiE/VPOcOUH+xOh/Cki01IRwYqVobEoq/1cPgHKVAGtvglFvKTxbygxj5H2d
r1/QXkrMawUs0c7uIkYvqHJ7XidENCiZlEoCynlxUmY9aoxH+iArrnV5EUYiD2CgR1tmJyF4ImNh
Rk9BoWJ6GydeWZOln2Ed4EQEPE33zY386TPI+IYdyhadPnJI4VjjoANt9VhMjbW5dwV7wCNP7Dou
CQs5XNoB/tuvGbQGRPZg2Wjm4RQKAp0LLblwj23B1NOe5YHtYfkx2XAK/GtNzTLVHRk2u8M99OG9
pAkFVst+GFbeG5IRmH/Jw64XKjbvZNRKutPECJzG2wkLh7YF4oSez0HypMzoT/5ZHVOkAQyHHMtj
r0eHKWfLn5MraSqUQPh70btW9DurIA3rlxyCqaFOKqO3Eow1K5wnxrGyG6mno2OAqXIBAxnZSG0z
92kRJGXNAJvESNBRXtZvXuSlcPopMd+a1/m8cjLYMZ4jd4NGISw/trKk0oyh45hF/xFtvi9LCy2L
dir4JYG1P6AhC20pr2+a5CJUkk6hWNoYd/msqJroem+Fmx14fIeBZStySVYD7yWMMi1vE1QoujcX
Kame52yYj8CvLVSCA9gW8laC6DolXHHcdm6zXYh/6iFXeZK7ajPcYRy0SFE18mnDhOVGIXu4PiL3
3/eeyPM77aUKBDYJXRA0zp4n6fHsfJrEEhtR1OaelB9XDvJKObpaWSE0OU9GEiqD4wWijREkcahn
p9v7YDmi3ZJ0Q0/QUBTwSSO0WH6UISGDmgacayAtAzSYrIGufh8snt13PLElUVeVVgsHG8jbMHnd
ODK2QFkEyPIcb9fcrJ7lPwAA1L61vIPLUXyT8K7ivHEAwm5iFEFli7b+RR67QmBCG/PCHrCF4MY8
jaN8Ve6/SOLiVv+ByrTh61xw+Rolr770zZblWweMQbDocQrMSHefK+Bbx7+Ia3n8fzZVhJnPYO0J
yQxKL5FmX94SNjqObKmnTf8hu8fqafdiomGGiibA5SzoDxRJ6pw9kyDhJU5x2rj63glIunoEc34P
MqosHZ3zsYbrLuxOMJ7UVSph300e3w363Rc7RpDWGnN7iOXm2eCTFhRPMdVr/CRtGU8SqFlU1NJS
r1rvlwO7/zWHjDdf0W444vk9N34lwAsyeLhnwQRm/IYiY4eYI6tH+D/bNhVu0fM0aoMdOU7xrQiF
QMuWlg8eAwuIFgdQ+TpyApOaR5b0eWrH9bo7GDMEgHf5gSNs4rS6K1Jj24h+FO8fgO0KEeEb5rc9
rM47MAmqxUb25dqx9Pt1fW/eQupx7oZEUXO5ttWKXk9cBdjqU/biSLqt2WBCv6o4QnW13AbwPW/w
YHQaYaIg7BRrIs/xx57JsmHMMCj4cu7e6Rv+A6/EravwO1wyh1kV9N3LJyLD5HJvHnLtkrLntu1l
fdp5tEyLY4fdMX6xbMS77JT8QQ+lSRAjqFD+JroQCtCzRNipFHR4x6Silu+uCNZ44e2FsQlim0Pt
zhSGWQgLscc4qwwgD8fb3hjN6IwtoMN30CQo9ON2KU8Ck2HwnbfsCMmMPoetueZGYacyjRhlSykc
RE2t84BYlv/CHttTpH0Lqwp63P8M5HQiCC+5DJMDZjh1UNDKhdpWkkkhT81j/Px3109d4+1zv9vz
AyG61TaRd8OlBBVxJAwurIDqc8jcPNmiViesQYuZFXx9b4+t+Xqqy/F6RViiT+F3k6b1GjopMjbQ
nvWL93c7x0QIYbtz0vJnxeu6fsesY/LyJqDUhSd2YB03N2Eu+aVUGjBN0wW6vayKV67NDA8wRGup
102b+Z2iATZ3Lw5QTG8WUrQmRdYRKMSNSWVmOhnU9CRTTGkdprLNrzhUT6WtwcIZEDm7eCjvCjta
thB4A71mUOBUe0LR91GsVdNihFdY8BdmO4BgePG4Bb0zC7pm0kYeHLjeBz0gTkDk8xjQhaTNUwHs
ie1EfUFsQbF/QwSs4OYhisEGjDI9GsQTUJJharyovQKfG7kxk62zHZ4cd//Su2idoP/d3NdT0GWz
rsDwtjU7E3+97Urs37TKlL57fn0nDckQ+/wd6giMRShLromyoex87zfwOi3UiV7iLyP01PSiYAwr
5m7hw3j4yZyZdLk9P1U9aQfJ1NNkisQntgSZD1FLOycsQiNLHPI6IG0ON9B8CjpuMuUoHd78tmet
Oai11uksN4Y3IhAX65eEZFoVbjbY87RyQuc0I9Zow16vsBLbt9BGAbkjXlWywvUlhQY+1JWcNhQU
YOLxYC/Zyx8vcAZLe86wIBhp3Ayx8BuQJ2fo3rlK801AFhLGIIoRiOzB+bRyZb/f4qHQg5zuDZ0J
wKYXW7sHOty0/K/37+fVGsG7i1+bPhya2Yun8Rb73osrjZ9ALxfJ53IXO/Gsd7pzPIcGXrEc/dJU
9MafinC2CmzVQ7koOcL4Iu5LrnB+5HKYeIRlnybz6TF6FYGCyk3XGzGLLW0kEdoO2gxEV859erqx
Cuiae9b0X2/QOAR6mz4UQ8Lx9GKjdVJxxYmpjNMgb5SB6OcpxrAC+MEwuLBRhQgboDLnJ+5Oy1Ga
fXnQX4oiS406BiZyD8nY0y/e6BeB+YBBEwGwT0273VZ+BAGGFuIBl734qnbXj8z3pSGVFeiSHiFq
qytC9IU0Crc4RV0iSxbrnmrPoQAwu2rVgjlL0GBTIkSJOfjZsHJb6Ejvy6swY8qO8d7HiodKSUV3
WI0kxeryPaEfWAKOLhtQZNdtSbgFXtOOno+InYVR3rXUZF5l+6hF2Vh9MaXs1148cqyg9IZLTmHr
twSoG/w/eMIsRTNkR7K4o/FK6JczlZvMTSjdVsqfZkgyjkxVnfK09Gw5MRFND0bm+MZLAf/2iDwf
7PGDdogcqQ86ZZN/MAGuX2YHYxOf0rWsZKUAwLS1hQCkOHn73ScGmOHQzL2Cd8H5+k65DxXlo3db
xVyXScqsz0DsPble+clKTNZ5SY6TRstLU1ZMXnuE9ccJbh+n+hETBO+OHc0BU5sueUIwObwtyvTr
vpOMaqgfE480/jbIlWGOFE56AUUF1LB/o0X4nomnMkfUCPkQCD+JV7MWTRy7DdFgRkz0eOprMV56
Ot9KdMyqZpQh0znx+ABhWfFElB0h5GYFAUt1r/jy/xBHp1r/PPf0mqhUgPhwhrFPoFdD43wMFA9T
cB5Bj48MfBGqP2jmgAaf4kv5fL16Z0zmSqnv8eEil0US3lldqXVZtYhuqKS9izZVmVzXWjC6PQUo
H7g37NG1wJUwpY6Lo5baUSdWT2rI+eCfSwcSO4ZoYSIklmnf6rWzpx8Wu+q+vzJfqOlqDWvSJWAf
UVYzgxIqLaJTu9ABl/zAGdNI0icQl+4Ok5pyhHGndi07ezUWAlvZBxN2wAXkuSS6F30EmI1/i34c
2Z5dSTWWonGvA64NHTrbjpTRytq5mGYquxVFDjvFK+nQLe3glzbJAApeb30I9kA2GQuC7W3HYJI2
LT5jIyE5mZWbilAlr1QDfzcAC/6chUTndnVSjxEKE4yhHB0RBUesrexORKUsNFAbJPkNgmf1ReE+
ESKERGF1jEyRgFzpSytpgM3f+z83X84BIfgTKjpa+dMItPwlf03AiLP/Q4SbQpw3nddp0QvGHjlr
vNLGyJleqnD7KBf+KVwrgvwruvZL8d+nMVE35M893p8B6XuknjEMj4oUXiNw2pMPNfCezsV8qVpo
q3Fb3LzItJMWVaK7XP5rQFGsRpayA/qLmSw3DqGxlNHp+FgWU/LK0beCDoY/ClS8AhUF5oErIZv9
2uQJ6pMCMDe6L1pvJj5LAKBxB+hfdtpACO6Nme8Q3ccAv45Lft4aOHJHY+6GKHGMIbZ6jSY7Nsvc
c6evfEpeGx1bLbP/dyFKsuuJkO51StqDhaem+t+HY4HkyzKKLQ3uNfbpdGjuZ2qJa+BPOZHIgCtw
SLcpjhjfcAWY939xXUVS08YPIQ1i45d76fFuyyPn632WY6N/1/xvgUJpLD1iX7fRvBjwu86O/PQ7
bOq57t+c4HFCaFt3Npq0NCXWeda+y29K0fhTzMU6yDj3NgC73vlyRrS4Makmz7ok1OOsI37cHCCX
bwWWT8AnH/0Z74wc2hkx6VlQXvLajxt4vTq/kjaDe5i88ePJuZSXh1HOwQc9rLomTarc2JIwC+wl
ME0G2PFA0rfBLe2JazTJRfo+Lh8RjSIhAClauF8Ft9zwmkx54XSkaQjE8AEzIs7ZW4R07Rx9t3+B
l64cEPbswGIORQlvj0B/BruNpbqns+ZQI5UWnOZa8geYXCHkW744rGH0fqY27fl7+SEvAOUfAawC
NvVK5OFI7qsggGFOzX8fn56RlMaw0PAUSqNVnb4QzmA9Jq8cGBXxdk7nel5r7bTnnLeGkTzKL4Pc
QZdEHkZZUlGWFhZHgoP0MjIBdX1R31uwGUm026FkBLNMvxpfzuFiPgF2696bIPTg5vMDu0yTa7KV
R0BakXbKfSGya1YRihmUWr0atGkjs+zuV/ggG9Gkn6UT199RjmI7rzzYASP4Vc4+I498n8+tYse1
NNf7ykaNY/Jc8ZV458agcXL9YRFLMegaNCMFuzxejO3ZYQHUGzsYFyvpz3yfshccenEyDh1mYq60
nFv/i9QQo7SnHJvSNwhm8p8J+SleIqmMFrArghmUcQIehCczDNSweIZMYVyX48llAWRkH9HeEJxT
S9zkEQBq/1iYpC4Z+q2mPs4rUu1/f/CKbrosz29Rbjcjta+EVJs9HQu6ukgbMZjlv4Ik9j+4uq6f
0b9GC0HyTwvfDYuq+Y0U1lwShSUgaliR5icV/q6tNLNAXEk8FL7Z1JaiI4j9pzle6Nu/wgjtgMQD
Ux7K4/IEPdrp8TTcbBWJa/RTUjYNUFLeFh0uMgGQko2Xej0/zSeJy4DHRNUpoCbHTTyzG8WzLjk8
+E1owJAHSTfkuVIpS+CzIWO6mRh0IEWdCJNoT6fNBQchWTEFfwu3KdCoDNwKjZNbbJWK5Z54tlr3
+foicJOQks0dwk9tNPJm253vtnABM3jD7Qi042CR7NmGc7tzzdIwOtRkNvxogL3/NWOQTLtIWw5l
br7psEfnbmYyrJ2PDUuJg9L6nEenwBMOKCKTgmR50iRj8qzEIr5i/SJiCyepeqhM5c+KAB4YeVaM
zIJWNpkfN9KfAUbGtfIHgFB3cqIssUn23xo9VWtfP095a9CYsELDU5ODzFe/ZxIwKjK4idRAQxYt
oyqJy1MdA9G6eM7L34En4o8n18SH2FELhp4uJx/qR36k8g6on5rm/QE4mcyTrzmDilRqSH1QQh3V
K//A0go+YdsNAu+RU8mLIm2hBI0Svr6F120VfY9Zvhasdp/AufHJXAYQ35notw/HquYcpuRYORVT
dEQCBjwFrnp2jYC2opCIpN1+yE8IUtiu7XVVQUrtcbsTpN2wBa1GB3wXn8d1OTrGH4a7uxykyk0h
fkWaIE5pOJU33NtOVi8gm0tEfQransgOLliqAVSWRXFK9olq6aDsaScvP68e31+QhmPl8XsRB97f
oQTPYT81g4DUP2g/sqmHeYxyK5cD+4ohjbwODJNLI1BM72Omy3sKomixDCh81tVKGBfonz5D7bkH
frEtHWzffYFqBMTvtT30MhWmCh6xokO2e3uBnXV+gOA/IlBuA/zVMwtHxXYF+uWOiAehiXmDZ1GT
t1g75S0Ry5XCJparPhmhfhITvWuv519Tb1Q/EN4KIJWy8LF7VSJaq2H4RiitbSX7x1B09JImVBv6
SiVhE6cdtGVjV5Z85IDwYUdpuRJiwe1m0r59s//8Zx2emNo8F6Sg/WpChJVL6nEXhDNx6+ryc8le
hsAj0GhUOuUK5G6trgBteFqQeEDge49xzSzUBh0dzxtLETObE/oI0p5hrsT00nn+oCoEkjaT6oFp
pKNwlmeaviqAGY+gJm/Uxz+/W3Ra7vdsJ1x6bdKXAKYcVTulCPPHwBSO8Da2RpSd5MsF9qTaYOYC
rCQSdj2dI6Mu326euWtAVc8UMtmiAxDGx1Jgq9VOgXDWaH4+p3uZdD0qR9g7K4sRNQN7e8dxphdn
b0mHK1RrBB8tsiXQHlIp2FPMcrF2o3oodgFH16T7JacRivWynLBj1KzSD/96udzMnry/+hmD9geP
uH2eDT7L6YVwn4DUfTcJcLKquxueHWKPqdab4oh8ZLeWyXdbq9XmsVEaam619iFwgayH7fe38bUa
3Icwy5zIYhd1ZDQcceYbfb1cBk+ecnw0Iml5ddSnvSe/Jqx9AKHsHJuKm/jeVjv/EJThC8Bitshs
NaHd53BnqsRoTyf4RSkMpFEaMO7/C6xh6EyV59xGzOi7a16wY2R7sos9keIWxociLp7FN9kWrZgM
SBlZ5/rt5FaH+d7c7yUrupOkXVpmYYDZmwRDKFBYXOnGRPmhjHndoPZsoyI38IsT2eOdjhJyKEw9
BrtlpIy2xezlIOp9+At4vJJe+S4H1lkHNa2hNeokreJ3SCn0ySdOOF2HXlyQgWSRRuMjRdEE8t4L
QWJEFTOPqs+JpjyO7JRI2XeHG/Ioa8NDcSSPLy2wOOf9QBm3BUOAK8IPdvFkab9S+a+pyujWIN3h
yD7c0eWqxFsxeIFh5hWIGYRL3sloMJFCITU09cd8ga3X+bEaQBXg/jcXowD8TgkIAxiflQjLTDGG
mdVcRddN9Vb8MwZj0omiadNuuMCfjZzZG6BMddyrZiaL+Ha/sHQmjQ/g/ibEpdAkS1pgynK9WPLd
HkI2WomrW60qrW7gjD2G6e+WZQNZoLXZInKcZJErdEGQaeen0qWQsLrXsQFpU0IAswSFmgD2WptX
arlyMG15S4gLjxaIAX5Xg3/Ii44Zq63NjXm6p6Quvis9bwKUNk+BMzMlA3NP2XcHJWvaYz44cWnU
fQjpwKZB08PHjE727SWtjhXQzR3ahJ93rgzulff1Ime/3GFHUqTarXutdVqaNcuORtXj5Jod6Fjw
LrPSsQty1TFIAJ1NrE47OUj8Yr3oGe/phqxmz9IyokisnX64vplWVV45Guic69bEJuCTMm27eu9w
bzEkKhrXhSXrMuGo/7+LEA1f9rcMgec/0ModOnIeDp3cde22ivoFGKSAnPfHqTJnaAdUkv43zrhH
fJvTZwlVfd/XuS+fg8d+6517fx8mjfqxcaurTMV13FOEK7IdUtZUJk1nirFTzGkzeLw9tJzNMQfT
C1QFQFzDbQZKO9DUQFZADxyvwVZTKj0uMb5WDLZIyLSO8rQ+xSniqqaLLBu/U6i9VF/Z9h9KfYN6
OoQTyQu4ZRo3aEk+8t52c+b3UdqmtOWKyGZJJf6Z1TLGoSOS0B8Qy910+xAwHaLAaemoMB9CG3Je
prTuEqA6eIRkCLvdbgyhdhY8I4byRb+HdYA1kAFWudvuB7IkXzbxkbf30MyEwrgLVIpQqWifuOxV
ev4/dfZ4vspbf4BaLvgAi4IpA0aYzEHCCw4tpJqf55S1A2A6w+GUMWF17U2cL/22EehQTzrvn1i5
qf4JUxQxGjHgGluWWgRuJAs5HG9bWUhzT2F6+h+3/41t8f7zO3e/VqEf8bSQcxexWWgsOBl0+gye
OEAZjh3sGdFWBlI8EYeim2F/7X4JLpZYr4wJQOCNJ5vgjoiz/GiJOSAhjTbzWjLZcixSR9GC5V6i
tsP/oPBz6hAZxGXIeq5R9dFdoU/XzZXphB1ScycpXwgDcOyk7GL/JfX8cCi1Ci77yUZN9wirjSag
l4dnmtTIDhNhsiR6yL6poeBmT/clwzT91J6DFemi75gDvhIURrxSYs9g+nxIueYFAUHjo4YuYtHz
OREvAUHGhgmjvtWzR0ZgJ4z805ANAD2BLkPZ/mPawCtlONjWimORXl3dwDQVNza5YV7RahDJGJ/V
QY3zgSgbFeIhkFg3K1h9HGur8TG22MrVtl//4GjJcLHRi5i+KAEXZAqZu0sNXBZCDs1P1jiXu9DT
x5/BZx5e9hENwllTP/jPpLDSY6ulZZyW1hPGaglOshxv9PdXZpyz6Jf30eoqtrHy9a/KEmtoJDZ7
3IxIzBd9EBPQeQKxrj0IVzDzKnhM7+sCwsED1LR554qP4ildtsNk8jaOgvd9rhZtDAGKy9WIbF9E
BjF7gLtpRrLLmUeAgnLb9TAKRLLyqrVY2+Vr7EKC30B/qa2DwP8Ahe4U1IwgnVMFVCYhxZjTg3wE
y5ZO0qGfQqQnADZhB9VVHqZjFSXtsrEj+CTbsUTyrg6rpj/gNs4JtqSCQKP8qIRcoV9ujeqFmQLY
Uexcmp/ifmXFeET/9h2nGrXZ2qHO4P25tbRMwl0UfmmamNlSVW9OaeMwrbv4U0J8ZIksMS3af4Cp
qANY2tj1CRlcZ5Un3edM8j3RwdZwbFs95Wx62MeioXbuIwF+nE/rs+A7GxakKwZDXOZh41eXKOwA
FN1MbgpMj3gPlhARNgjWuWKibgHc8KSdD/X9N476s0c39O9A0LcVsn0040+PDtVway78a3v9Mjp6
OyIK1FgG6rRCDGWIROB0F1k7TbCrSjUiNdtx0u1Vcf64tf3FAnz31ynMo0JRq4kLcAmNgNoFOZju
z4uLTnIaDIsnXtgI6xRXtHkz8wjtdQMxiVI4BTi5RrEt4kLnAUlXySYKGwvMlnDSmvK/ulwnbVrP
hHyLKn9qwWdsZmHwjbQdpItJYN0iLNrfY63J91WgGtSnaSH9lCz5ubjq3W6g5TCqvGp8dyU9sFSh
/FOY95/EGIFqI43SoKCcXLAjcYApZfqULonb9dJivK0EQHDWusziVTPqR887oK1vSQoy3CzVlQzZ
G2Xszdv7rKHVQlCKbx4bISXfrLGcLnoQKvUO/ERJKFvpg1mxQWokH6K48VwHWp4/BHt5qQ/BkLxt
/zlLIuIAg84eRRSfqlqiK5Kp41Kpvf5DM1sNgez+5tCQfgrUFEgRCX+4uz3Te5EakXRVYUquuWsw
s0xiDQzV/dUUTAPKhxBu/Oy8zJBseSUCEaCJEa505bxee1IOugl0sytbarYoLq9w61G7XMXt1mG2
CClW6LO+JeEmERKcSZaW/pO7Dv0sqBXML1C56px3OCpdESUR4NCa7VRZhl6/hoNxOjGhE2tmDvPJ
M0AA/BMUp5quQYJX3nxy4QUIJOd4ZiqtOolebSZa4Y5DlCUVTYw8T1MRxXxHATs8TPsDEzXpTupb
N/Koe0VevgGcaf2ujzGbKlv3VC+Ifz5qSt851MpeAm1F1A9u2KzyiPTwcji0RecyVhlmcP57u1na
CowQbSDoPKORbPBi/4gjPGHyGnq5SFueE+MgNy/oOjmCqSMqTBFIzAmYzhgHYoQBHvSohU3lQjfm
M/HDZUX5jZbcmUfeRs4nOj1KnNe78PDA7JiBaMZrdjR2eWxS/GPD5zQs0IsqmXH21ayY4x4lwdkT
cgdwWg7pZIUq5ljpbKe+nfd3QwCciimlwyI07BIcKLbPlHnu+iSHod5gZJTYghf6SHuuKWd7B1gP
zK7Z8p/OLFvI+Ts1BJs/CaQxIP8k1fwX4cIjbH6xmCcpu9xN7H58bQZbRMoJHPGZCRV+s7tovOKo
js+R+BOc+xMyYcujY63eICkc8RQQkJO0nM9bDaNn+QkyYOOPumpxESqlSoKuH1h+P7oaQwiK7aL0
eBLsw7Cu8s8u8NU979LfH9RpeQp+ZFvAr1MF9Sp5UfX1WM71bVKcSOCS5prGrTuXD5X2RFtSaZZd
A6CumAlbY+88vQyEL7dG0TjROFawSlrSkBnJIgj6+ubIJXqgNcnDqen+xojAggCh/rZrO2zWXs1/
wUMgcPhhDfBNXPqAiSz8Pcptiytaw79mnBec8gaYZvVtG80sjDsbpqFR0kGmh39wdjA7Itrgm1+V
4jY+loTn7gZlf/a8rgMBXTY8H4XTY9iCkASvhoquzmB8cjztega/sIPC63hCe5lkRVf4XdhU4gf9
MpABxAkQm03S1bgt4qGKDelgVKhv8BdPnOr+U1IeTjDG+ZIsDus8CY8aSaPQAvRgLuo9tYK5OxMk
w/yF5lcH43xa1PaD+7RZBlWPfQwkPU+Gwhhhbq/L04V04I+d+JOzW9X/zg/fpZ+MV+PLdYCNnnf7
0EZ9u07M9K6Xn3suGQm9rgxntPdyRXMJhoMqqDWdUB+e2yUztrjOccYsoBphrPRB7W3O0VLeL7VE
0idMP++7XVULIOQAY4Yb9zF5cnraP7wAc5l7SE05Vu9DchJAhzcNkNzA2m30Fo3nPqHKsoZ4vPyK
XX6DTvMLD5TeL1iHPTkNq1/jfUIGprbywcaa8+h2bMXs8XCilXimu30hQzDoy5/7P9boZtPPUPRZ
l6OPdvW8tPOgRzuYO22WFfz1BgfBpXWBUhUQ/wMvZOUHlkrFKKZzdVUud5CQe8caofIobNBU/OMo
0rnOxPadXp2VkmOi4jJo1177m7voBmB9tH7nRcMSLkxJSwgVjGtUHMbpr3Dr5/soGwGtd56ivvQ9
UKmS8k+Rq39c6q06Z2eyopijUtKpcWorNHhSNaJNsPlhd+cTHb5zN86CiTCk+GIZbaFaY/yVq+uV
3IX0ihdW7kUO/N8rpN55PeblrN6nUgkgCYg/OjNa51cKKEi2pm8Z7CkX213lfK+qPcjbKDgGoTbs
fF78GNWbOUqJUd6OVA3b5GuC/ncsi0RbhBzFCI6Gp+8JPdo3pzOAIaDsr4hOhecdxDAv9aSiGw0s
8L6HYrQhvGbDNSiIhw//jHZ5jyHvBqqYAt2iFQ/2jDiN5KoqoArMoLniCNWEMdzdz8M6JF2w6jqe
xhtalmlE73PTW/Jj5OU8nleIL45RjwH4S27y1z66/fgpBAq+lSIkyBAEHYC9uK21KP2UbnW/NKUR
wRHGiwDoKVg7WQ9tDpGCVy/44sqjehLk8PCfeqmoWVmJsqPBUarNCoo7ncTssSkKclZCO76cPLU/
EF5Vv7cNTwCyezQEx2/xoROVj+7miW9vvRfN3W3nYKDVsAYghc5GUzDXyHuc66UpxzIGBI2dXfum
PO2lPCWSlbDMjNbYtI2VcwEWCkaz3Hmj/FKKASwFJ0vc1V+HHhaLiKHlomgXhqN0l6jEnfRk2guB
Pkrj+l//Ga0s11eeMV4A/VUTtZvGb8CupB7Q68YJ1HZ9XAPNHp5vw1LUx2RTjaGMxOQ1FNjnosY5
ty5TpC+OI+BAkDKbko0q/wHp02iS0QYw0+MeJgEQzsIvL5uR+WtjQBEh+stvJQEATfB9/MpLZn2H
79vpDXdYMp/kQu72YUTMi5N2D2BvGlNsKZS5T+jeOIFwRMlnYONN224fqYQziTtlwBHj6PjKxNzR
rLSYPnmImpRBBVKq3rBaXXy0yuSSWwbIgM9mD3xSca1y9P40SlQ0hk/jDKppwHd1zZoRxvlijINQ
AbBd4AwusGNVSZhWQsUyK9rwk5jgZ3dYEDKEa0eD8oo1khSWf9/x6PnVwvvkfMOO7ItxCBJm9JXE
wkCPTTp+ex90x3LSYqbP75aY5gX1MbkbZRzHUk3/Yish/5Yih04vDHmraAudJcgBRKFSMx8+Wx6v
Cv6nGOvruEOw8oj428yacWhkPwdfNWDwag4wG5FVPI5feazqdyL05ALxVC7t82jH47TzZeEe+51k
URe3l7TjyQNeF9LYa/ila2CbX67JJiC/fOcPqFXj1KhGoe2misNZbSmHah28317R9NVCvIrpBvDP
fOyexuH5JOUzhe0jwONQtasz4WnaE3BNAh3w5pldzyGnzZ+dAsGWdv+npeEtVM5/YwthlueY428z
f2FnDTYKuArSCYligiNj2+ICC+wwxII9XkU3wbZtkrkmMMYmANy7LFXpgxP2/mnbE+WOJeY7t5s8
NFGlXhOipQosaFIuFR4VJENH26U+Y4fdMtUD+i3BJvxjb9D05X21HoWTa+C8pxsvQUUwUYi1EQOP
YDJNzXrGRpE7sWn56Avf5WKf4gt8YCAzpfS/AXjqKV1usnVBPLuNpuuaKQcROT5CvWWMqlc3VYCv
XNenOIYZ8pTRJlOX9WrsGmnDfNyBaXFfZvFx0u/YvG2a6u5x31WpBOikNCRBwlwgqjH7SvfBUKd4
Aei/DFDSvBZGaa0hOifDPuncDwb6J3MYRSJPirr4IpJLRGucxOtC4uN/bvSulhyvBV2P5yjVSYN2
owVsMbI1VvynAoWuMfGyuwqQfrBV/foDSeC5B3QLK9ej3WoLNk5KfuLOwTHwi1qzu0qbAmd9YAB8
XRKGajMsEaa27Do8buC6MDMEEOtaOZLNRS6oEiXjjokmK7hNLV1jXE0dTtgFBnjVI1wF8RLgsy4H
Yp6OsboxVHvOf69msBki7Vdkgp2mcix5LJFcWQvq9wLFmoSD82p5KtECPuMPzWJUu0VoFDxmT1iK
6flO+5wo0WFZPWNvtaUCXrqSETadK5ku9u5yPnYakrkVj4CcAIT0XhYaBn19hyX+dfk/napSN88j
64GEVbRUmpzk/jnha/1jUTSTevRLJFF9WMuFqjmtkQOUNyj7ZKonLKXKcC3P49d7ZDflbjH+rGuX
WrcrjaiT4KoyDAx3Joh13icmA6tDN32Ad/cFYGJhQTE8pUIqcOhrx1kjUu9R/qQJWjUH0I+UGXDF
dzVgJ6q97aqwM88B69PbTHY1sGDvJjnwSpY79xKXulOgR3IuhTpWIaU0mKxcBk6crQToHPoiZ3L6
jLup9rXoTcQ/q2spJCGVZ/9kkblW4fsSNoN37URil59CsUjXcmmZ6n3OT+FBtFas/b9JJjAPsVrk
W+1IbNYLaPnW1mzGLfmE716n8QayIGJB07bmZtOkT94jAU+1O59TWDYMJMq/WlWzOWfzmVKThciV
sYiT76+H0HM6Ot1rK2xMF98J0PHJDMK8DwlJJZW9xNDYCNpgVZbxkdFxxJwj1RT+iEbrFlIATn8M
BL5Lf5Vm+FN5P9iHdaUjb6k9oNBkv0VVQy5CzbL3rh9n8Ixt/l4mcnJmFIPg2ZAhxFEc8xwI/VfB
+k6aRK8v8IFB5ywxK2sTxDsBmwCMQI2WBGrn/ItP6wmI1kuapYf5L+z2kvaivxrwRqQpcLkR9uAG
VpDW6luHiufN9qTdhqGK9YJ9F1qi9DKcq2FDHEsbyCvu0aHIU60luMBbYiWoHWiv/GH5xBDnp3nU
XpGXUW958dS+6o1Uzx5VhjNAKr1MRQ0WQX+mgbO5+cr8JAogN8myp3+mMKgd9RwXwgvGqQJniywB
usu2NDy7XDOIyipYtybOhM9RJomnLL8wkxbQUn/4R21hv8HuQkRSEJQz93jGTFw7u/CsyR9LHboi
gwlr3507xXkNH/X5gCwUG8fB4yVQQX0Eoe/Et2dURb0Dl2ue+49flzL7vQMTp6uxprncS3esLSha
aNXNwmKY2GCHMO2iXbF+SrtBxyPDkedDKIYSLma854QyCP50VyzoG/IbE6cG5/hPNYXpkth7+4Ls
BdMair1pIAUN1nqI7lrXq6Ub2C75j2bBP+tECb174A6sImAGlVb3QSZsHuh2cX/pwoQoCnUqLOAc
v8hDaKX86Q5xyeofiH3icNHQI3icwfnMmeZm5K/bu9s28Yzj3gY4TXm8xD2yBzibLbR9a8BYn/oN
Wbp4lxeM8CGSwPwktbz6jk99B7cgCaemX/3x7Dhv0x4JNiyE1rmVxWM5Xhu2sL0pC6zRG57VrKXH
3slRUwoYMEXHth/v6e/tYAOHF2QLsJN4lkgHd/B9oJpq3NbbvnH7XYWNL2v536ELmptzPB1nx8qW
sRw67E4GBE6qbW4kR0pU9ws3dEGwTNawQnmg1xkjviGhUPYXXkmiWrLHuYl71pjVx0G/BnpIfl9d
DUeVyBcDawOmu772+zb3hxs9ipg0o5Md0pUXWHw9CxKBsOoV1SXsF5ZKyc3bKOfUqm9Mxud5wV6S
l4y8bDMN5jacskTW2oVOiWmd46eu5UMtdFckyadgQd04beCeFLJqVx51myAqrZ/Db6l3WZnbtShP
cdalcQsqbqBM7sjSFuqAs6ji5MsoLIZkmda3rJTA+joxCb8NYOVZc3D1xCX4BMptpas8nMEnIjZV
WFZkMcqd3tD1xd4Btnwy6MvSUL/2MqO67gfE5KZerbs3zKgHJgI5QW4UKyqY8QNEh6lIXdtTuFlJ
bWfX2yPHRJgIJTbIK+CpOgbXRJ87nTN3bRHMaX+uye9g/dSdZqOwrLE5+vP5BKZ9YIkCeCr1M8pn
6+QxugzXB+wB/x2o/RhyB14doFrJxdSgDFJz+nht0nkdiIzJzfx8m2ZDkvsUK5WuhN/RKGZJO9wr
yJw35ap2jbjkfHspAT9LgoS2Ifz8YeB4+L3wP40oczusmNrrzVlUIBL56LZdfjYTcFyk9aTo93hB
LS02oNo7439uNs6j3fdmZ3WLINF92pPTJLweGDVpzcAiMKhfU2vdOgzUA/+aC9KFpch+KeTU0iI2
gxz2sU6Q5r/mQv9sW7U4KmtxFkig/UlkBu7SEGva/OYeNQ7oOpu6eWs89ieE3rjvqyYuuTNxY0Ur
MSnZ2eCiGgni55lEL6+m3GMmgh22sO/QUsvZdOB/6TqSUTfoZAE4FOhslGP8u5j7eKWfdLtLQI3D
Kr20ubuBkoxTh5rclSK1loe8TURGZHhmuNlzoqJ9bcAlXDwuYm0hzGPi/QsRDURlgS9Lbsf88T1E
MKHJbxRiispEOjKQkp6HTMCWzfYKmUNRNCPx1YpkEL8zVaauuLmN5Wg1duTHZxZz5zZ7mL5n6gOa
OY7Ny7kA5WSODN4i4Irsr7SuCw86R1fMHOf1jgeP1lPGg4iaxK3lsskafVB60bdMrl1NVjitLTmK
8Eq83e64ghENpy2iduEhB0G1ysE8VO4ESTWAXZyDx6TBBDab3Fhb5edTlJykihOfmLDWyk1ML/Pf
hbq/WhVSjSk6aMUopEK9hLL8KUJwsuM7zZQ8ln7Ja7iofaxXH5Pq3di61B2OkvzHaPnskrJUGItE
pfddFFcE/Cp9bIpS+rOToxn7G85HbGXIJpJ7iHhmLYRMX9cA+XE/tVozl7aSpBOw4T1/2QSa3H8H
ZCXbMb6XWxP7bC10LnSLEuBKi+h8eyavtC9So9KhmhXIi4WCIuEGdHWwgWoVudS5DvWqNelmVgd8
NL+Q8X2gu8EUxY0faib7RTdiwif/OXa3KwtXv0+B3aGIVjX6p+7sx+fEiJOrCDHEza5jOLL/rM/o
s9gMORz44USYRDGUeNNBU668kUi4Zyt1Pmo/WpnmlTn6b/L4AzOHD4L2yMymLMBIxti0wrVCw+lV
dvI4dRiJQuTiSsWT7th5Zf3qtAYfVq69zb2Gz5Qb21/KcZ4B/0BiCsEZh6A75n13X5bcjrr4IhX7
kanN7PWVp9+EfRZic3yZuTCjXERyGgkG1o3OH/XexCbgOGi5cwhEEI4TehZ/Dag2fjdeXXSfTLGQ
c7jDHsMlWXVJajvojwhN0Bc28EXMAv7aPyE0rLx7NwnFVeCL6rMzNEkzr7jdqGhr2KtmH550s374
Fb12VgXYDhw5Xw+clCr4u2ESpNnme0eIIVtAC5yhFXydos/XDtSMWlazSpMLmZhljr+hLiEnPgLe
af3GvNjVUvhMdUY0GbO+gNxRowN0XUh2w9y04yXS/C5eACcZd7hInLY4bUNUMttFtOiY0TgIJvJI
M0nYTBAGdXAyhO6RO7LIMmrlLELVBZILvnjsXMVCuP1ZbNhFhJM8yfNR9XDCghj2ZBviRf65Vb6n
z6XyNh4h790NjEpoZ1b0CtOU9ickoj5V8MBV7UABBH3xDI97uGDtC+RH8aLv9BJOVgZokoUw3WN3
oaxe0MdAg44tZqtQ1lTUc2LLlRrlP98w3w6iyvObMsyi/2g1qg/Fr8GbtK3vjPH7XTwDh3mvRuwi
Ze5A4QCCpqIRWEMsuWVleruxbxb+ukeM0Pbsj7K9/Ywtso3dCWgq0kM2m0vTmqkityWUs4ozHAAU
YaBRR20mi+h+9NjEC7eh5QWhIBep0EK4PJeA6A2/+G0SsZOUQVvIE3wcAKfBYr3CRigufQSJP9rJ
OfgNUzrlZbfeY8I51vxnh7cIUANmsNmu74QafhDBHpEm+olk5Cs7BCab3KR1PEsn9/CfIuP2qX2W
CvtUnUv9/tMb7w1Jxb8nYUU5CcozJFYsNAt3ZpK1I5vPUaXjs+5XVHiGGy6ms+i0ZvA94FHtMU7h
qkk2/xPRYcSna4WldPEr46mgAGSCLDd7mlTsRgBZ4kOr4VXtwtIF5oFLbSqeaqS43O2Rs23HF0Lz
A4f2g9GNM1KCkKTls4sGzbpf4IGN88e3o7l9pzqi1odGGyEv4ZElI4S9+2+mfsjhiXT4fFMpNkv7
KVDBKntT8YPTA8sRj9AD7f2G8Hc4OWWyjrTSvm34LMDGfo50fcKEOJb6BxuG3EVUvzZ1cGFmadU/
B/l93nyNuPPtKsQAZe3V3bLWENgZokvfxocor7DTYbqAajnCa4FcjWynMT/ZS/v2AADVm3sdOAzw
oRoWUXrXpjmoNud1rC30MB2ikIyVMBh+Dh85uQcszaB52JMaHS2pwv9GGOnRQ3+SZgfXPOftww5Q
6q8qcFDLE+oKUUXX4OLPp1nXK8FMVraMg2XIL+RwTLGEvI+Z/6PedpbyROq/jsND8fe5G22k85uy
u+fLndU5+UdEaknS0Qt0lfo679eJg311bRAYIMFyj4L+nS4llSYxQ9dbWjP7MoGkOYaw/v1sq2Ll
f9BYZhvcPbkLVL5UGz/4No6mb/OcN2wQ6Dbg8pRzN+2yKeY5gKSCSwGPMerdEpwpDUZ4usw3Hvu7
cuLlZzw4ETjCTSoBBGCCD+IqLo3Jxya+Pnp/gnyI5jdUqa2NwVxRI96a1+EFfcfG1kTte8S+njZt
RsSHNpN+iZxt2PHEJyiI5h0a+0FE5INReJNYBV7WX4kgZpjTkApDT0bHcYxBCYQfFGEFObIC/8p8
Fy5ZT8yTgu1IJe6RVuTFinzZ67bXnxdqX/T9St/IhGITTABDAjO0D+vKfq3qlNEW5H8t28DJxxWF
OKVb59efUxM2J+x1a4M81Clxib1tPw4zqdDPIkju5ry+mGQKx5tMhuFKVi14yq4NjMq/JqUqsfSm
xLSGO73uGJImEAD0pBFyVCE1EmPmXwpg4yzHyzhsQOaXDsbxQ03kscOLmt92UVWy7M7a+KwET6p/
EpqA034lOyBPurTTjKarZ+NJm+lpJGXD0KrC6PB2ED+RP0z0CPefzRQYRQgiOchB1UvD/oyrJV/7
t6ce9u/6A9EjTVKyc572pIIr+UvUlvZUpxoPURE1TG2K5J2LLxAECJAhfyNCAJSmnMCZYtq0vJAt
EaQts6ucJIs60BeoVthAMfeMhdLVIsXpZXc52IjWny/ltw5ziRV/ZMMHpGs+fJLCLmJNqBA1Hnob
iZB18Q4TL55y+tOVYOHIIOlijeU/bD+1LYW2QpctOPLU+0VYtXZo5DDvAZWv/zzMyajF2exceYoc
Y4nG3fpGvCCcwaStyN7B8gbB3jWiDvUtjJ0K35mobVgUwsPxcrb14gsjbZEEyn44lT/dtoOxxI7X
ctKssgBPyb6YV2nulmbl0ACdEmDZaMrxqvzCpaP/0I5eaE9qMtTaUFGWaOOlN2D5IcEeASTztZz5
6JTpEM9p4fZ2s4rBpNP5O4cb7ViBK1GZsbgt5Anu8ycB3b6XX9mPVXYlnTiRwjQm/r6cjVBjAcZH
Ok4SgwOCM0C0TETUFaN+eJlAPezVWYE0dfxZopS/OEYLzNaFK6ROPvEe1jZTSmB/j6xWpvZzU2zx
Ar2g1WGc7RpddqROt1HQx8NTNavjO0F62AsnR/0RUvz/97ZQifg6vKU7dZ6za3dhm6NATRVgf7BJ
CLYOmlgGSmaUQR1bY+AJPvWL9Ew/GZUpcAlho0KvjlA9lpYOV7b3XjoYrRgQCoR05Q3SjsiZamW9
H3JU24lWTCCYhTagF1FNFCyRhiMpfmsL1Mwplm1DiHqJPmDMPQMPSzNPe1pTDoE4HlGlpYuJEwGX
Spo120pubrWURxuPgFk+Mg/8uyUm6DqJPNQ3JEv0nEgQAchSnogvgP0VbmFS1BwJkxBa/rNARaZa
G5NtMo2kOU/o6lWg6yjZxU8IPlZkUM2UWy3Zt5sa6wfx3xz+YIXKQHUooEZZyZitSzZ/Oppkxyof
25JNfb6nq+LMSkD6lce4UfuDz3mjaqx/bDpUXUb7T7t1ad1NCEUuGQ754Mre9FdcVgI7QTv8JLZC
teV4j2TFbROMoJpJmHPZ8oXxvMfh5Wqaah3aZ/BprZjbXoJc4XDPTTVNnzTAyER82h3X1fSRQVfc
waestHQbf3gdG5CXcfIJQNUsx6obFMR4jnEcOlU5+oFoSU6S5bzC2yjcAp5Hst5pwuI6psQYXISt
43JuWvSnTTEr97b3iq975NyJJy75dx0Zg4pEmL4Pr0bnMiZAYw5unBaaHtr0s7CSQpiiyit6lGqT
CLG1PMv3tVEDkTBYNk6u21XCHv8BLi4F2tE4Hclx+X1qa7+tlK6YBVP7tpBHJRZyulx5euwzWZra
xPdWSZoIo6My2+YiRRAlFEjvBzzCvzjSv/PfeAGvZUkaQGdOE/2ge3oJq7/8LANqaDvk+rpQgg10
zpkA/DMKMuEc8L7UU6xh77oElEWEjf6Wvg6BkvXhJosyAioZC8NVh2DXBIy2ewMvdOla4r+DLVIe
tRIpop7lNvzSNtoNwOvph9OGoOGiJ4JDYNqv/MajssDnpOxdx0HJ/9F+lkX9zS4/RiuLBmO2WpD9
RBGKpVFxpT3vfuDiqiVCCjap5KIVyUTbo7WjEeXe05sW3XKJ0J3aBDtkUzYk+TM7aXFETrdmBDyk
t/SNQWpi4NFUygyewJl8pI5HjBSbV4NWamISOA6Nfx6jdsoldFb8ibxIy1/G0TQm0XZv9iFUc5IF
nRdD1zx0GsM/9G2cjzDQ2fk31wCEGyexsNTYT4DhwLsrCWLhbNa93FUKLBAS0Y+dpKRWpFewguEW
/InCIQqNwbO8E8EiOd+zdOPpcuD9x+Q3jlPAseNYZ2DK07dLIrelFIQS/Mzz+8iPi4FVlP7Vv6mT
BvdjGtzmW9XjjJ9kkMbl6kE1ZNmINrAQ2UQanPQDR8baKvjQpR5d7uecWiCVIm39FnyxstrPtxAG
By6HxGJyjEL0VsghkjQj1/loeT4SDsGwMdvNq4pAW1DU/obZVVIBMPJcrOoPh3s6iaJXPgfjGbZC
C3d4lntC/9ROuYCF+iq7wWNLgxAvDY+6MwunSgZlr0Go4+ietNZkX9zXLJ7F7+dnS/GpXYhoSed9
GlBmuC53o2+RDVJTf2nntw/IbJYhDf73D4RdfqnpZpSXIOynH5wU67Uoh6zyqbTH7vxo0KjU98GP
sD5hH28UHQQJaiJVKzgu/6mB4Mu9UvznFsFlljQpY/rg7LtAzLEhwEsgV8hnbpijRi286ZaobuZp
hmN5Gqv3lGjDdldTmCsVdFNZWfuqejK3GBpviqeqrH/8oWoYUoPH4LBgl5V+SojT/KowgQCiN1fW
6id6OKgwT4L9FljaQK+vkV7w/vXHQn+aM3rG/WuPp6eugwXSBUQjgwgrDLxSh0IzFChGJ3hVc7DD
ndvuQ6G0pf8HqAFQtqnqJOpMUxE24VAKrnjbM4HzGLcwNN5hhw57yxmIPiqUXUCK6yWBx5hShjkS
NJcLDUhXdyjr/tQAzKBTLIplju+MLyhiES7qRL/Qow0K+N/vqvxG6ySOP3nf7+jend6ju65k2KDM
YH18N5tEAmdwE8WV0gn0FQyh3EFfZGmMXJIR/Gzym1T4U3BDarmQg2CxJVtbmhJLunCVKj+XOyeJ
DpX0RkuYOl41jUDjftFmLa41q7F3t23zkh3iUs0FTRQy3CfW45GobxV0yLcZUaQZz6FBmv0Iaa1s
/esbO7MXv5WvetJhO1mY2lP6eLx57aFTuFTNujNMkDsJpyE148hrhyWus0TKc/8dOjEPRyZGcJct
yCkoj1i2PBgHVo85BWBtHOknaJ0vlOUlinCcif7ky/SJtHYmBV53jWW6b89aEZjH2QtZPkfe0qKv
a7c9xM4Rxv1hGIxl/AZ+oZJYogeEScy/uRzt/FbckJpD7rwoapijHfd/P6/0M35TrqNz7Ifz/NL9
qvIryVs1zf43x6eNE9Fwco1fR8kmqcTyhmjrsTuaGTtsedfKh6U1r98KmNsdAaPJF2IUhKP69Lo0
eXmZUpV4EI+5jmdZSTidZ915FbPky+tKhGi8Y56lCTS5W+M5YQoNibjKmcqNqRqjRMUF1tS76MzK
fKxns2FBayqHiq83eBSGdxgZfZTcfpE3EUynFgxBfrQ/h7fTCI4Lu/F83i3nYhStRyLPuIuDkYZB
u+BMCEJ8OhYbLLlyMVTne/BJ7yt2awTBuISAdrFb0H1FZbYLh3ddeujSrOwrYZoCQ/05AgOzgUGw
eKBvrnu5WmWOSKpCb3POVMq85LlEX/zQne7sKB/NHgdc25AL81fgj5L5Z9SvEY4mP/03XGJt/H+J
T6j05KPrgbhPRVunsXLiQFw7XgKxJ0FlSN5LS3qtQlXQGr7nf1pZRVIdMteRS+h232OnnW3dJtsL
OtYH3ERu5/gCDI4oA1cRwpJ349HU5lvaIyxq6crLVEVQLmaYi1i+W3nlPQOld2TDOuIeOdjNDJ9/
giuytXN0obU5QtcpwJyxrcmyOKpIbGIBeDdA92Js2YmSpwpJ0xwVP5h8KOovZOSNDT3Ozd4tPXzV
DlEQPV9xSJ2d/rMhoLazD0hO2IucgUH17ZtaKJ/j4lcI9Io3dlVO2SrYrqRrYZdX76D+XIbfeaxn
7o726yMp5hHOYieHfF57D0pqjcmNPUN7LereR5WOhek+/A68s5bG8O7+OvPttFSfjn81ePpoZMg4
3fIJTDzV8OEn0FjtxrEYxZrEK/JffmX7d7I8x+/gF3iT4YLJIKdkoG4s1xmp0JnxqUA3v6QgWp9d
9wbHsSmhF30iFRuhs11lCcteVsuY8UVTrULcKpiK/UbOEr+hW4lJt143ee3XWZ0C7xBoF4LzdxeI
vrp/lJ/r4Yt5frl7nfpFwLEb+hKjtWK9Z3uHLwTMz+5FASdSugIaCr7f3AlK6idhWkeigFSAsF0c
Co255oUyw8ug6a+c4EEPTkUurzrR+T2zvGs2urAi11jQsZn/i+1ppKcN7O3SaZLCdGpcIzWW6MdA
fdkMnNmtIFFiHgWdhTUYSwt01jyvZX0Rw1PvAXUXGwj8ihMzblCBWUdA1i07wmekrjhjtjyU0A78
sDtU5TwRxP7uh7S+lzgPKzQ8u3MnuwcIVhP+/MhXqD49LxfMdh8G9HJUoP5EBbFzHtAPFbVvka2M
kiVZKaRvMDWeP3HizejT2cDBlgS5pwG2Y/yYijk6Aex6DIuBbg7+4EEVIEFkFIxpA960YfJImtYp
GeBy1wQWmn+ie6ECWJUTPjMMaM7jzgCWcZ+IZ3LVrQ4a3Kcrbsun6WShvDXgbThSSfImB1nOBc7m
Tk/+9LSELUlpfstBWAK8ctL54wT3mVT3/gzcx6u82iFLUZKqR0AfOjvMO9zwNZr7rqtJGmibeCWc
yetTAf8iSMpin/Ujq7szG82xCg/fuv0ew+C+EtMfxEDRcWd4yB0UPHn9BJyCPKOOzMGbf7LMrRpg
DfKGrrtaRjWZyFkO9n6yUnNSDrO0N6QoJZgt3md6bdXhyRqOLIg8tMNcSlHZGa6kigvcB+1ZugQ2
Gn4a+amkGpTtTUlw6DWi4m6k0MQVu2dGqVIjKEjzl2v/QR8C2gROkQyD/QgkalTsC37VsktP/uc8
pFmgD2aGONjmp2+qBGbamcmb+y67YUCRf/Fzwb6qYGqM2Y1gCMTOKoVxNw/yrbWvAYHNPP7Ye+6W
OGZHnikTFoDLoir3BwyYcqki/HDHbGTP84eKcByt/tKpbsjQySO0IsZqK0mK/gQgMx01QEVWVx1h
NKvXJYSP33x6rzxi1ixcvatot2oM+N7iQQnqz40FSFRiFKxKno2D8mJEyfXbLSh/BMlozbtSP5wv
TwLaIlgbjYIy2xfra2YZQ/NxRiLAHlYRUdTksTPpJP3mmWKOn7YGxTyuAoiCmhwq+KTLJRlSi+wZ
gZ5aguQflkIMDgOzJuHsx1NDzK+jsRHrEAtrGJCxcfT3XsZlniRgx/bvgMZgMQnndTb67x6KOF1y
wwXP8GlJU8wNRQH0wbWwubSSoX5LvFhtIqnowvaZKgipb4dX2bjHoV/nsCN72pksiyvamm4p0Fz1
w+R8LDwmeAu/ZGAQNf/H1sIp93aHs44D1Vb7bskUgDCZ8zA498ovX5B6K47ovYtSMK4HZbI03eQW
7gOk7PVmBqxfIDFENfGgxDAx7qyNzyXXOd6kFXfGpBTA8LRrUUmatvVSSeseh1NfCOTQoIdRXSD9
+VoE3mxuTxPIVxARiTdWHTqOKlIp5m8vMsW7rh2pPIYvXo40TkXaBC1ep6kKpyFXQToIy0Qotcwo
t10fD1kEsyBi/z3m9+Y+joDYPzKi3qZ7snf2rui6hZtR9kaD50VU5chS1HU0mRcRxhGOlYDImBBy
HofETITb01obMfGdkjZyF8ikBllq2PE5/+qSc7Nx1RGH9v/7xU9sTNGYypW58G6H9G2KFMaewOP0
K+keH8O12JrGrP5JEJcjiA0fdBAngiAnokAp2Y6FsgHebCcOsG+dj75mQQl1Q6OhbR4vaXXprMBM
SuCSP5RorT7FVH5ODd/TilCY24bkwiTuJ4TzG+W2lHVhjYw63Zb72ilLYx82vtSMvF9691qCSIgh
E5llJNyKOuNzk9P9pK9xeLcMfM1UQ2CLuGUQq9RTcTaQ54NMXQoSBX3yZ7YpasuI6r32wTCMdrnC
8NGRQI8JpAwDW7hohWRgiHkSiQVBWE/wJ2Offpbw/vIJaEn/kmN0y4uIaWsbdq/xIwh4ErJfRCUZ
MrAs61voS0CBhzCRABfKMoFPQrVQXyiBqyORlDyJi0MmH9Rrtu7VR9f4zQrL6z0g0KAmnY7iBMOw
SXIA8oc8uTxO27ZtJvs7ewXI7eOO0noh6iV8/7+La3FhsSearTZvefs7OUzfZqbphXDjVN96CMjT
nOClAjxEG217wteaftrFhNnf9FAmJBG5WlhRt+c+a3oHeYyl7WmdEBe29K20d1JBAy0dpuP/xEkV
2gC7jK22iabgfyoJIRzso1U6SaX8neljJoXDOTiTS/vhRIW6cTokmilLvipprxMKxuZe3kD97Oav
jAVpmDpM3MCTQbGPIO/P8qQorM7RwrLZvg5ougPpoHRCkH683jcdpfOthBkaqoAhQ0zqAfBszSw4
ytuPSjyn/fOExLfGlR22rSB7x2vLyt6k66V/zXhRnWmymzRrGOtXIf8Gv+G7tpNhP6c3TCCJFGAI
7pYrSCOAoZwfQ6vgB2arP/suhywnZGus4m3kgriwFF+zTsW+thv2rQnLLh2v4Njj08Lvkb7zeJB9
BEmwO0iw3Muufs9Luo2rtsJcTgduuRlhxBVIqfG/FE9R5RW/UyGX5gokeLhQPUUNXBmh1po1fu9Y
InuZoB7dnYpR9C4JLPKLZY25Id2vbXjDbzuhCCr06EDJOQGAfhDdUlHE+TxBvaBqvw9CXxnXcgZS
KNrywvoEsah07/bdMDF3TaccXRtAW/isHe8pmCjRJwGyT5/YFveCnK8nHEuFU+AJrb/QIIlXkzUT
m7Q01b23UDXo/gL+TXlV0/JHcY4U6LNBiG7ZIopWAXREyi1cxusUGp/ttrTP0JxQeUfwRMd4azpX
qSzQgZzI5LyWKo1plJYBAP/Q+GZsnukd/BPxF2aGktTNkq/rN+EsBuFfr85GVoeMqiZd18VgmJWQ
TxFagqaeZW0fdi3bwF5/8Ujd3TalDsV5nASPS48Q1gU0UGkQZSsQkM0LY2/kh8zw3Ox05Y0Bztnc
zep7ygY6xRHsbXpYWuMFC4zO3+w2UmkifUz7X4mTYSPILSghD6cCM9IrR2K6mVBpvYMWHNYYobxU
VcfXKm9iWuVYLJZPL2wJb/oitdp+7LSH/TjrVuX2rrqXq6EeEwjKz0dg9qsk9sBLciSAr/5VQ5dc
vWArFSP0y+4BRf1yCBSrqzNtY0ydZSoUszEiSk5P5FvkiXFdxUhq1PDpbEUf7TrBLBxRuf3qUz0p
BTSJJeouXgDWHlKLWUdN8dWkHFIOw6T4zsAsUkYuY+4nsU/9203uVvL3kPGoM6EogUIF+xF57lfy
tLS7a7MUM0asGI8Rij4UZdO8V3/Rv8XSwS2XBVk/n24+ySto4TWCJoDTD0kRqgVbwbAET+Wt66JJ
kZ+8JVfb59Hi1e1wLHlALKIA63BySbjXCAk6ITWQUOKVCveoxb4XVrZf0bzxXhk3aLEF7EuiWocZ
e+8sgFmwN9u1peFz6IDAig8AlImaN30sllK4iwRLBsXIgGlp7AzrYXhOjmhYzjOHYHqJB2pWSPD7
BY9tDEIFBvkGL9gcDlcvhFJBmV4hgN+XUTa3x+FdYX43VbaeBspNbdDYHEbsmuK0ZdxK2rJGTVep
Sv0VEJLDOfxvY3q7Qmujd65rQuum4xLHpigm4EuZaIZw8EQySy71Ln3tEF/lTHDpMPwZCgjRJ2zh
FBGksnck0AZIxtVEbtJLYGpxn2EZMhDYpHMRfcJY8JOSi8WLWHGxdb3gKf1dRpLZiL6qQuyMDsuG
7kxvy1XoAGaclOrdqWTaVPz/o3CFo94hhnYuugQ/1X79Cx3kx5EDfwxx1aE1vDHqntdSEHVOkR7f
koL+1HwZpLqGpVGag69bgwkOryJbbahVUhKzxx7Fy7G5KCN1v7RkhFEPdtwBixbuWVnq1O+85RWb
SgN192gvdUU3SeOFbHQbq4Zl0/pN/fc0mc4RLSPPHSKHkpA23ZlKP5cHAa8Zszm7EOPFMYHov2zj
C4x3SgQBp2zmfMSoHZBzx2DAChll18ij5DLc1Asz/lmgcNLJf+9jamzZ+GnP89vZ8bR0VOdYwBvR
Jnxe8PXav1zXPR/Ubs6Cp3+Zmjm/W17WeOvh9NbjnxkRJJXxBCqXhkFANScd6vmveLRO2A1XwlSH
6Wgtve/EPGjyVGHLOTzxNVkPpcCRNc2SFbLTMP/0LlVyM1H90aLR94gy3cM9rGyJWU1ts9vvuBoN
u6kurq6xMC758pJ9ozRV8SbOAxNv2Yt/ON4FLDGmNptWCIs2CGBzk8PqXirC/HakDJ0szU8StN8p
D1g8yWptSltfJBFvk308taxddTC25nJxyGtEsSmC2zxfZhJR2+Wbd5bsRxK2FbELKSMoImsmN7Xg
L3lezauvFArdx34cf7GHfPqCZmlo6C4S66ekyGQBy17yGjz5Uf95fjYVM73XeRX05HcIEN3s3pAD
eLqpuf76rzHtLjeMWShh+O3bmMK/OxSjnXeyBfZebznmS2SXTbGCGNe4SJh/kti7tQVHrEJPaNJ6
E/JoMw6ledS7bRhkx/rguDGURXdvYtm+uOSR84eYpDZAbVhjKxptcSiTUJGxZIsodYEBX0LN8Y3D
qe0Vg+0lUpOQQlyYbqkcCguaKV0/4yY2CGclZAUsAYExHa7ki1llrj3F7tk6RH/ZZhHvdHCWjQGt
C9rq75EQN8ityTZ8jiKPoZ3FhlD+qZRZCEz/kss+XuZI4zFhEk5kURntEpQa+JwVZ9aNZcnv7ou6
F5gPRdMmQ4U/pbpCHVrnwFhaThJ6N0M1CO4jhKuqxGKgp5MNzbxu8CA36oGCgWkSXgalgOMwTR1j
gc9mxFKBUXgVyEeYjSm6d4rMxcAC/9e2h9HFFQGbiav3n0zc/tCGD2OLw5ADpIhoFKdD66HlpLeF
inKHt2ym2kyx4m6z94aKQVVUpqe79uCFXamrZoDJN/wvizevKpGtHGNyTAaXtRDd4x4dGDMJsQ+7
knPk/FJrfNTSpgMK7zOt2kpinJZxDjAZH6B4jCYH1NHpvn+uLGLxtXPuEfSMLmQornYWkcf2Cqfn
Xoaf6gGvwq3J4SMM8mi294FRFZ55LKvnfI+tKwMvR7Pp3nKl3GeWpEFaanXWJ4obWZ9rLV09Ad4B
FyRwFx/Xx+V/wjBki5//oMZrpGiXLSI3ZEDAXyinuwqV5rg6y7e/+uf4/EquG7ZyXI5JqFVx/lhg
8mJT7ZXchhfqsUOwMaPFI0W2k4NgHm3ehFX7ibzOLuDQv3o7WBWWGKAVWzukxc3HSBfWUZ/CYgED
JSDjVLHSZmZiQby1tRQ/pKsonnkD4wkhNykCYW5JYRAN7qBiayipOIMFd7WUQoy8uZzahFTOTaCk
nvPieUOQb76Ke+SBrn9KnImE5Fw8dP+EagY6tTVoWcTr3E4eg6ySjUkH3RwXn8vjT5//pXnWj8C3
dDP5+WV62FjVAtZKmfh3gfRQg8oS/4niY34Bk4WpMIPskD7pUD5VZeZUOIzZSOwVgbW9esRRw5g6
msG8RDcoWqsJrqtZunyiNCav0XZanEQ+4Nn/JICBXuVVj2l6VLUatbpH09F9yH18/9ax43WHrGf7
ucczSr3uuHXNiwpTsrlml1KAndnaU1V3oKOB9KX1TpClcqVF33+igJLI2+n+xo7f4Z2+CpzzmOTJ
DNAnheOliBNlZua51ltwWVv49kQVFAm6+Bstk3G73w7gRZ1S1EhIX1KsXu+O0vypOpmxHOEoUaB7
g04fObpnmgWYcJLBVwkc7lmq0zFIXEY1QuwxcxTiDjR+UIgndXsYztnQ4GVjdzBqGAurfN1BPYSg
ikevCx3T3Oqcg455VRqoXFPKMUTuZOyjrDDdxoP5ovbm7tHD/w8jGtdPOJS4TrswVfw5O9k+2q7O
1I21Dlto/ThSKoM5i5q5DtMW6u69QXRuZXFAMB+jv2Gl2VXzNyXVb+pf5YHCCHTEwBjQ0VWDq3hF
vqjn9G4C5HQrClhWJrTcPLKsE3VdXgYB9U4A5rRL6t1WQpd3MIQ5n6L7wvFa7g7zBydmlUNq1rPb
Y5RKGRKJACXQRtRimTEDrLxeQPmY9ofnUm+xj/Qo7AdmNneqCaHBFb1Rbvs/HjUgEgvl/ICVmp83
SbU3/uDa2jr57Tz/d1ckg/6ENlLIjj437e5MC/uwaKCi9Y94/GoYGMj4huXj2lgRaMIwRVXY8tdE
gd6IuDEBfaLRXdjm2XGVnnqDt7ifBGdEyHLZNPvoEapFDsE6tK1s/2zANiAMpURpRd4cX7cGhR7q
eV7CX9Rgy6FrZ8TvrHoS+o7+K9yTHI5vYVoGC8xzPK3sm2hZYDIkbJGBpIRusHanxV0hXZ7E9xVC
Z37UxqLZg3V47r4UKY14Xy1RtQ6ooytR+vmRLb8lM/H883eIabQkuVIHGGpQUm6UuRfe8sRf7+xs
UK9Va55+GboSGAXKua6Ay7BvLc31AAPYOZFgIoqBD+t7Y7+O2AcxWmxb4hHnjah/1grCC0duYFMi
a12zmKMpWoRjzsDvPUsoZ+TkdhuCSm5Zgpk5/T+hQ/vNHc39/OHVTkqhAhAdBYGrHK5SILLiLyj8
99RXqdtiZoKuntGRhUATqOGfzZ2+NHdZ/ZtYxNgjY8w2+WOzPFu2UswzO1NITJa1PY6e8hs0eAJw
fC22BGOl2HYnY1G4v9NXCD4FdDjI8YjhpJlKxXjg2mdMudOtGGkjpDUxDLgQieyubDXXelS8PEyR
b+Vb3awsCW/IvGY4XkPeENKF0upG9jv6SA2UStxocRZruY4VGWzBUUeN7kw6ynzkgQ4KlNNV8Oo3
sVt9q7SH34xqHDqbyb+V3R7oddPvk1MzWzffMuaVyVeUJm/inu3Oe/c+4pIzAr+bYUnKpHlFLax2
zzACIHBKPReoxr8SGyH1tDYWgM0ut+JZbExBXOryO5YC77q8NoqXURogm9Q6GX0Ecz8Xsou6/L+6
MDcEaAQmhG5aAKZSn9KqJybX/CQjdPXjh3ipOzNLmvpgD5WdyXhiWUPnLoWp43Ed5TWRDXfzMrgD
Bgd3326FVZ3KbQ07L23HEzMBHuUIo97IzFJSTTShop937F9fv/nSs1xtor+J5r3SaM83AuumFRVh
lZb8cKTr75xvAmY4zV4J0UW5a8sNNGiUM1Moins07WKp8KSe1SpDZEK5qjIj3EwNv0r7KGZDIPIc
1IicVjiSDcJhU+KsCef2BY2wQ5UBXDCAbDDvQGf6ZjZAnpKN5yc39M8pR4nddlMypCBTR4X03y1C
BFxHF5DVNHodjmiNIFpvLft+bXd0pnsBz4cRfHerSmBG6dXTOqFOYNGXXI+dwbwHRJTS53n0igQ6
HLV4FuQWYh/+CGNTMFM7kp0uOWf9PvCoMJCgRJfLE2CDZihkeoTbioZWyBG7KcWzVvY1lT8v/VPR
FlKsTT+zjT2hORjYDlhCrwXfPraCL+Lr0y6LQyz3sV5bNQoeFI61Jwx30934hdH8LnD8nrRC1Irj
1hNpx6OxjYbmp6GSpK8mL6QaNbFUsw7MT0fm54iXL8W49czgntttCk9VOK9uixosWZmciMN4zEWn
DrAs92L0YXfEtiqR2iyvvbe/oh6ifANH7sMv8cUCU5FMU6G8Nj2t+3sGmOK2E5nysTQJPGgeAyLO
NzZFyXlcpl+iIR8l4zrMVr1ENVjMD2f8TpfTUpFWoH9p6qJ+DIrzYlgoMAk3KExp4tabNocpOqLn
efaIorDySthgBgF9JNVZ6lr96GsVkOy0x6mwX6TNPdRtKgS9RyT1z1tjlSu6bXg0/2V78e/qaLYT
kHIEL5C+7injIFJP6HNFCOV4vl3hJc8wvfeOy/ybguGAHLaiEa0nDH9hODHhmFe8XhfcTNN8gba7
H91zezMkS6+5dHOTiTZY8zMq0nOTQbjaQrVA9EEU/CEoEpyX8TlPW2ClmG9R+m/rlDjF4Bw+VoyZ
mgBaJQvpAHqjmM4oUQJWFDOLHySPli7vSmlZ/ewsARv0G/pzbTglXIWgiPK14k/NunoClS8Ru+u0
Rkv6XvlJQpiQYvKVIhwtO5f/R1GTtSUzHCa/xwheVXUY+PKBvhObANdC7AG0R9M+02WT+xtOgv1j
VHDpkEEL5Dy2mvhgq+BpP7HzBBDnohPZvaqCO6L9jtLRcQj1z3C+BsjzGmp9Yiba2P7VIxhiC+kj
7TK1rNj3a7nvolxrJSKOFuZcEmS7leZV07BsBjeuttnTlwqNr1szLtt03WPN6tldrkqmbHMAkD3H
rwz4MQTl/TA+CDWbnwKgr6YcqZPz9Fw7foVQI0aOIWjEZbs2zwJpuEahghR3tvFonL8ZrHLc0Jst
RxsMVikZuoUOsRZ335081r75GynBzC2szBzZQ5O7ouTN9z7ocLzlOvmXrqpS1r8QUhEzWU/2r5To
GGUNCKJ8KaisGCKeBjqunz2H08qsr57mOone/SSgSffkRUR17ZnEpL+zTQTK+MoHgTEd/XuHznnr
NrjGkN9S+7S8bQ9ZKy3cuPCkG/c27mtUuOZdtory1b+1kQFanZLv80Ug2WpCV/hKY0AZ2K2GEMbw
S3opf2rivHfzkxx6y6kw6bzYhXdOfwgmCynmZmuXsFfiEFkS4D9/uu5FnWMXvaaLp5CjxtVRb3bc
A2bEaYOR5JfyA1Gz+3HoCUDKgcRxbqwmZ9jCijE/tIQxHaWjQ7lJj80Pz1O11n/RqvRboBjq8/a4
yeLDxLCotjCCZrCiSTFqpeGpeGx98LOtOnkT9ZShswtzi8vuqTpXSAciwuLWFt1DTInJ6EOaC72A
sJZwoRxNQgO1nw/suQLXIiYAqXwOAfVkLXqfAnHEHvJUnqWHfnlRZL6ujAwics6HW1aPLweMU1O/
Lf43GYHbjEGH166D5qdKruAZjvBH1J24i6HiXeS9UNPU72zjYVwwU+q/PuhJG9skD/q9qlR3L1so
/+/OWFkaaW2uurIT9G170kmaNMDskD0oFA/PYKMUegG+KMni4YrKMxnUsK3R05r/rMRDUd85xSi5
eyV70TFA0k2uXNni2yf+OdNZw7kU+XR/PtFhlMXH7NLzBz4WXGDF8kCPtpF6NiSad05+V6CG2IUu
8oMjfIzDD+PdWn5RrnR2PEJcTp4kirNoB/oS2jbVgAIstMnZ6BPYvHfxNMryrQc2wXD/PP0oY6Gf
Fouwvw1KGYyL2lpU+sk6IrxSngqmlzt4qxGLmzxoc8/e9VD4olOSJkqThfProfcBrpXC8Y9CQF0H
YNqEr/0srHBXZ4bSCUpmVSsnzeK3CNCsRaWOJ/nEtwhy/3RxqzMADl21HoiqPwuO9BYAR5xsvMfM
f6l0vLHn7VEe2rIVc0EmycsxDIMm+eTyXCBpojg1UHp6GwJZIomWiFqoJvGTrTgvvoOC1PmdRXZs
gpVEQXbV4std2X9BovIE3wqWyiRNGzMv1XZ+v1S2FmC+TRjP+xYyNeqcH24+65YuJXscfcWHItry
EzTOxny0rzM8D2xMeXZFI32hI5iqPRb2+A9OuKvGjLa2kwF7efSAEwgBlJHhyr02ab8mS65Vd/6t
jiR9djcQZBixuGSoX1EfRP8JfRyuiPi4iIv2xlkqMaH3msA+cis9FkLuJRGjXOCit/AyFTzhnco0
zSuv26rSlR7vVhcRWKu471qPOBPWFvY2ZpDNmhG6y1JRC5bR+FViu5Bm3OLLRzYFw68WOpdESAIq
GtzJ1vbTp1A/AWwIa0DJP2xu/mYqfFBNf3NKTxo3FJDGL3CsPv1JjnKVzxXBmySHTymSfXQQevJ2
cn9grMc4B7mgP9Q4fxcfY4y3K0YqU9JdWCja65g6dDaSLsadC7M/RELvdYt5w7rY3BPik8zOlQNC
sWxLWllxIZzmxEEc6lFVE7+eQpiy56D1xAe1yUJRoXcfFfra13g0a0Rtll9VYkXe0CGyRrPF1Uj8
PhXArSBOUUSy0y05SQE4oagoO4R6b2lXRIiD59ks8LKDnnsvRnUsHVHsVUCFWQhDyi3/CK8w+D+1
Pa/1uaR68dFNC4fQhQbD9YSdW8Ii+U7YKAOPp7at8Ia0zeEjAcyu7O3/a4gV1yVSItQe41GVDU8W
3IXyBtzmAGzLY5q5iuGHUj/VAFT3fLWcRYTI6EcAUlauWpKQbukNDBhJkcxhE9s/ZcGoEh11v+Tb
tAGAL437/Jy4TBJKxc1lAfdIAKmyzjD2pXNZWCLGKTuq5K34VhwqjKbSroRHB7CI5gGlYE94OzCk
a7qtjl5xr/06lNY0hKLMKVzUYdpVMzP9SZJn1wFIsNq4oamd7eAqJhpSctSYf/Wr1HeSCrqsSg5F
SaxDa0un5r0dCvuT1PIov5+9Rs3I2o4YRcsJthdYwIyoQEfKPuKo7iaNbgCGU18t2VeJf9QBWgjL
k1gwQh0xqgbSliNCEGYHevXzxTsXHj5iBiRB90BOizMQRe7C1gAB58jpjeM3/o43EWZZKBCFz6nW
q7IX8DPFxf7+kV5ECezIXqwRhfl0cthp29T5zJp2r6BKIzQXgrMaC3ouaMsUNpouktLtwMLVibU5
aaXGr/AbalUzi9qDfB3RGaoj4ONNmfycMIMT/be0pMzsfS016a8W0bkY0isr4tUj7pHWrb6Q6noD
Tu/J2a7mSwq4y6j8u5ZboiV3xlauLLLNAwGfmQJg/Oaf9D0DR5c2C41vWrX8rZZhCIy8qUh0c0dh
2QG/wZF6M77e+x4hqI7OLFKDFuTsN0Xg8JuJGQ0pLypMH49mWOux3dKM9ghOxy/Ie7K/yg9hxsYj
nryjQeRBcFbaGbEsx5ty3muD/rg4GZXrJIwY05CsdilN5hYqFdkDU+L1tZoCx3rrGxVu0PHcN3De
N2Wpul8B6V655ESa778Yt9ANUP2LamL6raArUHlI2Ki1+/UnsebZd6A6wdCea0AliFzTxttUIOrz
nnlYwidLwNXmC7+ib6BFR2FC65j/Ydzd9f84ur4UWUfdU/sr/BKv+q7wEeqNW/+e8J1MuwVYoxuO
B1ctxtlgZWyQp/e1gDMSlRV3nS7U8q7q4/a9tNRf4GK/hiovKu/h0KxH/oMT3M7SISaN15/YSsyr
1d9BS8dV1Jboc1/EsEqnaL4urfPO7WR2XNHzVBqqOyxoTzH7ZnU1V0N7+ehJ9Ey+d8Tat/KAVwKA
kZFk9qxF2j8taKqUmh5zBDsBvUsZ0OgoYcj+DP0GDhw7yIbrNKo7XIu/1b9IimYmBuEQSwqX75xE
aZQ9Ckhji26MRqDokLd2Yf8C/KNv+/b/xiHE7illRONYuqO7suMzdbgieEXDNGwv3KecsM3B7rjN
P9MwoLRjBR9DLkI+ToR/L7gTZ9XYSBww4r6FpJSkEx7D9YZtGLwyhLdNuk6kZ3aupgAwUxQjcnGD
zQsaf6boSBkqCGPtfnzQa/GLKy/oqBAeoUA1AzDZDL3Lj9vHp9Fg71mPwuFGPyWkflMsB0jlE2zF
JwMG8DbmB8eFDV+gDIQ+S1d3mn66KIj3cPBpR6+3xfl4TWubGNVo2xrQQOaHsYj7cM70SToyI0Bb
c0b0SAFxwbOUh2PaAUU8JLi6k6T1LXi5jU2bblsgkgdjbXzteUiiChRf7NPxd5BpJseNW6PhGTLP
7T/0nrx3LyFob7iBHOD/459VzuGV1jzuiPhy6HCL3h5guT//wDEly31ilIXH/93L0VUJ0lK6IZGQ
snkiTXe51x+RiSPHaWpFB2VIxHeGvHpj7aiyZ6OSbuyIPymyNgDKWYQjRzALs06uQow7mEoQiln6
2sIag7oi9qTh8dCfjSQGw4J/v/Dab2jA8trAfxrS1UDBrY5aNRKNJ1s0lc0kUlrr0k9b+ocNjQSp
JagEzcD9YEDji4PfFPyKSe809Ho0um7MIKj7CxFC8uCnV46ltulPIIB0YWjtDaWidopTxTJ2Nnol
IV8cUpIE59UbOoCtdIg2c6k3/IIzsdtOpJhAe1a0QI+T/hTsrfV9hsyBfqODPCN7XbhS81Zr/i1o
zhFWHC24gOidjvJcVkOApDnziYy6+pcSmQePqnJ7bnvXXp0R3pdPPITBFhK1pKiF+b6IHtUwCD1b
U9x4gM60TBTAzD+pqY9MTBsKC+GvRLo3A4HtvGoaGcrO1zEJNMErWFD73FjVkoLm+YDsUTnpd6w5
1CYzUly37ObbOMP5V6xRzgE3ZI5y4zAkqM6lvTKRL/3XQnXOrUCKeGQpGWcHTv1qib2KVGCIlA9Y
+uYzgJxiP+JTwy1746CopM20TJGiAM0PposueaxspDJU5QpVfgdA/Luxy9Te8mLo0OTZIH1TEbOV
V+hifgS1DZV3don5A1ttLXJEfkNiKvWg30AV8Kwjv2lvEOKWKsasg71faG0yj4TVO9UUAfqzz2Gt
wwoUmjAhlLaicX44rGxuNcIJ/MvOJw7DpldJczdnOBbMlLnUXAWq4LLWU4F7FSic2mZUc5p1qjkD
03IQuqEDJ20NoKei59dCE4epNyvIlDIkjxMej+JTyzerfC6DDZiK9BMm8vXZbdiA+yDRAozRSSO2
TFBRbd4AY7GR3Y/Yo7zacCoQwMZi7HFdUwXjAhCvPcifE7YCpRGBeARz+3aDUBj194qvJqcg5JVi
iFVvO6tjEMR0pAnFVEdEr7wRoaM0OuDfsPQsUJ7U6P/SKw/lG0/TgAJjpsE6fhdjBRFe2LzO7ymK
3KtWzn/IC+MvikaHAbJQRqM3GinOmtJ8l7iuEzGE7jX39+vdf3pgfOhZ0vs8XSEcADL0gNgp1qAa
2HzHmP9mrCM0L17W6QQ49xkLT5uhtQNQdbY4fnOTnoNnsiilXV6mlTpqFQYM9WnGpE1Sh8RKaPxR
Lkbz9SLAW5O3tVkRM2olvqr/T2c9kzxJYmTbnp2dL8GvZXq+IVTQNBHYXOOTkMDBDwAx++giLhhS
DWTk9Fwyktl1B8z5+m/o9ZxXLXCqGoQU22X/8HLi+efdThP9hRud7o+jN5QoCQQQerwzWQYjJfoV
IT885MHdqr3XwaM2+K8lCUhYpYQOTVqn6PtteLtADZewMbmEDqZwg2LpboCEfcgALTowKlDB14ko
XYPM53mNaUvZnxONoD6DomygxYugZz1AG213Tdt+J+yIhqq/FIaemlMiRr9ZsEP6mYZIk0dqlOqM
y7ef78yHbGE6cYeYjrOkxBWgzbWhR8S/IWDygauVy5W/IeX6l1jz0JjKKKkrA30m/aiURrJDxa8O
ssTpjJzwzrzTXx0FhOUT30wkz9YbMQjVE8ttSQkIdXHiHO56yXgVIDisERxSC8qBgNfqZLJ+3sAb
AiG/l13SeUgz2bclPHZ9GS5AotfDcjQ2Q8MWasqOrgjRkt8Aib9chje4ESteRH7ZPvlAI/Unn5pJ
cfE4TIBpsjWj3Ck3kZMkY7IlG3sCK6kvns5CNneo5LUdMrIfW8ub4G0Ir41Idw3QGUP2tdWH5FVT
KKn1zashF6WSi5F9hi1vBre7BWxWnZoPAi0PzZbzcjy3LNKJWOIRjon0tkiroC5CEc0C7ndKNI0Y
CvZ/7jphEghSUvUhy4ZfxXYkZQDENVmzyqewZA1lTjHsyDQKeXpejdvTfNQINgW2gFmUgsBJis1P
DHSzQzqSFVAHd7B4VznusInrDsWnj5gGFzxiGXXawSpK588gLJqLkZ1ntCH3rTRTo8WeLhC5Nl9O
80XAErN46Gx9PpC4NhbxJw3h1Rm/eJHeTu8ALzAygq54nVRSTLBmdtT76amXwwbH/zdgrumAJxOS
wk5twxRG35cF4CaRtfFBRN2kF6C8l1+npCoPXFxBb3eMEVFWtARiTC35BUsl9SXLczaP/MfOtIfM
Nzeh/jaxY6GuGqFaLH+T0jBC34JeCF/3L3JGu11IeT0sZ5UpbfvF6Fw8gMQHLd7d/P0iY7Kt5qv3
pNYmRATLHZEHjAQ2k4UEqBtxnnkCQ5KO74liawT6jUqvz/NU5pHDPhQL4ioG12oTLhRTYbrjhqio
Fu+JQO5t0RgYdMFZC3Xfu7oDBAHAMUe7dEPvjM0wJ4WHhG/Wim/1IyrY6kfU+QioWsR6o38pnSic
HAU1n9qhkVE44Os1+tIgSCXcLzMKVW9FdbZh5TKD87A85HX/CB217XUopfwyHIa4EFAUSESqff5P
jfJqK7hbrfw9ykYkhitdNf8R+6h8ek4amOo/4YKezX4N1Enk3xsnt3q+gUoIKU1gb4ExDB7V8nuW
OfQOYTQaen9DgGAD8NFdAqKV+08+iQLAw/ObfiDuNW5YF2jDmcpiPInIjXU4ERL7ULaBzeOOvq0o
vsHrnqdWlyWEUilW1ZJ3Pg/MQePf0wgG4mOtpwVLQLiUm0TOYXUE8yIlRXB426k4j1HpBs6u+3Ln
MvaLJYJiL2ADpWzncDefToXT/3r75Jxxs2kXGMo/Ta4vpP+z5t9R1AXBPUu17LQybf9bAIlrsDa7
BN2/cuPFcqulhGFnfu5xVwEGtcx8174rsCls7EWl43TcS1rOkxEypsagQyIUItSxcpgcwlLojrRH
2P4kXNh8WCqPZUf57r8Ie8fR0HSC/8lRHD0fPiHMr3+Rpzot9boF36l8Ooy2X/8SadkAjtRMQrBB
JbKe3S2teOfIOXUq5Fc/wxo+2ow3kLG6wymK1Ke9PedxfwyfTuuBBoOc8zB7RIjQLXsrb4eTFt3B
Sd7R/Rd81wqIU5usUETuwq7iAqKgy8V5WY+bx3SMCdrktGIOq+XduGPz4BwzPM0nT7cexmhq343p
IgwLsOYsm+0BUrt0lUYCb7DZSFvn7Pk5FFoKMR40O0RGTlq9PfZJSfCWaX0hFdAb5xGbHDKY28Bu
G9v5d2sfkggCFwSeM4tIV3TV1UCckAsYsa/BourNG5DpgtFZK7Lj2vrUM5LAPPhuFPIgukFuVxit
EX8C0wL3PUVpYZfIEQTfd5C6wmRIl6B/PVbMxzCOUYA8Q8LJShUAjUQIXguZz6lzzB2EmO5JuogB
NCkIWZtwXC1sCHkfQ+IoPFd8tc1FkNIOUtsEnZ6Zkh0+md3YwYFybz3OmcBKZleybukLOzB8y1lj
0O5J1KVJ/H188m6ZMrp1jNa0/PBUG04A6lgEhn+t2ySkkMSt5NoDfaA02BFGkEb/UDmLD6Yapvct
zRxPO9byo7oUhuSr0t3TBxpT2OtepQ9sH+y+3WIj5i2fjk56rxSZL6o27KsMjKsoBrgbsAFCAJ3V
4oxlqxZ7usjrgWlbJTYxMfMZykchyH21LpID/ZOJFNvo3/YUzCAZz3gd/AaWyz19T8mM0LBNg7lG
MgtGAWIYvgjUpRIFDBSpwW2mUMId2KDuIyITtNvTtBWQBGDJmN0cwsz/oTLZFZP+83cGzP04ZP4e
8Y+KhBmUa5M3diFlFqvQpA8e6VD/Nwg4Pmzs2ftmiqDOXK/t9gfoFkn8106MXVxR6sTrUDpv/wsp
8Vg7gE8Q08b/jL3nCILyhrTSNSXhYARruWkQ7t1V8oG3ggbkE6O+hTxbKkrLJNzDv5t4DwFZf1Zm
A9wSVHhQJA9ufJ1aIs9schJ4f4cMZNlR8csgOaYTjWEK4pVLdW08O2HxY17rm1LdAIbKBCmOGVfq
F+If0PbUqcHhLIEkO3Onm7BZg1JHmXD3Y54kE2Gqv//DFgBOVZDiMxKAQmAUGwYQV3jpZU/sZgKP
HEghRpmvG3FtYvjv8IolV2v5SZeMb/G9zUJD9ptvy+oqQ6o1qrNElEcrk9Z0OBwBlovbAaBOxzzL
QnTsJij1YUAdvL0RD4S+Y+QJyuny3AbOR5pbGzLRoMGOy2rns7Bw9sGid9iORj5xGpTtyv8xq/qr
I5h0IBx3s9fcDqolAJjZy/E60OAP4ejA1UWiO26fBNfVWGHkmMQt2xk7mWRmJt0bWBqyzh3eCOz1
HrWv+xRca0Ro76aPeXMYypypXDqvsUqNLNWqapS16nof6Vjrg29sr1tSBc9WdX+PuExf4rzPH6dj
hBAzYRhPBbvr7OQHYx+Pi05n+OKRZ4F/0+pCZJiyy1ci4iwcN0b4rTPsJzgkQRKDjjEPW5kj2Aj/
u/FT9AmFgw1APsEcVjc9MOyQFc+sPZcEDXhI07i6ox+PsUtxxz12QTJ8T/fizfjwbRPGkERJRQ/+
kctZ3fJWZPuCkJpZieL+rAsiyrgfIjjTZPiYdMsaIAj9YEdGUkJKUmSkl9s4E3ieKauS+tiKitkd
b95yKLHg/c7U5ER0eKJ/l5rXxqST0I+dL7SbqYc8rK7klqAfq3OfQVL3uVp7CWENI5vZrfBWhn8N
vLTihlx5vAb3C2pF6dIU0cw9eOam50xJ3fhi/IVZObQZpQtfhD21hCUPYrp8qLDB8+iTZLEbfSkL
yyhHVlmxC3vq+bDTkh+Z+x74KC9Pie3Tqf6llmWDIJdNHDDA3X4xgPX2usRuLOr31yazWouQyoSL
hbs46BMJIoJyIoECxE7BHHXrv7SPe1rrNt/V7+dHWGAIwsU+gW9ANyN+Ss27zOi2sHk9+AVBkRZL
mKlOI9kviXNOynTAXkHUEjfF/KS+oHVJFdubpOOZKG/egvWSu8I4gQoXQlCEtrEd8iZ3Qn4xp4WP
NclfcJG7UBKiTB+tsidVNZkIvgzPJEoyPTJ3xPppQQC9YNONihTjDCndU98nmOCjZcfholWN1veE
DWZ8Dl1hIZ2q3SnnHl+hC5bMoM5X6L/qiVKUoX0oX3qc2KclwVjxU8J3NJZSz3o5o4fgVqxz5xYP
MIKp46T08ZHZO+Z4IuWF9QiDc4iZNFBbdZ7p+SYLtFDqQVkpS7JfnwVph/Q/POi/kP4qFWOschU7
0Xc88DUKECqP3UGvy6qjJTbJdKS1I8NP1mFQUsM2myVb9CD5Lp8F6J6uakYzE75poLqjOeNtQulv
9QgLYH7TbSSzuQWVFpmazXG7R0siBpeQM4CNmKTkMlVlGfGU2OH9b8tZh4fZwA7C7+4svZyJMFhU
Zl2Hi/SuGi8g1MpRCMQMgMTv0DxHWYdz6DgQhOXecFSLArmGN/VvZC6ZVenydof2yO2nZPOm7Wpx
qNAg51Chajv7oXdNO2aFMsBsu28L8BPnLt3NB2guRMIoS+VTbiiTq6ihaVjlSwjMSFx20L0B+HtK
mykDvMYS/4KF5MXECEde4bRG7GiEg8HcpCRmMrQCtnubn7aJN2CQukyrM9U5xubDClGWi9XqkHFS
rkLusu45kXQTQ7A5aoRoHs/bQTNVtuuWeKh6rDV467PuoXkyvxT6ssv7pFclUn9yzw3F22//CnVQ
Bmu0BEhSqSbLrSfql74iFmvTY6OkaA/y7RZQhPqNaiCff2eOsZ8hWyWJ3tr+5ICduec7dF9+lPyx
j+xfKjLLRx+weiTtoulgCoEZpkUZ1cgM2zB+Sur3qY4xaAcJ+9Eopp3uo//fo3tmFW4o/KLeMHWC
WZpvxlzNXwixDTRA4daKhkGd7dciHPACwkkjtUPPGNmtIXJnPk2FwdbWPffBsUPKFU4Tw6vNfNIc
qr+Cb4ACdUZ+ieDSQBCsSvtW9ODMsC8xeQOzNQMTutBokGunOXMia/3LNKbKWe+j0BIOJw8OYG8K
kPZy/NezroIerXnDZU3VMO66dx8sdIS8H2CwG+HrKR/XJJ+Pxe7Cy9J8fMfYpzSWmXQeqZGCKtmZ
PgXrC871GTllI5vwRoNUEbOMrmyc2zFGxnQiSiLQuRG4YCAIh1Y7uKUe5iHh67i/tn80o7IRSm6l
GDG4HpMsKs6kfiC3QIZflofaCOkqwYX5oY9NBJZO2bqzbd8y32SDAUprwv6A0zpqDBQjxrk0/pS5
yftwG3iA40fz30nnROdOZwfZWqu+bOgFZGAISf1ctu5JHoWR54KW/8dTbtZLRFLhc17yLu2+HRUF
dVyb5uKJsaiqQFXH/XApf6QSxYmevguVQasB8atigm/Zhic3hPf/OvzVwOH53ZXo5LqDem+7C40C
hTcSbsi7HMmEmpXzOEIGEn+MIgCYqoeUkswYfggdqof/NnZ2UuAJv1af8rDI0JCHssIINu+INC37
pyGmBexib8L7Vqtns5bMiYJlQuxVRmCVkZz2NZDkfL4up66g4iZ79JFRbK7Q1jN7Nplmh/mLWT1z
ztz2PYiHugW3kixFUJq2PdVJnbNuY3sYxWJLiEVl+2iGl8QWaxE44xB/7Z5QpGPJHwXpiRKI79NB
tzFeWaZ8T89mlG8OBSTNCJyYJZClv9S+BAS31OcEYIPQV8VBrWKm7JURGDXiPUd6YCM+c2MzSByG
8GBec9RlpB1YMXjqMLDfFKPT6dyFShXbvPL+FvD6KWKU0msVqymgbFtCq4qMHUl2z2BFGImMp4lX
38YfP8wopvsNqVTxPouYY8LWcKpA4LnVp+dH+5yklhjAPlK/JCl0pT0SzmgKUH/BLniM7PfIll30
A4TlHfsRP0SSgR/GfvQ/SkGPEHxHgcExRDbF0oHKJD2SavY+KbMtr3rnDO9LOWSaUfV18yUWF5J3
6jQZFZqQHTV/kSTvNupI07tYrdkvfCGhuNhtUTvTsNeCyfQhVbUcnEj0l0Gt+8Yge/U7RBUfg2rS
IDq4pUGwaqBZWKKIwLsSswQZA2QAWdnt3Zp3hLRJsYDrQ8Fvls8pt2BFdyyxd/Jz1IoU3zcAKJMw
hF281xjogOWhU01CKuS2dI6/2s78LCIBD4k9c4rVoX9UxhdELLNsLAy2zIkRoI8YljmOgz4OKNrp
M1vf8e13ZPJmNEWmHPYOGkTmSnI5epC/dxuWYSpJfRe2RwvCBbHNa/vi82Ws1G6c2da6qFiOxJFi
ZoixBij1Iz221okVfjOWi2KYnJz4XgamEnnaY+G76tiguUvdk7oy8c6pWJsJViFg4oLCMfJU7COC
FO26ah8tHr1R9S4SiHOSWwPuJKYvXNQwuh+C8nFCMZLs0OpD6PLb/ixhhXvNlZx6S3h3FKv7zyIX
EEc87YbXKyUgPRqSVu9ju0VaeebDGBCAlpu/7WUmwVsLKLuZXPy0OkhBje0+MEMeh8ef5tBsBGc1
UFMZvW36F9i031uZr0A8ekdIeUYd/fy3ykDJ1wVEye676pTo6U8C8Zu4SaTzbCZ2fUyU3Rbthu9b
tpXy7gidBm5cOQkGuXTy78kjTaRqQUCeiP3QYellkdyd0xkKVO7gS2/2yMM7YhePf0LglOLg9tMd
H0HFCSSVr808fToh0O0cXs82d/JBJzHVwbxTaX35j0kRZJu9bRUskjwEz06Vl5gUzgo2D72circi
hcWAvxM/fRj+w/v1rxEliJuTM+0GzvQep7+OzMP31zv3ui65mTY8l3gNhQM65/fIJSaqdFpPhRPi
X4FORz3zSwA5mYzALMLeWnjVL+1wu8qVsXofMjApZEKlnV0JtYpCwwuoE4RJz4etrmXMWubs9igq
zR0h4lDpvMXT1YsX8LrvBuGcBmc3UKLrSgArHdS/4VYcsreZ61pi5y8XtkFlUTF3F21fMQgvOfZN
e/PbxDb7I30fkyySppEpRIIGsRlqDUvPuprfIVW9/5hAUQLyiO2aTX0urKc6cRkqiYXDVkbPy92T
7kT1sqtBEfNgaKKRW4kw70fQ7PHpQj/3QW3KpBFZIPw9coF/cOA3jZDYA31WGID3k1feLRW20y7f
cGvEt4jfw8Ygowj1YP1US3TP6e9RxU6XiFfLQEhvO6hFEUMzDw2us0XCZcCCZ00K2Sc8jtQwydbu
H9rJNZ+pQ/9VC/gp8eKhccODJdl/3LhtSFnryKmoIpkBuH5O1FpiLY/+FtisniRoNpQtfZgttYd3
29CwhIBWNOhuJqjeg83UDlJYY+LdrRdeA8LbGVZCCigGoTBzkpKuMFvc6L5acq6l8+XDoBmQmNjJ
hlfzKbUZ2D67GDz/ds/8MaBbQpGETuqSkTUxUVL7zw4DKMl2wU9euPSmaLYm+jAtl9VCh44ewbqJ
f9+NvSZi4IIfobN2hzGbXUVoGJ3hnOOxtcYKGtjPCJW8coeORIahyYjVOSz7szXBv8iW6lQZf79W
tvRFMez4KGvQBDw06LVGrM/++jpz7ChzpeH7sJyaVkwN+mMA6vUmrYJ12qxL6yi3AbCD+Rbt9dTA
yNBpvYw07y2tk7ikS5okMxgLPiScOcWGWAKmR26VKsLUkpeoPOHPcy6bqxc0Do99MKBkyersvZpN
jkHys0jnQ6/HEKuM7PcV3rFwtYsr8cMruWymH5fZJUcKO1INd0bE2GJM7SjmkCvfCM8tmH+ehnDE
h//CF2pwnHHjwQy1FJ1pMsRGEAeCwgQGjoqxZ+zO6uunwWVCr2RQjoCPSKEqfB0VDJRTS1YY/yQ7
K9NU+qz5aPXdtllxrd45Yw/6a/KlJ1L7dOdrUqId1SlfriYHa0iBr6g6fHvjCv47+q/H4KMO/0A9
ZXMP/BVxz4dOTb9ragea8UZFlMXfpzgNRJYd4eStLhxZV6fXJmXKmsZylkS9Kk1TWJ7iC06BCouX
A/HDCab2qpODTT+EiakzVFuJTezqF6jw1N6lOMyB0SLf0kOQDUpzx/wQjHAVh4ysWLwdPVYUz3mR
zT4sgF+72RV/8W0wdGYu0XC8lecgaSFL21ZsXml5SjtUByg9W8wcgPfVs34s4qW55ebhNSHGEdA2
3u3vjhd2zqKqRjvtLFJQk3NfvHaLCybK+4XfJWRPTKEFHqDu7B/NsY+IieS+wWW6bTs0nI4JLuKF
8hQE0VVen1jiAapxri7ormSpqPhuhgABpVSZUOcJSbnBHuExfi2Da4NUbMLEJFjitMwTwLf6L39C
BW/+AtfNIfmiPlM/eU5nAaoRa7fWf4OJfBLhBqF/nLRidcYRhvDJWDncYbs1+WQrmZmfBZxoA9JU
eTTOrHMf46QuI76VYIUOE1sL4osmipRl7mK9BbDqgmpSeMzL215elYCjLY+bx3RxqhRYelv09tUp
PJC1AsugH0pxWcrXP08XADyeNKBgc9xpG4Pfa//u1ISFV4B43UAG37cxYCy1+aEmmODjyuKsLtdu
XiUVgDzBNXF8SgsrHtviUivABNk1RRtVtCR4+W7CQgfalNtlcUN75DfOkYgKo6G6RehzdnKDGJNG
9n7xixn+xiAUL3LoDIjbv/xgQoo0Uqg0Y0HOZ4UfUGjxGaZBa7lPNiD1pvcxf2SrKGTtU3Vqhjko
yASsrzbw8n60MbnoqLNzVAkSfpKFXM8/tZKon0wnXhXAr93yzB7zpPVXlObfplupbGqClVTS2Bxg
VXdj2YlBuPXKOdiia+4/lLSiKyOOODXWyaMqYEEFDG29FSuMdEZPLqGuDJIifbODGvQinACpt4pe
LytzekzqqC2TNV+89p05v7ghx07BKpRMBAIlz6nxOPNWFJlrQqlm11vQ3Fo1btS7shCV5rF7InAV
BR9/vjf0NUHUGIa9oS/uBtp+TDbEsp9Oty8PLrgK3qcPB+hChXP98oT3iPwcdo0X318iZww61B6l
thytPEyZO0NnZUW1jQ9PsW7Ox1TnGDD50lOVcrdHUBBaE3O5YGrC8UfMnzbcGZkECsjae5aVDJl2
wdyJA26ISJ6xy1bB0Hg59qBaDC3SuiZvbguHzpdH857eRKLVpwqsvoBumOwpNWTLshdwJYZq+eAl
5LbMJKKy4M8wFtL7qta1lXGz+MgBoGFwsM6Uw+AbE8E1OkNdKuYwnPT7oQU1V6l3Pfh+3HRXUfZJ
48E1nETR5Rn1cilp4oOjdpttoa6G1cDr2+Zghz7+AQdk+jepNaQdOX8WztBdxVBbRUDo1W9rAGYb
ofpo08R/2w8E9Ouqn2zsdpKWPUyzEe52DvGFb2bG+sj3eAsX6MwIZjiVE7T97ot0u9qyHvGhak6o
2vPA8XBHoZDDPm0M9cEtsee/oupz0GR4lsoFkhRTR4yVTTPq6Tio7/vEsA8pdeUQEo5cmbw41sN+
fw/43LufbQxktKNNx/uQT8fPKMkcmeXBMb8aUziwR94XVKjz/2Ro5GAFLhz7PbOg70L3hv43a7bZ
4FTKxR0vcTU6LhXuyIES+QBFcuQ0M2l+a5ZtbzQ9m33kkCmCWc/ft8svCsOKkl3js704nwwcEUgN
Xc79AMQ7lP3B08n1nTaOvJeBLKCt/ENIg6WUNoBEBE0iX3sSHBO+eFeS8hmOr2cRDk7VbPLW6fGS
QxF4mcoWMsnXNnVS1w09qzOSIYgjNQPyx7IiwWgncA3Mldxfuq6fMIDGVzkh7J8JSc41YWzktApY
Vaj5B0EhivH6JL0d8bL5O/frvUdjCLsA16GEfIaqJ8DHTUYEpCCDy7JhpYr6Q66IJ8AvV5G/edED
EaeGC4V4HQ4s4MqSWNYvb/wac44EL97u30U8upjxK/Q89moq4GTGQ/8KFhdJYyyprxiOQAkH23xJ
juQMdPcGHUKCz4Z/011tLt1v1xW93Wp7Elm/IySZKlsQG56rOfPtAOLdFkUixhVVLEccvEc37iSa
rHV2xXG5LkxfG/+dnFHXRG4PA+mnDF2Ls4pm08z1A8u4ij8ZsiMkHOwA3OsCUM7JAmsiw0ZgRltw
moffzOsCkxr0j6TsR+Sjox9nbA5zapuy6pFzcaLbLWgxEWmXg3sd+N/65+61rqplL2ZD/wBYEHRc
2gDKW91o1B7bDF04MSP/CU6adXtrHoSCQFBz+JSL55K0rx2jSPeLxZjw6AYckaRPUGiV5b2cZIqR
+GLlOPI6Ko1IA+p5CaMt75wMQ5P9Ol0EWxV/KsuMO0AhLnGHMcWCxfFkHXW1LcZq3TiiRmgCOHet
R/g0zdejTBlZf3iXS/LQzdEGFiaydWJ/4Ai7rcXE+TJCzJHyjgLLe2iW2jTGb6Tt8Jj1VllYoVke
XqXT6VbDZYTkXbcXUeCeR2Rjfh7VpYF9uWlO1QAKh0u/RNW6tgCW8EhBR3nk1qWunIlG7fRVOlKV
mDyKItbRCC3COvaAi4i38eZ7jJh6u+wXryg8I/fXad/obmv1kneH9Bui11dhaPyMIGreLo1fKOUT
NkcBLbVZX9ITTQTVRx6FOQR3/PNlGTTuCRFCC8tdav6wQ5WDfcNXVbvNJd6vUhGtdYPjcVOsOT1n
0KMqrDnVEyBlxt9A1YPQOZE3BviU/i3h70+3Sn+UYJ/qo3ZQozJ5U6QKe/jYkxeg6f8waJo8qVRs
N6ID/+ttDzKgS/88CnIx3VS7HqOM2WniU0KLp/QqF8ulgCZGZMbRtrjlHdQ1E/6YOpcGSxEQEL3G
LH5vUztkNILNonaMQs6ePXLdmBHA0zL0TdQFLRv6+IpB0N+si09Vav0HuInQcaTGjoKqGhlQDRDR
W0esPeLyb95veRX9K1UNmWIzccKGyMoSNY2HLidpAa8FX4vYvGFcDjCu5srCF+QJqdbfykpbR4zt
DNWrO/SGvbp0DlRKmngi8yub9GtS6YhwsXJaWE6vIZz45fpsbnCfhT40k2CIs8K5bjYfQJQSXjyB
m+Lbvpe+mgj3zaUelo9/iofw70NL0lTIay0a4XsRWbL65EW+JUOS3KqWWcpxrYbGB9FqyvP2Yx4E
gvr2r9accL4OuTi/BxkPl2KwOEj8W5V+48CJl7EaoCXW1OUG+mDLjqyGCc/BbiN0Qqs0CQzEBGVT
mpYwKoFSNVhwPTNHPt8WmItB7A9C6ks9lqZtHdPOvcpL/J810k3KO6UQVfH1Z2ddQl/GlAFok8Gr
28qK36vi0OAeiRNKv2YiTKzCQu7paiEK5anmBvgHjCbNfYDnJDhvbSik2wLzEFUVTTDvHDqdaCtw
H2DZ6K/kdfWuNFFAR3qP02ndxPdXwONY8eFYnsyDyZjZ9pq8N5o5GcRtTKzOnXimWQ+jN2p6qHiL
sk/9C2bOtdJrSSMAUJ6D6HxbIEyWBwsj1n+5y9I26EwOJkRkOUgyDBu5ZBPOgIyTZh+Mmn5WAEPC
7Crkrw+JqVxN2UJiPxCBcYe2IRe7Mxvs3sb4V/aq35jvrxEnW18sbOqWsQkFPEQMWSADAUT7DJlh
GC9Wf/K8bWCG6Ao0UWvvMY7o0H0CHIK4yme2gFYlTQ3xyv/GQlym9AAlsG+RnLN2ADRJEYT5qU0V
d3gd2h7BRTCohNQrE1zgeG1uDJMFYZbS/S+iZD7V+8oeHb/SBhVyQmVuFdPmqCr5/EyHtE+qo1km
og7EFsduk8TC9FGZYYKBJSqyt+uPHc5md2LnQ57n7jEZfqKTAR24i9IlU3SW4AMTN5vyckM9aPdu
YdENyaxLuc2O6najApiYgX81AsyQDqZGgPMhJBkFouWskWEQpccvh8WoxFOFJPmPKcP5cmP0nli6
MwEWr0H/vnXEHLYJ6KaUPHPQsaZ0DqC93CDb+i1IttAX9hBVAGnNzji3zSQuJxpZHNNTCHdltrX5
HNM0LQ1xNkCWgM6+uH6SXVniOr4A+DByN2YH766T1YQKFQcCz9HB6F0+MibvsvPkUCmCeKEFx8zk
quRJO1h63Zz7HMvfU+U2Fl/5TK45SCy0KttxQH6ZPZm/z1xXMN2ibLVKZj+2RIBg3hnLkYO+wqgK
exlPwEVT38a3wT6fMgIeQYqQ4GDcLsH2+s44k46qxJSKsHHBSnJiThS0ntvBbwRJek3Ua6YikO8r
boPASCl7/dYGsraFmvtyOktbPbqL82rfpSDByafQQ7l9DpoexOd8ig2eILzisluCrXgNnm4/f7IP
qKuqEiKGnyj9nq3BPx/EhwJ4JnbEzix1MDeHde5DdvZzBo437shld22tViUfDYKgzUUPnCCjEXdZ
zLJA8I/dI354oI8xK0RDaV8z1RA9VAzFhKBjI71f0Ck7mh7RtI7Zcm2OPCwF+35jHBJhKdb+ayP4
9BEpGMb9meKtsc7M2SM4zutBrlpkmGnhSAejMWJYhozwHy9/2fRwIVNRRNPUe4ayTxJ/hfCb10dq
fCrttEL+v5LK7qZMoiESFTcNS9BSdF7XmgB5g4mAcUWBEPWPuwkl2Q6XHcQ70WDGKKVigi5H0V2Y
eAzkC8bmqOvkwSySbYS4c5O1x8+qRPthTH8wLQrP7GAsDTpaRBkq3KZvQ4Qp607xxsaqkLMQFYmu
qwY+Np6LgLqaBdH9zdxZas6+xizImXbF97780XrLoAT0pRHoVIwHSnOectnysNPB96rCCmtf9wxZ
gI2iaC4720fhdQHyqivgi5OMNsO5Fbl0PgiKErRThGKINCw9K5f9zfO6enYbln7+GhAzPImct9xp
MgwSgw1a3FEq5hkMizOtchTP9oXd9IMMFyRuzxIJ+vx/P3+l8hAPJHp7qc6JEJIxlIbctL1eNTdr
0toLY4impDQmkZ5QEoiO9R4haJ/jZDizB1EE6Rcy4gE8Y0Jp/wJ3Jn5eBwmkF75mLueZpZJSR4FB
1lUkSqXuPyb4ZoIo4fWx8eoh2fRWA1niXIWDl9Z2Z434Mw7XzHz3v1I8Fy1aZ13yvkXCM8vjtwKY
W3k9KPm18SzuAAY/iIgV7IM3fJZuKWTo5L1Cyr8SG7AzErtUcGqYav8zBFLZ/+jsWcyy7tGDaA2x
OXhkeTj9DQsWBG1rp5SCgHDyENkRXVCx8MUYBpXh8bNGIGIPD33zDB0wW3PFGi9Lxzpeab6cO/ui
IOYK53ZlPjlC6OmBrVxKLfvjJjnXd8PbS6yXWNW9otWpRriOvTJqa3vzu76MQWUX2wAPCuErO2df
ZimrnARfiApfMauk8irp1iP4cyD8VfJTnJE5AKcgOsej4+eoVON7S6qGl9TycL7zjfDkVmiCtimq
Y/iWVRGLtvu52pabuyOWXYJD6nuvrIWyj5sSWjAVjuD8jPi8rmAP7AI01zIfPudCUDFj5h/O4zLn
73VsoEAg4MxYdF8WLr6khmTvK5C08Vmy7jy6OunxIpIpWU1lHypjHZPwWAOYqhL1PrtBPlxyHokL
ySlAKVsO4bf06BjYVp2qCncDIKR6qmI78gPtgMMHR0i9Tc/0jznFnKN5lYkpYRvyxFRsB9EsOeiz
ltgH429klaoiWwICbsskvW7Hz2f21kAYpoGYtHkfw0l3XyjRJhRBCahgJzzhemTad7WfcoEuQ2Oz
6XXryc2HKD0FB0o+n1rlGIKKul7ArugO1k6te+OCNJlqjCkLgNekXEzIvX9LrD+gW3xDQDfXsNi3
b2q4dSDrJuoJ2ARz/WrWnT0lvvWdbbS5R142zPAr9qZkrB8LCa2fGWrr7JB85OcggRdVCfi3J+A5
t5onFKESQY33RC8X0y/qd7nGq19iiw7gElLVvJh6+fB2Fc1XpP5wakVMk2c8k7CvuhYd0H0sIpCC
OWG99fyELECyabI6nI7odfAfBJSMPZaH6VFPMUkrSaUqxE8Zuv/qmoF1HZEqf38TN6E57jW0wNqU
ZsutMccNegMxvJM55vV5tjY0eJkszvuBzIbKWgZ/2Fg0aYgKV7jAygi0yNC82Y7p1ewQuaG1Lchd
74LMtQRthELPFBkDoR2oXCgQ7x7e+5TN+FhbdLIst+k8UinCmaxSl/k7DprTkIzA7BQF6m8a98zI
B9VZoKLhapHuCeFKFrTE/zxAU1kg06b7sCAOCVfVJutYZwjOUnlhrghyDMh/nLYdL5smYhtEjp0M
p8t1u80QToUWCgPHcN2jTiRvwsNV5xVCAjIsfnoTvv3xWRDwqbR5WpqIsmHZ3bJyw4tlTJ0iKGyv
YFmx9/kpMn7QQVzyJM0eyLbAgItVEPgnXJfR9m3phezS3WR9W1SmKz0OBAfMvFoR2IVqMfCHB1I6
QqzAbnE2Hr3pOrhf3w9yjozEmr6HWLC6/l6lJCzsB8aqh1JztF1Bndyo0Aod7SFTfn72QI9OCYJr
HJyek7qfmcuhIUDR+F+Ke7/XuIEYZuL8W9b+I6651nkxKLcJn22VKZ9m21apk1/umglo7Oy+9I1T
iO9fEjc1q33Tnepke6/pCSlf08U4UPYZwfIM9CwrwCvTajafKF88wGUgwOhsdlnCZsWnBgnYiDkz
vTfgjXVUpDwkvtiAj6Ugi0+p2Q2uMm3Q9cNlsTUx3gdgmnGSIcfjToFyLkiI8sxbPtsVRPfFGbjr
N2Uby6Rz2j00dqJaBZJu8LJsvkEmbLy1loTWRXVNPCd9ZYZ+rpzgX2sosnKLXmGIZNgknfkLBYDV
uJu+kFaR+Zh3iVOf71NxUqXHA+pXEenIOOB9WjwjWbMr1/jjKi3FZO1Hfk9uwnd63CUw6y41hCjP
vhhct64XyFSUQoWA4wXphW5DmXKRnOwilYY/c60cuzJ/I50CoCo/gA8wtdo7ZQsAxDziBPrmxlmX
hV9w7gEdzasec1hDM+jG5kUX93psVLvVfUwkzYTAWsfVNfbYoEssu90TD0efjZbHfVHl4tRaZiyB
QpW3zOT0lJwM1QGlapodotFw/VobuosNHUCZ0Zq6+nD4MFrRH5RxwyVr/GUBHK5/5aqBqCuQMXkC
G29hmJFqpRkPBs9c5RqmB3TOz3n/nIK3KHVZBDDYMU7XYtXnM05RRYfTFW47bvlmaViL/VxJPUV8
XREoPiiZ2P38O1RoboJZwvpCJnyzU4rXTaoQyrNy0nd63yKlFUYEPd/ND5aa884fM3HNsVnm7lCb
2q7YjMsl2F9KJX/wzvjq3cFRP4z77C2n4xN+Zz6bPPf6n4M1BuUrfn9SsQZ0/piI6etfRptTZb2Y
eqL+gGmkGYanJwNO3MpM0AWJ0p/zLCx12I8qBWK54FyC2bnyGnAOCykAxgFXa4/Gq5lafvEzKCQJ
UWLl3s1Uo8bpc62hVUXiVvsYzwVCHfdLv2r+I0a040tRYtsDtkRWEjlph00LDp7hl0ouSJDVA3Br
GJ30U1oPVdpCecpgqTQPyDHFqy4TyaP626+ywFhrBZtGgnHIKxwntht58Z5ucG/JCA5vaPtGElza
b1UYCw/Q0Jq9HQJUEGgboK95zIVBn4j18yizecgZHLygZNrDtaHTIyheCEbVln3ePxmPlOlQ7ZSl
YTSmfx5AIFEiy9TXZFzBzDr5qvXsYHwS+WMyYxEFMYpILOFSAtUeqb5QVm4eMuLJHJNIpz27Hu2E
HSYt6XK0Bh3N3ba8751ws3wMHUUYmE7djS3tEXJMN2w5P+xd4eUYcOti5i+zADHewspWOXQ1EzoR
y17zyPxXRty0LOR2Pm5hc4qgDalA7TnUSYjDvfnzUH7FVUSrOg/RhqJWaPDBXva1UcSqgWTZR6na
3DZlBHhDYw/cK1b63biBjuK+3Js9I0o8z+hT2Awd6hrmtuenaJlCnPfISvAU8y5d7OohpthSQr2e
TrN9bzfPmFsnM6luUikapn/SU0/nGlSGMRy+e5dCDG0wqEFdzQgG8pClJ/0/JkEZuH3oKciiT+LB
MJT9x91+hZKmnp6GMABOGJb/DL3gNlrlA45QiVxi5pQbaD+RtCmkyWsvPvvkSHUEjI+/w4C4S4Jp
fxkX/0WsudNV693wPXGlQhvOA9SW6IXhjH979PIIYe9ensR5ikb/PbRp8MIe9uPutia3thVbTeKd
TBqcw6sp6O1bPLx5q7YPVRY0GKKdEJBVm8nZrqcGichdkUXjId+MqZuRmWuF4vkH1qJZZhiI4T5i
OF91adRW2Q+RXjR3yco3KF4OpNEWZHet/OH3jh4lyXBHhBz0uLqlPBqYFJ0OQSzS2dNYAOKZU1jb
kudQbe7+i72bjMgv/lgOcHf1kX6m95ur7eMsW1nTne3l+sUdT96MWNnrMbUds0+X4xlV+WEXXuGO
C9xyG8mrBdfoR98C7tHEmAwJM/VJDC3tNu4z40EjbcJMhIhLCyBue+Wf1GlxcdrHeO873iRPcCeE
pZSqvIXmggr7Lv1Choed+FUjHkNRdrEwen83O13teNicn1EGWKVLlfiulmkGxCAEhTxiPegvWJJU
PA9TrkHHDDiUpoVP4OXxgMy5jy2i4gm7m/V4YcF8uBy+EfwdVkl+26g0n1w0sh1IMNPU5FEp8oUS
yRc6R1eWeb8z3sK5pLKNe8XAJwJPgS7X/fLm6WzCHuU4lvj7JAZ6Lb3K5FdtswWCDui9tuWbffaE
tzKMZR4+9B2UZXq5fkqrkGbs4ENWDXBv5PrD+qc+vLnrgjQqVtX/5bzD/PUaF+BBsXne66L4P+5d
mtk2MtqeicsryLmyXBAw4X/ShCjUVmPRD0QdBwANtgOiO9WZyXN+KUz8Y6tixgrgtOeHX/dxShdD
309zGnIUQ3tquBxvY/5Ngo4JP3nndiCtJ/zQSNJwqApy9PMl6MNK3Mv4GKjragSx2b/odr8fepfp
XQRC93WCMa8tREKQUkcL1+FRpygR6KKP/UDS4kJESZDF3e3xgMLxZE1Wlwczm+/kz5dgUZuXRbeP
hggRKHdj+OD5NLqtqLcU0//IFtWIfrXweSO6NPl7PE83sLvs+77FC8uprfN6Tl053Ee8iLx5cg1g
pEsfARF/1LFvxXMjY89v5gu5w21KdkVvVqewVN5cO2X0Av4bQnHakd9ZiP4gWMn04GKrBGeSoS7n
hig97QIFn5dPJDn7OafTpKWcx4Djajd4Cq95EwBgVCDcsM3Rsj5qKLP0m/Do82goliU9hAK6tTX6
OiInApJTN88wgkqDfewx4IBP82OfRRIL1LrE9L+x4dKg5LWIAsr1D+28TrngJdiFrW5i3kGttrfw
ZCmDlrIcuwXxaom7G7DHKTeneBTNnODqrKVKeb6tk15pEMz6V7v2lJPJ+xm1eplW2u/yhwnKC2Ix
Jow6MoqyUGoNhkLAluzdFXHZRsBdOqZ9lg1vwNvZ083Q2q23M9zGzy37JfU4ZD05brPmCjZqNLSi
oLSOX+ewH2oF8PkYRxP9KvZdKn+fhHCdxdvHCTiOUNf59bd7Sq7007io9A+FveGX8rRMWksDP1Jr
pI8v7oAFOG/6JFwF93ABlldxL9y9PIsxQTziOsv9bq9vnqLn5rFlRgcfau8D2VCKNTD0HGeUSqHS
cFP3vTGBfuZEAqtgYahWLV2JnMIs7rQnM+crGXn8YzFhWAkDR08Q83Jpw12OUd9wx3my4BQE09R+
gJ9IRtyzupLYg/pYwSJpMETKg5XUOSKFvOHqnuUXstwf1xuFrNS4x/CjgoqkrgjjAz9BdBSgnFUd
m/tmGXSROSsCLKmiJR9IJED3dV/42ZHueEQBu7lpwZGqsbbfuXUgwAzEtCxkMjUEflPffC6UhBpZ
giZtKPfVdzc5GKLhDE2cT/1mhH15+UtelWXysroNJJS4ICBh8esWbKq3hF9RtyQTZ68HAhSdhE9+
R8spWKOeBpgePPYjSJNSSutFXgr8p65+GAZpA2JhgKpHauE0+GQyVh7VN2Wr94TYefr2/M9oAFgZ
B87PMLb7kJhGaczTS47ooSiDnSNWuyzeS/Jeng9tLvgWBvV9USHyN3Aem/kZT8jtGMv9nKW7HlP6
+qgKbC8EHTH8qti2Hdpam5L5PpA77qZ1lnCh65SLyzzWGnMNw2nlRBC+mUxYLonKeigrpqEizq4t
7evunY5IyGb7KWTXiuhnqWZUzpLkYURpviuIum65EzGNkNpD9fiFA+jv0iiyn+E8Tr5w7VEl50px
0JDNKYsIzL5NvDjWOyiJ4H+9YfFBwkTx+xlZEPFUlq5UFqCYXXs/Lj/tAqsuiPrjfQKsS0bWLJ7u
p1Z7APc5GMcUFLe4bmLFKMmFrZzVI8okPLmQvosPydgzhqLec4WTPNjXF3nAyOPumlPDI3/7Fcs7
tfsxWrFaHFATd3Dcz1BalgpzNcPg04bhxisa+Gxod5A3bnO32vRmG61n3AbFR5ShruFlU+fAJGV7
7saJcP5Vl7oukGUQw5p24s4IE+r6yJSeJKHU2Wjszbm3Re4f/qx7+fJXw6WUhuY0+t5OTZkEEJq/
7CDTzPNmxbq2BH2JNJnP1Mbhb4hwg/6IJl6fgPC49OWLIr9+P1VXwjrubSgTbpK67nIs0wrqhSHj
S2x6Yhgv9Tl15O5LKhZdocs4mOfWGdRc7xrryJ2QL7290OmiSLJnhEUS1WK2z7KbhIKXQJaQ7Kv0
bvVXrnxrwf+Djk1YhvgCdIsXK5rkg7cbOwSfsxWRnGt5m7IAXifi+ZsxOCWVTIQ5Cykrcv2Lj/eH
NxjRiPyiZRicrc481/sSK57Yf4GoWu08V9zZJlom4lc2Gnw+Mv/lA/WkhziJK/f8+vJKaZdfTESD
nw1s2okSnBoAkufs4k2FeGsz6By2fqljxnrXwvsc53U+R358YGrPSgLivEwDL+WmAnHZJrL4SdS6
TyNldOv6DzCuvnmpyK4b2RxS8+nx1lR3xmbKJlA+HnnesCFaQat60fqpKIjpfLTMfMv5aUEtHnf0
a/UN2txWzT5OZHNILYNRLOufxckVVO7oc07l39T8iKZTDEqnP91kFhSYlQUod/ciZnS/IShFlHee
jvSGKuLZHPIdbsOtjF5KgLm+MPvYavXrucHkb8LYSqjyNJjAT5oidRGgGLNS3ebzPBjAG3+QNRVi
YNt/5jwUvl7lbZioEMLn+ZhMi+aewO4o7n4UUlE5vF0so5KHK3CTBLKNj46+D7htB+4o/K7VkeUh
IZXq6eXCvkD1+lcSWP8qxb2WehHe0KfnfiDu60mXKRViV4QLc+L0Q3f9LiJ06u19FeVvxYm2WaZc
XXkp++lE0BsyoK3Ud4ZfhIHQ2p77BgIjxhmJKa0fuHL7nI6ozncWSNJn3NO7GRwln4yssiLhFuwk
S+JhauQjUBLpb5sajdmtyGSwWA80HAh168tfWr+r0cUjwvYV3pK7PvriO1DOYWA1qhi2GCeGUN9E
YZXaP6vXLnIn3ULCgqMCcPZ20WxtFTiIiNSC3WUQCsSRatPitCQntRMu8l/8HPbVy36vjuMYGWQc
gDR01OfLmNKDmLJGPN9s3DZVjm6qBnq9b3Fmt/VcNysHra25KlnaOgiaeLvcbF7hnkudKnYrM0s3
9bJhYmMoLbOPd+zibHg1Z5zsp4bmROErlAjDLLblJPh8DJpMcFnqJRv6iFvhNzmsMYhz1m/Y1yu2
0tMKALowMcxET3Uk0dlqaAw1bbxi7YDkZGR8zzSmOxUw9/Af4MgCbRs9lb3vFQEBq4Y/CG2FbcLL
nRWQO+mSZp1hfe/VE0i76YG9D9q7ZMZ5cEfhLVqssMS4FYUj0/P9FywVi3XG7lj/4Fr7hy69ku7t
SCm1eT5gszJgGY+jE3+iNDT8TZbv6afIzsKjiXiF8jobdImz90RU+Rx8Lz5PKLnMKEZjr36qbu9K
fXln+A8nwo2t68J4Ipcx1lBqOP5z3MlWemu/uG3rua/OKW9BcU5xCpLEKboqT+dfWb05AkOuxia2
5YCFGb+GbCuiSm4Lq9gaaWp2/fqsyskcVSNPrlhO4XnWTxAYpBMQNFJv2J1DqHu1fnE0sHGVTgXn
pcT/IkdR+yYkHyG74bJ+p20wsJToRrakFv4DUnLSBB5cucJXzzjQ0SoMDc7cTbXCna+RVA6n9NZk
YtYUGhxANydy+DL25w8gHwnJ3pzIbEzPQOlBaU9Q0Zvlfmsa1E/gxXKSlJLvLjTRTAg9pxlGx56i
lbUqwL5Vm56m/Q6j/vmA0V/65SbOVP8kg1cDpe5zbzmIOZwKYR2fOsTLQpXELHRivLiFLFLcpUo3
Em/ddfqg24G+7YeaSRDZK8CIKWya/NrKJJYpwnKbmLRMtLEnQrPwzmRj/mi7fEUxXBCBxOGVTSch
cjHezh+4IrEzswTLXvSYlYUXw+6TkaVbeFBcwrlZghfXrsJJiEYdtrjx+XsyPCg1VYP69LXpTsv1
TpStKhCA8Y71nQuRUabgOGQ+Nl8esNRQdOrw4mSwJ8nV/DgN+kGg2LWC3muW0p+TffdTh2h9wdnC
HCVV6QZB3gLMaLJa/gqCPVYTHpyB6G4mtk+aOp7LAb4ifRDzikR6KQNzMk/vngR+uju4UBOWJCAJ
eXyIXFZGWFjlePVNVCFh5GfzrgiLLxuJOEGnoDx5vit0GrzlZVsf8XNaZ5d41raDvPxfXRlf17Ip
eNFm8S8qw8w12mTcHQkzPjnAdmOLP24amIbhNBI/xZLqLcCRETHxP1Zq/Cihd/Av6J9IOu60XoMP
VOjqKIPz/wZ8CDyR7cfjPjYrvdp4s7UU+9UAHrve3vSjyTSy0/Xb/SQobJ6yjEfe5bWUwemwMeuv
MpjM4aupGVRkfiKEVwlj3GuEgcYWE1lx8xobKo/voeu2BsBecUcOIP43nSwyL6T1Msxa0rsUNOIP
l90VSlgMWOPHmi79bB2mpl8KluLAEypwI//OnteVe9B3XWnrC8VehM471SVxU7RHmMAkT1L3EOZ0
e9+GDrJCAsEDWXLQX//HjGJ4gpQMPki9K3SMejl+L2rWcQh2+yKFpWstb5C3LgYeJODM+3bq+6FP
0COmnGqVKtnhTyf4deiaCmaR9bZP6sbOTuTdFg/Pl3Cvgu2Jh7Tl4VSr2xr3w0MuchQRMSnktT1V
4LX/44T13MioFN282WYDAAohZ6aorVi7dV+y+YCvlrNmtxVxj2rBEuh585W1GtdN7gqGCCl1knLH
wfK6QLQgWfvrLUVtTN31EcLFaLfjZ6B+bfH4Q5Mi0Bmn+dce2NH2R49DjrIQMMKA+o4xdBWv5iF9
sMWlji5hJ+hp4PlX3ssJ8GeZ8s4xjDEB5Whz0uFqkbFeVrLDwE6rTs3GiCfcJE0ax/H+GftdooRq
tC6hhdobF1RM9/ImmGg9TQ3QLnIjVKjglKV8U6EY4j+LF1MMIStLffgdsE8bEYnBKuJR86j3urfa
eQ/NHySYtkFtkq48AG9I/BCzoZj9v1mTGmJKy9NofgvTf1c/Qf+QHuCDSUQwwUC5Uof8xq7ZdP3Y
Dkyyz3/F47JrIE5nB3zB3DcM1AYKqK08zyRN8JNAxcMp/XTaJbudO7RdCMYrSTb6DDwD63ViwvTV
MNmH76OdZC8fxLVNwap6RGbYBQRZWSC4jMJvUcOm+hVT7+53OsSqJHv75rHbPzKxZ9bN887754ZX
0UvfmZXTdw9+FJukpcAxBTm/ACtbfrkjxvBz83iFWsNeJc49W4kLgyJYTrvQijjsz+UJJHIg1+0/
EmMOTnN9RP2IUa019AipBpt/5ojdy13ea+PJhoD7jedh4AiHF9vREXIcFjevBfG3gbk32HuYM9TL
dqtdQ2gAN1cOITjvpu8FObLMMaNLov4PZziLHYz4Q1eOpZ2hSzOUK8t2K29yuThDtNPQvIZhoIL2
RztX+MkubOIM/VeF87FpnVdsQLB/rXfr4AgXHmxbh1T9Xs62xOAUJ9taL7HJ5NV9FZvcfiuxw0XE
DZyFF8HvDvROoAzMubWsZdhaj5tEsjwpILI4xbFdVDxXKNKyYK7xxBL3xV30W8NzEp2v+YBYS/WK
Y5KLvNykO9HvkT+UfryIPc4dLclz3PPK1ljVShHAeeLnElRZvdvjMI+iiKtWFt/PJ2LYRD93gPxa
DrrtIx50WmNQ+UbTCHnPZziV9SW8jxX/X8c4t/t/AuF+EXCkdG/feoX/FMCwkDLbHN+9+mlxLs4L
DCEEmaf18YeB0XFxaLMjCqO8ONU6bt0ttBnsKIgC1jL/7Kw2Mup5nRhbHpU2MJ1P5H9JqtJoNaTj
ZXg6CgHDUp+rEQZsuEXIOjhZGT/5gvBL733SMWwWO7OMSKKYdy7qmqnl44V6QIO/hcgiYTjymo6M
f+x+jT0Yid2vPR4oa8yoHuxeiyv48/NQxxq6QgL2whzz2bJ/EeoqbLz5y9qmg2aJKUBFD5tfuIA8
JZMipUPG1eMy52PUDp3qNg8NWdF+9B4zKqsyLnrRU2scnNKDifom6hMfuE7pDtbLIRL+uC3RQxnp
gghGT4sTHJUDsGHWSZYHtgImU5VWTi4naw5IdcpY9UYGf4dr3G3LUvaKx61SdvNCeLfk8lgSUfxy
Tnx8DHlM/bsQsNK43osraHB3N2VslASqKiLDl6DB+xZl+278Z93vpP1XRW2aXb35KtaGLmnllvZL
SMFz5jYTi8TMeKVsBIZGyLd+vcZsIP4do+a/h+S++ugQYE5FyrcMIU0HqqArM09uztGS8uCodsHV
avNZChqBFms/o8J2iMZuvcty0wRGozWHOfX+VaipedSvYZgqGPDrbJxbNAZirtHe7ttOrX8pbWjI
ESd+JGqBkrrEELh7Bjq7JpLRu3sBukHdwffiT++SSoFCnw2Dr4y3ixtRM14nTLNGAkqpyVF8a0PW
SGNoXY+YgYZ9qusgWAh4IjIckt1QBIeei3OU/uPwOSQhAoSqVlGrLfCP/YKsXRhhCciAm62avzt8
d/I6/gWT2MyykMG9V0fnJzwJzcrRxUVA65JSoaqjJ14VOZUL5goNOwdszvbh7n/1v8nubdcpE/4J
j04DVuxjPn/0Lj2wwpKyYZkMqUna/90IHi101FAqWtiQxwFn57p7v7Mvt7Nw2DOfYJhZvgGETdSn
/rZl7p2uCCoj97zyp3xxZ0Z+Y3zrM8PRR0tB6NSocgIaFshq0sFHOWjqTWH3Bo2wpvuN8q+ddbP7
aDs9pgOBEC/fY7AxNkFm3N8mz8EPaus/9TT/R7TPtrjvueS2/7U+ebHUnmMCVUsWhN2wnMyoH3Mg
JmO0gN7oZqx4zhH5R/DkU2oKG7Ty6KXEHQzotHo6CMOLuMfIwRnL+Zg108V1kwq+MeC475t9vCM/
YsLFWyqdB4vvILgq2ZSLvOEl9fXRODZwybAXobhNtJpoteProHzuZzXbdkUJAmgv5gRUUfcol45H
h7Fr9cQbOM3rM6TPUfIqEIt1e4llyzVHz24sfxhLUkyxJibPXuuUUxGfanctiH0+PPWA7UnMXd/V
HEQ5ae3gtSj5Q6Vq34xTE1ncFDSYG3/8CDl2RM2R50kSbzqZthy7tdVKGPPeL8q9thTVnxYoHF0z
Z499FdRvvumE1DpO+4Xh79jZVzfe0T/VmsYXXGgPyhtE1UOuzsnwJLxFcdjLNlmV6r1orz5nfhqK
+9ouktA0Y4Z3Ki76SXEo+sDp1gU2hmJ1X+yIZsK5iNzgUvIourze0Nzu3ikeLl3GFpm0/bswvT6L
leOTSvMVwUyKQ0enlf8ezsSH0qLnWCLbaHVzkDNFH/pC6jhJDlGh3bCEgb9W5BBPOUD6z1nll9Q/
PFuygCux1KdeSPZzzKibsRkJha4Ax6MFZisMVl2jHMbRdjyvsRNYZjjxj7Hx/a4tLUZt/I615nze
7SAl9L+xda1UOOKohNSYshtVRZtD1IpYju9/S7t/V3wEN+h8/Y9lO9xHPjp4jDUcNCONWbrXUXme
4GOvg0KPXGI0XrEqPc8VUWNyiWWkABhQXUtTk9riSFnpWVINpLxQZOMZ0Qwlv8zF+y0iXsvOG/hY
+hhrjnTJ7np2ibRka93o7wWsZfagXo/eNIKduM5nWltbMVU1Cp+A9ejM+998MFpxMaMnQZaeqe2P
lYiBtzMnglLtOrXcpaP6AKJOyS6z0kCGWVNpBAu6RBMANR/lcKgVmHeBBwjtNjvPQTZtRnkTAAbB
ET0AGF58B3yw3e3ipqiGIAhuh4fSvypyJ6cPERHBYEdWUtJnZGj9ku50XvObzcrP9CdaUu9w8g+I
8iMMKiTbfspYZXm3mq7A98PBEi4ecSM0gbhUakDhhtle0kUUIhMWfGJfdmNkPUNfvoGzxTL95uTo
w/vZIRbfYLPrEktdtGAqwUJSeEewig70HnJa+Nw6ZKEdNpi7bVerjSbhjTIC2OHEN2EXzeWhKRW4
G38lbwqAyPZfjJb9KkLKGXucSms+eRQImwWNZsogtxmxGzhvtjqukMbvUx54uWBhSDkbBo/y9ijg
oskb4eLE3VfdSuyVxZLF/XJWv9+II53or5/ZVVrGr0aH5c9T2terCJV6c7IeZ2KBZQTYVj5L9Yr9
kCRdJCyv0z/NmuwGvcZk13XK9sXdg3NDnfasDPhHf44gUhs9fWJsUxGTxsNzZdPXMiC/A1hoRpnd
duyWjD456Cn/+lqxag/3KapZ9idmga3AEUrxAbzZKWxp+1QJJuFlbXHuyTDyPefHiCsMN8TY4Ldc
pcD+D0ha4Pvs+ZVcGpP/wW54IYn1IPkD9NAhbdAmYDr8aJoRvesItmBWSoWmbnL3WCx+cRnGdClJ
xhNJurAy5cOMeLlO0jXMSo/tvpBtY6icbwrHDu93o8/sKQgNnYFiMlmlJ5Hw/+c6s4Xqxady9TZp
4T3Mou2WdsH6I8M26j4vp8k9hfCIUSdhQh1K3jOlt43gCcLjiQkkUa4o1lbLc0eWu+cx1w2BfchZ
dNQxwXJ8n0IxwNkC9hwCTALNrfL3ilHT/AvzWj6DmwQXahYdYDVSSdv0jwMgE0mMAH+3VFoCd0fc
hgmNu7Cbvn0Pyig/dexvYPN8fbZpZrIwOgOHvLLowROp8C19St+EPCczF5aHDHiNu4il8yTCzxOM
ITO+0zMpJUWFMaD1lMclL9W7tlTT0OhXIUmGAiA/tMMOidk8IS4RGCGvrhQ/da9LHCRZQaVUnbzJ
LtTcmawm3b7DVM829jdbo9/Qm3jZxag4x7BvgAIcx9b81YwyJuRGrTPWqE5XJf+IwVOWSGZ7VRX0
V20t9tLfBiZdTVlG+fPh+J1sXF2IJElKP1N51lpMf8Seo5tUoOeKysgbGHyT4/P3p8bEp797M1gk
Bwuq4R7jHJFT4fz1SYdPh16FjbLd5XR+y0DqD+NIu5JLBcSJdusBDYBSxM3O0SyPIm2IdOv/WL9s
VltAYRspoHKfkF5VsIFccE3usN8wnUeCJooB1aBDOXEgueJsRNPMFB/vaBrADFPj5tmc50iFDal7
h5H1D+Ews7p31MPlqr5zxWHfRnP1bwMQqXGiVvivPsbpOlsIIcgr52biZ2KfRR8gC38qXpmr3c5H
tJAz1WLrentek8ViELebpca7t9drbr8AGvxWBM1eXgvbVW4zJUKpvliaibY7lyf1aVcdlZYIuA+v
G2dwX0Nimb/K6e/QOZDYBLF+NZVnpe7R+P0JXF8Vi/Nh5q0PeCHpt4LSs3AJh4XORE3QIq57hvq/
mBzxfgjsVp/kNrh0x+1qVNTSX1VPNKz3IbPHNZ7lrf7NGe1uniyUs9pbd173mbgKjicwN59zzvAn
2n0g4Xn3QtheM8IDLj7+zfiaIyO1BMNugTFC5yntfQyfsKct6by4L3ZsIN02UiEKhoi8Od69BBEr
lpOgDgYWEkorceHm99XcB3nLcrX9P0jd3jTOKyH/AxAW9P0kfCT4k7NYxGQ2ULd8RR6iS9VY2CHS
xgL9gVazdNsETomiIG5kjO1KNCCTNl0mPfUGor3AYUDXEQP+k01EA0hxB/brvGmsYHJEWbczrhwU
1wclvjQHLZBaQEm3g186sVrH54jn5PK11eLWuUlpb/lMRwpZlN2MB60vcOXBKU51ZkHS3yUfPsjA
eCoRL5zcs+Bn4f2QfYrE5Uf2FcW6zaQmOBWcMPlcntZ4+UnRGW31FMrNS/CvK8ZqgwutCw9ptyvr
TRt0hhOeSxaILO/XngBT+4RbHMbO/TBOjqJkiPLi82xzFmqUImuJA7Z08ukQlMGiOScBBhbN8oJ3
pwNVjH1andyfQqeWIvgi7b7jO20qThp3TRvZo7Lka1GpN1df42O84sI3QSUFRD3Z3yE56qoJqJ4N
al7O5MGDCfTMccj9pdXPODIgy1aGJpW05l7Ul3ZwiLKmhoI0cZQFG7Upbvt6egJueFLdnS6iJqOf
EWphcD0P0hzWXN1oyKgSQ9UqVgKSVlowV/labYnylMl13XbwzNBH6oyVOYDPqrNBvNuXEzTvnH4K
L/AvaYxDj+ZeZOmTXwDThMGkL3JLqAkpouJwpd2EqPZgphs0qyN0VLx9dxbuBt/JtnyIBK26wRp6
4eltJgpN1alb3gAZtcRsnYKWpoiZMkayVnAmvkugtW55fTUWiyRbdmWBORxl/bzIAGJ9RVSukGUr
ReuOmy5igrilXRGLNguCQyPdDyHH5h36NhGzH1NOdkb2KHhgrl2JMg43iRoVUWHDBny/ljQhE/Hk
cxo4zpwhMKguVQssXA0MEI6OWT6mstda71KkPCHQqLxUrSBaWNXgNsHZ9NxwEB4rC/SDCe6/+4gw
QrNiGmlRfdigZDToDdxQOT1SJzQ6onfYxGj/Yr5d0xJ01W6Uqy9tGQTol58kO6PWZlqFB74Lz4gm
G8lcUwG8mh+cmN6PQKaxROcFS3warwLtXazqSKekdb5HN1R2h4v10krLIXYQW1ARnOLPFqXYHm4z
b3UPqYke3XA0xyRrhWouzgqkCatnr9cNG9Otglv7rjQ2m4rG1rvCdF+KhiZIpTEd953Jx+fk85eD
h87z8n/QxtiL2LtE6AtsmYioPUTQyGqF/oiagFTnlJJjh9sQpdv4ymuR2KisK1Plv0CaFs1ggvFA
g0dYiuTc3pf+txxlt6apCX3C6Rs0DrnQbUeCqqvBrpNxpr9yZ7BNwCITmZKxH27BiElzQKvSTBlN
+3J31vp9aHe7kr8ddmIKbhzbCZI6t7MPqWN6Z21k+Cgr5nnwEfa5yHf/q3sDMgIzeiuXRsF4K07P
jK3tUIYLRu0gZ5phZsMzIwNlxTxFYmLhtlqy4I0c07lJEwKFvc3GTuhVXZ2PehFMHTLmFZusdQHn
YaGTm9QA0bSqZYuuYuVj2jkc1LKOHpPl6WxG15g+rLhjfYgMZko+5bVKCYOAu8ii9SrAi5077OKM
TtbmswbPE35BuxoI0cPy+Pzd68/hXOtdLmN+cnK6BF/jYX0Ncun707aN8hKtvkQ8vauS0ZLwnGN5
UQfNNAi9M2o9yvYXEh8ECj/VOhtBxjJzmAXVJs8UD41Knwd+n1lLzoWK78AuQZYGuuc0h/p7g6AD
gMtLGfPGeKDKGvMw1jkkSll40uIZMo63DDigq1qLtBksHZNvsg4wQf6TClR5YiZ6e84d0Ir9bZB7
8dFqc8rgbnaJH8ksq9I97Bbz4IHYBsL3FAjXOkI+ARsd9gjrmW346+oL+IeU5k1uWjcRZWEtl4x1
nvEwIvPYhD0EVGhkJ0/hhXLafH8tdawUc2BChEu/Fd5XWogjRno4E1C//8voKpEj2ZDoLxOVlDbr
kSu8wh69mf1/DYqR5ZeDJW1M9Vuo7Ty2j2q5OhHdqBUAcrY8xJSh2OWSM29uZjY1+BjQPPmYMEiw
prCeufnDxsWZV7wQ3Q4vGq/f31zZ/+2ZHrajvtCiIcdus5/55Lb/gB+oHIVSSthprzn87HVmdci7
SddAvDX7GOIC6mMVm89lWI03zy1KjhkpNupoXQ2ZFcpsYTOS6EAARxVDQDabNF84kASVVjEwrXp4
2H0b2NFWSDANJ7v9+tjxVwKdOUgf83bq2UEo9PuANb4gXB9zxVLlQYEGCEVNQ+6ZowmXG61rp5qn
rkDuLK2T5ju/3n7vda6N6jB/s06oXP/Y8HRkwOJ+iygKoboZeOwFMOmUGTVqVpT6NkelQIKRRh9u
KzNXJubUK7MwmxmhCZS1saUmwTOvFt/h45Bkvp1TFlSSmeFHkdxrB7kMDCMCcx+5V6fJ9BEXeBS6
ty3lKZETEqhyJGiWnJudhPWXW2f4AeBjCnC2FyqitB2wzDxreRp7lHK2qhNzR/CFLcPAPnfyYeXX
Q0yzoytkTklscbbr+2eEH65W8ri+VxM+RiB1+4epprdSCLRqEKyKLWTMKhLgg7eLzAFC8nz9lpX0
QqxYl8C3ZLRfdYY9SzFzg5atG4IxoHyecZpS7DgzAFut+ZDU//MPVlge102BJB6lA0kpFLRaMJEk
kgak+NhCB//HnxDL/r0m+d1/QS2TKeRKd3Ff7ihI+pVsYWGroQWEQDUjRC1XnTYIxDx/0Fgylnop
l8PttcJsg9q2P7WjHLKRKeqWDaTYMjbbCq286qX3H2Gom7Kt3ZZpwlgpJsQguDXiKnIng3zF32mj
DrS4zxZs0bbbaOUasw3BZdepnEO7L9wC9j46LxxMFC9t8M3NtFNsSv8Pdle/bYZu9Y3fYNHXkTTI
sriMAhut3cWnaFCrBasHQP3sqC+xsCUSmGI3TAZzuj/664HNfYrA/u9QqIxcZe4lQJ/1L41cKHqy
L9ja+cBV5rOPfzPc5NwKYuX4y1Xmz2pPGhBkuGIkjnbnTLimDUsg7R5sGpStUnF/e+GYzbsdsUkT
ZjAGpcYKkrwWMtpC25Uy3sQyrUMzBIk3NmLwvXmWXAq9FnqtnWKPOAodKlMLE+8kryXpxGxyujSJ
/TcMb+EwKnyQt2Y7jY/XcKyQPb2/qozWNXGzpJJSaSQQsdKQNJHyqUqNqirWaaUMvKUV8VaWF+Wp
Xi2U7JT7z6jlHJ45EfUsIGxaIFDsB6Q87eXefagTPSJggr+hfbPNrs/JHJP2cNj+zP29Up2cfZxF
bFB0KFrMQPl5q44I9PtyI68LVBdhFsgnEAl+dikdzmNQe2XTfwu9OpLWugRDQ4q0TnkGVi0hmevD
x9w2E1bmLtt3cbFUPDtXmWsHYg1Ica6rvRVgETAIzCakIJBd6YfPAy3ZCDG6gXxN2x2HW0YGegny
zRz7pmvVO2EqyGzIodjcDQlUrLPMAVpWfAG1WDOqbf7fN7GJYvmqUInp5T6xmcM6IX21SU3E3w2P
Rg/tJ4Qqabcsx84kcGUHNzspKIustK1X2pcFzYeCXGxlckw9Il0o1Js8e30vLAwFN1tB91+MU8TU
IAyih5bbxquNo22aHWCQlBntszUYCYPakhZyQgpL234SVqrPF2upga0TGrPO8XesT7F10v14rzTt
3QUOg0FxzswCq/uQ3bQGBToILmsLfzW0VkSjR+UpxvhnZaHtAOGaM/ykUW+9d/TuGCPLikSOSroi
h38kNozRhnRAFzaHM2llwbt4zbGdGQdC7pqI9MkamOgM3edym5BRII8ATAsqZ+ESbzA/UMCXaSfB
jWPxridtdPAmdNlqG46lBnleTgax243AEchL/cGODRMNFCP6mc4LQqQohNtLZRx2Nz2rYm6HkhtY
ZthCf1XtnTgaejcd8XwZie/To/zAtsQ/V3Hpd7dG1+CxbEjvUcL7IMmFelVHCu24Xam5N7VReF+U
ik+Ko1ME1jQ3sSwkaT1tEuXYAMusgffIe/yMCmCp5+piotSMFizp6bGmE9jJU3fZhuCsadXgtFps
XxAe1rJ0M1R0qyIwvn5SI2pg0/xIFJUvmsvhB+Opuw3Js3QchS2I+LPB+qrNgWUavAC/4eyzdrme
kkmA7uEqlB0dLb3sZHFflhXd2tFVELsr0COtJxlzaovMl922tIpOxk4x2TudKKkl1e09c4lkQzdp
qafLQGQ+frp2V3TXJxgRCBYhBTDdF5xn2Y0NhEfoYfDBnKsUjeLk2pJXF1IIRtgEhDo9Tt7GykGb
oEoxdxDy5mLr+VB6HUYgU0CNagVb3Q7cYKq/vB7RFgRf9l8lCFtV3EZsI4SGIQoYthyuUTrj5qtQ
35BxnrlEN40cYvO8OUFrY7N2Rz3evvSArXL+Uy2DaAPvigMGqwuWbL3p3td/8AMxeQRcDxrRHjBB
FPJNkThJ6pBhNkwWHATAMVYprCQDDbK69I/wJN/ybK85tlqj+FvHIoU/vr0GMBGsKifybh0U9yxk
sJCgBl1E+/jrftkn3hkc3HtGE4bxBRyUfOMBMmfBJpOmgjvfkL5O2dshYSCHogX8a+WzDQmakMPU
fwDmhPpKnvP55IMdxhX52cM4xMSqL7xdtcp8FKQ2vH6Y55TgH9p/ZAgjvTfleteJIw9AA5sZ+CjZ
AN8ax0LuCX/wYZHFWDEda/t++bcTzkbpD/lMW0d15JXkZHGOnzRQT5uxTw8Ach1U2rj5u22HNCUt
8ql78qIRldn/6GKINjPQZzsQNnPAFRFKD3SKKMCgSy+JFTLEfs8eAOOirHz19w7nZiyfoIo/KTXJ
vmZsEjgVT54VSoWv2Lndg8/TopzE+u5n79LMl3DS+HMio2hwLla9Vsx0znT8ACm3QT0gj/nt0h+6
VX9lss+1IeKmWfknCB1DInZj7uzxTYnB9oJoIJLaCLoXksdSDFF7TU/naod72FCnyAqug3ge2jeK
yKUa7rAt7SBaDAI20qaJTgmnrT17dFi8CMxvFswUDpetmjUf95AgK3Nk4UHUYHT2BEPkRnqL8i0k
b9c5M4NYUP0LbjnvGTNPRXyYld3zu0y/xWr8LVmTE7ZC8HTkvW0ow/moBZCoB/8Xq5yT62dbkmVV
IHPKIYDEcTd1aIoRtNu9AdOOrzbEmnWgjOKewKUaDGfs6gXxNK7zX2YwO26DWs4iryVytOYMB2DX
Q0RfhIZgs+NtNLypHxeJeWd4AFNe+FWV4Etiv94QqB3u6eLV5AbdJ9F7ayeVyO8bHHe0kVZFEA29
KifyH+aJ83mRxphkJy+WzQdGoaAmLjK04imfadB941kc6wIUXZ4feQI8iVeXHfoZhie8UO/MjNQv
FEqCJXpRAxDwur0P/5/SNGr3v5lZASAisXw4JNEiXBYCJXsjk8Z1G83Uz6/ymr2oGl0Gdwt5u7T8
RjMGcWkn2NyPrkc6IeckeYZkZWdXUoW+8V5uj/9cRoyc+BFQ7syXJC8ThnfBBIyLoyo23zHJw0W3
NRFd4mOGokECTehpp++7lXcskJ3x8Zfcp7V0bmZoQ6vWrgqEyvpXZKgOBJJti+4sUAv8sk26fUCw
NJyR0ZCGtbJ4delBpQb5Sszhh+I3ichdqRDp1F5G62Vxpv/QGunMvjwJljTpfjN5SJ22fcekDR1e
liwhoiEorleMSY2hczb8Pvzmod388FZUI2lW48XZeHAmL+zsBubQCNG9Ea99rMdWnF9YZInYJkHO
7c0Dh2opZw2MymUkXL1ZnpqvjcKOLLNi3KeyrS0/U//og1WNuQfsBg9IE4UZP+6QALtJY5ahg/Ok
AiSsxFEaZCOx7Dw8ASjaCM35TF6Be5z6vg4eMX8vHEQMey7KMR0rTzcs6AAzYq9qVNnzkAl8wfmI
dsY9bDA74+ZK3t2DTkAyIxfGt5EUyN03rDAbhE40ri+SGz7Xcy7pmdBLkbuVXb5Fiar2xYW5bJgj
uY9iWLaFJaoYMsC0fTRSMuaDMRtlCqqprfWFdiD9Qan1hLGfdwMWhEhLndVfC8qS+3hJIWBt3MT9
8Nm4Er75X/WhX/OU/tjAa/zG7ik015ttVJn1/ggDQphbP5BxImwh2IHOe8Nk1CnCSQJ5HRd7lEEj
yOrlEhXjMjFIIwMV1UsG1k0qMv5tXpHqe+lROdA/oC1ldsZDnmW5WMwaDoHGC5GkFFHEqhkwTxYD
TFEB2CRCpD42VgQ2/W8+ixSmitOT+bvMt1W+gj4CPRVWjBlbUOcR8INbZicy+wmxT8thgOZeVvUc
bOjDE/Otbu4PeGm7E0wLjYQjSCL0q1x8M4FvLSOYxQ1eEwK2UGTVY2foJS61xibI45O2YlHaQUog
ZDJ32yE/1VhjsQpQ1cpg9CB/QB0IWP+Un55vvAIcRXgNdY350RsMbfRunigKqLOdw5l3a8BcDjbu
E2M8pUlvfwC+9jQjUwpEXNL2gkRqTyrFIo6EYmngEwwz90YuXHO8cZ6d1Z3hxeKoE/XORyhr8Nwj
NFXU/MSUDMdI7tmQGTMZx1fthpWgPSfTRpbGXFabInQYbUZjryIIE5eJjW7hu+EF9pUi6qebTHX2
6AmiMscI1OnyxBPhYvJa67a/Su1kCV0mhorz+wuSRhtIvrrkDKsIf+TkP+lxD2Nj3ho6XXtBvkBP
L+oo80cOvwjmjmXCahST7U4KaxTutOPqiwPw7z/uUICyq3k+lOXnu0KbLU9CTN9/5ywoEruwjIVW
alvM+vD1NP2MO0qIS9ctfEI5Jx1T0cO7GjRhyq+LmJvhDm0Dr4uIjaJj7RDTpsKFiAQwcmng3mAk
yNDm3kucdhAcK4pUuMvRtnTCarottAD3jCsfP0vWkGGuQKKKsAImmt+vgBvvO0wlJJE4EDc2nxj7
zykSqohRKCYg4FT5zSzIty9HCHECZ1EqF90zjDoYG1Yzh9XF5XL4yJ8yvZTDr38g/sqWnBvLJdoE
E9carSQMRnuQJPeqxPPnDzBhY2ocl62YNZ5PQv+BRHrGy/WKeACFV0yfDG5K07j6uhtyPfrWeS1y
qQpZCdZ1lBlFVccJdRxHo1BAHnsqYmAUS3DJa6/nG181hpeU/vFbh4cJMvUEUt++mEVAoaF4HYlf
iVwzlskIH5zgDc/mgfus5mIQnfPCswd2CT9PChHOUvjPmXbp2UknpFIfXixUFiD+oEj98Qsd9+T4
jzK5I2kvhEWD/7zn2wjATqTLidrD1Qc38JLKAhtcnWEEStZmbHkNS4CccrnLv8O7o1gEZONLEj4C
7e2t8oF2opEO/mwJWe7BbV2xfHmxNCYfkXpDSuYVAoGxooxk8P20Iiz9M14fT7zwlVCeTg0YNpPI
ik++vsPvF8XIYyFVQaOi54yf+X7htdNkX79lVZtr9UNx/yb9IBqkD/kKEuwPPNedmOoC639jJ5ru
HF6MGRPWWj6hKcPdnATeGHgHuZ731AfwmY4JqHut9W+0UhnpqwoAx7fDTmp+bC/oqitouXbjboPN
LtGhgJvq64F06lJ+DcXB4oqmAaGqZRpaT/dK3Pb9W2EhCM1XWxiW/vV4wPtPtOKMD5S7VUZ+fPNZ
LPRls1OYyaMNLwG4Os9WC1+8uNqGJNnXJ9XdNfPC4aYmEUqagbc63Tq3YJ2N3Y/Vv3qWmqpUk3ra
+N982DIvByz4ZeV2RDs06t7GLED5i07I1rm+E4Qfg+jEre08sg2nEpeMVINunBozTpUC/YDRmc71
Wd4NqA/m5UlDywlc4U8VaFdRxO6pyerwg400MlY/0fGaRodgq711iCtTSzV4sPo2Y0EPRuou+BSJ
tUYqLJmMopcWOGOSHgVZ5OX7EfxxMY4909Eim0ycjOytjaLCDQ3/nM0yOByty4Mq3dgy3evZm1Du
z8avVhA2Q07qvRo2MPQ17M88FMfZ+Fufg5ErgKz3/QHZJi+/pb6akMqdB+kYcJYjnPwhFoOFd6DQ
2vY4+ZtcVC9xD0HyJb+Fz5Xu3Q1CDCRxURUuHBWaAgc10vbZy6O3a7TarSWLxQdTRSLvI9apNtEq
tBcwdJ37s/nN4ZdBsG2jVbg7lpP+PfYTnLEnxxIeBbFhpXEZu8Q4rvmA/wLoqufFxug7XXbZRAk3
S6UUerkU+43lrTbt8EhuqoTZ0PZmrEHKQ0wCwBtXkh/KlHVB3MTV9uUspGezyQz7w0lj301vqqdl
20EF3cHQiZeT6cb8gk1ndTqZfgjnPzC8V3ASrmUHZsoows8XqCzImY3gGstKBlIIgTFfP+/b0S1W
441nelNgzJyGkSEXmBB+Au/bDy88IiglLIsaWWbf2bDttwIdibcqJlgPHPabo1oML/boA0jZL2dX
pjfUcAv0xivyTSuq/ClQJiplbYNhAR4R1oPdKNSEgy9exyqWn6wNnnKaR0qk7FCiiPzi+zvIbFXO
sytKK3ZfjTAo7SzLH6/qlq45HKRpeDGT1w0RuGP4jI73zn8nAm10RfGyQudz6S3Qbl17g1L8yn9d
hiJCReF5Bkci/J6z01o6gZ5UvRNXZs0LzZ2OhX7giKHV374NSYZBHiGMPV9tg0xbKTinSxNvPc37
rVCkKjxWAeurtd0Y7Jz+EwvBjd3WWBFQFlrqafXoIgu8AZawOmAhJWYAdPMt5M30wfpgJq8UfE/Z
/nCGxLTeuaSJoXgUZLzZrvhVRn8JRi3Hxb0t5J9AGp2F+NzB4pCLec+JSbLzAOLOZa1+jS+BkLsJ
PQzoVhkP/ABHwyx6K54IE5ICWYujayifcM1xeJ2jH+NCtxzknt6Sw2nIKU7Qa1KReOjwTucwT1jU
7JnJsfMarDFN2KUfS6pPHYyJpwBs76XU5Quyj0iqOeh5YylMCP+U+9RZYq8OUydPuNOXCnot6g6i
EJmNCdkiIMyUdWcOCFy/32gjmrug0gWwnwSbRTNrtFaVqayRHCbc3JJisIV5kzHKrug20hH94DOw
YfVUoKiuzYpVgmsAdcUzTTx34bD9muRqnZK8orVR0wNikdFgIB3i5sG9DwptPddPuFAYvhTLJTMk
sjffZG14t9aUkeBMEptxOfSNPwbm+OmbBJFqhvvLJlzN6gtA38phTiHdglrp0hqG5+50leA0ckR4
X16qQJtyc2dX91xQh4DqSlSCgoA+Ail+WbloLrDH8A6NfsQSzVEhAicrUv1RZJ497BnzCwEv4SW2
elMrtRWYfb+hivn6AuBzoRg0CCBu/JDnRA7IgqcNzbXkDJIf0LtNr8Arv2TibmQWkdLij1W9lZTv
NFIKXiirgF3EYCMZbQySQ5ZEGu9cKTYIEQsj8XryUrrs3f1Rjrl8S6TfBV9z8b7hiOgLWHOnGAa5
vbdaWe9NMH9FP+IuAo+EUMqDDjqsKPkwTqxOGiJuiDBmDPxLjtm30yio7nN25J5jd/RY2gH80+nA
sRPjyExqZ9ORekPsjhL1pBhRVPK1xhCpjIOksmyJ8AKa7YQhuIf59P+sLc8iFH3EOj8fYvDWckeS
EWPSg79TTGES9ZNMKcZrQDKiHXjw5ANhC5y8fG/mQr9tnAwUlE0fkMkSHtH5HZgIp+xCjj7IHGZk
lOrG/wY4tw4h50JhHrcmmNYSaROWpltw+jWHkvyGFOZ7eNHb/3XrqtccHHwEoGULtjSGO+9Jm4pY
n/Ar4ypTRrcF8i04mUopfvjtkxlvYcHeXxcjN3GkTzl69uF8FYnkrELuK4pIRiCI874gGGIkZAk5
agoi0GpyrDEBESaVJDzCtp/f/JgHBluZxCN+9SGEBn40GS2COeKEHa/Jz+DoBgM5xouyf/HgumYS
MUI1DeWLqrb7fDOnLkl11FdUCVYD/0wSTAGYE5baItm6NLI6AzSDcMnnEeLYqpERRj2weyhFFwm8
byWePw/phJNnP0GAV6rKqHpS63Ax1rKeZrAPhza0JnfM9B3lAP/30v3MPvLYhDSWqRQOcVXfmJGO
dAGw+7R0wM1+n8Ikj5N8D2e9TDynSHnEUGe0/goULXLmG5Fdf4OjA+ISFbUwpo4KCPaJi3qWoaHY
oKg8Rvyuj2eS1dd0VFkm5VO1+g4fI5d3TqbvTz6YsLTuiFX+uDWcyoxFqPSY8cMN6UfMUM9xEGYZ
UYk1ZnsmUcXeQmm/4IB03FDJhStSs7K26CBqLr2GBLLwV5EnfoaBpI7JeYSPFsW+V1Vz55ir8iwJ
UOeio7hReA4GD7fRNthAjPc8JE285uin0DAMBMkIXQAnCzCBVh+7YufP896qUrXb20gU1pnerkiA
6YsgCwdUVWX07dEknBt3PYosM5pj6OaMtPOb9b6r5KEcz/WbW/7oa9ipUi70ICqc8F8/2dQfL6zJ
dUYndyWmYfY6h5BwWtUAVeJ0B27et3aKUkxbm4VcQ+ralu8aFP5v6mZ+WUkRA1VOHyIBLe2Lwd5G
JnUvKNFvMctqi9twuRDs4e1MZZGVsCrvXM5EXiBhwUGzvdaT3Fnk0Wa8y4Tw3AbAN+ECdGNaSQch
YmpVHjArbiR+FtQnAB8Moulq1T6ej6+lmlLOdUG9IDNA2MLKyUus7JiWigVESrrBHjUBM9IfLeDE
LIDNQ7/Kj1oz/7c6eDycYtH200y/bWvJqOfIIwaNaATcbsHUYyEj8GBscYvg0LZwNA/4kBb3wREQ
ZOnPPZGP2q4XGuq9bLsXRNRrThPQ0p1lMgpjskKtqfDSSX6idIuC+T6Xt3Dyu3T+ZG/egEcK3sGk
BJn0+iKqtUvviy2iErq4Rxjtd8RIA/sNsUV6AFFeqqeQ/CZtXPQ85bc0TQaoLQWjoJ70OepftfkF
q9trVbhcqvqch5GOIaSOH4S5v/rjwm2PHk3rBwqucau/5bhVhAq9JdOUsINNw5i8gsKh52sc0Azd
Km78zAnYS3qHPlF/ScV1Fp36RhvkL8gVNH7pIh6CCadS3GPlw7DoixlGYXPZsPmk3krZM7D85cNR
O+/aYmZWhzpwptw5BMiee2dvCdAmi6OiSfy3FUrFL7R0X/KGKOPQ9mtWc+j7vJWKMF6fFgdJMKXw
Es03QIbjuWqUW9q9YUuAoVxqxU6KGJj0hy61qOlHntJwhmfM61cLs1ue/uwrNwY6aIAQp5NgpIHT
Tx0bkQwwvaBm403Tle5YcyXSfTRdmJMOdNvn1teaxLbIS29pXy+HRnSzn1cQMNP9R5SrzEuAyIMT
+IYGIEj383rSpdCJb2iT7A5syyzW6Q0gvNi33/rojE4kA1ny1giH6TwWpgI/0KGVnINQAabkGwbw
qTgCdkH71DoIF3agr6EvRXmmtgGQKFNysH4ij7CZLHy4RGxBtQ9Ea6WOWEGKomrghqRSXlYE31o4
yVU69/NLppkRMMDHbHu62JTVxTviWtqXtAdFwfw0+BVo5le52Xij4KXki6d05ubCbipe0RkYXAvi
9jh9jkWLgtgJxU95dnmX2MgOI/WmYUyRu9zld6rrn0F09gSKXcg5RRD8ftvZ8J60oxP/rsYq4Lby
p3N+PgXBFpVeG/c3AYto4aEX4NQAKJriHpA301M6h8cEXUU+HrAbmyezq8gToTDfTy1w/q41abKp
Ijz6Vd2HLhF/kVGPVEoiJJSyZO0IADUdiqOmpDN8S675+9gugAkWpNbblc0qy7YsReT5sY5p7+Ko
6LV1quHqhgH308KkELi9d2b5nlg/pcASweoFJgD6cX1yX/zTFkqRZfjdiXppDOjA9ZUI+CljP8Ty
t+4anvC0e6705vERKz83eHFg+Tm+PXsyWmyVjjZsWvT/YruWwRUuuWDSdxXDRUgZbzNtmlDYp6yf
ZnjInkwlGVgPrv/Ex8Ib9xVWPGYGh53ksqc3DViv3JlztKSzLBfVrL5H8spPj+sPYSg7yHHlYf+n
z2hAvsnvYtptxMRINVsHAxR7phV3LEhMC8D0Q1Iy1aQ5eSQardWI+p4g0SKyCYE9vP0NzRy8NZia
htu6oTjpXyEVIgx50FRfVnYli/j59eHMN3l7ux1s5EkfAEHKXmzJp/v6sZIRYcieMPzlAUGJ4ebD
oh8Ad8gVGCOv/CUg5pAAdbl5GG155D+FujHlPB+QFpdAXJBwItmsj941njR0PfAQpDPNWiuem6K8
A0ccooOSO9s95QmhARH+6O/qD1s3zG4sS940zSXXBZKb84NXjlPhOPfXGLFycLqV3imdQqdSILHb
OppTLfYoiUzwy9H+ohP4Iqcbv4FZAgpCwqvsFtSL1R/LLhIyclGC54nb7PPoETxqUaiGmmYk0eQ6
GnEzTeymDKgtchA1A8pa68sZ0gSlJi33WZ5WKj5oYuVKk3Li+tbVYrw467ALLHa1R9BCBQIXz9Fu
gURlrPGGxTIh5GAXbD9UFaocRznvVZjrZAZ25sNCGOzpHX4gcqFew7q6ceOjlRGcmqpLCKaadMVx
1RuzZggJVwSWF4ko
`protect end_protected

