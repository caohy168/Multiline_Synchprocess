

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nwI9apodsxWnt8/qZ84l2L5r2ru1rYRvzH+cIiU2LZ7ZFrYGVhrKUku8GacxvPmk04mNLHGAUf3D
0KN1yrZ0UA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Sm1hR/bXnEX5hSLJC+m0q+qTo+GE1jW/bGh9GYODVR1B61WO0x3DI91rmMkLB3jXabqZYmZaVRnk
N8AiDf+w3tD5cTm9k3UfnHfkmqEgj8LBJAWCYHciLWzjmW7DKTQG5Copg5YaoAmLrkH/R11p2QBq
US3uTE+2f5z8QlQwimE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y/EngzI5VWuiEHV+TKhmZG2qH1QkzhsLqS3InhpMlNY6l/FsFenjJYgIcwfRB5cHNIe7FLSQt6Ne
y3HMmpsqF6xetN1AMKtt7yIa7k99d/5TC5vyU4dMYs9g27cqHYJzk93esgZCvjIZLHpcXw/tu9/b
4U5FbTjst4GUWQQ7e+FOVWa1BC4H7jo6ZOE8mZ1oMeTUDMRBFFBQWv4xUZFg+dKul2euXKFScShR
h6tknaycBcdNbA+6dQJo+VgrTTewvfrkpNyifPBwk9vIitRhFkJJJVGsR6T+AF/UJfY5dEYYFuu5
J288ggKjbjEUNQnIyNWOpZiuhpClTTay3laNkw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
htKUMvAlzdN4BbAAeNmEM6Yr1UUCORwvd6+1cV737AnX/e5QyMGFY1ZuaVzrrzfIKK+VWd/bFDYR
WeL3jKvGUsyl0cMQ9jcxLrsCI3RnUD8yDbbqyDu9KMj34D7UA/k879CbEg7mJQsE/OUuwmk5Rusa
S2E+UVp+HrYNnNymuLmmn6wOTCKRZjZEMW81xyRvJrDTTqf12SjMprM/ubdETBwwiEzoIwLeibWv
EE77NEiYVwYpzXElBkB+JN+riXCrervjpMbAzHbeomW24pwXmffMMvkj1nRzaEI2QRT19Hpc4iqq
tT7PSLFxC6iyyFn2bd5a57kSCEK5ZaaxszxEVg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ST+OORnrF+3QguD7AuqTgC907V9FPxT3xpP2TfPbwAQB2+m85/czQ7xrlMYLNRNl2qldRPC2JAtf
yRLJmvKEgyRtR6tv/9gg66CdnvMVGbBmprZnmsgKpHGXcIGIVm6FR+ifL/5pZcFZyTQCKYlbE6bz
YNrIQ8EskAk5YXNHRZU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Zz8HkbKk2BMn9pYqHdEWEMFHnKjJed8tZnBzajqsks1G6q0CzbV0FSYoWS1nKj84tIU1JkBaGDIt
9sdF4TFidxOJyhtrmpNfTChKxpMr41K8vo0yCOwdi29v/VShuI/rkIBCSgrdlmTBWBEgiBS9aabp
Jqqjo1ol263k6jlcp9rOjaoU+lcQMEXCkHoZu/V2+VWtTqhoSiWKgDQ0jJptGQig3wemEM16ctGQ
xX4urrzlEYCVTlr9g3mn6x8NgAjEFjJqmg1uE21AWGXfsNowkj2dYZLCXuVTF108ULXlOgx8TBHk
tPYc56T7eylPXV3Y05Z7agtvOLTYldGNSnm7qQ==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VHzNHo3jyVixjpbjlcbNuO7IrIjCuYoXTAjRb06/SIYnbUS1pXATLQwryf5S2ETq0CYvThlIAGS0
xbNOLpEIhHMaY4VNrUdhUPBHXcXHWUCHudYKaUCB/Pk28QZKLuHYt3FqZh6wdzI6AFJdP/pykVJb
M/Pyyc+uLtqsAqyWqtJ0puNrBSpFPSM5259v7Gum4dwYGluRNUyJPq0CnQOQDcjaKw42cmf2DAtX
CSJb79mvoLdsFiW5ePQbcfrrcT/FhIkNj4/DqMVl2EB85zQgcPJw5Up3lLGw0Qd2Cd1jeq3A4qcf
LraHhfdfhy6tS33yDqFUeXlzvLfkicvxivScIw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ir7vg+6icGbLB3CLLO2WEVH7p5OyaYzRs27g9ktjlLGEA8UZWJVD/LEebYJEdrotzhB8SWmHZMDV
/tU66bmEBeBvDhzPDFffP8JEne90WI2d4WsOz8gc/qUmQrWkWWpKaGeRzRKobk6HEaC+nXg3PqfM
0b03fbE0S205+4xE/rEnuHBIRBfZd3xmeVaB0HKBt0SGPD5SSQQZpPD38QOtCELjuuuA4RtmpS90
kaKEHc7Je6wpd85YQOJtbSfSfwms8QmBrV2vuYX5vgvFoWdrKhFu6ei5xOtYRK3gX3JKdEXLebbV
49uISo0iQ96Wfdc+51UDQD4Z2sSmPF/BKuQ5nQ==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LpdRmMYH4gdKs52wqPlK6TsP8t36Rz9etYG+uFXIxoYPOw77GvCpHTnPEq4wgKvtHfjSBYM58T8o
VFR+rx+dgG80Vv61h2/ALXu7WMVNRnj432YN7jUfiNGlmdGjYf7j5bb6jDSZd9SGg9hOG322ua8w
FL0iNhZ1+8bqOC5DHZhVoYhtH7wentMTqEBB4I+Xy3zK2H07hbY20A+hZ5iviyCzHMtmQ5LCJzAb
8LeBnGRdOv8ntIJz3n1voQKFpamiYGRWqDwIHC+A3vf0VlEiw8M53hPC9SjoIQqQxSnkzTditbkH
fDStRcfPfMIOJ9yoREe7QoWlh0XCwpflnMvnNg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
JWNKbdkTWBruQSySiq/T3NjP/iwubNc56E3ZAdy/+JqVklbPP5VJY7wz+2UK0TEIE4c0XSdFwBF2
FnRiEfd6mQjMLP2xZAEA5CuZrfTMWb/xJEO5VMZr/Mje385XYvu8KS6d7mNA2gEItGizvqITCSPw
lA5ktYy5hBewCbVy4vGeb6D+C0P/IvcxajYSwUrt8kBC98NuSMBghmYZH2yu2lDgr6hZRLSN2aqh
iV4l0Ge5+kPBlXa64RR+O2ZUjHTxJTaJNepQ7rm1bjyPrS+9kHR7NLrKeV3r45YmNEBUfZLLRBy+
CAtnZVTvmTKNgJ/mUW5icoSCAd/3+HJZXLFxVheKGeMDmpxYOLwAJvr7YoHIjubIMhO0iqvi0kn+
I5fjzcOiMeSGzO2egsQ54Do9k5N6gE9EXaDmDOqd92UckKxJyhLP6RcAneTrTxAkmZe1C5s3goC8
esyXifmEkKiLg8cIYUu5+6sSjsHy/3v/GJMehbPSwAV++Hg+ELj31/4E07eaxh1f+MoCqyjJWtWI
FTf7anMeH/Mc4TGck3iVXlMoLazz/EhFD72bFCf+m5GVAv2SncXlTm/TTbl/SkE5wGT5UGUMiF5f
sAvUtpmw2KsbeNJvXR7rl0iUBlSkNsQaP9V+z8eM0nfBUsABk7rNHtBJsXoy9HfNKTSreJfo1UF9
nKhD/kILzKszT83j4JvdvT6bC2xLN4hPgcVS6s3Oc4Okk2d2qPSiKTil62we8X1Ae2covPsQTIX7
4l+P2Y9JrBTNteQRw8+KDBG/ZsPrcyU7dAydM4DRDpy2Af5GwB3j6/o1RCwRDbyjMa0iUBOd0R7Z
PhqURyzn/YHGqqSgdr+NDOIZEcgXn7FMJy3mpHjU9leiab3D0Bn134XwLa00ChUr73+kjPDzlxDf
JU/wbzZPuK7eNQGd9V7DgvQRuyqaADQQHIXv3+tBrwuIY6eeNac02igGrBovxeEbOkgbTSWsBpPl
cfbAwc3e76Z9iCMyyzMHoNnc/NyfUKo9KAC4/X7jqrT3IIe4rKT7WJTtrBLQiNfZo1+6ZsRCtNvg
eaRMuGSigrTgk96PaveLRx2hwgF1cXGV3n2b92J0qgJVVNKUmXOGfe4p6uq/5jEB8crdUEwI6xCS
imaYrd7UgudgnWagPR4EDRlq8trNtujepo/2dD2uZO7yUs/CKAeEehr66Ht3AgIujUBYwmTeYxmb
GY8oBW6hu6mQbmFIWau8y5W/tL99PVJqTQzMtMNWEAjQ8+2bAVI0MY4Fh1ubwI001tiZV6tET5tB
B3gBNLRMwLFC2Ue7w3zVN8XEBbnvQw8SYtcZPwI7m/A5iUewc1eUEqEnDCc2rApyxeCEViD71+Ng
8INjTH8xObY7B5Und7X4xxf7eBMOJza4+tWS39Oorciz9sSV1F6D4UiJTnN7te9tvqBR+UkkANNV
yaXLG7jyf/fF/fbPMwKAeiLxHAlKxa8IbN8ulXyFsmzlIVR/thaY7P+dQE9mt+cEZNDqTQRBHdXL
1Aj2aqFgvRjDBlqj9MuSpCQ/kBbitUvf7aTiXunHm9YCtPaB0Wv0WVLIyGYbdCj8EIw6h26UJ1/E
hBGdr/OoFDKZbXCB6Qy1FBg173B9xup9YTYeAGIROlndXgcx9KwTjtLx69O6usTW6BPXzLgvXtsh
fHCFtIyM7GuR4AnVHM9v3e+dxkwLMIdRsK2OVtqTNz2oT/5JWAez1Kuu3ix7Ypf2WX/mmrhMSNL4
lE/ceA3aJPqxvbFf/y25ZsioaiZmVAvXIQGTgdQHe6swx18aDDjKe1lSzHtJEwpr3YtGaP1nwc7P
AvPhVsFMrVwGSKQpGQjEvncCprqqVlFpiAyJ/9OcwS6zwAUyGADNiaw4aEq+9iP3B8mggaOGK4VH
PGC75ym8YbCxNxB1/Ty+Dar6qgobP4KdWL4zuGI5TwdFoFXvBzlayZ72V7ltWHQhBkStP844Kl6m
PzDKCav/9nFK14QfV+9fO/n99BukJgPZKD2E5u2qk2FiEbmr47qgKufn5fgwJZAcueaMOLWvt+UR
PHtnlBxpYDckEIpFazhlslaOxmyNWvUpinSBCopQ0NhOTniWiFPzBJMFuhD0d6jz3NZqoocifR8P
loiPPNi4krF2aLQFW0XM1lQfDq7D79/JTCIUa8Yf6GO8ylx1vMNIbuMJBjHSy6mTAL3vlCvMmvzA
8j5pyA4V2zBeDEKz9i+cHimJGLsC8q5mSTIegR4EY2F4xyW7gqPvhS1+AFnR7nv8R3uLS58UG7zL
13MjJDnPoO8lsMigYFFUFXNezgkHqtOVEV5aGtmOpjL7Cx9G1GacpLOyjFU4e9QwtzCUgODfYpOI
R5sxevptsRFLu0eezMU3mdEsZ0+ns5uRb9ODhRrxt19/oqsQ4MQrXBNdWIChDBVb/j9+StHNvjKd
7arnnwoHjcYJ5Y3iOFL30cA2R9MVczPKRc6o9jyt81xwJM2+bmbxPvffb3jqWwCozASIPO/hj+vy
AEy4NBP4YFbHzglTj1SA9rEb7XhMon45L/2nixXRHhn/1hhaaSvylcJPyjtGGJXeRPkGwwkA4u1p
HtlcLjcm/MlyQrs2LJ6HYVkA4V6Z57gbquhnUTMOMoo9F7r/dOCM/e6nVZVuDMQD0qlPvuIgIsDa
Ff1IMLzB8CSg0Mdm48E/QXBHJdliAplpLOA3UUdp/hyy9ieax38CyulVjJYbvT5GmjKHPgOfz/c9
m0k5YbwRR6TKvtSnVgxyqd8BkTJ0sJZ5j5b7usZ6WGkgsjP9aREBD6ysEUIO5W7eUqHET5u72JcJ
E12cypuh/8M6CmmRmLk2vTnorpkZrPsHa5eIY8q+hAjJx1uxEUD5UH9TCJmYp8OhSmX5ZdVmHFBp
5hQhCn2pd0+6jcFyA2JOcWTbOsz6zEhq7thwsrEaKMRMup/NaR/g1zLn5HIbsKFw9e+YJXpzRYJ0
B/ly7J98XyuBC/IpxPNdG6ZTeMWD72vcvz7hNqPsNt3c2wSlNFRBKECrqQdUa7QEA5TUez5V07uk
MLI9Yt/cnJ62GOvBdHZYfWWKQje8hQ4F/w4TtW3/dNvycE86hOwR2f1rohiMdOZ+hmnR8Jd0h7x4
4UgEZ0qG8GtuTNA+BrJjY54Kqia8MfrIsEFcpp9hYDKEY8fCq5W7yT2K4zm6Njbs8OpVaj5VyI1x
/vSdcJ6EsqllFaKXTz2egbDnumguYmo8YLm5Tk/j6d+jqy7D19AD63RyeqwzsCXgsXD2OZ3O3lrt
zYCH+dBxAUwP0LH9Gp0YCqBBOIoqPm/HvgQiynRLrThJuO05h0PABiV+U8xQq/2rLKsjzqvew5Q3
2+ePDcLhW5AzAZCDq2so7o9JcJKadQpM7g/3tcm80DhCxSODmT4GxSX0/s+upNx+4O2llWPpcM1z
auSiZndaEXTHJKy275edR0KT66jLqxDZS//DBUXdWDHkXMsUXjCsOYd6+DG2tcwU+UCRPERzmQyo
YH8bqYJDZnmDC7CWaxiGTHKRYtbu9KsCaLKbn63WK0r/1CDwfbS7LAq+JF8hr62+J5ibV6uWX3mf
UPe6C6qLyTFR2sRJGE7/r9rGOwYwr2Em5cZt41LdhVS8jhyGFkGBgKyhUTTyM1qxSvIZ7Ok+/l52
zBWQUAgdpiZJcG7x7wmwgUTj0EZ3G6PDth05jiuXX5+DFT4zzOtZLXbUmZjb1BSrKb1pAbx8ghi/
HBo4GoqJsa54yj2hUECF5Hu4w19y0fE3N7gaxPpBabswooUhE0FPQvy2W6TY34CTGVAfKaLcOfuB
WpCzoE6spFMsHWNkzzFf2mw8AgEIfcTIOv43sKmQZZwNloY5x0erXlUg6jcQL+Xf3k2Br9onxrMX
cScRkYaElmgbCJR5H51l8nImxEUKTTquYnkNIfSJqa4kI64YovRl5SiIWVMysVdsU5T9BHTpvnxv
psid6aXPGx6q0Reqx6oIed/h10Yqz791E4i1VpdLfFibbdnI80aVrsbxjqmbzIcN5ft0R5K6Mfla
+32yC/vmzN4BGLoTtreYfNfY0YEXY3ssQzwkU4ou8zK4pB6WtQFbLCDW7V548SRE6sgSuTDlhcSz
dKfy+Cj7B9EmN1LLQ9I/IN+OL+V4NZBMlU2iDFx0/PkOE/uu78Z2hrWF5DLKN3k7L7F7btbXN8Gx
AyIMChTQfW1kdMPbUCJSCK0zeJT/GJRyfyqvqpKT/3kxatfrQXfEC4BX8kXkqhDaWE28CW2TrtLK
o0L7VNyI+w7Wf/eZiFzCpA4eGw6PlODuCbO9BQAnPk8XAxZ+2qgTqRX7qnnMV4M/YyWNJrrBnuRu
kQO5F+EM2EpIlOgoQoid3iH8sQrr+wR9sNwy83CzrL9otXdBP0MbPpVH057A/FmQcWKzoCNvlmRy
6H4v3rziT1bswgQKWhIRIsoNP2aqSYlju7UbCQj6UTewtfjGQqtmMVz13lEAYy4vTSUSPINXyNJD
O7dqrMJ3tn8q5ICa62/2bAIKjdCyIu5TpzlTsR267euqP6awUg3PH95wfQCGtSlQLC83g8EXy+Hr
NuEz9kqZO28yUjouasr77sljkmtbCFGSQ3wpzki2c7r2cCfQhc9ke+cyIBu7FCO0GEUh+etCpJKo
+Fu+YguliWpwpOonZpRIcJ4AHhteSW1aQoAucR+B66MT/LdMsQdTZnwIeYvL6QwCR/bAUnSTLGIJ
agLPR3DW9noNetqTV2ABFmN45mRMlLs7kpcfeROZzHe6Eh6RsvUBY4vG3A1G284slv/Rxo2f4xoG
qNqGp/rH9ZMy2l3Zp7deVDXXqqx66AYm2IbB6HsiXI6L4k6Z6Db9Af/c9+hFxA5kcjdP/VcZFumq
+cVTukW5FaikB2VQETDpB83ySQ0WybRIdg+7MjVqr3szmY1ClAKBr6WQwbnpkJGIiZME1TtY0nO3
odlsBfDEXbGyNkD4DQNVyxCogLSGXbIAi8Tb8+lINaEHUaWp4DmqdslOW/s2bV707N6788giCKPz
KzmihzlP9UJ2BcDbq9V4ptE+P+wLveUSllp6TabQr95ZPqxLd9cSnZPSmGRUGixONefoq3E6YM7X
Q6EJ2qpEPaZRgOeDYpoK+2WS56njkf7mys5wJGuJulfoMzdEiCcus5lUyNtyuR+DduTimxX2Fvs3
QuQ1geqcq82flQ8aoF+69qsbYAGC9lue6iy3L3531p7YUVOmXvNdlTp/KG++DsmslVF9guRzCB9n
8M+Ho9uUGTyUhCA6ZffRLZFA3ojiF7DcjjZdvYxawtvnI+JnW24ShuCIcn+/qbFOyaLqlv19/6bL
584PBtvVgEAKGiTCEDPGQNmeSUaGbnHc0mQQJFheJm8u03gyXg+/uQafVhVlg0dH5l+iYa+C3CPH
BaOReyQwHp7FeDk0NUl8lETUdWJH0waqlHAE/kQ4yrhZBa/P0FsC5Yt5mV/LzgUjvi7O2T3DZud2
Jp8nhKlRa6xe/+UdfOc5vV1r0OTHhmUU8PnPyQSKsbQt1Ug3IfFeaWeiqi+KQqG67dwGXpw1ZWz2
2EmMAv8Hq2wo34pSQiAjv/cLPrXyvdn5x0qz/9jzHk/THk6qBEfkfAxAEg7E/CyZ9O+DgXslCjvT
VwE0m8MGgyvHq9CUhqN1l4137s3i/Hgq5IOmnvI5UH87s8d5U9PEO+dv3I86BfJqmgb8QoZNj0qp
kB4xrvYwrN7zwtBy/WZHaBkiCN1RQHNFkX1seFTiM1fwYV1ILKEUPqa4Hqp+cqVoCLD59G855OOW
61T2ivHbWnYO/mUK83OLu6AkBboECN9TTJrzkRWiujL8x3J6aY6wCw2UiMv5iASqsPM80Qu4xToW
yL0s8dfsJB4HdFsUhWaiPUAaNcG6J5JmTsxCUwsrBx6oEFznbSLCmkC5xNz7a/6cjrfNidCTJzAp
HDciZU+HeR7jBKlAyf7lS5MbSxGKAj6nwbwGZF3PulitOs+tBOa5VH/kfamioDtHQUio9HylOkWc
Fn0XUtmBnU6VZ97FLEQqhEEsOs/s816qwhOz8gu/bCtcX1ZabOGZAQrkugb4SoU5rzWHDH8JSqDj
EJyvBehm+aYOaLqh9KThtvk+Jgb2imgeAKgJ7x5SSZB2nch6FVnL52NgmvUuX8Q6SdnWWZ7TKxGU
j7dLyR2lj1xWdCqEY26zvuaY8IrFHEuO7KtQrsw5NS/0/c36S/Lkv8iEbadhSdD2tOrrdy5e76g7
w+iii8JFTn0/LO2gnp6TucXESaBcSTtOKnRYfBMGoyz7NMTWYuA6MkJRsVz3nBZP5bmnZoKbD68N
CHIjJq59ZOPeRODifh66OC6VnT53I7m3V5ON0UvWxaYfw1h8soZfY9Q+n3ZPvQip8azjFuTGO8wC
uQ9iGunK/46PiwsIP1xooIRXyCuU5/SVr5vwzk1s1uo62QVlMN0Cp2NpUaeyaR+wMhP3HY/OdX6/
RvyJa85SWZhPGjZEIi8G49O20OcIhYyfkb6Ckxj3/L/bGdE0TfODOhZpr996/IUK+cWtT6ujLD1q
T+uDlzi1POespy3HdFSi4jd/S73hwScViuvhPyjr2z7LSTuxIyr/dm7fD5IhbQGchJoWc/BPboAf
4T7tuA2a97QxCf5WyE23KkIZYisjyF/C6+amS+vtXfbzVNcJHrwdO/KjHBmpxVEsweZTTrBQHRIA
xZoU6OESSB/pBWlH8jne4QZ7FD9Pk9S04Ope0ayZ2sPmenwFk+KPzE0aSQiy7MK2d5QIxv5cIAqR
PCMafvn9BYFtp+3NTjnFMsc9volVN9Jxuph1t/pMeTZOCOIssEzvREiD4ln3miIVduT1b9pFN4Ny
ciP//IL5AiG2siXDfcQjQC19Ksaq+YA3rv1qAT1XW+pFAtX6uFIeH4IkrkU5kab7+Q0ptAnUsIgI
fYplLrRvRLQGPoqTl8vPuNBHJfWj5mAtYts51ukAllHrwi9cewHDaqwyzAtCxa9EftGdh4FqzRu5
2T8K0tvWOSBESmEABeL1lgn3qieVeUVGeQYj6WjD4pGRfTMfbBkqYrHEW9UBpBwcxvkgvFOxiwcC
XTUKLCla4xRwSFtn3DZZfgPKdgVyegJHzqfWmIm4skgTkwAFIzLkZ8LwyybjS3yca7xEtMu5dj0S
utoga77zORJJte0iTZX0nn+1tswoeJU8Pd2TFXgxg1hIKvjv8c//Rk9ZUKrrhRlI0LFhKwnypPEU
R0nTI+Ps8/FgECdses/V2/gdmRaSDFytsg6RQuYNyS0VwVLxWBhyk4XyZQLKLAwAuXLdc7c8wRB5
GL95s62v+damQ/1suaJVUWE9EXOr/SSWKDzL3UJUG5aQp6bL+MuZT+KXU/mjC4haag1ctyAubLge
mJmIkky/D6tZw9enwuZRrm7A1BPZHGO+AFayZmfaYTs7Wsnict3lccBehCWGSIAvE58OALWYfxfK
BKqcp4m0gPYK19Fgm5yF3/dhiPYdmB16GLL9O6IYydZOukCEZzqmiHr71LigB/iBDEmDjpgD+Oc8
sYSmfgu0EKddnz9XdCNdzih/3pLoZqzmGfj1PE4EeLqiPND5hz3b+qzbLmq75b5df+DDiF28t4HL
6fbMAZ9wbyA21WcwTY6VMufq9WvaEVCMPUvbwrjsctyNjA5HbgIm9xyrjT94ShvO6oaX9i39qmX/
ZhbsTiwdYTwYZ9iQrVIgSFstdrdhPt0IITkMn9FF30axBHTw5702LjmbFaFB9g0k4AyBExn/DdGF
MBLYtBmvpSvlQ7TQUwl5Xu2PSK2zqHKT1NuAajFl0Nx/9RofCtZxufi7OkRcNxWc54R5EEHTx5ZQ
EY+Syk0p0aiN8TFBpJU/rq3yMuMYRempQVLBsf8/tof03ox4BYbakFSg5KP8Q9SKhXlxo3P9j56F
JTMn4mSak/V047a/SiiR2quGsfq4BnyzeLFBlt0dmWQSYusa8qBDGjWgUSXCHk69xJBSYb16IATC
j4HumlUDDvNxYyJS+fu0lE77DLssnFNUJYejQ/emQJTL2Do6SdqqP1eF01WdGUGXXrRAKy6ltC0q
BF30F7A2PKtBta6FPZU6Jc+fDfYjhGX/50J0iWAC6EPhNpapkimnwWpgUvE5eam7iL2ZOJ9GWfB2
e4xBiAK8YYlty7Zis4luIwIc7XUmrJjH7v5XiJ0IV7QRY1A2Aw7S/qm4RDbAGkLlA8szlE8ysMWq
InLdlfgkYT7ChBXNbcXYl+R9j4VFPvkD5bZJHQaIEDq8gQ6JgryFUalAx03nmSjrABrd/KAs5mBR
avm18kMUVE9YIRphQEnIAvp8JRspfSldZWZeBBuQO7IVVikp8ij3AEnHGlptW2dzFHusuF4IyIhn
wkfPJXVBcK/o5PusWj9U98WVKV+SBPFWapyHoYzsBh4YmVAMHeD+RAQ+nWcT2qg0s3FHOmc1RL1d
1iPlxytBnMuToE+xkfr6U7gR48y8Au8L+O5XytuHM9wXV77bvN7OLwD/8/Nq3mzSHdrGvCFDDE9+
mKzljN665IdRJnw4dm0jNs/dulyi+feapQGJNglujEwXzfbf1i/sXEqUt35EL5jRYkc6ed1sFdxz
FpzdHv5A3FWZxxYFy31Ktde3kLv3zOXTXfhW0UhKTt99Mkfinmi0/GHVMa5vCeYLm7ND/tLVyvEX
KUYfIoZxwYdb2FWLdioZKJF6gh9VMfWJLNtCLxYQFhYyONqOqTHm0MYI0XgHNGb4X4VJJrtxVfbI
2YESA65zIzWXoQ+Zk6uhBuXmG0/xFUBaQ/6zDqn2W48sW4vliFQG4a63emrjh/DbnDADS/r0Th4A
HJzTARBZyuXmwujIAxWhc/XJYswQSKi35vsC1bd+xnZ5V8xKQp/y2x5zjeJeL4OsVU1m+suMkytg
OMDf2/oBpZRdyOXvcG4gyYMJxXSav/LcMn+mT0Dpwr5K277Z4ppMjY30eagtApUhhogPQiihkJbs
B6Z4BdlwbdzXk7W9wyqPXS1t3jiOBac5/8b/mS/L2zWB8MRLM4KlXi0GomEeGfktvmCKV8epyobr
Fs1e02nneAewVDXOwrHBUW2gWRvL20jp1nVwGAwI6fTPLtGUuyey8za37Glia14fsTGy29EcCIOb
7l7FZAwNDIwcMxg/yxRfSeH9Givk0xidpTJ6rNm2HHFRFRDDtXZ7gR1yT9DL57hLCQ9e+tVsE3tn
ZsSDbXyA+uJwuzmPe973FwXP5MwjLzYgNOUGLiQ4sK6mlosjN31Yj41ug0s0Wgr0QPReAVGFEzJG
X3um50jYBJ0N0/QgBqi1cCr7wTsdol/G1KRfz2w52Q1cfVXrRrzx+xLpNFxx95dw7HcFJokQx308
lGQQmZ1jrzAJWYLRrhGKZTtAVhkH+/1fzA9o8wZvXJC0iAW+7rqn1/7flV0GqG5bTLQvNsMX94u7
+VVAG2Gu29HerwZNAgdVOVghZejhea1FWxIMLIDfjcwcvwAbCYiMZWiTXjfx/3ThfGZAkppzhGf+
OSagz/RdDXBnt9CI4BB31Mbtx7Lr/mjWwNrqZIQVUUrOTQlkTRR7gfDQwZ4pJTW30K7qxuNYO9EI
gx2mPdolAKFPndZThgrQw6kBKSwuwFdgpYEKkyypSMRDX/isktJe1cJtIdisJdbLDEYAcjqvT4NH
XOReSy4Gh231d2h5GDO8ynQCVOxnv/0j6znitYjX6b06PMTUR6k1vYz44XY9IKZnI4EQX+IWsXNR
i9DHBct32TjYdwVNC0ehIkgV0o5GjIXTOIVkHTs6sJ5gRHCCwSYMqS5VNKsVYT1t0J4H1U37L/xK
VUXSb+/OCVHOFxFLG9uzFgoNUb9apohjlLdxhX9JbZq5hn0ApDZ6ht/V4S4QDr1ZxWlNdo3iTlET
Qy+BwqBdSp1DSXJFglGvlmSMmd1Ieg9MF0He7189cbhF1nppUo/boyYxdIZkwqu8zV8lG611AV+l
g5vLXORV9VMLfpMn0cOpvgZwZuQl+ZLfPwNetS9t4fpTtfCan4phe+YZIBFRI4SxQbiNddFl5LCc
Ikerx8Y01q+7k2lchzZ8pnpodG8RxhLx5UCjE21Qq1v9F6j3o6hWg8wYtbjovyClpdy+8NTvj0iW
yVmmwZh1OsLpOrFGKsLFt0SG/YMkIP+HCB82OvAgpCew0bK+HkBm9F8QFdcT89C1DwthuYWe7CW1
v3cDBXtNYlcYtI1cNXNjtNIc4tbmRUEBq0MmMRMPpt8G5jYdRRkVx66I+NiJ2UbvAY2MT/2IluEe
UjCGePfJFvIPQjm856Qoa8ASU5edbaKK6nqMBWzg3UCLhLNN2wz2SUwinwJaG3N+pnBtMQMoKliz
LJsOtem3pSiwSwnD0DTrltxasljX5tAljHMIr8krr0IQIlekqlpRM/k3rs45eAPNRC5e8idP2lGd
XNj1AiQcjkSxLN9xtPebN7QDBro6lgofxdYeChph35HWCWaC88kJWgtG1Zv5Wc5wVcMzt+MhufT0
jcVWxgpg9ZPIujSzrGK7qmNjr8o2ka0naWoEgX2rVgqEccudtk6iL+ZIvU1ZlY3osF/V/NHfDvoj
562Irx6DGRKfRRpG7O6AnjJHU8N6p6r/3x4J64T+Y34sGiux56J89A4GrAaNeamX5oOvW9q7eEoU
qgwDE6Y7Wv4yAQVJcYq3AF1urRAmXSvL8dStz1xOhnNDkQsPEfS00y/flQMqX9EWEKHUtgBkzfM3
wDxKn/38ibOXX0O7SJNtOUHloOo3U5fIT0TCMICaYDzIITbgBrvTTXC1xD48P7DZhc0l3xMMBT0s
76J3yIE/C11YoS55FwfDOlOVV0uyeh67deTwSF0dtjPSBVC1/uGvimyzv1LlVvmplubTZiTVk6Pv
KP1Zlc4jR7UhWGfk4S9/1QZxIYVjIhKRSEdmF1CiUb8OvJXXDaCk8B4+LMyjo1tdIuug0uU5tQUP
GeRSe83LPKU1VG7qtYOrIHmgBLb/cd0NBpC8kQ9vGv++a6/weVvmUeeD6OMja1VvT+3+eIU7XoeL
9EY+jJP5XqqwlGTvRKHdc0TiMHeOIhPzm0BFa3/4HahUS59l9er3VD4dXCPVFSxGo0IgTUUK7XA+
ML3cFaF4GTNxkbsmwdOq8euU21kUY0PADVZ4+NXF1RAUiTuuaqMg4tOXLDecLmGKHeLuNp1IZ0oN
zjFVO8Q81aCkcs4DjbSFaEdkTHE3EyYCvv1gaqOTt1Exq51DCFsGhFufZmTHexEPWmJy3ukgtfuc
Rwii0sSo6riGd1cy4lGqmXqTGwVSs0sFlKl2AEOfrEce5wJG+j0nN3bDiT46EAOlFTgLq+YVl5ws
zCMcg79ZqfNTnE7ysjl4hsTG2Gmum+xGIkgGSmY67D3QxTSKO8Tq10TajUOYxgnyVNtIeGlbQCFM
oHpOynr6etY5ALirtvcChBAtRpXlaDb76Rkh6UrmOkqpJbFnA6fXOMpB8qwkeQuyhQR4+9V0CGEW
NTi/16P0d391JLzQq0v//s45munWnWHf58zl4SrFL8yrn+rS1JEHl+UCtASGO9Dwb1+clm++i5k8
6UM/lkHcqELncCRNe/FIV7BGLD5GY9y+BjbS4vFzwM1nxJ7O9QYP/6jBcKzn3HNLxVLtF/JAyclH
LhlizKW0TpjZsYi/EBfMJexrX5ExTr6HWOQZJNbnA0LE0pyGgaYg00A3iUKrRg4fKR0AMIFBnhWz
uP7Q4Vh8XipI1VAFLWk+nvT2tAWlt2JMcs8U4dSKZ6A5Oj6Sh2UmR6RaeJiP2AzkHWoZ+q7RuANT
enaqATzw2X5RaWGruEhV2tGAETLRsekdTZEFv5mEKOMJ7bx9J2azwdk5qIW+6Zo5sTrLFo0ndir7
to7MzsCOncQ3ZO4dytQDc3o8fbzhmFptjcauDYaDHm5mF2rstH+pbydkQGUv3l//FB+G3pzEHJik
oAkXVNvhRy52UEsmZaPUOw4cCmJ2niaR54fIPuGYR4a6yTg66CsZI4GKFIfGfN7+4dGa4qwMREY/
uAg/qwydYZHkiupRwbfnSsphOOOfV3ITg8rlAgcVL4c6iq6NW2Y4v6+0mezcxEoE8+1JBWpGCqGG
+WZjJS8IqtOFwR2wrwUFJFQDJ9eXjaH32HPJBXJSiMz3b+FNeNBjunG9nN+OU4pWIXkUPptYgSGL
rj3Cpvi/x49iYQE7E93WbOvmOoKbFhrkR6qcys3/piXGpKNA4WnvHNpoDmGkio1XIyw+sjrMAcjL
zR5vI0VfCK6rFhjQHbvKLeA4wluWedAIBVov5Q/B8HfP0eTFSuLKImQyrvFd9E+O55ShmNqyujA9
NmXjJAIe2Hl8NjoNTHA25EnH+eu+h+SDjadO9StjE5qu77Z1FSzPZ4chk7tcgGqeo4vJ+j4ohQ5t
vs+2s+IQQsIJXsyRFy/HEeD2D86JoSHXq6sfVB7He61CprZG92c9Suzto1NK7cIA1MQ/Z7O1HDPa
uCrX7V3CsGPsvfQkFQQF18iDgpWdbFIkjp4BoFAbEiZJleO/Y0FSVWsy77RYldhG0eqzsS+G7Hxu
+4o1/LC/rki0fGYJq9iDJEvXrFcQ+Md3/apt/o2SNGZGbngHanijq78aAL7BGL5euWKPraZTEZU4
tI4q2lcsMTMiMChnvTUcIr4rg6u+RwI15jg4/h02DrZDFoVcoSswjHnIe9aki/0x9jVf3U8Asq1s
paZneIzzh+d1nHJ70dgbusPyzpOJ3c8vQHv1gy3gaByg0hival/yPGkDKtC17JVF6z6i3+EL0nBQ
3gp50D7IjATybj2orhDlDr0Br8JsJCV+TFbs51HeuytszANoOs0NqiS3jTqwkE9kWHa3w4zIn4Dr
BWAJlpmIoDbXpNFbPuTZKPxBIr5K/q4d5Gc+ntVkh0j3UL4M5HhUzoqvaU3LtIuO8v04T/80ma3m
NWnPQNfzo0skDhSaW5YfmojcARQPl5inWpaLSlKRFo1gjdsii6sOt21/EiSf11LAznvtIZoHwfTj
BUbdty1ldkdS8Vd7kEw/Kt8wyZgkTXtmIKfUC5YFAHZztYN29g0unCSZ1T7RKO3Tj5MDgCPWo9vj
5oz5T9f970XA63HG0vZiNq7wkhgKLnO7NzvQgD0el6DklyOp7huVU1/cMifJZsC69JgHKZoGppJb
bv998qfnfBWDIzHq0WGTbFcmgfF8ajAaySnuKkPR9MUfM+kKInmpqi21iW1ZeIecK61s36fVu+Q9
VCvKb2riznt3d+lTDTVtHmNKUsTEhpNZgBrmYmfOOuslIWQUvmFf4qVokIAyeeR4TsMexOvl/ePI
NYmjtsbMEVyGG4qR83AhFTyqg1fhYB4qW5SG3NvLNIOL4yFQDaGj9s7A4h7ds542sKcm9hcQybLy
y5V0ifUodLj23Xe5BdbXtX2pkWQfm7Pj7Mf5ykPWSZawk2WtMW85XRZoMmr6KsF3g4n1K7xSJlm3
T9FZLp9ju3WGCQNGhHoxa2HKDN9QPmkhp8pO8KSkKrLJ+TED//ifPciAl/Q4kzKsJaOIJPCnFbME
ORSFxCeIZG9nZgRJ+dAXLTYlZ9wIw/9MXI+LkkCs4vftcRCZbcmFfHx8CxfxmtDOnw1P8ej1Wjh9
7lSjUvgzSEbgjRwLI1+/lrTGv3ztqeuBlZ5LevRoVbbC2P09dLmrcZpKv9LSCllqf8bz7itkwlqW
Hp2uDux+EGfPhPHSE5ZxLJiGvXJo4q3IZVxo/uvLQeGsNWAC6wB0UnCOglpuN3f3XWnVvuQk4VOr
u62fHL42z7eLodL/c0E9mBu2WvF1GpMqaRkH/RFEgXR4sxaKQsTuxMPaLYslS9pimVEsthp8/due
iG2K9Hl8S4SWIDq8dTsNgOk7xRk7VRe2DXk5kr3R3/7tvFZCHehr/O36iZNfc7NC1YID1dXjQB6J
POjTOmfF5T+UJGcDqP+nHhrJypr+ZbYHk5iXrzHqwUdAPrwDngqSZgkrN386lUlxbVWiQSLzRmWo
/uWNnqCyUYDftgVS6Pzk6oLdeAcGuq1tO2Gye8hTJ89VArt8ZoUahzCMUn6LVAxKU2bkHDZD6JLs
6pG56EfSOvXnZlNcYIldqkmCEGrf5itI+OoVkKBNliZCfFPW1bOCJpG5O8qEol0YIXyOTLyZ8QDz
A7tThHbtLTAnAWnuhihF/HEcSvvK5pvc11bbT3QJGB2PN14zAEvBOPjjv03+l1RV+5y6ksYqo6iZ
xQV7bzxEUovdHXPqdIpFm/Mu431aettyI+ZyRVXTCfM8Cs+fIu/k1Zuc6vQpxxSroCHd3rlVtMqS
x1mJP4OYoNuzs3ADfC17qc5wvwIF2UH0Ugb8ITxCh49xFfaxk4qCBSww1yFXybzPSFTAwY8MsL41
J6fm9cY1n5CF8n/BpysOiSFrqLG7pE/+pFQtAaH8QEyki/9H/PtOnS8H+dagImLzQ597xBjLgdou
C8xDl5JL+6P+l2pu+3PECuu4nXTuahNuy7hvR+4IIyfAapZ5h0F4xqFuWYq7jjJwC/6g2zsiwcif
cgVnIRs6lo8mfmRt7FNZwvBPUfiDbqmuMwLh8ecokJCnoub13M2S6c/IqJql0Ky1N62IxabqfZ5+
+gmt2HVnjw/80YZk+dGQjb9qVQOIsHR+MvjHpeIuSJeCqmoGFeNNuITIvTNRQTzvu2pQ38jTC13U
DoE4+Fu05heyV8ewl9ro4k9N9i+DNpFyhmC1sLfMmpj8mBpFHB703HsdX47U/+opyUebEOlJ/irh
N3eLPj1SgGwDhg4pJphjzphjzUQ+CAUsSKIdCyOIGl6VmZhEoXI5DIOpm9tHTuPSnkFoJ6CYY164
qmIqqeDKPTQjJvMvQ5TyTbrgLrYB8+r5ansf0bLhO5gCL1uoxT0glpag9BX+pudwovH9/TLpTPju
LzGm1BHB0clj5yJXq99zAoIN7lmjqYJ5a1Z63DJhRt9HdfCmYDW+vpCDlulg/zMiQuWSKwS5fFwo
Wd1hjW0CFgUcLgJDRSeQLMgRDtLi5D58hSPc6swxXjARWxuiyRWmDjbd5ykEt6dwqSl/07k95Wz0
yLpGIvWQvz4lpGEHVBR9cPQPayoa20agIJ80hMtetiyKZ6XCpM2UKXtHT2wWFEx4t4mkcGtDN7wq
fbKTvWDxKRbHdNeT/GYAFBcdImoVLtuyPK0aG2v+Rn2SoM/zplcvY8hgILLkfIFhBZlHPWKc/U13
scBKiAD6Af4yW3sEz+2fWO4MXICWM5PdCxnkKYeYFfhIj8pKGYWmCTA/xWLeuktlYQpZc+hQQwcy
vW4VB0nX1aLByhOB7ttuKvzEzJ1KjG9b37GSKH9aqu1hV5SIafTyRVA/gOafRQG9Jdo8P7CsZRIJ
f6HMXtLNTlEjA6QNcAIdBv0cBcFzJFfgUTERVEIKrioNw+a1ictzRO3HKP/3RVTIaEE35ksLY7nL
Hu3RbiDl7xNznUpKs2kRlTOolACRTofBQ9k6r7nJdtABoiiVXPTUNaJ9kozT1dBsDNulrjtlFGIu
bBMmpaCE9/4RI/JPZeSnRHWG4Z95DsKVkMVTlAKZXqKHIF7/smuEr0ZfeVvBA6YCdCxgvU1lnT+l
s6EimD0jJJP1ylRxT6FNA0bt6/NQmHLlpli6ylq8baFVXHds57u/EEvElTC89VvQAZuQ/wZ9CFE0
drouz6Dg4pfRthCVKXcWExI4/VGKMTa78udfxQlZdVand9JuUcxg+oBPoLRzSs2JVytFAx9G3706
uKJIag3GGXa7Zs21ugCm+fEbInyg5vD++qGorgzs4QKnC31OzZEitzGu1f936FrOA4OZoFiyMBH3
OtXQdW2ntwe4q4xabFmpJS4N3UzxYvJnNIC9P/ny96u3WUc0wn/lFaH0NBixrnXivC/FpvAzG+V0
ZoBzY1C3bPtPZ6OHBEJ1MEJUdiFprSTiFz4T+SYLtUiNo9Pw4ywY2uioKlqY0hd++ykwdw+Z2Cm4
1aDYmlDWL4Qqrm0JEcEaiy60h/8WgQWraqmQcftouAu9CrAxc4U+qV7+PO/hrKQOAxD7VuZVRcHb
t33YTHqkr7FmF099l8SvElFREmVINTyDEZgiD2Cguj7feS1inrO2pl0PGgobXcea584b5zkOOuw2
r2DkmddPD9RbL21TC7R0Oj6UVWysDvjTIjC03f+f2EVdkwCl5My+LMKkO7P9AAniKkVxrwyZqVTw
Li6PlKPK/EnpAm9UEy9VUJBCfffqQ2FcoDJZjXE6zXKYeS9jN9A17VXxJe2ij6J5zQbkKpkUYGWi
BHtVpJPhToYGSRQKhzqYNJURI0yZbwb//pG8QQ+AXslssWCawK+XQ1bZD9j0f3QmjnxRJ//SQLo2
RFbDigiX5GcN1Jh7gbbJq905wwJsGpvniAEKeLYbcswFSmOX1XoB8euT17Og53bigGyoUWkKSXHm
PzlsB4GjUyp+3TpkrMEi2TGLJaBIaLutEzI8ZWZoHwgN+swGMu433K6swaMriqvQdjv3crZcZLj4
4zsVW1IV/Rn1FAHPZc2cz+M4qp7BYjF6iX49Jup0sMW3bkZyHBgAAEya9vKOC4KZhKlI+XYiYDu1
zVyKUuyPpHCLrMvvFAhd3ZhMWRRwxPpHn2mLfYTDvNauwwDErmkhUXDtu42/XD7qmGQZ92d6xOM8
9NFCV8InqB6LekYXx0E1rrYUqlJgGCyTTSpSJ5GQqylsr2LYKbaeqHbID+k52gvWg75iPMsI1UVW
b7Ov0o+48fTo4XIMivVClTL6PcvDgatotUihF6oLFa6kT4QKZrozqABfZbDWZCLJa8pSr+6XzmjC
aouw72jgjTOjGvwe/OoQCEXj3CXgED3DNJvtVMsbu+XccTZByyhgs5TDfectrFfkst+9INvYD/ql
jtpKKdrYLYdAvLH4tsK6fVtIioV8E2otpQK4/yvoErdFlqnK76pwO+oFdVTVDUKMumelR9KehDYr
dYcaD7QACvl6r+vuguj724a/BNR4GqSEvQKGkN/0nsIaIzftqT5OTvQPes4pnglAsmDnBqJbh+RQ
wnkebRm3ps+cO5TliA8sbDPLpPPMa16QjkJHAMPcHmnf7ir6dc12o8XQ9ydEOQJ5wmLuVReAZg5M
u9oVs510VVqJT5CjqI3M/D3X3Cs/rlb+tMI0ICVihZH0JT5eLBtuxHNdGhl1gdz4UXppIRXFV9dM
8SHXxmQh5uA/hlpME5lhhh9KoLNa6VUPte7+bSjHdXbeh+64OfL8UiRurHA3WySOiwna2zczMqQW
AcggStbB5XVrzJ+mmxm2iXpXZPvdGempBCNHV8VFdRHBeBOz3hOA4u/xWWGI+TS4F70CSeum8xox
MrCls06xoDPcTzrqyHTIhLH3G7pXToUBEK4/Y5DaSoEc6LdftbwAwi3ap04Ty1+mgqyvYFHmVUhI
RVp0TzCG18djG+TqEtVYyZ54Ywtpc9rh/L20txuu6zWfxgfzuDZ7J2wLMPWTaUKhGYtGHXzx6XpG
d9qY4jDuUpXUgoyfwFg80uFF6wkZWWrsUeCMWqzlz2fEKVh95WRxw+Y2JxVdotGCSPmkEH30sO9H
ihG6rimaNk7Mi9o6SNZ1iHiWyBQAdtYo4uX4SF848Bgykbb6np59LxNzLN0Wg3flrZm4YlEDXZ1z
H7YSzZ+83+DGRZZvUJmjZn2pTvaLUnYYYT/Nk8UCu/iJnkzrC3jSfov+XIIW6DFWNVDswH6E0wI+
1RLlADwptIdYLAzeS3pN8AJU4beyX6rv0G3WrnW+KU2G+1LeTo5tvohP8RiHXBCWWjSeczDuMfzJ
q2MLPGOf4eVlly4EEQ9A79mLKyoAoOOkAJ0jXV4xDFJ/Bm8TXC9xBb6Fog2+zHHYNNvmanBWjfx+
Fey/ohbMdL6B5WzGFRNHK2l00aq9SKNVK8LM3Swzp5E0a2bUlIZHkVnbiaEDTpe5ojOfNUi1QUA+
ZFGSQfwsV1ZFopSxknBDTqMkN32mXZj3JNW+D3sn8FByEWkHQfJA5ZqRlV727lmovqOHbyr9jSTE
HT4x9o/a6mTg6J3Hao6HlbnLgPWTrFAwtB+IUJDalmONWtBrkkLvTN2nAFattAumKPKucKszHAW8
v55lLFJ5U6R3G1UjsyPrqU/crbQimLyMypJLe/qR2NBOQqLrZJxOtsi+BhErNH+Ug7iWkWwZkNAq
YkJp2l22hoLGiFONrtj1zeMeXOBkxU/JxzNnoV0usZE2BeefrbMO7gDMoNE6xf5GuljtOU/X4T6J
EwXbsU73YUQieLsQe+zZZKFloKOXKGci2JFl+R+mx9ytv+0m4xqe51HjLaJR9HxQol/2M2DvlIK4
h4ZZuXLy8PU62WxYuBHe6Tr0Q26WWwhLWN3ZIBlRXeXzarhB9+ivCK3URy3qAhodBzpgqJAM+U4r
tAPpsBLNx3mQ7m3/UhL1wHZsHEkLuLhHkoB1ADiAY4OOC83C74hXkLH03wpns6UQ/w/jbONo5232
B7eXBGAcNLOj5BDP/ahr3TXn4vvN7ZKE1kQuOYZWXA15fRCTZtQpya3Xr6CJBRgA/WrYURho6l6r
Oq2VjWcGdnNhBEGKc8tefwtW3MIB+ewgufWhMABAAJ6fjyjuEbFndMpPv/mdY7cmnqv7eRIijfQC
//2tTv6VFhpBzf75GILb6uZmuMrVse0nEpDvXcTffQDN3BisXaS4QsL7QpWzhfZTUtsd76lvPhJX
roWlLpfrI7MbQjiG/g9Y1xvjc7y6UCOGIUvXU3dHJtT1nbBWfchXtsrSE0JOgIMAZC8UP9WYwBJq
O93VLigPf+QShUePhbQ7dhvrwwMDOHTA1lG6KIqVFluOZYe/ORpu7TvQiinoBEW7UDT5kSN5+tsS
9ZVGC0h63whnTmmSvxLBBqYTauvae5uMBlU/3hm3g+DXTzZ1EKqpjnvi8/oee7hjZZRd1Xs2pq2X
fcCirop8QL7K1o/Mzny4Mk/dt+3ZPt9KKi7Z+VZYqg09dXkfAAOwkcPuLrDRSkv0iraMsVHwVU2U
A4W8+igsgmgAQ7LAbmh1vfPRljd5Tni70EhfM11DiWa7ajBWo2l2e/sefzNFY5mmtslODxo4JpZI
SOiQWj/X2eDLpnaf21T5g6iBwyxKHht2haMJqzbCkivgkHOMcBzdG++n2EeBJlhR7WB+pQDpk5E4
j81ysx3qMZe/UTsCNJrpiZVDMtBvHHy/I6fTlwc5KxKPR0v7P10ynjksi5aEcZUEkgbFAv5aVewN
kUcIVaL9WD4/zT/ZogVIGBWNqKewcadtU1Lu+38Oc4/uwZkCjSzqOvbsxJYIFlsFfQX/cya0wAgD
rZ02yQl2HHQSpm2MGCYdLMXCmi1uD7pKb+A9U5qgPRYDHtobaEGc1bQH6wBsaYy3imHvVogjEA1q
2tS487/LfLLj6YHCd9JxqvLeTR8icRQVtBofVL9Ar7C1yuPmPNE7cvLDNl0eeLu6xP01yoSQkD3k
1BNE560LNfEJKWANpbccXfR0B/rGqE8JKKK2A78tUSo6Kia7nAxadk7rBZMFcJ96awfd/pgnH02w
FeGERTF9wjFvNlAr+mkBpBAXL016im/mYTLURDwy9y7u18HHjhQ3gz6fkpVrBtPiB5/JrsZUiVrd
S3MFx71gxu3wUVIF8RW0xhAobbBLvl7G6vqyuPSX+mEbgTSlACJoqUgW3IfaG89pp93FPFdOo+xd
rpJRoMTmxyCTPxSZ0fy1VaMqGNfHoBJlSqIV0gz5OOJC5zfn7DkKOew8Ogimnp+zdBpasEdfVouf
S6PtaOxl+nmK0wyuQ8RBwyNC0JJfMm1SMIHDEMZUeXedh12dTyQvhvzcVjVHWzXLSSPxJaf2AqlZ
PZ4u7crYKthUpm3gqMWkRUOyzMrWXWaunEjmCHtb8TxmNr7LKUr0tgzSkcit/U75Otx4NBGhQLy2
p7bJDC7bp4t+QE+3z0EQU5OuxQ3FPYRKj37Hrcyj5TSS77Kp7/W8rfIEDJHA+HMGzMMyxJqIspdU
DLfRlbURvSu3hBRqJfytDgOSpZwmvE1GPdFQoTNE1Efx7VTtn/PXxOQWv8CoMlNr57PdcIW4vZc/
98zsPbKIShqR7y/v9Lc2/cJXN+XuM0TmJsgfbjYah4iqg24NOeRcTMgAFnxe4usvQNIeWEmOG/Z3
6JwFVhLh+8R9LspqVj46fs3Y5D0H3q/pG31vcpvz1v5W9mePsFkD9qdrOCt0Hu9xZ3PXLTDR2Zw1
VIs7Kj2PQ5zpzKQ40EBUGDHUUHnPMkQRce8rP+4NokNVHJP8NfU5NYAKcsNf82lIGcD2PHurUeGs
M4Jgm1HRv6mt2iF9Tx8uYDyMDtWcPnv5d6V66N8Zro2VAy6ItRouXk223h1W1R4a6EZI2jqmqyy4
h3cEBMtlASuoIvoYhqjt/qkOlBiYcpa+snEbKBWGFFGQZXwWVEC56zfjxkux/v2LNhIcm7tu6DJb
GdiD6rARFqeoD9SK1B8TGRnmWGQQIMgooN3St7hdrMDv3VO4nJDqfnORMF/cZv8cdwuWPu5Te2TD
zodxPxGXbHIz0SAE9m7xnClPKWJnvV6Ud+7J3sFt2rlmRMJszfjTAeCQReX3L1c0sM+qXWjotOCv
enFaQpgsCmdkPburzrL86XTxLRsVbrwZxZqWsFl3MdyHpUt9hiZ8CXgzfybkWOg6tr1mkq057lk3
K4RFScND9NCHR/CIwOflk+30LwDhHIuhfjB65H0Zt3o3i2SReaMBk4EE0ZlOxNDizcsLI1jQPUfi
gYnydpE8aECIaqOgAvU49aqblTPR19fbTxnPgC8d2tPQU/O9CaamOY3aosueKZEmHZTAMiY1c8H1
IoJ7GVGrBED3MUwmg/OXB0uLRidLSLzHIctS+1Y9Ps1EAXImETeDjcn0ZC7qBoNVN5DdnZB0TY+o
snMWzUG1FdBej1sD4JPEaZ98+9E/vjN0eyMnk2V25PqJs5MRX3pbWUTBAc+UGDmhhsoyM1DHaHwp
QBo5vcOfRdRUGpmV4gH17l+HxgPdahOpwLfzrheagoOuLfaRaI63bpiKhBEjjsrkG4Su8Ue+ymoI
76Y0kqigQBGu/1uvD5UmRtasqnlE6Yb+LOZO8OsRXrfYcy6l2zcxrjr2EymgFgPpLJNleC2xHtK2
hOHArL+dlorQLryiPhXPSbiKKUsy07KC6ycOFZ5O1YyhoJZVy1e/Pp10IJOeWA8VmrPJdW7+Uvze
Ep3lrFWkHpxWMkKMEMJSXZhaqYdZ6l3gXcXCEIuluIavfpx/Gu7q0ail7stE8Wkils3uiKw/TpjX
NENTlnU8ywLusnmlmRyX7YZr1CpB/wSFxAHg8zWaGQJJNT3iOByqKYUvj9yntZAAUSw4YSfevbdM
NSo53p4a7fO/xklXeJrD+0IXBT3OQ0y2OovYUKQyIWyCc5ANiCy+MFNCs1wvJTn4DlWE/msNeT6I
9WGYY5xN/S4yZeaTjGaaJ7cMrkIe69y6nFZnd6oKUihSp7WY067bxwrISiSTEMPxUCXUMNeB3y0z
M+dcbQ1S6ZIc304hMkaSGXFqraMXp7u0eHZiIXY8o6WQoFnfu+56ia5YjlAtiV3QXM/u0NHeTkuK
+zKNF7UBrK/1icBfCxHb9gNw0KYZXZE4pyhuxKI/164NCpTXFcXuXYgS9E7cwk3kBIpt7ldxc1zY
sn1VW58O9ZY92hLQVXdiKdOFaXFrkIdzBO0KcmGdWmHX3eNucmOfwlpMdgd/kKEhkZku5+l3Okcd
Ei/jctUPwfCicgTZLtowF8uZlDynna0BmqmRzn2y+IDYe0d8x054QzymMPtuTytQ9XNJv9Qbkse4
OBhAqrNdvcH2iYNjMYkbMF9BlcNSk46OLQgX+XH+TIE453Ql1JJN/kCAYotWr5oY3WohUOfIuyhF
ypG0g/nfrUpMd1dw+YCdl+Z6jGrg+RblNNcQuuu31uUlaMTdypEKF5WBI1ZysFlB4guCDYcuUelJ
qNPic9hsQGVUIcYqjpjMb99qfQE1Vtr0T6kGAfLK+8IPT3Vo51zlAuDqgzPzqXTaEEvaZN3C8NY8
sr9zrjaNsN16y8e4ZuPPue1tmLyQ+uW1R40CZ1ThmrggXscxUrQk6nT1aZg/K8F3f4pxzjS3S6el
alHIlZvWrwJJGJH+TOCIDwzWvwRYwGQlTyDTFSfMm2ofxd4y4twkUq3y2w7oeB9K32QnXNQhziGu
aPa4nfjQae50kjAp6kk9d8hZboD5oJlZcYapexAFJk1eoHg3w6wNcusWb3WRJjVL+vQfVCUvr3py
t8b/b8o2IR/RuGYEJ/dSjWghNP47asZEirOElVFuRoQj5ZqRGwEDIll1n0Qu2vkjir7sQf5z7CqU
ppdPZl8MjAx5AhwG6KovkDVPBzaXNfDaxzdyZF8xICV4EKc8FZzqfK9UMYT4cFHh0NFhTBAMnHT2
IMkKCYyvUuSxPiFYWw5JQouhTNVdvlMuvmNzdEQzRhDC1gD9rLOYuL8cdeg2shrpDfCMb/SPDpVG
vYlO6ekeX2NliRAygqEjKoXMFuOxDzoDSN92b+fzKDZ44m26lHAnr7MB3BCsRxx+EC5UrzfOBSJo
4tbnqO1YpfSTlXBBnGYBK8rfD7r7fbd8ZdSfWs57hUOadVMXS3H6/51DvYgzTy5udp8WrOYHZz0x
xpMmS62wWe85y9UEwt4YTYQXRIakAKVx/xQke5ULoBdrQw95E+SWECl39uC2lUspTIsa/ktmsRRb
Q8+z8UfOE62mXxHEG3lbY3fP75MZl6DX2rM3cFkw05QQU5N/HQvLxBxblWoXXcw3w8zU8VRH3uEF
ihMGfWTCWOqnydGLF2/oBwo+qAS1fvn32kcFPtmDcuIHFpEoNizLQW2q7Y9sJxcKSL+OgXPbaZWf
gvLekMJFCqsaYFDaD47k97tPrd3zJypR8HjcWOnqSK6Af1wwPt8J84ivqMZ7png8kqbeCuSFx8jT
G80va3NSYZnq6D88YD0L7u1Aw/HmEXmGzoTaaGvDZTaHkEmCvbIyVRLhDWY4U0uhihGJ6sgEQYuL
f0Vxju2Z654JvEKjs3ASRCvPY1dDr3Bq0IMEOqQhxkM58H4wNZse+vswpu7VYxM3UX/1w/lH16TV
aTPKwPYUQ1Axkue3kIJ0Jzpb9f8b90Pf4jEUFvW6NdaRyNM4k8nfhxM+yfREBfiTem4LRKj6Kago
vWFhsed9GyotI+f7zEfCyzLcO3dSCMpTa3A6CniqLTJb1Iu4ESO/gHHymyoEm0Jh4Ai9gHp9RTPY
erjQbefoSr3JLKhoaQIwdZk88H04n5ljJRKxG8hTLnPc53AWdD0robEQ1P8KqwB5iuRciQ1EVG+i
QZDaBJs6fKMhEzVHkYlePbIV5a2PLsNULj8FyLcyMglgC/kGv4BDwKlbmrDqy3FB5uaMM+LQHp42
29eZDGDt9SemKRtnWXESWcs1Sbnhx50ooEiRI73Sc49yNcAxkbgzwMHhqzgdicu2w51DkxfuYIrg
gyQKudD2eSiU5p2GV2qXkt1nNEVndBrXTsTjHMtVDpUBO5R588d/bAU9odjoy8gOkUxWJLntecJI
EyRI420PzoOwUd7twY227S6URoLIEw82TeRuGa9SBcYLCbNIeYw7dpbOcr3Kr9X1cBQbC3qR1LPo
tD7sb49TfwJQQb2jrkpnfgHXF57d3SpnON4iDRXpZBN+Zcqj32c6WzLWJeVovStfVbf1MRQjDnoG
dA1NmHizNviCRQeNMRk0Nk00UptCXJYAsf6nTc+wv9AwYn9BRS9+/HjswwBhSSEtg6W1sdl4TYYv
dWRXiBkElLcdGbTW/E7ehDPAJDqnZ70ooQDMI88xjo1ooIDpa5b+kwVGwxUw5l91qNjsuIrJd5lK
Lg56zLp9J//zdveIqJH7seqU3zye4zQiedxdipazL2qRVY743WWAU+KHKDY54DOKS6frroXWGyf0
HGHS8OFjq4E7SOSdkxkY42AxsqOyA2YMeSMT7iDl7SVVpkZzLJRNALFalVKrv7K9tFddrtrv6XjK
LoAR2d+rz94JF+yw3JFcQmxNsG3I9GaNwnU2eYxXfEdlwN+kXP4lem3g1zapZkk3qocFja2VlRjj
4b5yoFt12EaMUelZfYnYE/IGXylnNOOPxnToT5457aBXZfjff62FW5/+B8B8dcJZk3v6/ZIh9ora
9Xnta89/dJEsyHQ0lBM8Al/VJv45FwOpf1wN5Mf22kbuUh5lit7WsZYbpK8Msl7NY6GfViyK3F21
73x3OaP6aYqs2kp/INkKaySxSRIlYgbEQp37j6evj3pNWNiIpWgBtJ4EIhIH1Ev988Oli4/WcmFz
nYBgHQLEimiOKjXSm7gSELLmq0fZYKGWT3qznCsBzu/2f/unDSQ3Hcyf1HwjTNPFieG9iYr9kyH6
2X64295wRNqK/nbeMFzSDlhPhPxE7xw/ygc0qXYnqdqqvvcVd2ZIP5V0cz8h3OEHVR8GZMq9NfsQ
sA+JENhgrM6wP6ncAmmlt5026YKbsoujgXJe1zzYMdxIg2RKB/mbifgWLqD7WIgSvfbNeOR/3QxV
nUnyfpeK4Pfn3an+EH0FYcpkNeqXw0vBR6KjbXjWib1BsBwVAvY+Dgj5IQhoPYqse5kE88D+lS/+
9nY1IyZQoV7iUsAHPSbsOkNLUFCIZ5tf/6jL4tsK64ZAsbvLt8EzyzSFO0z+yemHOuufyeXlfzKH
Muhn/L55rZQSlKp2ohJEc005wOFH60hj05IK3TuHzTfP+f3qO9RUk5930pctus5r7ZFO6B218T1P
l5/JLl1dSREvmxpYSnlJl9ZILjW2+WZTdaFIb0+82U6lWk7qxhJX2K0yUxFsp6g2OzUdDg9ySzZz
k3NPSuCHBoCX/jPYWAlfqrSpQMz0ZNUN4B02WDn4cup8LWmJ9EfChseH1NhgD2D8fkTSh1iQ1/oI
pLAetZ6spW+G9MQlXKNJeNsgGSpZql3nbqvcxPFSg7TuTRDwY9Y+Jlihp/u0R7Z6Dx3ni5aT/coO
rnnGBb9lVX67MsOwFrFxVNsolR4WJMbC6JtX21E4NKfVQ+BVWFpKKiA6zW4JRx4Tbe5ol16VssAC
jb6KyQxTv9SNF5OSSREDF9dBOuuX9OFW3VDO+tlXKv3wrBMUE5CXLzDRsHrDoy2Y2FWYWlF0BIkO
fZ4XBV9wiyvmAUf+TIVxalFTcteD36MxI04JK9+0J6hx7iUDkWz/k663Dv4DbzylMwGh8nxbfV2D
h6nRbLjhV9cKxL5/HPIT1EuDu8LhXGGogasmkjnqez0qHPcMbeoRY9RGjSuwTz01Qnt43XD7SuK4
f0CwPTTcL2WkHYs86LcEZkK+V40FwCZpH7pLeezfD9Zc9J/nIlUmfgTg45zgLwXAtZATwSGPAkQg
TuedB/TItu8To1KkrvpACxYc/x3BF3WcIo+ANbbxstJmAgEB/Uah/xA+C008grXZW0Q9nl32387f
MeAfy5LvxSFq9tCERt9HOHcV1gcw0SHH5nz+AUin7PciWtMCDlGuf6vpkYaK4gXirT8XbSIW6jjU
miJvH72N/Z1O9hUAJjMUCnUmvMz5QF2VbQ3unpKD6JIIq+w99WzrzL31ewCzb6HFqRgH+zjUsrMc
fk3G4Q3wptvQnj3yRheaIKaeQPJdZltVJKEjxSEb1arS1GdPV646F511ofaVk/m28Ld0iLqba8gi
Ht9LVhVVBJgD/BVA08GrvOI0NTn2cFoJVr7hcRhqyU8VgDXm4eX6uo6TR4gZWX1qpR5Ppzta64Bz
8lMGggCcu2t9kX9ud6iMJN3S1WwHqy7aeV4SNe5+o7k9MZWrypd7URet9d2TrPrjxth/jzpZIfGT
J68Bx8UKN0vEbzVSUABIOCgbnYFtMCeias/o0koJ0KxsROmPeIGFHz5nyk6D9ayRA/iby/ZFYZOV
3dAJhHczh2oMV3st8viYw47Z2XkIpugO1VFXbhTlgSMIlylZLeravxmQl5om39iJor5N/NQ2poT2
KkOU/p6+wFWOGUdACAiOHvp09m6qHBxSEwHzK3+vBf/rk0HXOwec++gA9ej/ayjEChA8I5fK6WXF
M1Fd8wkZplkiPRMox8lF2lodSe+h6mLV+ABDl7qqS7o8aIcGrOpQjYXQaf2moUdurNHO+isHSNib
oA18i4Y2jNsZSmjyba18lokPWJ/0P7PpSvYPrjhRDgN8ZRzE2p0MJv4qisJ8oe/3yzQMEvTL0Z4r
xSDFKlTnz4dhqGWytYogmRls8fYeEFRVPNWCb2kIZT0FmpjXffIbWdtduteSzpBcJ2Xi4CuHRrHg
2C15EDger1l09N00aeBmeBZ5kFrgkT8bnJKm22n0f3ztSk8sNKtEKUghcq3j2Z6Ti3fJyEcFMONz
dvrXAOHHklQAC8IGGH4qHwm49phrRtrIU//kL1O1bEzUeQ2tKaUZpcJKk4Ez6AizrMRtTToYXK1o
Bc4kP3nYXVFGJQQz3G2yRwIOA0sJmRne7LjuBz8SW0k6+Rll3HKofmtArFDLfvjOegIdRNRQWvX2
Kzr8SHBMvwuglNuozlpJJwPKTG3//SZuSgqqCqnExtbS5ViKQK9Yx0FUngBKDFWEs+AaGx5MUl+N
vl5iA7OXZMBeVgfEg5KcUsoLNiUbMuShpbmXWakMTLQMNlecETIOsMaIOSz8vPZqCTX+meSKw1pP
wi29CQ1S++QHRKN/Ek8p7lu9iCNr0bNL4tfzbdycSQW588UvWVMPLR1ncyLhWAu94GfRnbGUqGlS
z5KHNdesp6LSZ+Bm+YFsjWEJWcSw3sfBwgMd290pTBaunrVnLxlsYXfeJcjtMfooxmsPhqkUsRho
6gfo2gfvPIBoMgFF3bp6gVta6rvx4SVqWyJMRh55f+WbbtaxPNgiSbROjFvrSkJP3zNSt4s1yw+g
i+91hO4Bbp6UjYe10J5dmtk3NMjqgM/VHL+d0JYhvIEMS2dZdOwo6rZ/Aj4C27Pzr12xW41B0UBE
dYrQ4m96gsMBDP/aft33HunWX7P00o9Jic1MNFYYTZ7Qnz7dARUNWxY8QQlDyENgLqxzCXLvJNRT
kPYWqPikdnJ7oAn3aC0oSjHQjVwb40pGzO3l+CQFYbLAxv5AUGzqXlWkxcnQc5GjdPlMAPTGZUGb
kobCF23PXBo/pDU+250cHT1Cz9e7QTzBHugv5l1rBDfEMDjyyf7x1GRCIuZTEWkOxWRvhwtk9BtX
NslNpol+a+IAHKHjOlRJB9rvF+19uK86GscuKxqataVjmQ6SpyJ8FO5cTgobxLy/7zidfS+ca5VJ
xEPEJ/QFIHNQvDr3iXDmmpxxOmmFUQ/cWwgawXmAPbjeNIHFrfmNrhNFUP+aDSJHLOx90aW4WByt
dg8Clx2/4xg92oq0v9Aousac1P+COdMZGJL8Bvp3O7RDgpVIBktuKWMfeBS37Eo1k8Qv95l9+pNo
0lk8ZpJouayIsxoglqPcExWXU8fgioDeKkUZQ+h785DyHoAlQ+8hl9L0VyuA0t3bNmEVtO2nI/lf
CQqxKfAOIla2ii+sDpoYdb6T9T5HSLm/MdcDN8hloSa9ngdw534lJsTJRMBI8f6onxa7sHW5lfK7
KJqKVf2H6kLq0sHJb4+yegcp3MOzmPxu6r0DRI1kYCpjGuZot5bETB5g2nbGy90KM8wOaUUcjZ1j
8zRdhKkTZ29J5Dy0TYHm4obRzdbhR1UVOuH0l8sNJ0wN4vuEBWd5IOPH6tWzLXcwLK1fY9v+yUkg
ASCLIISxZVU67dBzXR2VhYBxt2zLgl/3xp5cHxK0SqSeT/obI5MOu0WURHj8x4UYVeEU/ANtAxYf
ggeCNCv8J2iZO5OCaCxOcQ5M1Pf2Dse4FyCnrl1e2+N0LE09z28MqkgJqZCjprUh7MVOj2T5peUC
Xpr/J667ZHMiSqxbhc55OcPtVn/+Fgk297y56haqzeMbMxpnFiDQtk21tYWnZb+43YAlF3cNrl9t
jO922cYqiaLgjKtMccJxzXFf/Icrvl7lbOn6Yag1lIIu/JGI3J70orduB8A3joARLTC3YBdK7d8D
hD6x4BWCUdegah0ahlZruW2RM2KsTZoTBGk71mIMWkqpnpovQ5Cd6ZRdFO3GXHWCy+nPue/oZD6w
wq5Q1Ep+wFDgNIYfZ0dTLiREKDQDTmhIQJGPENAwmnmCDQqeAJMc0+ZCY+c/LPnV/ZlLWicx95xM
eHfHF7R1T7tz95bk+z/1JI6zCpAHTnai5ga24+XZ+iim4/rZvNNzlAlhLn2WQ3r3KZwc4mKP7CxX
f//mXrtgLTAEThCRjS/c/AgkWH1v2Xr0aW8mKxSXaA7SzXAWk8Dlw8X84UQd21RYkdbLB6Q5ZJU8
AYqUNt8IVi3BPp5+Q/xVqWD5jH7WGuWbh5/lCu9iFLrdoAAhVCtSnguvMhD+++BKwjkgzmb3fRT0
SIBflplRw2X+VRqGKAjbWTcp15sbFOcAP1taOLVTpnvpYl0Ui1qKqUKYB5LDl+WgY+kVbSjUXQ3c
LcoQTD/rxltDGt9vTsz80MAIQS1Ob/xHEY1cn5GUlN7GlokywxyibGE5PwqURXl6gBPx5OLo0lzl
VN0FgeQwfV9AhFc0JPwmfSOC3R20443F5CllnEIqJ1zqd7PUENgzyS1Ot81YpCOu0Al36nH/L60n
2jW8sPH65kYO+zbVuOYeZEzPyeBqb4Ik02xTPPFFhL/2oU5Bgja85H9G40BJevXZ0wlPO5pjPIwn
906nPWi/Wv18Zcm9ZNAsbX74saNDxgCGkfS8ryjxQQESvZK9vNrjmriTWKmf4LXdyS90HyXakBeu
gPdfmVv1j3ovbW4bc4OeUzPhmD+VBsNtLd8IrjNY0YRjcWdZ23Wyq7SjoeUr99IhH8XSkxtM2dCa
P+E02q3CdBl66DsrkTyvW0GaocWnfyztXbH4SlGXvcgi1NPhwEJ7cXQoZAuDnsjP9kKAOJULlH0Q
g9ZaSVnrWeAN9i5FlozxXA4NVNEU60mx8rwJhPjnWvMmH2Fly3hqVJd3tv8Oezy1wLcN03ijKRl+
TZ56HagwGVNYwjPtd05VQDDcYeQcmkpIzmS2BqCWU0V4lOpP9MIcM3qeOpDYFvvZkV6o83Ty9cth
L0Fs09DisyOacshkXZCj/Ly9x14uLm6WMlzl/qHClPkN10bkQFdhaNZwzG46mAWU4BViilT5RZYg
ZfFSrXhRrgHFoQUcXrq21rBhQXpFPKuVj/boKd0FEn7/jHo3PSJ3ym4B1hFzxp0p1OZu2yKtr6bw
VvcdsY3z7hUClM2uMVsVvC7LLsrJZcrIvjwB4uB10dEoOljFXF7FxL7hPlb3Gz4tcBk8WQOVxqV6
qMqBJJpubxo57VKM0qqI+GzIV8jSC+rpZegY/R4KEHhgKwjUNEOzBCPEhPmIn3UkDh6NmP+EXbC+
fRWUro03oDL99waWPYfNthH0PAcZI1b5WDNZOY7269RcXu5dLefw9GuS0vubLuauBA3bS3m7bd5j
w/blPiChtF2d1zrPZaG6dlym74bqeykpfXl7YfA+FKaoXbz2LGRYGg5Cjrrwgegy05+hTSmq8UW8
ojGUsD0OaFR+M/ylFak/6WRXO02r6xZ4AKPOTUHHoQuEQqKSs3BzwQ5vvx1xqCVkjodL2a5UiuRr
x5sJ8hqjY8ETt7NBXEq+El9QtAgVoKWZQbEZz/79d0Flrap8LIpJvy7QwJnwDrlreJsazrRTLjjD
EM4XNTbWA+Y0fDvbBnEuR2E2BkoorXvoIp7fkAviDKiAO6P+8wBlpsxplfdVJufdwdJIT2B3o4ZR
J1MRC3pf6pEn5LLB8xP5YyzVy6GD47glACqQNAB0LELX62Z6YISdEmsif7yk/Hi6Rfq61cHzFOgK
3Y3064eZMSCQjNB4AOMS3esMfnnqk6BFscSHcQ7nGSQ5D09B/1Rkvyv4nwokVgRVBNdTlElwprnl
L6D3BzvnQ95ruve6AtuONZKEHopHbt86DFxLYZCLS21CE04wiP1GaNKhs1Wz7ZC6jJahUp6nzVzF
SaJWg1JGfWjMtGWz2emQmxCu8B1iEh5Ao0BlLaBOxRDhBWIGISHlE0ftD/fRISOo8n6Pmd8VSDNK
4WEXHOsUJ0kZlt4Vaibq8bKA1NFIIsqjmHp2Ouupvu0wNR2OWsW3PENz1kqmPTnKU1XQDVofn7Ek
gEqEN/Ag5zxZCAlSkQ2QlMzPUTzXjSxvHatqcnrjIgovjsv1vc3PjC1oKF3Z7q5vKAg0EYTmHyxh
y+Co/SM0oEe+rk11DR/VHa36iWOnw4XdDPXmInyiITF2fMpJ/7UGqC/5WXkgyhhFia47Y9kfnYu5
oIpomdb0QZ7sau6+q2Rir9X/YTfcOeJ3Ogr9ENmbr5SnBj8E/d/VyZLGcBOPl4H6/nGMQBE1sO18
HItEkNjUpl3Z55WTPfEeAOhPFQhxUzEoz5bk0K33EbFGUL+Y6NJuhxzNnSy5JTVBmcrv8s/G1eiR
N6G7Mmx1As8Rza9oliU2AO8gpRQo7DDYO5R9czk7MF+MprS6bRf7VHC7iasCddHzAmBWzyiJXFw2
7EwGAQmaNQUOKWCpwZoqxVNM+jh8su/53jAHCH2G9fsRhcnblkenHGW9GoE4XOP/SvYvA8loBrfy
TqAZNI33yz+CqfmFs6VbldVhABAbtCK9bitKKglaCBDLdVgdAhg4d/uQBBila+6BYpPi9eBexHBB
rlDuY14IDs4i1KD1vsM6tOGVXXO/JO06RV3oCbS0Y72/GUf45h0WE9tO754EyBHu+C/6s8QORDnM
CxFgqxlGJsoHTQDISp0GWyznyQZVIJFZJCr/BxHggW60wEXjxyy/YbUNRiTvxJaZ4K4tTaX4R3KA
3fz+cpLCt/ktQPmk8JdcYyIoHL+tThARJevI7C2fNuiWF3GhTb3KFKBXnum4w+QBf3TolXMYVxw9
iIZPYSEu8CVCIvsnYx7M7uNHosI1d0o+9wtJtnt5UkHrFwUT8wMYHXhIgTqqxBB5ue/cmAOnzhAz
fi7gqEDXBnAH8B3/OhwxFsEsd3eJYFSAIeybt7Bqc8S0azHngr2twCYzAfN6MpgfOKDIQgG3Ho0L
1uRm5H3zspJknTYn1sMlN3qUE1CvITYipX1OERkIkggR4Ge6G/Sn7iiJsbigts3ATp8RJWb5q/aq
IeUTbaPd2YaQemIZTAlCQf0x0LN6TK9w7BTtSEE1ECtRZjAXK1MX2CiteruCpOOKMmacNi1Nj5lo
9VKOINAKG+EpkCWawpTeZYdi5qMU1dhhflQSGrLea0F9Vh09rwip583vw22UxXNG+TgCo744vGgn
NDl7ne+HdlTR87woi6y/6iA7aO0ubLAWnvOT1p2fbwYfPH0mFKYiIGzPVUv442ewTIDQb9hxCwnQ
PlLnBJdCIQQvKvtSnJnHoSjxEq/jQiEPyT9qjatZ9KXsfFCzd5xFDQBrwMdpb/hzFriupF6SmUwB
PO7XAjofnt3abCLMOneqjRAge+Rn5pfZn9pbKYcMSzOgV6SMp4zDIj12SztOKVcoXgWQeS7a9HA9
NEL+ldZrhP/j4sAA1/dxeHOaehfj36jh/kKRx5GzbUKbnzfcF/HTEe78lmFIHKU1ixxYHmodli2Y
2+fPkyOzLpJE+yaucmrJKs2ivHmnzEd3zm44MgteKz71hEoD028WWl7Ase8mjbtKnXYYaItOj6CB
bTN6RSoiRcs6vHIX/B/rMT7WGjqU6Vf64agkvVkUxMn/HPDj6a/Yinm92ca+mGJolixRTgMTwv0u
Z6xZbRfwhVWNIUBIYFBrdTX0T/y31iDeo7TE7bSdRbvRkoyFnqysrerkUc5W3jD2N124RGhwsWQ1
iFND1ln4EUPHWzNpWBxVKx9hzBfgzD3JTn9weuTiMoB91+SpYTMG99tfpX+iUjkH/3/KhEoCw6+C
w5GdzYtuaapFQSFTOoI1L9typ3hAAshOsqAvFJnwxwuoreCJzsGcfpYkmtmv3aRMzyYGnzyadwpa
kk0kpNyEHabcrYm5tP5DKmtw5P9XN60VrZriJsmqY4N6W8C3Yr20bzwauB+XzhLEhjP/pnfXKQZI
nvj9Zv6fXP5iWyCtwT9KmXAXYcFelS7cUS7iEjwjPiGWCC+84dh7xR1bv9P8pICCgQUHmvTtNeEo
Y9d1F+DR3TlBttpEHezOTB0UJi6G6UzSYekCGh4PpQKZcVMXVUm32y2rfp3S7xiMlFVYbVzzNMJB
RkUnIjYgRULY4F4n0CmNy7YncvDHue8TIlSHbDI/WttCbuaCLcXhv9i9uXGz+1VNRrojxOPshU61
OzvFZGzPXLMciCo8xf+UzAVVcAhO6xKDYiVCHuA14u91XZbkWMUohoDMl9jBSbw2/P9aJK9PkW4D
gVDXpKgaC/VurwzY0MWCykPfafChlxmtZtmGkAiS7dVo7pIWnTeWfEhCUA+4YQLHb1bH6zs1C7H2
iMPn3GpZzi+htbiBorB43pTtICd3AKuKLOPUSgkic2a4rM3sGtn0uMER80Zz1b6ZjY8jZ6As5eET
iMbQVRM+Wc5FNVnuygkPe/39CB330oBGiEDQQYW40kbRBggFx3J0cxhtZqhcvGY2ZsdIfO4cK+UU
aIKUpmZoXFdfaxLcM3WsaMRGGUvzdG3hPr+Sk8r62gNTGnldxsCOJTQj5IMobAZ/Nl+kDcLm+x19
9jF4I21rAhNSKf1fN89pWSmnBr/gA4nov4L6gIyerUZt8BKnXrozRK4e21sl54/fWYvds8MEwAt6
1vSGWjY9UZY01I0VAm0VPNmkhrFQibkhUOHfWteRzJlmDc68/17A/Dg74KXBzIKJmxjjoBJwPKnT
E8Zc8kzvtg4WmrO73xAlN1nu5Q/QTw6cJSkj2EzFM1xiGFl/pXGOIT4apBGa9+r0tYOf+mhhqti9
PLMyMWEixAvvVCUGqGkNvUkumiA6A5Od4kDLNNFpyP0+DP4pmLrSqOmIzHYq+yyTB0D/i/1Tg+Dd
uk1z2qSFZ1fn1qrvriMDWI0vU6SEmhLbIglDoqWpu+SFiX1lC5n1PsWip4t+DfYy5mwlBUOdX7PM
fSh27kVqLsa6ezCM1EHSxkCUC17nBtD9tu6HDHaLXKeQZfmVAukCrXwn5R1KSdiPNxQjOAoivGKQ
qcqLmVccr6lQIHu0B3fbsj7gn+Rkxk3Ge6ecEnnqb8LP7og/WnFUtv/R4/ws4PtPjX/xPcPiKciD
drSTzaGmaqseIbNKCNTZlu6mEnRyS1QHyT3eAxDxpeyD4NZVdeVj59jqfks1E5+lYVhvqXJebqW6
y1qbzl+uJotXaPnGMDvv6zRNZnChmB9idsLQpHByGynXp+oCbihmdf+oklDL+HUjJyy+3beMH6kf
UR5rc34N7YC2zwyzzDMLC1xhDmmK4+6VwbxRbiLdXPsuizy8skStzTSKLmvsRiOMvBX4E+V/Z3An
VhEps0PLTIYpsaeU4RSGgbAA/NwcNRKXY08CijFbmsD/QhHfQ5NYRc6KFJ890+q09As4leleJg2J
n5G1s4S7HjhL5SM0+0jVWcuCaBzMYxmzBWXsj/Tz6MMGmB+Kq4+UFiaasZAgmgraaSfkerE83aJz
wLAsyvBKQvugmePAfIklvhz2tde+P++SiPvWVcmTo95eVYgiaMKRbwY2Of48NTbQ5QpGpK1kz3Wj
NW6dA4yExJWfEmMZpm03l35PL84ZSLXSUUROQQcv6jVlT/kpIvjEKcK8qyyxv/e7Ub1sBKcoLCmp
20uL7m0cW2hZu/tlgYdXMvvFWiX8/NFoIzuwRZ5GPGo09Xz3gEhHHyHxft1m188Nhd+00r630cUV
8S8pJS7Dkj7DlehmsePBpWrr3BaoHafMOhm7TScGOyXhW9s6gPnJValEBt5aQGJTX83EZGM7Scyl
h8aNi8AcvHLQp0cLHd+1RO4nL6WgyM89U8+4bMTYrN2N4Ilv2SezNSfR4oYygUEdteUIpK6G3pqB
v4KTKqNHoShOMvzZoo+MXqD8VCI+v53obRBuTVFYVGrYCyY4sD7hzzAV6wu97DNYXbi++AG+aXQ+
r1/v8JHmrSWdbnped9mZl/MFgeYJz3W3qAafpOj9thxN4lySK72dIgGCt4hoA1oYpTv5wrpa1UyF
d4D25n+a5II+6ph5Nwhf8Eo6FejQXCAeTLJx5zsGRrRNav4jfsG0yBV2LxQ3PnwGdh3Z/g0kfg2t
0Z2wzGP6SYHbOxlj4OZIW33abrQW050mUzahAjAHSemfFmWcD4waZ5kDlx/aSNDPRkDvkKw7FVt0
WeYgf/tPondjJanZySrmKTYA85hcFupqRCdbynN/AmAIBw1f3t6ktUL17bQcBXiQuvuYomfaRtpY
se1fbaytgWG65KQ+N0FFwOU/SPWNny0b1B/sD1edOJIqEnr6O4NLo7Aze9jSC+ayCPOf+DIlUtEm
j0P8Jg0CUNBbbgTYy2TInxzkw4E6e4aRVK9GevFjIV1IJ2867RTm6KKgLX6LseVqsVthdN4evOV4
qfs6c3Hq6cozhtzh2ZbfQjhIVDNavYOKyWPSUJTI9941y0ULY+m5Alw2l9VWUXXzIefvY2c7Qhzp
2TG1tspQVYpM3Nl0kPB3QfJfF9pI5ltxiV39ZGz8ac4SutxUTCcOhFUz+/ir2T4kdz/+vgWhvQBD
ocvabE6dZ7IrPjiv5v2sai5nHH1cjiy2usQ3LoXtQYEhMxEPWt+2gPkNMo4mVYEupY1RtV953xvy
X2FKdK4tvxi4OQo9wlW+uG4Dm83onxizSrnVIrlNJz9b/2p7YnlLaPmR8bY1MEcQSa31zypHQHRB
Ijk24AUGvW44U0QqBz9C+XYOMFAZHB4qmCTyhfE5SsszGghH/pKHa/y5xZNJUJ4lEQN4/fL4zs8O
pd/8IAhQT/F3fuMYIQrTERsYkvVG8Yr6pjnb+b77mq5107MNhAIx4504jgk8YLbHPAKfcoc6KTDn
2ekeRVrayYW549Xp9cfJ576yABVEJCBvuRxPEKkxdjFjoD+3q6bqNI9tML9UulqfBMkbBbSKGh9b
UhR4ACBErYvprBPABgaThbMuxuiTNkefLu3Nct+Qdc3gNjGN3YWxYQj5+ape61Uo3rBLvVOGP6CK
OhDworQSi6Mf4qZIw3eatAx5pr5Pl6SXUSB5DG0zwcRYVE4jfcd/4pTgjlN/D8eO78rlRvwlU/xK
G2NA/etjebgInOhtx32JcsT/o19gld9UgoNojzHmE+du4S+sXyYG8o97FAbvcB8+L/OU/J0aA5IQ
oDlIRezQMc/bpBQaOCTR/73dRV1KRkvknKGNCt9ByInGsXzLpbLS1JgzYkix5rSfGq0owmNVWOAh
rdqp5I/+GQ/Ryp5pbIQ4HpeUFeEzIcEIoyYmUHep8T+PXXnDqcmsbXV8913qB8ThWqJ9DdvL9FOk
Wf8puQjfPN/JS9yv1QzudCUdiORueayddSxK846uzCHokwFv6qhcR99sYEH9I2DIFJkqbkbk6KFg
6Yfslmc5++ISJOCshQPXehpk6HkoPTdFk8cDDzToH83FcUZi5duAJdLljPKK2KuRPwmvYpkTxYnU
VBukJCfZIJ61qi+o
`protect end_protected

