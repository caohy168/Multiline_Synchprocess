

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NS0UzMRfd15c96SOZUCS1fp6CRs8wjCMJONa5Nnv9aEx79OUbnyoXsYSo4CLFDR8jsi3YC4gTGTd
MyvJDWUn1Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hZnsHcJwARteBAJ9FOgdrtMNGawTGbjcJtHea5OVEQLpN/1E3UZeJQvMM5mnBKjJlNnIIddV8i9M
joJgNubZ4x/J+5MH3hTdxxm7F4LSVBkzCDCdKpy8cg6sRALdJlGCLBd5W3fL/N1Vm2mvnpWYOTAK
o/bvQTpb6ITD77LnrhY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R5vX6KxpkN/slhDNucavw1UjzKwMJVO51VdByoN947hhTDMG4hIQ816kJsxI8/j9YOe47a6kVgQX
KY5bGd+cKmc7Sj/0vw0+AaRUi0BUjWSzIKXTRnPH+tW2WtD0kJSh+7VgTuQBcqSoKv4d1hTuP5JL
M95KyED97q8kA8W6/tEFUdFDODI3RK1AjVcoiYvmLp1JHE6N+4xV9DMw8xy7xHVPnxKUVydXS9ZI
5Kpm5nLDhGrx0aFmATRDTNL/Iz8QjDkpAArYSnHBguJuoeYzuJ0J1ZlDWpswin87gylwAFb44HxZ
nqHKf/UUdwFz42xC+ufZ21dbt3dIGLJZuW/J3Q==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kkium7vGgI4mIKVYu5AQtLq7e+Mob05Zqln0+g6ZaWnlPFJRayAUb2TGgpLHS5PtaVScG6fp7jAK
hR3jUq/6kPviQVKWL2u/4LhcA4kKyI9Zdi+ehWy6Tnh028+egFThp5uoINPpEng8RwwI+6IV9naC
FSuUifTc2tuuLl762gUP/eM/n8VGC0/A2mW/JvUel9ur+8u3BftctCYCVxa4bDpRr5qOXJGA4o6c
E4X6LDHXzpiVoyMS5t2r3OL/9fPqkK0nufzJdd4SZTXUqjb/RszVSlGWdW+08kPsxUY8m1oqS2K5
TalFYT3jg5Mp+kYfDfW3qlQmAC3mJl2SAKU53g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CkQIlfatrQuDsmTnRTe2/gzxK2zxoe5Evnu6XsZZXur5sC8gZMQaMz//gFgUkCSJi6IZG2S72YwZ
/DWOIKI3TWXxND32Nx/hdK6B+9GNQNAe73NLPLq84cJZY++JigrKxnm4um/tNdK3g7KtL3maNF+M
YJxE5p+FssMep7I1eFA=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EmZX2JV5yuh7StMKg1MKBA95BI+QbntliTbj9Ha7iFw6mcWRe5/6CGQ4XD+IIBUvXHSt9N3dYoIo
PmKyvOD4ATYMfvlrtSTiU0NkY1vMMBoIgaVMYc4MWiOOqkLX5QCr1y4tP/2tYFT0XqOadBl7mSkX
zlFIafpoH/LOglrVSIoDeBEC6MfVsaj2w++XvX1XfB4Q+0amZMXDTJWJMAh/IXT47EhyGLO/yis9
ZfieIq6d9JNguG3rVoKcxXkthdipGLh78LhCJkQ8FEwwGSvTbhQ4zgHstrRwdAASUDa6gwXxPpIJ
qqbHLfsfv3nb3kTfiGn3wbY3N0IOKggKgCcBWg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AboF/gdXw5XFu8Y69yIdoJn8uAobuhjjThXr2RSoL7EztRuvDZOCvet+2p1rluDW2+roz8+34B1T
nJYCZlru6Io6ivyh9RLqrWtjUfgNAh5bdGa3criaFYVKBbO5WYESngDLA4l1SKsY/ml7jdn559js
3PXOVkZ5okByUMAkBY9xgMS74kRNZbbWOs56xv4nvKv9udRIBNg9MIWZs33CMGZ6na7v3KN5Epq2
xwDAxNEyc/aoA5g51oYouiXbJQ1Nb2HoUlG1XOtMFCdrUfxuR2W3ymUPchBgVYx0ewk6YjTKjYY0
kbo74o6VcLrA4RehB/+i6DYbsVtsYPvY8u+VhA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cHkeoE7Sw1d0LekbvMrcrlfDu0GfJ9HoUw8fLhpsruaH0GbjCq3dlMBTPam2ODYxDCkoL5KkHnCy
Flu1mhCehzsjfkPpA1Bys07dlEsLcToR1mbANOUTbGzOUIoxpQY/N59lhLSnhvL4bqEb4ULGmsMg
tL3bvdV1qKnitWWmXgHqMeP3UEX52+2ODqtxSE+9LvBE/H0u+tpADs1/2g0UDOWfjx6qgqWpxcE1
nIcDsMEzJaatCD0P8lIqpMMXPTupi6XX6Jd8cXWliFXKHXevMkzZ66K/E5YBzCuv6OKuPSXVAjmf
wZJsjo1WqZ3g1O7+v5Eqc+ekE52N3vpm+ZqqMQ==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z7DnkfqlpbYa10n4bpu9gzVCQdqPQvlWpZyyy52R1KXRRDMK3xAnodeq9EtR6ZOsmm5PN9SkQqQO
l/gjwQOcIVAi4fVzDz8+IKXpDCqkqUS9w/NOg/0X3cTIKaih76PLBtiilbrPCaQggu4V92QkzQZZ
Yi+k/NGNjn8AoxTCOPlc8dFEeQxWTPkno4pRRRAxB6EQGemCa3RxC7USFhUJwDWozHilTW9mQ1sU
Vbuqq0D8vs8lzgHCrzvSriyzzI7Ar30bNUJ6xjfWiDaBEkoY4lQuo15QVyvXbvhwZNz9EXXXNec9
GB7pUSwj/cmVIDuz7ortZFaKgl4hP9NzontE1g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71392)
`protect data_block
jeiOGRQBB3A6ltKHiJxa7ONI1JT6/6g32pnuoRjiCh3hI3hzpkn393TMWrK+JzWDdKw6keEvUbXN
geI6Dvoy+B9pPIvYX39CBzKGkYHht3xVmFk5qI/vWmjkTpjCeT/eLd7+7JcpEz7Ar+iFojKEbbKs
Td0Ch9PwuZ/4Zpim1YnOMZIvP8ckx9q21uSHE5rLfNH6cqQIdmbCbFPGWNTPpUwNkDaAwuyfY0WV
/isZIpBRKyxQbMuKncjM6jmx+n4xnQ8MqJXysS7TIOWZYyLZiZFP11oo3WwNj7jHaA8dIvbK5Q1l
B7oTaeq0nX+a3KminWTlExtLYyZTw/GILfjqnFFnRpvyPhdS8YkZ4qhu9aRhXhNZN2b4OfWa9nFH
GjFDUtKm+nEtYEAMsCC+2I9fh9SFJ1qQcFFiTLRKGuDpsZvP1bNP8hR1RASOQO6FGWa5IjrS8zzB
/gnBGAhI9kZrMBUJeHY2vB0swWhvLXCqoI8ouixO+qMRCcWkJxazGoLb94mMHREFYP724Rwdapw9
myXgIsmZxTkultygFUaKPNX1nSWar0z8zz1Ttcpn/+gek2fobn7rJn8y9ugcDDgGtpr8mF8tvz61
QQFQcMtXaVUyHhYsxVlIEFyYQfbdkvWrvKHKZYqLeYY5ptbxZDwL1rYiQMPb5j3gHGmrTPSGDrcv
OIzd6Yv983/pL7d0Y2Oe4DVd5/Id73nmfc/t9gTHLmVmqZh2o9qsN+3h/EGg8c4RtzzYHBRl/mLn
IlAf7EYb6JQ32GO+BhrMor/xdI/KM9rMiYWanKriUEp/oCi1bFwEcet/aLfUsYes7UV+hoAMe1f8
I/o0nxmLYkVrebr+bmiGMxrVpISRE6lwhPYc/hybINLMI3myxmT/ycOfDDJTXdTjh72ivzMJR6ea
wttbpg59yEe+/4GD+i5elUQ3z5FUnmdyoeMytQDG6LW3hKekcOa5uvQQ/Si7kaXndmBrcxEESZkX
E6fLJUvYtSy3mBt2zYmZZSxwsw8eTvO2PCILY0sjQUnoT3xYAB3OHM0Wwo81JJ32PKE1lEJcsoAb
CNUcmNI2jFVuKPN8xKlwadJtkpiwRCCNX0a1gknzuxIlLfy8YV84Te6jiQ81ze9HOUU6KetovcVv
lo/xX3VNF1u9+vzwe/mV2CIZy3NfmpgYBvtpFJUWKGE+mSfS7v3GkuAR6QbDr7EIvzRRwtriG2ZE
CO17iOnffLiyIrPqOtSPliHcxot7XGVgynaeXGDILHYSnmzEsMx6Kb/VNuNLq+9dL/uXRzjZAwO2
2xStL70HIwQsGM7AXg8W7QZJuQXQIbgqUYAjhXU80rLf24cGcB+aTU2sDaA26CDlZksnk1SnUluX
gluGzCR2SHKznfg5sIG3H7uOtI2wvTfl2n/7PNhc1WBlamY9RESruO5cDoumtDlcrIUW9mAqPRkZ
AMh7oNk83mqHFDDOykW6ccYK0Ng+zY9bFBqXDXyBtKTjW+cHZ0HlOUHHMqkQwGUX6OQ+InipEOLI
LG1LGc54l+tziVYdSrAQsL2rcGzmp4ooNjTOrB8Wm8+PowPOUcEmu4dpWwE6Ju9z5S8thMb3L5hq
cdzKRAKV7bH4CpOylZf2LhfaXkono+PMz8l6WIzZLMtugsZfxSTDxTfHd/pQEcRvsxmWPBNfUbgT
PRGD3/sCHCOOuW3ep09CB6Wria7auTQquCCxufw6Z5GoP1qzlQ7F2ZrLwBt+qS5x+z9i2z1BYs6i
NUTagwBJJOykgCbiPyh9veXbtzCFWBlp5McOpAcbAZqLIKwLT1Z5OvYV/S11TXiO9qfZQJOgdtrL
riEhhcmqll+u9XsNrvzOWEUcGDgjNO1j2L3Hd9czm/4EIwJX8oMgvk9iA9TTGxbyiAjUQvkGCzU/
f/MrUfe1CX8azV3rRjFn42dM/coARe1azmtVcCFAKllU7mJOr64ok2fvEkOYDQQ132gCAS0rQCUN
hogYJorjAGiUCl73UAqTP0Zt9dA+q0CgoBYH5bPXuO77MZEGg5+2F/xO/wgGB9emqT0LIrZv+p7z
nLWVov031evzLSuJ2ogtNCt72oZtQB50/Ca2nU/F00Yi3RHcdSNi8oViTsgehWVT8dsPl0Jl5Hzz
lolzfpbJkf2zmsSkb3D4rMTv9CI3qvL3+Fk+p0N758LnFyevKpXjSOZo6xJ0HhEArx+bR5QTq1EL
OUYBI6tHxr7fMfk3ztVOh/i4Qx27QJfMBYVzX+C+gckcqHlmSGh/UoNVtF7ZoEpM5pg0deHTxcJl
GZ+Dv1FQFxk3l+bA/0OFeojz4ZhESQ6NQsRW8/H4JFvoNpOvR1kixeXOnx7oHXdRu/O0bx1bcuN0
8jmno/W4jerBTLBz5vLRDvZoquIqfo6R5GhchMUNLo7y8iJ58N13qk6ty/iUwyRoCAaD8gyf3LP3
CQjuCdZ+FEBCmRoN99VPEoAIHUK6WCYr7IynNqFwm9uW++Y7kgv2t12hb+uLyLs02W6anUb9vSdj
F7c+WDwx+k413Vc205bPMLpZGgMWK9WOcV1x9GfQuZ0EM4s0/6nx1qLn3xtMRP5n9FcTsy/A2Iwj
HNrYY+ZmTLYRfaK/KttjGaLJIxf/DipTy+6hoUwjhVFbYVtbfBMYe3/xVqI8YU1vuGyANxnDOiOO
1p/e1OgLdljyvO1LgGrBjVWM8Rg2TYfpZawM9DbAS3UqmeN884nlPqtIyUVU44sPeovOtyP7k1BC
MBIQnUEE66of4V6bkzlbewepNeRHs7Qz3hBbSTlC6r4eY/+FNmjMqRHvOiFt8nQKz4AlDCtaAAQ9
o1SiBpI0Lp/HbaOV4OHQR8W6LlLWiuLZhwNtq/d7aneGWK6OaYk0TzuPwslJQJYv7U1ILG+BJPvS
yk2rU4HnBSDQX2HjUJTSKIhThZi+OaOnuU4Atylopxgx13nmJTqS1ekiP5W+SkSIZJj1TNbdV3i1
kWVWySwuCazfWSNOrGGPmMEt9n9NRRTGn5Y5VQjmRRruJHW0dvt7OWO2sw9J6WDhTZN+kNTOw9Kl
UYQ7zc+iw9UzkxAo8uUJVcNvEkYiM2ZAwQXexDIPntaafdYXIwD53e2s3qFzVCrI95CLQPty895w
R/hXYFhuixFr8SddRb19vUJ6KgnxhUYc6/F56nzI5+AaQ6NSdxrCci0UW7eeLfnoQEKz21Hwf/mf
CvNRUsEXZUZhEzNQfAKsKDJ1VYQrkvKwShRXXKV3PxwxOf9+AxvWHnCgtQL6tNaT5iplGVUhr3jr
yi5zKU92l017FZbSfugo08RiLX435eZuG74M2v4YwUyVPenbSAv4CbMmBRl+cW4reZzAM3OuwOjD
zy/3J3sZODeAkD81F0xj5D4MRBVI314qAdR5kbQm2IcHqgG4SYt6/Wk+THlyyRF8AJp6AqF/54QU
ZbePrD3wTi/WSHRIaoLKKiZdJ400WnaFfTcQLEbCY24/JjatHmq/aXN+OTTvPv950aLFT+EfwJ9D
uGJJnT+faqKh/QK+Jznzez8WM5qPp/mOrRhyffJX/Dh8Up0M+1H6/ywtqZdq7pppYgYqZRLEcxAI
RJcFKLQq2HyPIfyTb2u3I9aEmG9lg4nhxpWGythkMgOCNCkBn2j4lC13UqBaUnmPzI4r866VBnkk
NZG7PNF0r4NolizDQ6qDRdgFoEZLwE7jvAVwS3cTjMWoXZDBQA3aoKtuF6kIEa5X6XbgCxQeFcFM
oINv3++qn6kNExs5/TgXHfQqKp5QWwL73cv/QG8Jh10hBKwmgFYCiVbuluXp59ZNzcFx8PjEwxDC
ET78v+iXP3QkYOeyepE3AqZeAFwOaBIZtzG7CXeNUMieN4532N+j4hBLSOT2sT+rsC9d6NiUrLvO
t4wXtKcyz4a4KDTQNL5RlFsKplxqYXKgrg5tCDrCa7CLg+8MHJVZJRcMYRIeQukjuERKU02NhKuV
sTbx8u7GmkcHdmFsc0wBACHxWrpnuAwDeR/zQmcFTIvWQo7O2wPrKj0RmYBt5OiZewpP0h9vvNEl
f3UW6PKiWSu8ekt7SAFgIbj1plXEQdw3Of2e6XTlaBbnFsZQ8OneJM7LuhrAicbTcYqGJlBw+bNH
beu/POHBe/hLeTHj3o3Jb5yoDeffitU53QTXFJiKQWyb2Rgmz/KzfAa/vf5FO626VuUpRK/lTx0L
+H0aBbNl88iN8s8B3nClnQWBY27NaodKiH+7D5diEb63XKddvQYsXGA/tBthFa30WJRXoPqRezPD
zvX+TuAb1XIcmBHqafLBfTKbSA6861ZS1MT1sUC2nx9VUGHH+40xkf/bbHVfLoo43R2nKb/LepIi
KKUh9GXaCmRfxvn3KthTcuWc8R68n745m71sBhCMt7AgRxylEAkfhUyNRE5xu5cjyGUnN/D0RQmk
I1P+PlTgrp4iTafQQAkeZLT9X/8MGjSMCVtHNBhyC2HqLvMUdlFoUedBb1V0lAaZbOd3IkSJl4EH
3c/QPkxDfMYNDqxkg5AxiO+2jjWcqrhrzf2PHYrAZorkfTwIL+qgzNd6SfS7I8bQUrpjKDGJikuA
d0Kc+P/get+M4dsSMBhud/H6qHg9xo3QwZ5gx4B3mgIwEx+bQNfjiwacEII7JFP7ZLcSEBp8UwuW
eYpMtvNVJFsUsbreGs9g9fANmf9nSZ+9jcG9b95dLLREQwoBAAZLjSodSjjnWaGunNh8v4ikDQPL
SFFrY9fTSYZBbUC3nXgaiYFCWASrmpfBG8D88hcry2DzVBRcGGLiWZMqgMV/W5oBcTSfN6ajMtyt
mwK5hJtL7AMtvCZRyrF1LksovdFm1n03FPwOF0UwO4A1VcUoW7ez9jpx87V0hkRz5AXuOzwBxvWq
RdCgGG/NX/OWYp2VKG9u2kWqcr7J+2EOOaRB2vUk1aLEyBcud3tIE3/P/en6AXKyxNEIUi3zsqkR
G7vsqSTClY493GX2c22x5VKYWpSbLoiFH3ow75Af5S3s6UwLeriNMJcuKJoKTObHlWC08H5X25MI
uz/ZKWc4snU4ohBioigihbtfldg/qv/d80XV1wSv4H33RMRBW/AEH8PxyoylRqhRUasAtiWbBEAl
74b2TryMTfE1Yp6mlzqx1zG8HtC5WQpDHady0pQDzmwOu+PladnrCZ2Rq0RFR9Ownw0nCqMWN5H3
jkKmaBinW1dWORyx9NIMkfOq4uQevXJKTg7RqObJokQIKTeTRegYVKtPwOMuIUwBvaIs2s2GF8Hu
ZvE/I19T4fKq7SQmgOiZKHGPWYUisyWFm1cIEubYGfygV441ag4zs0xoeFlCvmndhY3rQfTd60MR
Z9HVjwP1iHRwQMSI5zCvg2hhGt33fWuDRimTng8K6VLMAGz2bRL2hD6QDL6GwTvMvRdDNEQKMty1
u67rUMa9yWrWvPCY8rurFXC0CzqcFYL7aXdQfAHu+Lc9sU1KEISgSZZQirSla8H98ML1lB24Izuw
iQXFlOq9B5Rr9cgqLUaBSbnxrBFXgd/yhNB/riSLqvxVGqqASLn+yxkcJEdQ/OOPbSK8+dF7HdgV
U9o4faR1CpyY05Fbcb3H0g+Oq1Bffxzw040odjS9e5ZcvZb24xIIgC3p25cHkzr8su4oOW5bFHO/
dc92F6WB9cP3nIaWKwC2ZFccPNEIHLiXP4bEcDH/XO0Aj1W1GjZpouaP1R8r76f+SRguavnzySjr
SYbX5VFKiS39NwGiSoYcPzIq21UhJqyphi7FQISwH0+5iSJggdliEb3PuMjN0dy7TtI21a5s6Mo9
dxST1+CsdJYInZBbWtJw5NP5xCNWhNnR9bYDNKX6bLqxFMgbofdpRyW7Qwn3Oex2lLMlJcmjT9Wk
iupIRVa24NEJkTUf02FFiODnXhp6+off0KeXWtfKhcIMbNTK69c6K9XCsxy/9SbH50Ew4QhLoflv
6Izx7hB8hyaVNwH1CXY4CWFZR3IF9Wy3EjkhymbmTzLa39S7lw4x9QCnfmZ4BFVM2IBBRMPHSa3R
cVaMqpamoUZdkfFqsEOe7dSKkTZOappJWDZ3uITjlYbo39eTTPYASXbcpm7xWJ6RA3q4apytmqZD
7nY8pS97MXqOME7R7vqOAKgWrnckn4w0z4w6DlKkAPbBaQ55Tcjjziy5YtbBcH5aT2xRN4oSmBIy
AtRHdl+SeixI4TyqgvuT01tBAGlGBErzI5L8d5t6wHIlrI2BqvTp0IFqA5sKsyasC3j2vKpLnjMK
qPZ5jEZWg9R+jCJOCCUWg4jclzriYfy1QbuKh/vsqxfVJwSvi6Ck7u/dX492TjTeytRibGxYLVe3
R4rtfJ181RZpwQ0Q9guw9BjocxA1uYNNzHX1P/9Ad8Idg/KBeXhVuRpn6EVLdE6m0IvcOorN4JA7
osuWjogOZgP//7c2gEH9gFaUIurIt28sbEfyWOLMigH9InhnTSsgsq6+5T6Fl4874K1Iq9LJE4EQ
diJ9tutz82uA/Dgf9Cg9QG60MG72CAIZQa2uE9vKQL8UbJ58IroDX/tmv0dKzOmxsjEETEN1Wue3
ZhwDBjF+vKi8tmUaMWN6U/u7Qk+yVw4caSnM+nX2Be3ln7qnBrA0TgYSouotbN1BQKc9sExdplSt
FitcJzIU1G4lRFLIXEMyhOyNXUMi2EHHFwEaOhdMmVQuBsU1hjMSuqPrYfsWZtN4GDbKVBqsKNk7
37QFXYYvn/J5X1CpoVMWVojYbs1MTYEmo6gW/7jtxd9WMNHGd9rAv+IfLFdZFnB5wWHdF0G2bUV0
yw3bBcfcZNJ7k3m2vLpn89QYFEFvJs0T6SCm4twyze946yRZnjQNluaQMKdpNWAvZdE3TGFCHml/
7UIDlHrFAjZp6E4je+kMEeeVLfnRFoFLZgrnu2dhgNlicg+MfdIMmCeo9p2aBXz2QIh8pF57OVhx
XLqpZq9i6wwAXCLd6NiaVRQMZBtiFCpXXspEbi85GkyA0O3/K7E2qDTzg+WEaU9oH0pBL+YXvEE8
m6M8wUdo+y4VEqS3qutk7GcVo0qGSRJ6L2Ai100QKAOlv1qkz5we3mywKWVmtCZebhC11P7JB0Ch
SPyHqBaZdKbhOvy69qubmYGLefhDglQJiXDUE+3f4uLAgTYw0xKgPcf8WvFPMni4rGdI5jGvdrYa
/oggoe1hNXd+8exwY0YmoKDmNKNZ27c3cd9RY3Y1lXXot0k5IQku/BoFlP189JfbtNChJlaXNDnZ
+5aHDM97w7rHrBaAUKo8qOol2Dmr0gv/DaTx9GwTEtstRnXx3LaPe+c/ZSIto9AuROwZsOib3xQV
OuYz3pOasrgSa/SjOKPskj+tNlGyd6NphRRlOwHmPwtyZ4GG2wHn4pI1vgaJjog87h7lkou5i0gw
eCZGJsCfEEasHNNDptUuI9/6MZ7J9uqZ8OzvEj+Ntdv53FD9ofRB5TveLZmPK1fh5107f4uKH7AO
Zthy19xLrsjFkSRREhPLLldUwahiJARmqf196qtxN1bcrwN8wU8aiKtb4Bpy3fBz4bKCL+sQkB70
GurSceseOj36It8qlj3qKFGE22pXPQUrMmh8Bvf2s1Vj2s5SDQyrbRub+zXA4216dfndh70OlkB6
MZ8Zh4lMNyP7fgj4bSzCbskpfjqadFLZqSrFztgHdLJ4PpARH8/JjRMfUFIXgY3dAMksKZ+WUiNF
/IPTlx4hgL0ihtnwPX7ztTtt61GB/BENih46lLSuBYjO2EulbZ/sXsDKzQHNBYX/+PHlSkXamPYx
34j4O9DMEbkCWe1IjhvVHDYjX6sF6/bZnpv7fnWL3eEW2tTjaGIVRZHpIdkaAZVma9rJ8jqm8KZu
q6jP76eOYTra87Ja3PBscnqsg8SU1/U0wmYLx76PvAmN6xEKOPA7ineVTPd4j4rDCqUtxgDraK1C
CuVKx42p6p4oDigjChqlwXnYR7WDIhlpxbSecNbTcA9TaIny7n7gueYSYaIh4sjdIiviilXi4f8n
EW3njJr++HcTFskKy3yIdr+60WuL5zbhlz7FcAmA/ak8uDrchNht4ryOB6HJ481wGwb+MC/t/ArR
SLDc/2aHHWStpaZgz4yT1dgoKjgK5/bTjNgjBlVvF2EKtjmBLzI/v9v0A3/quuTMOHhLHE/t3EZL
3D91HdoBjBIcM5GFzVdk3C+UJoGYYAG1LEGeRCxC5R5Ezg9eoSI2L3lpxASbSziNMcytqncr71NS
rsbUfrkUevssstYyXs2a90aIFVd2p7HfpgugRcxvaYzRUg8pQM4OlqhfHApTemM9H3WbNY5NsQ94
wGiiyF41+BFxUMgLRFONEApGrY7pDO+qw5zZfn3S6o0GLPnKJ/AcMPum0uSLyRPLn2JtQbLn5Cub
imnBLjtqtKnLFUbpVe1i029QNX84dwr4tmj54cYS5S3DgG8ZU/sMo46j9p+Q2neNCWFBNluh4Qd4
PiUGuLAgzGW+MElXFGgK2QXb35JBhi+sJNZu5W10xRnXPUMmTl/bjSvu75aqktsSl20a9A3iG8VB
jlO49t2Nit5xWpJY4IR9zPqFnSyIXIiVZjL+cu3b+ocWa2XrQ9GoOWmYU1Sb14X5za1OUWJ+wiSz
/ITwjCTr3GKSppYMwQSi8k8QdNNGQ+norimcnXYYINdDrvZmT4PXsoEB1WbUL5F2yEFL5b92Jrbc
1+8yELd+dTesWiEOcWpDkwu6adZYogCbwI4APRFrzXYCJZJkEEjVu5bYaJuFjIVc0+kBJuSj9zF/
nYLvlQIBjKRrwttHxn/PMSV0LVQHUn/z2+bxUpeBStA3DeEl1e7rDEv776uBAz5YgjYxmQym6jPj
BGKQt3imLXoldIo2PYMhdakm82DscXH538hNpVZT8I/o2vaQtUFtcJQoHdEg0MDFZL9GJRw+hEqm
YOTWwcp+foyPU9edMpgEkDRKf4WxReGEFOKqaBsGynrMvx1GKRSQapvC/DFqo66jVJ/MZboguY4z
aMUuZ4HKqsFa9qoUiPNY9r4tdEuCNxuPyPE/+XXwaKahov8kvZ5WWRvP0nw7+T20gNqF9ITBdN7T
Md9o60rzfwrWPsD2AqY+dh5FnB0MxHoKrIbA3B4qDudU960iR2IBcqldbJRFGf3b/FEU0Wg2PXTd
dlb/LGj5cGC+YorpVriH/VGhPh166YLmgNShzPSdFcm+C4ooTePOY8/h5PwjSMQlHLc+9RFhkXfi
KftHZ1A0/Z93+9TAz/SQIB0TPcWBwOdgCXKE77zKhMLUO1X5xucAbf+xrdpWfotWiDKrDFGo6rmq
aXlcZyDfxph6C9VdaGxAe7HtSgM3fo+6IC1KLfKTgDW+xaRBYH2taoWwXkm2hoEwdCotbeDi8Ajp
CYa3AXVlFIp+dT8DFV84le6gyz6YY7+uKOrfRCzM/N44suqq9KYqFhjoRyxV7cYAqjapvQRhb5rQ
er7zMBnd7xjHN//lVChf3HkvytCRPeADYQw7/5FpJOYoWiks2f5ghIZbuPybj2X9h5LYfXWV2MMo
O2mhgKRpuspTk/A5ys7R2lOOva3Hns6jBEosxLVqxYuV+T8kMoUgne8wS2CiQAPUtF4p5Ajg4mzS
Zhb+Do7ZAao333PczqAxwV/+i6QyuJAAQro3eOj4yM6ZUGh2lx9Rz92f3Q+b+0uO59CYM1dPgQab
mSMTvvR30KaTYW/oh2uEu6nmtc830hSFrkBY1+m8I6XodDrfkN2hf6iu1BZb8+7cEQplSEwuVSSd
xSxUhfqmrv+igSl2M0T2ZrIaxpokXoBuDLJ520wXEYtNINA2/mNqGtKUnREKv/PQ6N+tAJKRyp4G
zqR4UJ8yYMvjisoAXhLwaK1vKMAlecf41DLdkcJOp3yVNKTIO++rs6J3+gTtpR2mVQKD3u7v9hFP
jMAxoGQ0W4FiZP/FvRz9RdOaIyt3I70l53lEoxCksChZRFHEbnyaNljz0dzoKDeZpkIOY5/VQTyY
z17hbsci996/lnVId8CQUHrRwJmNMjyjNeD2l+d+9z/Gi0uCg+LhTUKbFFtbipof7/vS6htBy35a
3nfduRdpgk1oyJbh4QMoHi+ohrpLjq5RM5ramXOIXTpjwYVPTpJDS1SiF4jsLN8vGtrmNqYTkFIA
ycRE1DSXLtJmH5NOuo6ekSJSxLL50rk1MK7jrnvaMw13PEnRD1aJD1hwjr4Xp4v9wvuK+EGOin2Q
zOQqV73wf22A5K+GDq4QJ4JBMsuFK7yaoxmNK4C6en8rCYPPCnjXT/fIS3vZ0IMzGx6p7StUqlo7
nYZJE0Qwh7D29n69seVyyWgmGnd96Py4Slb/VqIs/JTThL1pyHz9R31kqnA7IW9qw099TICECibl
LdO7FQdWY3R53EtINWsZORzqh2MXZCiyqhYq/kMto0wLy5tGjH5N+AfuyYBBS0Rxtk1fOLLwtMcB
gnANfwA+6Qi4ylJ4VYySs4OIm+4PUBnlgSEUka/44hueGB/mYu0e8YfPA3ZfiEvhr+tpcneaLbYP
bZ30/gyBDJyRm5tfr+XSUJsw0lWik1ldAQWWGH5NU33+jlxuA+8wp3V5iL9I/Xkp+tEcuVYomdeU
8FDfnUlzf6oUdczYFhSlBC0CL6t9b7Q+jEbJhUCWbGLEP91oc6dkUf0P/t3cgHRZ4oN7wpQOfr9t
UQkh00Komp69p2mavowrvj99pwyKWi47bqQaEXb5RLSHLX7JPforfcD5knAAXLBrLiEugC5I9YOU
Iw6kIbmaJydvID8AEByg7FOTKoueC5MZSBl6Fli7uMuPk82ACJty4VdEQkrF5t3Q+jicgG1lSC1Q
HxYFjjb64XaYhMk85yp+jFAY3IG40TOlFYm2lE//cNrId77f/lsPND9tu1tku6+mPh3XRETqCwJi
JDM8nis8sTP7eEc11KuAc/U4S0+0fr0u26RKy0hDfD2jPOEs39a3qL2pw6/jGwY6b4xP/cTLGkoF
52OofC26fOlPT/Hvt5yLimCCwW46zv3k3z7ZhATXm+UtDDDW4byjn9iSyahPNSQgojFjr2G1OXCf
mwtuO1Q1fz27BMJgZXrBVUGQiZCxZ+bH7kaLk85i+3DlMEARofNauNMUrw5t4TKIR+ZoOQK6eeYV
zSUcsqPDe8IXN7KI+xd9QhnUbtN+hG5f48FE0in8rNT9QDEwobx2btviba9Yb2XCHqM8yhsqHDyN
ZM4OKMTbZif0H2zocf6zRHNd/cdLMtTOugS8iyMU4wO5JuB5b6mExbwgFI5wfVBGd+oVYG/tvrJ4
r06udMMxuaxMfIaFwma46JdFFXZw01HsFf2WqoZ9J94Q4R2JU9cOPCHj7XZXaO2j2vJB56dcBpdY
RXUwy6dEjXsrlEtAXivKpMbJU+w/QtaAMsnSgzavaHRX9t/zj2rRwVHVj4Lj5PpAJbsqGl31lSSJ
NCT5fBCr1Q9X+xFQX5xvuy63sG2qJ67XMWpHVFJZl/K/cWrG0L8YThR3btuXH7vPZXqsl3Y+2Aou
An3INhW9eTTtBbckuSlAVhWOmByTyvU+jcTWCqd6bvisr77u4ZkDTh3LSgpqOoZ6UatbHo3BCaVH
8/N6hsUNPYThdsGg+ha+KPyY5pylQSPL7WS8//C899i1bsw8JssUhZmMn2fVCGCVIdjnEXXvpe73
lQ5tY3TIuxz82Y1RbRrNDszFUD11Dv0iBcFWlkl87seQe+CYljTGhLtuly5CkfBx5YXHTN+FJptc
4wGqnHv7O9W1dfCX3ecl2pym6/5Q4cfSTrXXHDlBFdlwyk4G7fBFDw4nDJTiMVweiIJgAzRYvZ5R
ZWXSEHgGDU5PCBxY6KuoYAd/+RxFWPN7wsK6/WI6R6ITYPQHx3n4b0z7sDWJq8u3w1q6slhpv/Tt
8xfLoioX9RM64oYf7jArNFfUpzvv1zgrFEGthGeuz9QRJ+JFowWXgeD/8ag3N3Aa/HkeKGYZpWPY
ilhmkuWEqBkZqzFWhQydlwjiNiWDWSd86qRMyLWNQ/RyUYdDpmaRPPh0zrBmrJ9vLVbp6j/nJ1eI
2PYBYFw42spjoHlMMJLHwR41AlBQawxwBorm5ZuWKaxNm7VmFRP+GfheobgEjkWpmsfAmvOVZ9qG
M9uaHnAF6UY49ix9qys1LGEq5x2QjuUDE8ZMJuHh7tNO4muni6hgKoNoM8zgs4txf9hBk7+t3S13
bPs6Y+TGg8uYnpSrod0AVwQtA9F1ZzWTz5VMn9OGHSA9DM63th0arOWdcwba1zMzprh9J3MWnRQx
sisc8EXPTGFF4g8GOmEXcXEuxglW5qt7LY2t3Tuvvm9t1AVZcKzvBvskCSsdtgzEYztvrCSvVMee
9roPaVhCQ373LzgCRgBuXmGrXpk8XMH3wV4z10g5k9iC52mRGM2zemgNuGb+XmQP+aM11AM2YxGr
cyUlGv6ZYCuMqdVuF/8MOxPpcdnswHa43L4X/vh/qarEYjRby7e7FNFudwEKwKDs9L+R9OB6WfOl
WlaQroVI+L9gFQrWE2ZGur/71tO847tNxUcbWrE2kp54Bp9l7wI43NviEXgT7YfXEOV4ROeJ/TL2
6twawjhEWxMh2TxJLiOga+8oS5eWGJ01FnLMqdXK+3o6gZNs+Pv0iM9YtWSPmcqFI36qjUXVL0Jq
IrbjYzV8UjI8wNbHNSixFrAmNqC8ZEefFdKE1oCyfgsULb0Cm7HiQp0Q0mEHOjvURg8QUZd6qCyO
6mBKBUfojRtzaY2p/bcMGiHcYfSDdg1+B/CljeX1PXypPfSdvDp5McFjrNo89kE8pNUkJl23seFL
atGh4VJFKe7pGggAjrkf4iYIdvHnP2Vwos5UDIrrxAwDCkhhp/ysczMMHwZL/8Anem4IE3zmafgl
Lb7K5MCCYydIq6zMDdiY9LM/A2fi80ci1j38cSytE2igbvSsUlgGjHTZOlZ+8vo6i/7qRiABMdta
dV1i7ueEUMEqIQhI97gFLxcCb4aM+tPRAaNlxTgsjnEiq9xIrJri4QW/oYEKXzBEgP9Ip0mcmSqj
mjCH5cYy4lCUJNErvBk7zZ8tDXJaH1xLB1HUbq/Twk+Q9XzBo6zEgVjADdfwnCC07ingAfBNX/Fz
03ex/o8ykhEz0E1EbYZB4nTE8s2+JNd5BjIv6uHntiRFoNiQHYBXKT6qeFP75sMOqph36aX8K9QR
Z2gdn5v9i7uffqIDYfhadAJJLBTNWR0paZDBIWztItaGx65klCB1xAYFdyCLfYcg0bO1DFt7RWYo
H6LTM9dYETC1Gdg+3jvL/UxECGelsVJgEbd9fxDw1g4L4c0QmSudaSUcD9y5KnG9wJNZLpnFChlZ
vlLDWPSDZBHMj87sVBVs3tfQlKaSGsDwkGAeIbVvJeMkfR/bV32LL7A98LyDVR00ZE6sOOknGH7o
NADQFgtwR/N3q7mHS8DDJNfHgkdZRYjWYJT3akYcFBcSj6qSXy6OWbluubKIdYpfjx3m4D4+1yIw
+MOWgpEUGR696CmpSODzUlpqWS1kDllKtbUpx0xi5ZpID5TcGuXAiAp6ZDTDaE2vZb8D/vfkdRdG
B3resHY/NbuNdyLLRuEJHopH90C9LWIGE3ybsXj5dWPkWlympV/Wb1sfJQ0oZvzSJIhNevKOcKGa
QPVIoanB06sTWWlWD9EHWZwclXjSVJx/RzBIXMQCq5kkHFaaOt2rdTDqy6GGKel8ZpeoonmBsr+x
Pm9FeieWYQL2J4vhFzfxDZlmcDr5CgG9WsJOB1tO51//z/DPXVHCGi4f7u5w69WTPuQxe0ixGhE2
epEi4mjLp4Lkw4ZCGl92b3vlvUN1GZEmnEcSyIIDUCioICSO8RD970XxvxpLEdzXkS0z7w8/dIDg
oOGwbYyk/XuHPtLdZFcRjNDKm7kIQWtaM7x7sbP3h6o4LZFX0pSU6lHS1mx7wsCIfUImAQpm5rbR
LxOiVWth4IZly/9axH/mrKRuP8N4VEWd0MpI8Ad3SQ2mdbZVPOFXDPmoL97off7J7oD2epS2pR4D
u4P2iAUWRX2GHpGiY5KMJEdLG7IYt6+92qwzVzFLXCphTbJnPeyq4qfCebc5hhsMNH910/m8qJYT
qbAAckPC5VfLkRxLDJfFN4KWMvpWtuqXivupqlETxdIqfIVvLWYuzpOjw8x+2G7sG+O6/GPv3mD8
WssV4GBmcHHWeO6JTY6n9tbxOQRu/kZJcTAQUEGrOjVNMSNEINFZEN69wDo6VJooJ6+qIIPPH3Qv
1Vc2xhHxJu1HFbDs02fCUOexsHZGhR3jMVh/H9aRQ5IFf1jbj1OnQV5T+rvbQndKuGuT7NdRQEzB
BTxKTtylc06lBNeHtYBxCdF35UKwf4S8Xrn0FsnNASaFHu/6AxY1maVnCOfG0srxgai717XXAfmG
lsdCyqCTJVEyoV7E0YzFirxrXBXooO1amg2HtdBa2GHumQgS2jfudlzMU5g6jqoIn/MvmF4QuQIk
YflmaXu0FgQaNzA9Dwal1HFYmp80j998eJk16IRqo1AX3U7Ui42dPfzcR4rfnYpA8kCVmuVFi0Vo
occWEL1aszCLzITa0wotD//SkMuPp5aWLgdgk2Z1fZnh3fhiOZwKfld9fayBaUVYE2WF1VfBz2SR
yguvVPB9hLYNr7WB/yW0twuboIgUMr4DLk3j3yWWMjgBXI56Cay59zpXxpjtw1/a+VR7sug9tCJU
t0YM/ENmPyVj9zGegzxk64kqoCQNj0+Coel8gMeI8ILFJBe/c93Ji75QRg7I21pTFFg/qBb2CJ+u
AixLP4G7WV/vZeC6BgrafKSy75lj1HPx174q9OfnNUJbSuGKgGMN5iA9714dBPVJb4yP7A63cOjS
efXOYvv/lLbO7g3sTyQuChNJqYS48pV/UjVbSmxPyQm1UX/NNa57XH5J0vOudh9dNhKcjCskhcKf
2KyEThcbSaA1FfFNwbDXcy5d8WTWA7WDpDy9iGSdwZbS0YqQ0FCO/ZtCNlI0T5T1EdavRMkNYDi2
ou08FOcILa3GkapoQwKO50t8nE7B8PaLcOscOiiRRYrBUkdTsf0Ox03RdPrM+kyVpfIpMps08It2
LmqrSEFTn9Z2ZrDoOE5njB7uEc0pKsC7h7iOxOgeqIXiizTzw+oNEMan4SZflb/QkDXYBorHdf6r
grB59O+QM9RM6MwbNvKsdKzDODjKL9FjMtJ7VLIjEB/ftj7WaD+ORYyaBw4B8z3AX4mcdErH95uL
n56VeEkRBUXSJxQnGmyhmBpEs5R7EXTz40UvxBDCd7UFaX1+0hyxEas6i/iVUUPfewP0nQFyUKFU
t1IQ5UKcXwXiHRvgHBzJFrI0RyJrfqlmGhhDDRRIo87uh4qGp9pfqpKKxVPnQOPgCGhOo/2wp7El
cj0AlbjDmOIErzcmgSsOYlhj+VHBCtPYieoR1+XLsllqMD5aft8/WSYK6vYFlUUqQwMPHrOlwZYi
f7Bgb+fqerK7V6KC1jFL1iwk492qTNcehb2HyeUo9XVUUft8HeF6lsvMHPyzHbsPlemANqsK233+
2xW8uc328YUuKY6PaLJgziytjl5wwj5FLmptIWjZ8oWVDIM2ISAmSDFRdpS8098+ITcGUHk4DG/L
VMGafiEFFuZ3f6TfHnOZibTvKhSwEwnRJOfZMySsH5YJoj4rB0pjKj6zVA+fm5hoGB/BgBbXlG6R
6G5Wn/tmMNIGeASy/nUT1LGJaBdAfBNf+TlSLA7UhF8QbwlBhtkKTuVKw+XnvWhoAaLuvThIHarE
6odRC63Xmpb8wHlY9eDzFqS95ESesZkwvkZ508ttBCbkh2ksllKNiQf5ukXj7c2G8RabDXcQiMfG
PEUF6T+yE97eVCmJkAhjEkGmK5xLoMRc3bOK8xNWCI8bBU0J4iqLyXHEydz3X5CLhHb2/ygddTy7
zHtQYzFCjKa8jKT0fapJdq4PsF3o9gWH2wLSTMdby8lWBQBr8ZebdnhvsJqLUTtprtGhEBl8LVrh
XL3iWsEYbaWGuVUzE7yccNhAET8eKlehSF5fb+DxbsC273vQNiqAzjmKGD9HCAZ0FJkZnyaBxZZr
hk6xN9KMF9eTLGEJqm5BqE42VwZPT2R8SBNlWRG6lMwG758Z9Pv1fEyx35Gv+KPRDKoQ2UCIMiFm
VWOX3rn41jk9B8ZRUZIJPsVWH2ahuQZk6vf2kllEmCr+kf7jyG5lMs50+WyQx1jSr166idc+K6J+
kLiAC3zDpDP6e88VpFqjgGIFLmADTVJ2VF9oW+6ANrKdDlU2FQO4N0wSQDvcWPypk95Gf+QhbhRR
JAan3UI4BYnhI5oRxKylT4/7Tilh7E1uTMVfvQ1pzUG/y8j/M2enmK74t4O5oKTSkaECOOMQmszM
Joj7D2iKKBcQfmaFh+1kKfJOn+crY5Hm99XCjNQMFtLPJJddcf+aZNA6qLlkm5Z9WRHXnfmmKTyI
CVLds0YYBwoOqoi5ca7Ti/yWAwES+MC/V2U+9Yhrj2aWVLVg8RIv1hkjzxbKaX40j5ClKGILnYlI
Pa7c8F+KhKZpzuwVW5VR7mMKf9ueWUT0U+q/+hOKGuDnzrvQx0UmB5Lr7xgaD7syPeqZQGvO5U39
DKHp1fHXXE9zFGr9virfVEBgGpJZ4s+PCroda3qZtGzOboFv7wPgvgdTM5wVfjfUZsSxCbrBknr8
q7RtC83hpYBHwFamP9bFobz8U6UiPXNW/CPZKn/LxF0i908P+21B1Mlm4GJLTJB+ZlRQILVRFCeD
Qx+OY+KCMjYRABrYVJVAqTt7ulmpFYra2BLen+JrqeA+4JdsljHkaycSRTB6ASpZdvx8tE58QrGa
sEHsyNJBhMFkaVGfe/utQoXOrimhlpeicbA2/x3bvG/frQrhXcZkvRKqPqTysxopHVUZL4f29xFU
OiWe6imLD3uzCqViD35UZ7f5BNz1TcBYNObqUTWKZ6zopkvVlHbr0YQNzTLINtNGn/r9r7cUyG3C
sJfx7sH6r4oicT2o/yHu9fmd29XozyygUQRMbeWwJemKp2QuDINDZoaNgtvpoInMtzpIekS6rScU
Abtlw8ud+MjVKsKNk/J3ZiJHTeCIESPGCgm//9AK05xQdvsg97nVp1GkWa55bjpl2/MqP4adVaaI
N9oPTUlu1O9th63c85vBk+d9s6lVwybGaNGhSb35rKVxKsTjoBavULL4iZtRKBlihVBqBdIFYk2G
0tLeGWTokmy/2tcMxsVOhFKgU7RVAKa1bnRvbtublruz3tlTACQJCnr+CTJ25mg04lMeVjMa50I2
jKuWp30KUmZxAWFxhCE5og8ZELZlQq5Fxtrt95KsoCVhHGlK9vpp3YMVUc1X6SbPn7+aCa9LUim/
ftHhQxFGNoXO4Ab6gLx4Xp3ENXj5MzUxCJevW84vxaJQbC1jTctFGPDHXJuDduxsPGnDhEIZgo0r
biyW7cnjvgw9UqkXPOZBFq9vPfcz/KPnO8peQ59zUGMKhLL+YbnL79LoesWp2VaiJZBjzxRTjzLx
fYurkPQS22x1KJH65A6uQutdXvw17mrVEQ3gSjToeWy84Q/KU+lFKZcLwA762gVBO8NaeMeqDY5E
VnBT5h5WatVm2dV415xZs+hmsDHPb2HNEsAWmxyvFM+9SLJFBpivdzpypR+MaK1YGv3X9HZyGb59
SY6gDzVQZ/fnDjupRxcbNP8CdRT+bFC960KAf7kDjk7wjI3JbxLVBXG6NhneQN5o0DRq1h1R3GvF
1K0XFmK++FOOmgWLXdW5e0EvXwfOQS9xilp8DTIH9aY1/c71FbcUjOc69VloUvp8gqoqz2Z4lgsC
GPdpquBWTCHazd6PQdV/AqSWygeJn6aG7XETD3VCnDUk/lGqkW7a/SodaOqm6IBl5ehnlExharuy
f7HldhOYzVDJEJVNtm5tT/9DVuGr/qZa2R0CQRT5w8JwQNYfFhMQAIQm4f8yL3bjqAj/ROqUAAx3
VQXFjcY3oHplLidlb41Sf/t6AuGZtTAofm8v2Jw+/qWvAogG7YXa34LLDeN004+oyhklLCqydZxb
ZSjPn8c2xLaRMVkdcy5ii9s3fH6DLY2bSIK+7EBX7GEzgRhxPwa6KMZ+qmzeIqB+K4Yy16UVBLJJ
Lh6R1FjEI5NmyWJ7b4mH+J61p0FP8TzU1SSyOZFiB1nsR2mLYcjJ2twq2W8bfsEgTdlB8gewUnBq
jZgX/gv1ZUj3SCcAAp8oxqwY2Tf4KDoORNBtm7IrksCgSPzWMKN5bpfdOoED4W28zZ5oI5tVOhc/
dot1wRVyZuoRw0HDuNSsLjn4kcqTYIxfDHAQxSZ4WXxGKpEb1vOCt+bFCldbBpVYyJRHiSZ8kj8G
uNOAeA3Pfxh5aecokDmU3ajDQWT5f9BghYTwGGyd9EDZ5rsvG2T1svBM0qq8Y5HG/RQQYH1zh1Ia
jTG1VX+Ej7IPwbaV9ofhddDBc+L7BOVPrxo11BbVjD83nWxxPWYa1CkjFRkustXUMdbbIwQGJzgC
LdV7yiVNt243fxq+V28dgnkssHKVyK+O8USxItuGE9TlHuLhGywFc7eLz1hwpUH+5PIqKLLe4CwZ
14qy3BvULAaUbfsQ1z0SXG3xQIgLU1XtOZiUGkjeFoSqBOs6L4fUXxjK03XDxmKbM81J007us/P0
Y3xkXvybj4d+AAnd1w5dsy+h+n440+/2wFaAuKzC4s6Q3r/zAi6pIlhCPn98NtU9sZ4h7UdDcjja
SVcVG1v0hcTU7BmKzsGYogO9KJ3j+RRLWabdeiUAbIPt2CGgahsVM5JNemK7mL5KIEqn7iEWk4oF
MKnZcEpm8YshqGq3D/PQWV7d8wV2sDkbk7KX8r7tZvqLVudFEXtdBul/2yQZ7hu1Znsf7yqziohj
5hxHbQRkTJuOgKhn91ofrfrVJzzz+NZZ0zHRMSIfPOzO816vxYNKzyefkB+y59hndS2TEgetMdJE
homQuiGHE4y/Br2rNArMciw4StHfsI84/FiIZwFUhdYdIZlVXWvhecJ4iuR5WZug2o/9OAoWfIgR
SRchdKXi9XcMGVGmf42zuVU/z0V21kBuydm/i62zLTIkP5VW7GhdLxDVVU4iWfyb5uJvAjdZSqUe
aNHluRNDvb2JZkBNyKVS8+dnZKKDg22OO/4lfzTQ8zBF/frw6LWZzpRBUWPTw3BAFyahGbBi5xb6
NtOoDEu4x12PGeMVv/GbwgsdAuEqlOtHnePIYQpF/ibRAsB48abqs9SRJTk0MoNzgBTi3NPSfFNQ
7nAcNZOtL6TxBEYFDY1p1UGKIjH9w8WtmpAW4dgKfWjVm+42MSZvYh2/aT8sg6VkNj2mjGY5K9Xf
L2WLfCNgUAZpRytjEFAydUWHh1rxAeMuh4wd8eskpaqI27DwTeRRDYzb8nF1Jx5FZgls0QUe4JG1
9he03tvxsfF+U84hbN9P8+ne95XvpA3iDFUUHYS7Vcf29yrNmR1morHwIAzrzKTsy2w26w155jnw
L/cDOAWy1vk8JZG3PWGfKWtX9XT794Rfz9SDmpE+B97YDxAy3dv5NWc3AR6ixzjMyswrnGfbHLlx
fUJAE2iPqmenoqJXYd1K7erEHLTWKnU8R/n3pq02j56Zt4ysxm/0Zw5tqyv/opO4ibUwvGBWgcJO
oZp6UF9lAxkTiTztuqxrpOJNDZ+Z64DshPlmWwZdTXMeTxBfi5N7BNvzFskro2QE6M4d7dkW0/V7
Az2FRWOS2k/Ns9VzUxurxt+zN6uj3ZHE8Dedy1zpU1mDfl7rkYy4fFxrXLoAOvKwHaELYkwEtnLG
SlloM5ZB9awH/YMtSm4E3k1+W4/4VqpozmemXk/kPnfNukzh7X1vpHm67pwdwWDNsNrOsQas8g6Z
hoQEps5lNiDr+s2ltKSCUMwEDV6BMgSVPRcRMP8xeKTZfpC2U82yXeGmBpUsMHMhNX4F5akaEDnS
tqmUWDLrFNHkgbpvvTbs4Pb7of55GrKiRFFeU5DQDPLDebbZs8c3XrfBCJgQHjfUhmHhdHTQa5Ua
cGymgxjUQ7W6BpGVoUbd0rrcLCABzpHWi1k7VlpREbgecEQXrJwyrpQRzBXIN97wMbc1rhb3AHIT
pl4hmgxbbePMFaS6xbzZ+2zRVbGav0w/ymLLR96xoehM3x/LHZO2JpozwXUmM3uI+Z0u42Seh635
kO/sEFD3EmRSkZDfLb3iKYkKH1RNQ+k8V2HtexbXQY8VLW4pGrpsklJJUdX+iJXLbbCY/+DxtU6x
aufSTpOodtwEA7d/F1Lpnt3IPweWHHq4uAjFQ5M1FXYASPx3s3GNsZ/knvvxrWnmJaNSqaqRHPj3
6mdzzCP3XP7NS9tkA07xEJGm18Gk2u8c66Ty/13B42lIEw6RqneDVhEJF87FR42rgXLPyw+e2MRC
2PZPWQOEYDA17QWIhv2CzJfgYvgrr81ZoaD4+zLE0hJux1cRYACZyeNNx1bEMJTsLbEaQnU69sWt
WmzQKALR6A7FwZW7FNJE1+O5HcfIoZ2j99fjJAdccdF/NUnPGvEKdNl+2sgKHtwESP0CGV2TYhni
QSs7X/zMQnyIic97oBnmZZKn/HE8He/4XB3lrNcDvnkPpQzHUqlcqkcapISPVHXXvFxc2LDSpQrt
aufJ8sEMJqaAKnjF4uL9+/kHwRuOq1gYixQoNOEQrHbw01HBKm8WhN9xm5CxLwwCOb52L7q5B9Nh
7g7VD9lbT+lQFYdKpb+JZzKj3DJ9sIKezQxRbpSISlpyoXhuEwwPXMIzhZwm+xShVaeAkmZ71laF
duK05ujv1iO9ZSm5cs0nA8PbYDz2g3E12Xnt6i8Xb6CcWdDBOakiPUXg+XrWZNiEUAbqfIX1U18t
yL0s0/mecRMqLOtUMpqs4KWyKKtWL2shr9gkULAoVkosmSf+INPNI/EoaxWU8vhcMxbL7W73+KF6
94LMwcNV/fLJEqaK2N59ZGZK38nrAtaul3PbJ7ykaCcHWL/CiEaKJ89GXYZnDPtdzs5hW838nugK
G5brfF+dBnLwgVEr+FDSplwm9lCNeY0LRxYPEYeXHOGKiBx3Z0d/pbru+rxViUJy5pAkKMerq+WW
OtyzZLQ7WumN7cdom4Ul0LtOyPUNeMnkoHsDjBWF2JyhmFgqLVNz408h8rPo3OyaSh1WERjcjFTb
BFoYsGikyzSe7zPZ71QGwVv9ugmIMgmmi9LCWRXGCXTOP9SQPExHU93VSojB6NWeLDlMZdt1hXY7
r6uPVkfpA3/IgNqPBCnp1BZu6pM0YMEegaTp4G1/tT6A7qDKcN2m4JaczGZjff+y5obuYXjZXESI
AfeUkmg1W/bRiAuWnGL0Pm/eQYVolWIkOfezJInBp7UN2o/9eaNX/Vw+7S6cijm/KQ+cypiiviUw
+wjyplpyX5rsC5fgYIy7D4/Kx+EwmZ0e2pKkMn8yvqQccvUdV9CjZNG0TSq9LEmGlze6P5+VkY1A
CgPjtfsvcUqGTMFV/dC4S3i2U6Z3ZtcEqVxtOS+x4LZbBgjCf9l4zk35r5R1iL1Htcj1OYaelntf
d7ddxmKYCV/YspjoE8nyH0g7tj2feGDEoWpuZOu9/sTgW5FgltTMHjj9cVECiF4u10UJPObX1/Vz
PbEgfRIkwS0psmGeTynIjgRzpyxXOefirHb4cEU1ZxvogH3/GtrCv9t6FF9c4N3PbJ+7uUEzTdRD
Z+rXQGmICFVafcghnJ4LUG5EAy/KZASBfLpoOICK9Go004hZVi7GsVY7iWY2BfhSHdcjSKvmodo/
i7DWonwXfc9SZBDBcM6wU1a8p/E29HnaNyYiegXNSaGZAz5yicVj5RohNOXmhZtp7g4D7gt/ZxQS
BjcWK/qq3w43OTQkCEdGHiiKAL4sjJ2z2GOHFnIKwgDLL4qlre/CPszXCnY7XQWqbbXGOmgS7Spx
YlBI+4ibrChb/mca1mMl0Nk6yZM+HEy6/67QIcql77oX0s2tHYETRVO9n8WVwfSc2vd3prBa+E9a
hqhEExLJ9qJmkROoGdrsfKzgXbcM9hSXbHV7DZTJgGyjzRCp5yITwdhJVzp0koqhPksUcqEHNa1N
f53xWWRH2C+2cHs1RGYuwy99aY7Mq9e0QG6rGqT5rvQBsRQrGl2eCf7jtcC7Y3phdxJ/EtMK47kj
Bz0nsSV3jKWbeEv1pkSvTwLKeIIJuPIGr58TLsTAiT15p8P4IRQ3olMf5ZTscJ5HSD6S8ZVtL2+Q
zdXtT3W9MKTne6aaHvLsC8t5+SXOlvQgh88Qlyp+U1loop5mxC3DblglUrAOtyGNkWWG8A5Ankis
I7lSOZ+GwF46M8Q6fE1OUhrX7N4cyxyA2mUYRIXnfFpCMBNwPG0wnHuiPYf77+CVce6f4qEC9vd2
TQURScA2827RRqbWzrOLAe6Kz+XA+dJDvQFH6UGVOLxxl5zQUxv5rZxe26fnB7XyDR5BPN5qSyI7
k1sctefH64e2erevzXNIPL3evf2xaRjQbiDRy4vq68WuDgIHUzY+f7V4Ar8NIJnF2yuxHwm/9Dlz
oAyxTf6rNazT7eJTdud65gyATaSZR7ZKkjsC4qjb2VrjEABK6sztRzDuqmzbeb9f76PsYVPx+nfW
D+7Q7bWo4zjpu2JXiK4b/9fIwwjeWRtCAq+qqUa8S5b1VWLVc2VhZ1Noat7MhCfg7eKHc6Ck6dFV
x+5fXDFZi26iu8td7DxxSMj17+bqElrG8cdSJnHqtjomSlJv/dHvGm95D/W/N7sLkiSJS5e1whA3
a0dFeQ4pKW5LzUz3P1LWxJCDvUcavPSvWCg/cle1An4PmNBLAyu8svUDLnafa3uOgCn9ayYxMDdL
ZumespyE/3fNKSr2zmjRDiJ0iwi0o+8s0EXgNgAaqUKFjYE9JLmi+FvZ4y9edS8xKEyNv5sprmwP
v2V/LLwgLjk3Sr7peZUB8z4q+LHEc4hZNWpEIQkfPRpA6DtK1Yb75Z9W0aDKQLsAul+7kZ1cYXCr
7UMBddO72dXjCELmGkaozol/rGDnp0ClDwCo6mGDEyiN+EugNgQmSuNQ5lQigaXhsVVburzZUT7s
3s6bE8AVswhdBCzuaHAEhIPLUZW7iF/Q8/IOCPkVd0la/c2PoHfAo0mOfQJWwqoSi08BkF3t9CYi
TzHEoQk9pi6R51fV/slc57nAtzPmLz/GhgIgPMQ6lKcllz5O9mB0QhDROS0YeD7cOpA8Bu3OhbwA
gRB4iYvOFLschFZT24R/AMXKEhDD4vT8AOsTpqNXsDRSPyy3w8klcBNHEDwcYx4LohHbZWwbeOU1
eae+vcWazRmOvmeJ7zyn57a06HTxTbbOmTao/rn0F0uNS9tKdZDGspGIl/rmg6502RhCErbbRB1+
7qjUS+PkYyO20HrgMblTaPM990IgCpfJonvpiR8CYvVoTIFv0EduyK7HgcYqIZK1dONhUcSI1THE
x4W+FhtMJ4mG1XWV9vL1VszRQ1GykMaI/MDmeJjPJtpHIHtlHhdOWJ1qhtDAhNUhlBUypp7DbKVL
E5EMJNJeh1uGVoE+x9EGDTqLUHHPToKulk0agJElrmnzS4p7C84YbkVH5K9ueb/SJ53eYS1hapwH
ypMvGmFAmuZQ2bml3hn3bR7GuTlRenwVp1fwqT8h8zAxDYfh2zEnjkeSWG5o2YexFFVCm+PEJppY
f35YH4L33Hpgs1y4ILa/V2hZiIU9ge+x9GQMVM91c2Z2XKzxbUAfNId1LAiDicmHrwUBNGuuzyQR
FTzDSAvqMCLoUK0mmKIQIa9BPT6Hm/lbs4TK8KrI8R29pQ5rYTIhRTktHG2iS9ZIO2LGVO+Tc0Gg
KeIJAqcKaV6voTMuSAHlKJpLh04syTA3aYolnTyFh3ROxF6dd3GdompWmFtEk7tymEkqUHqWm+Iy
iJJy0jfE3SUENK9fDQNoRBQN2RlJy4b3JheEDu7S8eB1nxLIV9r4hg3IynL2jwCvYgTUM3LWJTxT
x50Yz4OlW57vJFn8tUcC+LdaCOEsODT/hJK96NjFwTYhntqDtX6e1Z9QMqiPW2FqA+fuX/DCqEyZ
GnVvkpucN4Tes1FvnUkCt7//B+4U3iRfkeYqHkOqTO9miDgO7JdSO0r5uhqUmkLEsz0xoRlY60V9
LejLam1nrcCstGkumJ7MtR5uSNbI77Ummt9i7l5f3Y2pez0DQ47TJsZXSnFXJeblkVng5Y9/bl1r
52XKUwwiHi9ltU692tsCxM5At68OzddTsFDfXctDtvA+qFKOAGBEDS+7YGEH6I2lzDpm7nhdz91J
vJnOeyvOq/ZC202zIirv8EMWIxDMLxLJMdxyBdSUkbSwLAiCCOgPjTe1CDTOfFUm47oue901uuq9
7bQ6SxGQSPQ5lbZP3olqPBux/FtwfmAo6wNIq0SiaYUW5k2PLVe1D1su7WUkVFm3ePo8O7yu3zjW
B5VuRL/XxnnvWf7nOdlu7qqoF5F/qScTZ9hUaAm4g0tfRNjg35c5ufDOz9ts5ZGsATguMqUojghe
6c6xm2yVM1cJ9o38Vdyj7JC6iFHglM6Prgl6QesC6sh3D/st8a4/bFXcbzxxlQ69TUq8tpQX69Iy
wB7B/aq+V3pi43KJ8MuG8T4UtyGKY1rSynw0h6zyb9P3OwzCaMJeul19VEpA5pCtY8E7vUdD20MN
QZ30uTSVZpFmGGcINE3he5CCzGjIBo3QvuyrxYgFXnhzDQv1bJJQzPcdtN5i4PLU1h+S5llZmEDI
1XXP0vmiYt/9xvRntPBkwecahc/DVAHBCRhbP3hZ7++JCMEhMz/YVcCVNkEYSOcmpIJYhBi3DRUE
vQVg14Fd2+1iKhQWCH76nwjgGl16TqduEIE+MAZeLV8l2QyHRSAJgbTcNTg0UQvP3WODfpWdOmNH
YpDxv+jUATr/3Q6CcIaUJQ2nnxojdMopR5mho05MzISPNHBJM791xTOhrBxPYjVhEWZgR+fFLFuE
eSF19guIEhiKa8S39TpQ8sI4aKVrZZzHCkOUCmHdp/QLOh2G1Y8QUYA/hgueCAfLAQnjS/gx1/47
kWP8OP5VOqQGbmW+2i1VfkT7ahdsDOLYqPCiqA9SbO1MvOiNN81Vkkh623VJK+7JmVSh2o3bNdYW
6AdKAOlIKpeBj5Xv5JXxBJFyOHUsihYOXOOBBNYfqS6Z9dz/jr7bfbHIckvHArUvEYzUxjbawqDZ
nUZ+9MnkQ8HeTf/AXm7dQ3cZnclgtULqaiEn1zvxfnIEM1ODb9IhN/v7oT7Ry4+ryUcgDwpdoqX+
3ARHTiq+tN1lWInHCfo8MOO1xquFqUDPruoy0r+figbanFRRKysDIv+iw6Y23ZaILJQ3BpAu2YYb
Tnb7ms/DtmWaBR168yFhUIvckFsZBxCLdIK0eDap5VGmCYG3vdtdbipCrGI6dh9eE6gvNFKD6Wyz
CL0E3T9ceR8yEPfTKEMkq5lDrjPdEplwet1XWMzzqjWmcKW17OYoygwD5GaU8mw1f6I4Bolrzlha
nJzQZzbiJjS74nYCEYm1zDt1jabn35M9JQC4jDA7Bxj5J6Z03F0scnCVsRnkI0Ka1axDEOJGCT1t
/Il4QviyLzSQd12P8gJbRuvWhO9BivNLyx/7vzba/tYWQTIceRwV4C8pS3ZbQX7Nq2YbYJT2yU9Q
HPEgirBCflPVqkOsjNRTEUVMOlfd4Xf0URPvKjNlTnKlpOtI2AitJFOtt/VkXxxJd/fqk1IpmiWV
N0vM7qeRESWVK95I0DRTaZMV06LuUpR+qHp7S/+NycpFQoEH39inRYEqX55K3qT/Q4v9l+o0SQgO
XRQ/yjQtZ+yLoc0sYlB4ykYZxjxMLHq7xsfm8Vaj6orm1PAevtkn/eKCE2xzWZ9Y+/hR3p8oqFdW
Y5bT6zD7wii0Wj8kNfD5vEXuP9bip+PuwhauqXo9T+uFY7f+2MpFBMJtW7Ttdvlg7T+4Vcn3oHUc
IlI9YTEoLaLC/YilOazeRzbbkyjHHTj99CEZeJCRfn25++rVSy+ak2aOgA0rw87dXvxhmzg/DxZa
RngXX8P6o7y2Wd5Tz4rVW68aTO1xe0mB1spt/7X3mRlot3vqsGjTinbDLBV+Z3nT/9s7Siktb9iT
SLIQUcg9vQ4XZVkMDF5x6g68u68pi+yywQptig4fRU4FuwQ+j4gB2oRiufozE3O7vMUk1NdKpvQ8
cffmw+Lpufb2vKVEJw5csAEnxeamEXsPN2QXE6ZL0fioXelhA0cDDhyQ6KGXDNQubm675KMkNTtg
XNNBXmOqj9NsNpIzM8xGv9QjiB9ryvAMDo7UBlt5Srb8V2Q7cIlQzYeR8m3pMcgy5hVF1lGuoFv6
tQ+v3QxpyvuvTM3wTVnJMrdYgPJHW96cDzjqrKoQVodAB4PGMxJBBis40/GelRG4K7ZIgZtioAZJ
lSdJBoE+NNhPy27gsdpX9FO6PpOmnbkOnPb0sAOYKZ7u2vXbwIhtsftQXCRL1GJYZGw9b5QiAz5x
bUdbNePe5m9goluPD4774ywXoZkS8+5wvx2J5lTeOmzLYfBvblqnI1Vh600MNxtVmDD3AZmwplwa
DQz13smyGy3GcjPJxG+wVfwZW6ekINRtK3MYGoG+HaXNbV/BjsPEf4vsW/iXlDX+HFyVJzuthEuT
VHkyxjjdhmnKdtguPT3LCaYlW+dO9Jqv+tPqBFEstvA7oCdKB034F5YvsqD6T6QYe3fQq7iZlnsC
8HXzAuHBxQa3TCCIIEvW3SzOl6/j9adAOIyNXSoLIY9QxXzed3QCHPxaIqE3xjU3sTMbrobCAFXy
NcHgDIrQT7SR7TVs0VmVA/u0ClVr/pivjQHGP1QLR9p1OjG8A3+ylIw8Akq6UzKcfVb3vQleIUPS
QSRnuVec3SvUWt5XwGADAsPqmao/uz/Z/ACoKd4zsXkOFAOqa5Mjb2nQJ8MDxmKIXDZtDFof4r8g
H4zIlXYVqHymLsgctrVVJDLr01fmqa4a7eYE1NrTMZeQCcL6nBXMeOCVlAd4fBhYejt+2J6qAdK1
oJXBUGPPeF31aXYjyjqwDh5YlHKRPzsT1ZU1T1rHopiOZgiyVDUc70VZWD5F+1l3R61PZIBuJTnL
VLJ4KcCcsxgjqna42BA0tPObMybemcIOWtKs07Q17fO80L+vBcYxsbHH3rCJHPSp9g5tuUzuJOOG
oNBuo8qCzrHeXTiYCT3/LjK3FzEHWK+v+f3uz+q/8re/2tXjzFMItgw7re9ecHzdhsnU6tSlnCOW
gunK8o9lnuqnDq/axHXstRjsCMJ0p53fiLRqDoP7HsfkUcwSd0Gi1VrZx+jEED+vAdRZjsphkkkK
2RT0291+86eL/RtW6I59UNsSOcL9TGxN2kr9sjCkfaVNgh/SVn5lc0bibs3XlhnF46VA6hcOcRP/
1kZFxstk0gShoicwRVGVDfnoQYQd981UnwIa4Xwc3AsaBiHRntY3K09yLQydptdsxAZpWbqQwYZG
8+gUTf3JyYhr9/hS+rmljCv+5kbFg6041tqLKbUqsm06Y32q2nu7Mn2Sqrp4HOd+0tRW13pnBtKE
OTYMGVs7zDb9oEuR60TB+PgyoTuaKIoWfO5jZmgnRHY8kBxj2p5SBDgkt0HXM1evH8CNAboIEZrG
gWwZoK3cDjdaxQ5r6D/5VlLvofOIKK9NhDSdgQtGCM31ejfifnLFo2rkcRm2zhzc1hb9keQVGCvz
WaAnX3AR9ZLmQIjnNKZdaoHI3+P9luXJpkOX5vWAssvEtfGbwV7C6Uhcm8gir4OOlRurRfDFmHqw
oXmIz560RtbaX32RJt8jMS+Vnu0ndykFczbsFKHnBUrUdMFRaYVG0i9T5t2hbPceh5TfAoAv897x
XNA3ejF80YvNwvLLvd2z2jQXFd2ydMw8EeqsH9gkBtSYMmbNkK2dlyHAoPrI4Z7t+dVFDCcAlB4b
RW9aqiPZm9V/MJS106seDytaPt8+2DVhQiIirxufXbC3bqoChOocsMOrMj/+28M8cteIHVfd82e9
/6Ujwp9gSwkuz0ApWptKIdXF7efGbGoFZCZ9vWScEdjkaCAG5RtUYyWNoywFab8dJyNFMxTHxE5G
VGIwY68njWrRLCpUfb8Jk7W3/K3txqWyWeaNxB8YjGii5Vs/D6S+tB8mcLbIMO0obSgPTgXnJw4P
n67jIo+E1TjdfR4mpZfVlMtSzagokQSD8rCD9YzKv3MQirTp69ZrkHv6E35PWgdjVPw614/qlUDp
ZRslcuUy/GrKs7YJtABsBZptKxdOPuDEFxZ+ewC7AA+JpTo+bpc1Vx4gbWmPjkp69Y1IlSk1LdWm
R0tZhkmM8l3bCVN6zCzRRC8X022UjrZqScGDTrQ61m9cBmMHOCB6qCVFX8v+Tm9M4QvUFH8gsc+/
d0+BPbc68qCCWpS0v0Mzw27wKYXuBKhk/XbW6KOinC4GFlF8EsRKzABnI7mSwxDTzhH1KrAX3hUn
+4CcG8UsbRzw0DpA60Vir6T/DTJACPV3t1pItIlB1mfX5xp529rQC/hmDMv0iY4ouyNHZweddAAZ
nXrAzXTS1HG8thgnCHBiprYMdZP/tu0Ro6MCGPdwDtw05hzTeVCfCKQ2WzRFrv9vzcL9DepkmjCG
MnV74YCpADT1fWStP6mdO9vLO3M9+PAk2SSEZCws3sTgEKv6TsRw4vwL7dt9XefpoFjQVCmNP4Nv
g9XPHa2kPztMEWKK2b6PJ+DRZEIIV/PU2B9ToOmQwTG06XTkTUB7GS4SqnwvBOuF/BYShOddert+
63TZPIxsdH5ug52vBtJ2IU1J3iT3OoNGJ3ni3GpBVzDQFYHXTX11SxkuNTu+3MmG7v54I0r9u7EE
byugu7Ebzx20p7DAWRtQu9YadjIlH4rho+mZ8xsKyEitN5GGfwEUNuNYj7YLpGOb9AXFNV19vE4r
p5Ha1zXFcmLtoUhqvdB2Kd1n0yZDymzAjZxxwG7TrnK1kDq4QhiayBws8x7eog01/hxeHsM5pE9l
w8zCnpO7AvHPyHNugNPb/EwBSY1XyHSbsnOReez/SPWl0LwSMe3VJhBSJqD22SE90EegB1bGl/s0
wwKfE7dMdTXt//Ye/OCM53RtcKLATyGi2Bpq2Wt8eRZ96SmyqRR2bOGjZ95Om46by36KDdelEYe3
pC4m5fSuwcAPNQolPWhlsGrSnnu84iRS/WLL9+8b2bI4sN8fKpNp0ptf3FMgwX2SRdXZrvixscUg
MhbqPzINLL3TFExMTyTwcXzbBZWDaqHacrgWHz90RFQEFE3jhN12GOuHERrYkTh76S1clYqnGPSO
gWh8VYKRw/1R9HqT8Fb92XH6YC/1+LX2M9w2AaVhy8fNMoYA4QSzpzuDutnj7Dybavt1JPTEhOMB
NXNgegxsZXirQVT1heUXwtBrVmxDQKktIotgy9TQlmzJvZs3wP8OljeICz84TbzfEmBcylu73hSl
2t2iOuLW0S8uqCjlD638d+b0nG9tV2r5uhzGMiGL2K+y7aYmD3pHvqv8cKexz7E5+dFPla4cNzLk
oRrZCt7gHaremLJn27MddfQl3R4o3kBl4PSG6CAJveIiEUTmHCSVoSMtN8TOVEN23tQwPwilcCc0
lI32fSdKhgVmTg61anv1GT54Y/BhrbEwkmWbAW+fqQVpNT4+DqZgsulPptgOer0zKvk8JSa8LmNp
2YQzQkR01ZX8hGufzvKwDdM/8He1+EU7ExR/TsQkcfngIBEi631y/yjqEwwqCn/cq1krr4JV3UzH
kyhETliOAOBcimr9BHlxpSuTHTler6/mq2naRYW/4xHCG9XoK/Y2dFI99O5OokSMfvOgCPutQG/m
kbxX5pNx2eEmYpiZ05vv4VyGXNLJV8b7qJI7cycmUErrgWy/qS7xVDvfaZeYobhhj26FbmKi8odY
/gjIy5U0k0Uqb1w4BapIuVcQx/+6j48KbXDDYvqkBRYKuxCdIkDfdtC9VQ6Hm78kh8//ljqegGtA
Yw3FvOrUb1ZnetaLRGhXbblIu4i5zlinK16EY1N50Mzc7o+ENHN6AaWImiT/mgqB8tFW3/KOv/5t
xuKLDGhw29z8CDZj0+xKS34DYPV/Vn5j7EeUn8oqozCWJwd8YfEkC1wjMPKCenG1CpWLnM3SM+lv
t03QdTKGQu1SX0g2mdcXiqRrIBnA/g+JvU6gD8pQ+kbkTR4zBrY5OSqR8jmtJARUIbMFKbSitjE8
Ri8bl7zdWiJOfaMMANHnVjCi94dxRFfJpIzxaQi+pj2lHF8idH1AZLfGbqntQ++LE0lroJRA2BG/
l6lXh70O26/wxp3QXbh3SfW5PhMP5hOwcoKdmSelGEzSoq0CbHjqK/BA4RHDzP72hTghf+AuSCeg
+eJ2KNFRp5yk0IciSdo7PF3fuLBDeQEHwE70Hv4Zlkz6zduEtXO5vUIu7aoO4Srec9pLvHOUFw8o
m1KUYhw2PIevbgyeEN1NlXQr9uqUDrCaP/ARaNCZ/8PHMi4xBX62QIVxBn0pbVoxcFP+dGwFpY3e
eaRNXNMopPwTR3qLTcP/szN5E8L/5/KX22ZdHzPheYPn1ZuMKnCNq0FC2R/XM4ctLDs9sbl3ryQA
9kR4g5E+KGH6MiUDfq/pW8Da+4vzZVUABy/DNMRm+0pgws6IFDM0tnhironpK1IAc/OdxQJ+Dhbm
S851vUz2B4+9lNzp5cDb+GMyDzg+O8ceNVMdr6X9KpO/oGaDg6SImOCbcr/7V0OJAQJ9kLWiFLM1
ve0yF+/x/lph+ehLguVGGsK63JHGLVE0pLwfXIBEA9W2GgdOQwUEp5S8mOaPKHuYKyIeW5AjuK+x
BBiJIX5xFdtDG07ALun7inQWjDKopricDa4BbIk7EKz525LoS1l2uu34GENPjS9Mz+8ROu2rB0cD
s0Jpv6VewL72yQbNNSDMedN6WjAiF5cYM7eXdTr/iuy8ukalCO4Y9i1VsOOC2RWAyUWKj/sIaGKU
wCbg60lNs9JODJ/dzI1trXX0kk0x/og6DkXUY1a6zP850QYdLnkydGZ1PKLOK60ATF2Sx/+ip0Ur
IFq/24l0IcP9oBlWx3mqCn1B8OAE1KupPYyKasJpGrry+JtFhH6mLXo6+dqhkmuyI8AP/UOnUjcf
68pM+pXZ0F5xR1AhoZSeFQL0bkvnCKHkPqKMm3bs/daJZmcjuc/7Rbma4fXQogjvgBcsokDD9AIe
TsqyWZhJBLB2F+fJXmqlnpu9a+DLdEn1fhmQ4iAXH1rbaKgjWeo9DCUpBnYz3bIu1tP+dm/003U8
sXE+Uw4TRWdueWhkVmvhLt28JLLdWK7jP9LN6NO+pXxs3eRVC0IF3nAoRgNwOJtVyOJyb6clOsHy
Krgjzi64AnI7185FwOTPeL6lLhk7rnrjs6OBM8BQaA9WjhiYmEsWJwI5MvOHo0YqZG003csnLG6S
RPoNDphkmZvZyhY+NjhOg4BksRfH3lklgGywz4ul24291iOPr+tIX6uOZa+bqo1+B9Hk+94SwfmC
Q4Lu1tMRwRcNzZ6LFibHOPOh6eYr6Zut9tGCMIbygUt8atNh/iqbphN1aPJyLBljVRROVXBW0FMj
NQRm8nEp+TGonI/yq6BYPffN9TBw+9fGgXZinldr+pY9MeWfNGH9/0aaKGXSli0oOA84yPErpOmd
wBRnKtd48QvallyFJSfy9MoJRO/Z7r75xuisRvHyEW5JaWFxEHx3qywMK4TlF8i3y5a0TsigmdrX
cGQ4CcxBG3w7ULdhPayWY0yDdfE7CayAfiBBjtkFjxrul7uxFdd7uIxZc4f+ZiNyuFS/bWPB/L+X
+kxNF5JIceQiw51ek7RNKE5d+iwHO2CbJ+GrtASNHURGtLDqtcyNrfYEWg+/OpSmgsi6lyPRaZKy
gD8b0nztbjEhk7rfh3tjelzmHeSA9TeCpdfwzYuQu6cO82rJ243GXQsS2ItERMIfauQy8Bvf0jfG
situzCwCs0bkbVv+zCPvUkzVpv+6gkz5aXzq1Se8/ga+9ArFYaQOPeTNLWk4IUHSKc1tiY8+wIdh
GqqO4yGIYXk25vLt8YdAq8UxagM+TlgKdyFpdEBZx8wH6r2toYqnAgDQQblQlS2VqgEwgyGu+Bzi
l7pM0kn2H2D6RhjRQmHPRt+uR5OeNHk/EIcipDEdZXNoyXhWuNhriTMH5D+xAGYCX79m0Yz/qxgv
+wFE2Ts++ldOnDV9KWcxc9yyw5x+VlErLRejYRVOEHGE5MHkbMB8sAPEEMrsTa1+IDJr7iD3EtPF
iyMmVpymwomOT2IVGGRhQ0w7tFLtmaANhvO1Zd63/tc1lpFUfTcqdx5v9BEMBhp0WGFJDERkKM0f
bUPO2x52EqbKLravUBDT7iTnGIEXM+kUrcUvm6kbFUH2GlBQzvRICr7BtoaC8pwfUo9j46vj5ohX
uPhRVw97sWKj51o7RnOPQPQiQfVv0pqwCKxvP92Rr89EUTQHD/+aylavdK9ha+vkoAbLIGsTWpfn
9MMC9uPXEbsMbxYNV5F4wayjVSBe9KfWCt4Puzt7Y4qI2GzZYk+8tNQ5QojUDqJyxvtfZhLdC9GD
4HaldoNAL4FX9opL+lFr5cB2nNDXI97ggBGmj/WcTPjjLWWJm4tvFvib3rpkpOk7Sr/2rglVJbew
sPpTL0BzCmqyKjzaFgR4kcsoMBgznG5FZ9ojj4ZgXx1Wwu1ARdl4PNIMkgc0T7DSie4wl0p2H+52
fzmM9kAMztMCoDNrKz03UC3+3VG4i7znlIIGyT1uOwJricbwxA8K8SBxwq3YxmpgYloqxwS/O1mL
JnY7vj62pXtKaTBYEhjHn9D7rJlgQQ2hnITwbxt6drWNfa9te1wCm4k9R4l8SKPT0a4BK+vTSLyP
QTyVfrB/NpNHGYF5xziPW1Ap10Ms1kV7fFjvlZSRPWYfofoCsi8wjYBxE+35+wykbESmuxCc7hbI
g1aPBvkOaONgPqClbAYuM3ZUQJNzcKnSBkQ2Njg9Uoau3pnTJgvQ7jtJdn0CAr6OySgqAZ25ZjeU
YEkWkDOijgCfpurWpQqhKfodR7vNO0z3XxayF1Hg6ewicJ/2GjBWTWW9mu5/NNAfioqgqjIJWtJ/
I7At9VdLltogN4dEO+CJEviiVuojs3jf+zn1dnKkZt0XmZpOUynooeiL63+7w4gtB2RJdAzpIrVm
nCEIvAemOpg/ZwhwdeSV7rnK0F8AaRW2cmtu9tUkjVMayGsCry5kigZevO9/vAHO9PAiYKhdQMXx
gkFhqEXVvHVPDzjN921ouiA0gqMC7w2sS+wsCwyin5+iuTozKLp99PESDP0UnQa0SiOGYPg0f68h
gBXcfWDlEEaLu8KjzNOxWmZC29w/llMeKkcc2btwndarsWuCw4mB5A5WXVJAdGhUaHQgAhC1Z/+q
C2k/V9W8gaT5m2F2/w9SCqo9djeCaRKcSVtiHhqNhNIXI3Rc5inCeginh0pt/oOwCyCWjQdyt6/4
5az7wh3DoD4D52hSBAHOddRyXgi0uIFPuIb3SFN7TYlPKYqODumRAFrCeQ2gc/2kYWNbFJHeifIm
UtemtNkMNUqg6bFjvdhGAXJeqah5tzhACCDfjvVfovJu5GV6a/M2FKfUccAuDZ1YXT4VpWQ3ikxn
pxdW6mCutF1RvUs7VdYelGNzgTfQZrkUohZ/ehA88twk9cZaln8F59t6BaRL28PQo4RAAjBQ5y3C
AWDywwP5e8VSJdSWYYYjSNAtx2og2FBpkey+x4bbNqX5dr6o2txOH68qKclpchbsUAjgvBZKjBvs
pVWgsQnkhxkiDFv00015IYkks0gYUWuwwhgw6hekcKlZvqe1chlB3xpwI5SHvYzJBc+FDWfCAiI8
N+3XWQSmvpNEtWVFcOoAbCPtZeR9GO8L7lhQPPAEpeiGI+naqvJMu4O0SwAOTM1wvAi1aEnza0fu
hu+ZfsvnQT60nYimVHv65sFazGXxugTAUJSyWMa9YAz+vXb1sDtEF/ZxgWD4HR26Lf8YKzB0HRzx
USeQezu+eb6W/WZTRfyUFeLCZboxNKtzAiz8zb9oM/5874A3jD14j1mM1iiewAQGoeK28JJT6JRj
Jp2KgDBp4F8wGY3yjR1rKCgMToYchxhFn9k/hRDA6Xtt+3hnckADb09VjyS0GoXu3EW1vCiYZj2K
mLwwA7KqxkDJ11v7juhaCfpE2AbYSHOL6OwazI3CvOa7QZzDJ9qg7qDIHoiitIPOqAYKc4LrMXia
VtMRnJGZw8pgutOV9CM0Ko0Ytn9h/cdZnfvb50WR8mg2aUNi9ki8Hw0RJlw0VoNbFy/aFZToHeZw
R4gyVm1lcg0+TR78zr0JgetVbsbRf8r7Xl8ZeNrshUV56a9zJ5Cok5MSx/Zxh0+ZYN8Oh03Q16ry
1Ze4SnVWVNR5boRNCgXzv6YMBPuflE4FpjU4EE/vhETRKQ8dTzV9aniAD9LAR/E+5nD2ejTsxMiH
UuIEYFqKPVAyMnUh9QPzkKh4eYhJYP/2OTHet/eAgkOK94QxtGfx5QIq5XqTOOKZ/3c9g1I5H+zI
uC52F4HJR0kefWQmCw0a4EEiZgzgrOoVzQYSrFQTi1xVicSQ2GzM5CRX2G/Lt9h95+HmZWj/WwCA
MLAqL66juY81i8FxLr6dscUQUvVOCINcDBRK05zmZ6WJzvtfaAZse9G05NQolP9tCVOTyslaQLBn
EmisT/nbLcVR1bduNb4kblQJm/Xr8D8JXIiccjXfVm5vp9TadkjnJKWkfcaDHRBmI7LXqXtgxP9y
6NJ77l79LBbUPnkE1XIK+mH7Cvb8kHQmVBxNwzFf5gvZ6BkCwAF1e67MVJq112RfWfKxd90EGHjX
cNXCyXo0oEF2dmc6zke7Sa397lhaZdQFeQf+FNYDLcEGmBnRtZytG0lCBfiTVCWpUBRWRMCTymnT
+Jan0OzbB0+4eAhXM+996ydan1+ZC3/2TW+Ued4CC/eDnZNRrz4AAqrGhriK0N3GVvuehYHhaMSa
+Epe+tx1ds+mkhTBJ32bic9n0bR5HN3fXtiZELC8FlOQmrfqQTDnupz+H0upGc4QVuAeKkfnBtAl
qv79r1f2YrJwH6Nuxc1ASRHdYD9fd6DV/hOG8o+bRquhj00Nf7hFdKdMyxuCZOXX472xE9W7CrRD
AzZ0ByIEVibIHRGUsYs3SRxNls8aPT/WvntsrGERsbACXRcZsz7/vrk+Clblo4zCvMv183bDnRlM
41qNW4DKD68tYRwPfbtawsufJJZLSCVo97d1MMx0REXE/20JwqjPqgMOukuRlCweDT0aw40ud5p8
yHTxljco58D21AZ7BKhgjpMqw5j3KiL7ZrnREMt4pfFlya9ETPYtUiSHowjwj49XNCQFflidgMfX
oPSwcOUSN2KGZpTSCvQH8JKraIL1j+IQgaYoHsBvqu1RRwq21cLZWNzS4D61TDGY/SLwOzXORXMV
e+oKF+ko9X/Xg5CzD+eEgbA/bnBOSoIzogSteP2mp2JnkFSobfmxhs+3+bcsy+O9Dy6S8VWb9kFp
Aybjo9j85KM9bHixVgi8NPmfwy3mt3CNc+GrvOcgOCtsw9i7X1cWO11DiDIr8LUuhplNCqNXw4lU
/J0S8r/2YltwlzUPZJto2+a7Z5XxTC6geTVJxjE4IZ07x3qry3Yz9HvPkHm8fYGNMpU7V/XjNts+
znyyDo6twcsHrIZ1UlLfFq4RdhPd+KKmHNkZR6J767R51kryXRmgibhxrwob6WyGU8aWI20QfwDI
XFfnGhsXRN1H605UOSv9ap+xXepozQ0wkXxFQuhhYhCG74jE23d+yWFSUjnf5qVj1Zf6JzjommBy
4AdlXQi6II2tBpcxDxJpYUpRvrk1oTHxjXAtFnybNk9/vM06fW1Ho/PaRryCX06i8xaqQk93sqq4
vh4s8jwh4YqRBWizZHApuPikZyMJtgBCDKrBdaxIIG0ivnYwOlmbzk0IBwtttn6iOnn1Tbr302Fz
26rv2KXXcSFtWvC1QntfgnAyWokWsD7Ou/fH/xc0Gr74blVHTy2vpzisNlmrM32gzHjyZsrCFnU8
aKg0wEcQQQ6196kughzprvHs0+yyYQ6GH+QBrTNoPqpltshF7HJctrmTJNy3HvgfDDgu/Dzj6nfT
BgRKm5qe41GEDynmhZnLDF4RpjCBxNzAUU6zHhuvo6OasVqWJ/d7QzEWsxBnnIKjTyVu6Biei7+y
3s8Rc7QDC3eWyvFSQHVU5YJWkj/BFPHTCtgf3QEQfnXVJmy3GDhcq1y2X7bh4n6/5Rs+vMB9mDwK
1ADKFgnTGCJZ9VRfjm5vLNT/p7iwmvezHT4pfaDpjETxo+ILu5cHd+hl0HK6jRkGBBeHIWVQFqnd
NDGQ5+yRD/22/tat1R7ANSQQCoFebLrJkdEbnV5DRW6ytRGW8eXUPZa9sMJ9oqeCWtusexp2hfD5
YlbySWOhJ69BreCcI9QpC0uAvpRYFAcStc46Tv+yX+ayV0XAn1DOOEJ1Z8D7al137r0bq+mQEbmH
jDszJUfXC0ERtcEmWON/vjD9hbIBz8Ul++5MRrhw/go3u5GtMF95km8Ft1SxB7cTVG9kauhic3xe
Ce3zRXMBj0FZEZ8Y4Yn+AFRtJRAjBKDubNU6MdQ/ePmO/YPtuw6sKnqPTXypjmVTAPLtjK8Z7OMp
2j/C2NUY0yHooZ4K7d49M/zl4keeFrClwKojFJsG3e9TkEjXlY9eBUuSMM6O03iQBbAAek9SI7ER
FINChUL/IS1Rw92RMACoPD3ZEiNDTU9Yvu91S4IzvS+458SSKgZqAx2+HETJwxbNfoI+8R/8nuiy
JQAjfBCkCJ5qh4fmEf6SyESTtvS46Mc0ydEfS0dYVqVH5gMdeo1aXap82mQ9S2JUbi/40TuKHbyh
CgJpVfWSE08yKWFm0xrIAmuvdT7/dNm3S10cEfv9GW7q0oGJHzkDTqVvxrAyOCxAfDAmHGCYDryd
9tEig1vH3CNwMqYfzaTci1ab66FnIgbpO0She6ORC/v7ACvs5bhePSi5rllY8MZsHas9SH9aZKUi
HML0c62iPNBnRusTYyqxmXF+ctb/QJp7mkxxX/yJxQ5EQZez8MP810M+Z/EANcjEuPcC9UQudlye
t9He9TE6VxEa/Ut/CmyZg4T2SWnh5cDlJNcsWLuyu+GNv0ab4jTUTYmgatV9XIieluU2NIfdB7AM
bS6BOmFRLiB47cPYe2edSqP7moNU25Qc1eHCjPh81qYzgkq7GRey7pxgaxib9GGEMjSH4a3TLzVg
Lb1XV1LL+YZQu5Elo747J2yC7Fpil0t4t8zhAn4xniq15LEIC7Snzei3KiYfas+0RVMe7U4Ufoq0
gxaBkmEtzhdPBu/Zr2MLZYY0un+rMPDCs1xDukR5q0qoARyh1crSj0NJ4ByKcfoAValFGxAP73lj
ecuPc2CaMACWvIKawA8qKs3DWk9C6Oy6mNK9qOZ2AFe/whuPstsN/YSHW0YqLie0PvN+oNR1mt8R
VVFBLMm9+InR0kNzPkCvxij5MbyaFkHTulW+qOxvaN9GCCbGgSatIY2Il34ZFwE9LjR6VFfczXkV
BZXAO9kBxhoT6UnDt/VhcGpKsb2crZ3unNruIzMUqZepgDJ+9bqu8F4HeUX/hU7NqIxnHERcC35a
O0TSJjGBbvKiheEQLGOUYzS0fXe8XZO9QDIVCVB6tSUBmvZN7X61r6aqRQvbYMB6JvZBmz0OEjyh
VkbXyjhf0cc1gHwZtgnTUh4BLjbmvIKHnRxc6jVFZnGlq6IeIPksF9fb85YRDS+PdAxysaOe+5/C
TdkI5P+DXgfgGsowhpp/QcNrA8Qx1jI55sQGbAP+XK7GekKs7gMaceYe6YeWJt3jNF8lzoM//CeR
sXb1UXlw31izmSkDg/j+JCCIJul3yyuTIBX3rpKj5wrNaKGh9OI2KlUF2ifDCPC/nW9VIzdYlXRL
S/qJIYMf5liJBKtAKfSe96XMiqBJy336LSS8+s3DeD6F4kw1FmpvNHeRsOuvvDTa5m+XnVtNc7U4
JlFwic5CL+qXxysgyLM82Mj9n03arj2GF4igZMS5TdssjDthOyuj+A6laWEq+QJZ9BPyvWQpMZHU
Q6J9G2nHODaFVLLIP4QzojGHwlZVaZl7STqS/oDOKse6nh8cl24O97tx9XSwIxG48oGBNmjVnVZ0
0Zh//w/7mfa9RLkjvhLfJGa+hU86ZsdDYq7asi2iSuYaadP50ksxdq1zxAXsNJiKbrHBw7+f5A8h
YNwoEIvellKX8nUyWYC8ib9mSfS7gVN5NZBQkcjzn5J6/Ri3H6x1gBfQ3r15P8myydufJVvISMeA
DaTRYOS4XES1NT71ZfLAgzCXstKSZNs1HWTHdnxlJQRTdfva/u+VinOgOAxC/7LRcvdX2+YR4ayU
KqG/apfzeXYziUHoOJpp4cy4lFUSo7i687Ifah00Nqm9yXlkZE2prGaGpkvfHi8u2d9Sp8N0+ph2
cCGexppIMy2IkO3/ExbdKq/K5Xqsu0a+7fv4B9hQy09bhJULLimb+fQzBSMVFY7eFADQrnxaD278
WRDfPYJVdQHIthVXP8zoTM81DE5cLUS5709HXGLSeJXjy3ZssuYGkb55rHgk1QvaiP2UMMujFlSn
nCrcpmxBJGg/Y4s0PzRS1Ze0jg/CgBP3l2CBCwnU/CrIGSdptK0NCDeEiJIT8FW2HiadEh65avHH
1dbdrJQyPyvC9uPVvgd8t5VxhOU+WzNj40T4QlBjMBODN4ViA+oBAr91Xe7WC7rDnoJJuclPSyvr
xOhzP7Ib5d2rZTeQ8wJGqXZMxfbGTOeXGvoDN6ExmJbKrOPcXiO+J+u5vSvZ1LhKaJc37BOQPhez
5AlOeEgh2fTCMzIBUoguxsLmeNXGfIhKAkWtxoHDwm/j194atp0SEOkGfnxPf1VDEucjIOYysTOQ
0asUNvtZ+6eUIMKFglxVMH22qn7ZfE8H9ntMV6b+MhsafI8f7052J/IpmQkhPYM6mrHwWzNZslK1
Gg/ALZhfdbdqpNN/1aNSM0lXglnng0dNUso2c8QWZ7NEVagWA0BmMdpPJaJ22f+WNIyeAZTUKqHo
3MbmZ61dyU9ut/uEp21vTH/54ccyxi1K2/uopDaKB4BRjlmdPtsGSy0y5GCkKL7jpJYGojUEv9WF
HM22D2/Iqi1UQnDDp8XsTqOsmOCSpggWTJFlWoOKHv1/gSk49W9U8ydJY0vRhSqwDC1aQskxPDn0
mLMRRiaO+dA1ZSq1x7OVb7OOJw2pVAGfuuGeHdjlyenzAhSJw3eMzVECjFeH3dPZY0jqfq1N7AcO
mU3jeQb2ABQ5EeVLoY/MsNPa55ZlNc6GkGLm2AOE8B7WN1wb+BCKr0GwXpmbc5RX62mCLgDtoHEd
t86I4K4wiCkN9fJDM5JcY2QdVeAm4xizg/8DhE7giqMcgXtLylzRO9iWh226orn1sEvq4PvWwD9u
uYDz/fQDxGThTD3+A6ju+k9HMQZcvdvxaQTq7IDOtnZRB1a/yiCcEeHU5vwfm0fj+fabXINiCeQA
CBhyQ4XrhspKTnBb11KXRBYPnBUDpORy8I3ZrIqDYqmJYASLt2mriUe6tunva3CnmZjL+0kRHShS
uEGgPO7MjnNIgFYxh0e+3jfeJkVBVugZkoyWsnlqKAe5mBRTVa4sBZ1+JqVjRQQyZi9gbZimUXp5
aDgog9HLl53ufyhgXB0z7lAGnKtkG7S8/MIbGyW3Bi8mMmxVAzhdUHLuD1+3ug8s1v4EihsSUcI+
p8Mb9ZA25HHlioShX9nO47u4o6nqcETr5c4xhrL12LxYr11TVtIcWNU1AEa7Ni2ozRsptOsTu60Z
1IEaW2uhUB+/SDFRIgXo0732kCPC3NyqpBiR0WZwf8yuIcyojHgHjPSB59FESi4R1soAvcRfbMXH
m2b7G1rEJA/vZliwZZj7H3nzffznxYL7LLLDP1un5VM/8b2utsiYju6pd1Mb3E8pgUlHTynSRLil
6YDrVrjoHbuSHGMbRYAtdhqXz5eHgqZahZtmNRoYYm1lx4R+q7VsC6NbHHilvtifxvUyg9mDXmxJ
0Y8JUrSN5X9dLtlmEtY/ju+G9oSNwhk4fnNEAGn+fDyr+f4ET68LXY7EJ0FtfW/9VseHTVFdQ767
9rrvDi6nLZPdmo1tL+IAtzlcDiRbCtr7w+8FukrdTH+VM8SuC4qDszk+pOjHk3DPAd2nOJOE0Wd4
AsPQ12GzR4JdXvHTVLQivoU7oTFqhB945K37Wp1DQPd2GOrN0WGn+Q77Ge4QB+IT2WyCRDu+ACmK
6ZkRqoMltGcP9cUWhzeSf7V1EGo2W+Q2BgSAPNjc2imGMNa2CEd2B+tudExo4LiHl+lQzZn1+v4/
2mnC+6KhQz355PRgn4cK6MQnMV5NO7RRlXmTFHccWTaVbXJX0bU7/W2Lgis2KV4L0V62m5RpnlgZ
Jkz6tZfyywYS+b6r2yBalTgdR4xtXPPjWWyeBSR70kf12zUTmDTw0rK7y4GZ1y5s+YUXHRAmzay+
F3WxzUhJGYBjPZO5NKULh7c7JnojZpBxRFIyxCE26Hu3jUIBCBSuqAa0TCJOc7UtJJYlHKMmbooe
8+/Spv2SgosE1bZJi+atXdUCn2mw/cT4zRu/ylIsM4UfuHafgfTebmNNrzbHxJpSLh3fid05ZS7r
DcoCbEgCC5Ag5oZFRMvsdrvmAKL5JZRYDiOPbzdyIjzdQqp9W79g/75ycrhXVNROMJ/kaT4Mz9Yb
x6ttowgCXhHs1T8u1DcpEkDali+xnBDTx9kTJ3ngGR71qJapTyXW3dcsnAo08wTYJOcpr9W3le6U
YgN/LCIaj5esbXqz/0YB49zdJ49ER86xIsvxEXOG0sYkbiJKTUNRvf/bpYMdB3Hq+L9REnppz19p
EsRMv+PsZvnGepOxS/dkps6q1ZgIlJ1TageNe2DMyJpejqWSZPLE9TCO8+SLGDw0+1uFRGEdrJol
N0lS13X4a2G72vbANB8f2m2Nm1EDtjb6Jt8aiMwJZ9lMm5sp/xQG3lwPd5+W7ylkVfcckWSAbZPT
6aHl1DIU/q/JTLAsPZOVzzHwm2rq9YcmRS3Tb6+6gRZ3TPJgbx90Dmz8cmPg6iCXCI3gbAecDlNy
nuwJELb12HH3S6nhGpdhRh4PWIfCYe6NUHENhdpyg1/4nIOk1JOcAgJMmkGIqux9hYkVvF6e6Vuz
KyWtPQcs6XqIUodxKV+ZwMdBsiCW3JpQRmTRW14OrKfRUlhsI8Ckyf7q2Sv5usuaP6kWYptmxcBr
DRbsYwHi8B1TpFQdLygnpYWWsC8OSFb+BtVxXRVZQwn3K1o8SIWjruTPPw7qPKLt8BoARzJZh2zW
kR/kmu5L3DpYCxy6j/yhdJY2e938miOtWJnW05yFPjRR33dHv0y0YUjfHJFCKhyEg/rUaGp3/bg6
8WL1Ukn4Z9Sz8OM2bkVImZOYRhCiceN6rj3zuzOvl19quU4t2sMNJkLJf9WHrgbRYQSAvLsJ+sc5
VoWjaPO3/KnfDc5sfkVDDifEI45l4IECWyJnCsFMs0KnEtmy/as0LOV2MqvJ2MZT4rkZo7Yg65P8
KD4m16fE0rDJkYFvXOqap9KNKrITQqtiDi8Tehl3C6ce7oPhVwq42+t4z9c1qYrwq795zEaQW58U
q+hcYHx6SAQanrL9fKy7ClCsqXcmnjIMnUeTPFpE6BncZ6DolUl3ahPWAzy+tFnM2DmIR3zJK0XC
qjCo9pkuqn23G2zDojyd5I2pU3LmTfJRbvucgVM/mL92gkC4OrokUAhhYLfhHHZmZgpH3YsGhVyb
oAt8aFb+mqcfl7r/LMSGM0OE0Nks1RnkqZc/Kku3p7queXZTZmp0/dDAVGFtLMv1D0Go1XBX41cO
a0QVGGavo8Vb6qEN8jtlRijLP/DPE0LAau+lbl8FfvYGMUS7NMoyYx3y4D0vV0dHez5tqt1/k/FD
NaMMF/nS11D/DFzLAkpAiLAukpNfS+sEEzxPLjD6d114J8sAQDJsGCq9ksVHzU9M6X6udpt30LCX
lQdBvtM88HVyJJX6yOOUp0bPdcJyqCtO3wYFLXEyIDRuIeroS99zz5vWBtuO0Gi0ydnVfbpOUkfH
e6ETenPDD3fLdcIgkUU5sg7InfOvHDavuZHxFuws1kWIIUJgTeqm9gYBjQX9ucLMFkneM+vVuF8h
nyq8s5OGdrSfAQkfRnfaSpWCtcGKIXR3UwXDI8nWPanvlo+aS634c8VSeEZmCa1UWld6+hbr0+RF
ZPefjZ6gdEpz7XJvcpaX36rvlBD0PEBGjT2O8DFVMbhTQDji2ctEZcWUdo+OYKVP1PE8mkjau6PE
pK1wAHIIFCgsiJxOkVS0dAjA2mF67zt6U/Ke+midO/s2WmBDqfmpULZpJ+7ONlJxgrTfHsrv4iZz
YbqNy2Qk8Aa3BIe8IPZqxAIMyXLrNfCoKdxtuX8NexQZlRAmoS6sDdXJbebf3e1BWJa8sQwOXcmv
mOxwC9Vpqe4yatfNdbfxgD7YkHPK0roFB5uQdMr3mXmIxo3xxFp2R7DiHSKcLhQVKCTvdKq+LnGQ
2m6vxCrOClDCEoWfaHUKNza9K35fy2oa9rqIejWGmeGg66S0KlKUoXbf0qEVGZ1wGEVMWJOjhGr8
d3Ty5Je1QxbLjN6Swymh049Naz+Ggm2bzE/h32tHrzQ44Xv+h1nBQHL9y/WN9jtuEBu5++zrgQ3q
PLEr9WVTyiJCA2T5gg4jy5Ga6Ai4BZeOXLxPqNCNDR3auivAomJ53utb5bLMH61dlfmhh83ZBySG
eo2mfLuXxB26jZFbFZrrT2fn/UHi6MgKUp/MOsCtiMMmFz9DDvoWhliDYyChYqyWVbx99NYO9Dt6
UgPCq7yx2PbxAQSMkhxsUCZ5YnRcgQBpM5wIyZ6JXsJKVWiLa0ejjtxxUXfd1gr0IT4qlP1Xa8Fg
uysTEJn9r43wJ/YS8tyG/lY9R0M9H6Wl/5oAG9j3SvfggyaQE+/s8n8299i9pmjiNPmFsfWprMLS
jSwvlBe3IPqRde77f5zZTGkcukQP/41HzlkBBuIk/vfLYA4vGtcyEf5n4BME7xyIHM5SdCDTDIfU
nBu0DLpOv5LvW77KC7eh4IIX3xb+CVDJj5sybLqW+4O+0kWfgfpWcOkfSmzI7yp1GOssmXtGQ5Uc
76q9L5Fmo/4PV/VBPkEKL4R98OqJF8j9ecTwjyweqwQ3iURxCcO6vR+n50RUz18gQzDnH+8m0sCg
2LoQsERFsA/UIStFDFruClsMZA4wtoiTazubGpu09Zl0RTZljhIipnI0N0XVdUIPXRuaGbvyOP0S
83K4CnyENkvmOWkJeVJRc26yjIi4b4PqpaxZ3YiRv8dkEntoejZcn2ethfWJC8sfF2T9YvnUX+cM
htnm8uJ6+3y9NfedZbY7M9f94srYLzmPjy459Rq4qCFSaIvTbaDeF48tRNHasMZBx20acZFwPSAi
8VbC5a5aBn+Yi1lGpgPMqkwFhd68FUDjo5qxfcnqtO0qpF3rHtKvh5pD176JbIPQYSg1Wvb+o414
if00ojBkTKlFIjlLU2kF7MfPn7mTLVf5LkXs2utl8N3aAcJ/8lGmJk6ZZc9HTGzUhD32ZtClSeoX
VKFn3cheT1CjlkrtcLKo2x9B5LT+olsaQZuTTeJ6KcQ1x5agmsHPHWawArhlPziTeKeLngKsJ1Lh
u02lpgoDCQvkUkRg3qvH/V8ydNZHRbCyn+Rdmn8bmP/eLHiqPIt2lmZR7wug3Nzepb8+Pqw1oRXf
nhXxz/yWYBuwkCdQiCl9frjbrfzwttbZ6xHho1J3vVpIgZLRJWLyIQ7gB2SDjSc0TWo9nVlNdwtg
oHLCtkeJE3u7x6Okgg3oYmOOt3Dz9hsHu/lY3Woga9yvRBR+6oZujKmEs9++ro51oYlveQyMOSuD
vsLUKq1HFKt97xHEZvTU3wpYrlTKsnk7x9qkTJcHGf/Z+SurivRRQluy9/jxq2FmyuR7Xb8Cqn82
VuriGaISnWqZnnqhtGT8QxQI7+ojv7qmmSLjtZUk0N7VMzdDlQqeFf/OoESoEqmMQF499FnLXIy2
1P72uh8Z7R909L76fJ0eLYbQUKMHYvRRMHvC/bTVxbDGASCrh6bPiIOOCMxAZH13RgZ3XiS8xK/O
blwbLfo7enxmJcDpzjObWKKB28mTA8iJQYeFQfN7IhIWtf2bga48pL34AhgmWlM/7TR2opdG+eVr
l8UpLR34yhQ93mCjPBWmbMj+AATjvfRj9bOXnvBIc6DejRYWXy4aso4gEjlotF1FocKyncTqtzeF
o5tLc3sZtYUpHf47TJ2eBP/8h2AB3FEu47IUnIIgrBaEQdjBBQO381BuLrp4j3dPsz7N4Wywjn4T
e8bPM1xugFpkZIoSIUYEa33tUm6RQgs7JPmOBbLmXo76bA8A9bXN6/gwrBREdTCRg6zWMgRz4+OT
5+GW0tnZLx9zd4045PPOBV+EajM88arqdpLlIFiNlKiimXKRLleuSpuxOiGJ7wHTk7yRVpRCFZ2X
kFsDiK0tRx4s0CqO9IWSD3ZAhM2xofw6uFq7yE4g/DiIZYnEldEmpSCfjPZLR+aW6A61tvSFMYrw
aJnv3C1jJklSG9SB2CAI1935mKKnh838mgZn3ksEvwmNhLXWhqjrg8iQ8sOqGN17NUpfqp1KBsRR
ycrdjgEHEyKQwJrZDRtZcJ+yFkNzkgFoHuZ1AXiCUOPBfUvtYeJLbRP6T90oCB+zddCEmzAvq3Au
5ttOohpAmqKmr14zJKnXXoIUQTzI7cos0gcivs6tZR7F6aUsbURPSGPNYpZN0oKGoYWAgxDZCwWX
su9IdlTEL0jErInSvgB5NujXHlrF7fzWLEEv+pXqFrjlyn/6p2ANrtcgJLYQ9zrJWQ/oaxcmUloj
uz0sEKNfHNA81eFkgpYV8mMOhuFbqzEdv0N6PYVcjktxpBzuyA5iZzeO2wCzgnf5RX6KSxAR5V/N
tWHqMsO6XaM9T3C4Es8EPQzBLw3raui2VLWX3iR6ryWPo9xU1W3A3w2DA0jWXUOS+wO2F3r9W148
3oppvueMfvLS5fivZmEHD+zMnPiRoKJGxObPKNaLEkBsGl3hZbCU19jEXcChFxBz1TaKNElH7jxs
J44QVEleCtQybUsGQig/L2jwDma+VEwvXzMmkRNr7KP/hjUGBWHZCCEcHC2FLpS3cF/3WsDPzjAb
PLnQVOAHrRHW1TkQ0Ewqi7u55k1dGenCvZ6j0YBlQCyZHM7UN1oAxlU4qTVwlFW1aIm/JsQOyTnN
aqYRNTWDU1c2k74cpXPEQsguBwD2IkljSq6WqrNq2T9KztxGmTij/pb5NnwOBb/pgs8KzVB7STTP
yFhluzMcECK4vkzHTZYOpZ/emYD9UcGMVJB3G1WWNx6tnFvQq2D8GFArJ5oUO7Mfr3Yv3hhGQedK
qtKg9LuRxs4lWwHxULNsgP6NsjmnASe9t5fAqh+cSZwqvSz/H+kBedy0M75jHLcC6Nc/qufipTt/
lPRUq7TsUT07x3GRFmZgLaFeAynRdXf5knQmxZfiIG6C0cFBFHDj07D1/RUbGwudyNr94uNRvp38
IYs9kdojrU/Gb6mDRcb03X/PtN4IQumIUJJKsDLoGqBcoCI54ohj/bmlIBWGWlvAd4anrQagLgJM
Pb/3eSdftG+dKLk1CFIrMa9i1wTJlnxN9/PnW2gAje5d5WXkbKdchTu831gQaINvZTbFMezherBa
F3tl4yYRLn6Q1SEa43ZNRCfVIn6b4st39vjRL9wWVWsk+qdMWOe2QTDF8kNEgF4CMiPzrm4L5bYX
GyPQ9aJH9H5aFDE++6w1Hb4mAvYzDwSbX6Tvi/glwuCDp/8SdwQ0E8sLdt3HbsSzajLGUXNgOo3k
XXcPrPVMTDnmyxwx5ZASilHrkOcM7Lc+PdECc1oQAzGIKS9pIuFcN9FE3n57aKu/hhgGU2iJNdmp
g4Y2dOO/Tkr44DqW4BH1WR2YoIPhEG4wkYymZe8Qm2LOvmllSMzEy8XiaWkXboCFiIiEjcFlvMsn
5MYL2XF363RnwAr3xOlB4DBWOvupcCBWUIiL7oxFMenD5WSnjVy9O8dh6NT+Mk/DVXPaQg1sn08h
JIN+tV6Xh2qNmm2C3o6TWOCZq6q/mgSgyeW4187N6KLkW8c+v2oiMKytroTvakM7e1GwnMjsqrck
uehPt3ld4CWWfIJC6Vj2i/oBsRE6TM8LxxdxJMeqSvy79+EfvTShqqTbf1tDmicMyjsJKkd53eF+
yX1+JOVKQXu5lToGhmWFh3X5A+BU6kgPiU1qdjqYeWWdBwptjfRBkQqqNRcLk8SSbLkzH1yLwaug
Ktfun7avij13l02lOqPIMUF0/DK/U118r499GWC/5YHctBygM24FIRS3D68CeV5Ly5L1cqE9NVAa
h5G7PdsyKcj6v9CNIONO3A3p5eX5Nrg51e4TPXIIZ7fPsLInKaeN9AAMk2Hb1JkzaO12r/vYssTz
g/fdxw+qUN5T0G9DiPHTOQXYk6+jSURZQ5Vy+RC0pgDHUVjCHSHNO6zi+yXiRmjqSiSUWtVViqwd
5PhKFOIoCTQsOI9GxOzkdjig1jm54K++DZQOZr32ceVt7RGdZwoSULls/tyNZ9WTqRMA4zSB54Wh
NtiR3/1NspOE7Xn7W3XqSDWYl/qQT/i0ajwiK3XvJM8g1RSpgJybGa79bjcJc34kIUhh+o/kklkV
USX4lEb6UMTleH8RvV5MRB/UIYnuoP5JnbH8AdGsQKJqWMGe+l4Onx3tsqZVVqypj5LxAcuq+bEx
4W1eEYdNX4fxKsZibRqVJnbZSDOD4Zuy78zSqrU1yRr03sxRLpfJYNXmADPD9vdKLjvIol/SbSHy
7CNRubPOK/rVaRV4vAYMokcTB61RQ6Ex58S3QZ76Pn8A3ZpAEHRRAlHgK0rJwMeHprdxzkS4umhx
ex0wWuZ19Me6OTqBUyQwIKkcV6Q/B1GjAIswrUAseH3DvXb9PEJnAVvTmMxn4AMQOCqxWjrPrJpv
82aZRVkWE2OokXGGSgi28UD6is6ICiQJ+Z4Le038Ez9qGNFGDLMXoimCLyOj5FKMP1/RqM6gzbi5
rFzKK5C2a5mXrKXnd+YNewtGlxL786ge4NqCqemj6P7jSlo4YK6Pttvkq3ziZfLPXp07GfIxuQ98
8NwCksnCQJsqcpt5FSYSHvIbnsTMM6327J9u1sbC4hzsjU0Lc/tPdFG9ZrPVfFWd/uP39Rzb6TZ1
OL3DrARwOYukuHEIeiPWm+e2FJhBEQjxyVvg5+AbvkHpGQ7jGZCUo52bfKDpmxDLNUIca0cfxfEk
2qLFEGC6SpQdajSw8hKFHXEE8dveQ3LExfITeWE5jetDBQZKh6cH4Yh/UtF6SzTomcUua+C1i6Kd
3lLGp0xNdQoNZ1zpE2jX4uqDLaU/gP6bPysGBAmjF60JCEKHzNj+qk7mMFMhtNHEZKBZw4bHPST+
mPgWad898EbQpBZne58gEebqdh/vIP0c84LfyN4Y201GG+AtqooeYuiKIkCipLVTw6srOuzgeZJH
/Q24o0J+ea01h991ppGP3WWY2e821LUIghXAESI0uSm3YFNeHSTXKpctSu6Lp1DPN6x19TZOT6WF
a4P2K48revOn7o+ifcbt3J6mM7c78RVwvNVvarUgGtPJB5LdC2xBdiZx+uGjh2ZNDwPRkGvzf4dm
1gvi/aLOTJ2YF9Xu6YqMiX/wsRPtu7DghKcvTwHgARBwtmg3RJfLHBsH2Esu+h5vxV5jpADJYuNl
n0Cc87vOhCOoFg1qp0DsMeJ3KZWTS5Pdg4Zq4c4t9ShIz677YXagWjT1vWxT38k0Z2CPY4tv3unf
nKyGeQ7j3DQ39WXiK+rtN0Lh4co/gWbyKJtItR9L7tBulAFsy/HN5NS58zbQvZ/ZVT1WmPjlXp8W
GraVd9N+ay99ZK48J71UU9FG0TqqWWoZ/fvsqY7CoDVWK1+Kw/0AR9n633iwzg3SuDmBaTSNXQS0
uy64Rwgnm2py36VNSApPnQ9z0QUzSvXPlsAlep/VCCzHrOH5yssAXs1x0oQ5OMg6rEO9M+OHpJQ5
IcPZvUVbGrRZeenOcrRe/eNqCLilhB80bvnLW/g5KdViEbv+tUqZRu29mdXtDA3VL76+4fibs8yz
L3nLpC4fG85Ub4eOzYGAFLYjA1r1+9V5fMRa9K6PM/l02o2jKkMmcVHmuoeeR/cZjXk9zTJ1l/3A
qvtwVJDPVv3HpUwwQ5iGMauMiCQkKnq5VSzvUFHc1Mfo10IAUyckjQKNcyVcvjLQi/t0xDXqEwrH
x4PVcep8Zo4PmKSMZymqfK7Y8iy7fd7lX0loCIrhB5jycnS0VOAekSiJZMFSZQbHXo1yH/iHL5uy
iEpS8Wg+xPIOPx/jU+Fuk379sT5szxvosEvdprODlneXCdMlvjGJ7eWoUPPoOebVgjAPLJIkb/KB
X8aa68q/YZyh6aDEFOH2WNqCr4Jsl80p6Nj8MH3hIn9MmUwakCiVe+YUP1EavHYh3Wx265RPaGD4
hZeDSW2fNWvOsQ2ppDo0QQBOnDBfzXnwrplLB64hzHyWNqeZ2hLdDfd+0oQIZy8g5KXNgEX/2Tk/
BZ6ygjkmxpGnU3E6slgCtPCVs5Y+ANcazq0mpbJgXd5Y86ai517jimuWJsxAcIPd2rEDwsr82DBg
YDhi75vQ0OrZFjn2qC4L8AApa1gZcoqsTKXe7xrAE1fV1uETfBVTRPWUdotc2TkaWUBhjVVkoDM2
IOIAXi/tBUYI5rNEtnyeOgx5W5Fuo/+7MuNUAvAWUb5B7l/Yy2FARmZE+5yktGzfxyQc6NSu0jxp
/pa2twQTA8qEs9Pmua8cLWU1hHXH0wwi5OTWRp9PtYjGG2FfT6ejiQthufn5B3Etr6Kgn1SywYh+
3Shq0UEffXZXmTwJnLhGk/0o2WRdTk9+XuObdL8Pd8PGJj5w6S0JoZR0OTB3rF8iWYaSYzaeFIEa
N/gRlltCY5D8MMaSiMFqhw9sk8asPj8gk6FeSqUuiRf3oNn4/k4UKuzwlg+uFTOTCnK4UqzcJUAe
bfzQeNfsBdk0IuBIc5nHCgYXSxg7BEQeiNNVMxMlHJVDKq2DTY9DPVVv4tgHhcMINzo9HphJyDhE
sWTtxtvsxlLUQOjfk4IS3k5jC4Yh1ycpX7nmu3bSSoa0EUpWr19A5TbVbuaEgMLoLV6k+dNCOOjT
tNalJzcUGLC4j4kfLSZ7uGwzBC/lhHHuCXvECbMUXcYrRIfCkMXj5q13dmekhpLNjVoc3EuAtLO0
lCZURvGbykGfeKO1//YN1hRPASnwLmz6fi1YRtH9WEzvZkBYCTvyDQX7LQImOU6HCCowSyitwOaA
Lq7KVxtO5VJSLYo9CGlh2DMUoxnzkaz6nqbLY2v+dghxeIO6Dv/3jlDN1E3t+RyN3gS/5gXnf/Af
IWRvprZVCBxB/8Y2JEj4zQ5O9Gl1TBEA5QoKEfQCbCAbdgtbgK07vDke4apjT5CrAXkclsoHBmkZ
4EXB0rFNdh0SlzryrIXFknhOUxXW5kD/DHR8sCeYbwg1K3th0zCMkCTp26RfyIeNHhGqrgJEMlYD
aRogvG5V7bIF7XcHbpmPdEOXiqVY+HuohudRj08ug+tT0aUlQbGnXQTsJ3+DHmbPV+QaExZoVYhA
xVo7wJj31/2rFR/ABVDA9uuAoCry/3VBYBMOwqPtV6tXeocCbmb9a3b0Eh99kQvdOt6fOOKU+I/k
HI/YndfNvmj6ZAofX9rFBdnUPEfmM1uyWqMBjZCDmgQE5acFXt8GmRLQZvu86JeGvJ6LUwwliM/2
lg/vTt96i3Tls85FHydW1FJ8f/QLSmlPyYE514+EvPO3YoOmAPRlf2+TefUxo3L1oRtp+ysYxkUk
6CNUpux2jM/Y2Jf8PfrGgxmTqsTqWlGyLdCaJi6OmZsN4Q5GL88dhYVJkc5KWJw3+Fps/ZxutxVy
vyropA+Bul5SrPF4YW/Mvc6PwSlG8LU68qSUrZq22233hW4WoI/87qcy3Hkxp0LkFimCC4ZNAzKN
vBiAK5CanyA9Kc/5CHAzYnxJVz/sP8d78klMXz4gdcLTCbRaM7L0lVC8bz2l3iSgUBs0ocooRH30
Ajg1fpNoQpmXemNSPIE1CbNoleeFAjNUF5SoUmQQtvP96JM3+Hw2KyXlO/jCXukLIpnM6SVgPjuC
IAeUoNwkNSnyG86n4FC3fV2WI365djxMqkf5GZXcK2azdjS9R+LDyMQmwxWatT9+N3VFlFdLmtWW
L+vuru2j2vX6ngcmUl//fVDP0xuRYrUVFEdjSXGuZBLs4FopDLPGF5UdYbSLeUmejHCnWcnxZUcm
E5nCEyYSi6ngmcx3qPHgPH4gmsktruZ6EOpX22nRtLVPDng524VY2yixH1Q7+/u1qMHxWJA+N9HZ
Okx7o7iJsp975v0xF0NzPK9C5zPRJz89rE2NxHA3+eV7WXuVC958cOuQe/B9HsiatVcTTYO33q/u
CmYaERPWxUmmht1QaZN7HendmHoHlQb7eupx5g531aY+qu/g9SYf775Gg7hDCjX1jeCphWJYToeX
Pj8nygYJijtB2jHdnx4ZDhQNwTODRPIOtLyUOTCG7YYDTW28tMs0Ypg5F0yebEWSLFShtCq3349e
kNNBwRp0DSyDbv21EfESEQ1BkuuOEo/E2UbBKcn3qCUc+BUoPtRp2gDDzgR8+0Qe/i98wGqJWRhr
e7RecVAdzu5ck2PzyA9Qnm0VpxiHxBxQlq/nsw2eGHyaeG5KPrRBn6lDd3xkLGb4Qu6H4dtHe4bg
/CxXhmOmc07H8rFGM6TGWUBgq/j0tXhhPZpzLpQ4fY4N62OzkJ0tqxbY1f4NsmKeAznbyTE7ikQW
W7EM9bCOlFhefCWf93Fdkc0AWn0Fx66Vw9P/CyKiHpU6TgEUNCzqpP9e4bmjU+V/QgHJgsITSUaY
4xy5xLnp/T+PW0twH5+hdXu7jTgSBJl20ap96+R48ryZO+bn8FJOonQqRJi6SmjHEYL1SojK4JEb
iWRbWlMF8GQblpzQ3I6tJek1CsSoS3afReLtbVuMK4HvrLfPB49akxnBtmeKI2lyWwOz9MppITQn
VIzED2dN0aYpm1qcIoPWYELTrUfb+UwBHmTRuu+hIxf73OIpXwZTAUmJ964qicGPu/QwfBvETJ2B
kulaXDBi0tQK7f1uUdlogYPY+88dnrP93xR3WcUO5saSGs92chqfmgj/qYyIPlTI+NYx/VxGQCeb
pq6PR74Ph5iuqXsmHuugFUUkEJto9G9pyHIgcJXsgK3+kaMn7DZAX70peLo5yfRb/ldM4JoElwR7
6LpHVRLG76JVspiAl7u+QgnkmeLt1M4/sf1Cm9i9wY4hpy+8gnzRrebyTcEo7yxeBpz96ja6pIbD
Qs0c4W0Dk7RtgmnAf29IMVbBvWbzu0tUvYqRdA9uGBwZyM3rrBbTPDTcuVA3BWR9LFuKHnjUGUIw
8CMDWiXsE6O1fksYzw2S+84G/+1iZ19oAwAK/tI4ZLECRVT0mujmnyElPQJ0A/O/vyO/L+by/dvH
QvLJGuqJtYaRKPhmcw4lcl3CWcpEOZKENRS9+hNHpl3ETHvOjj4/fwdC3K9ovwANwLUT5HglK6Dn
22TzpZyDuewVEZmxHrqYhwqyHDSsEbvUcJmGHwm/okRbA5ZzsxabBc7zjFwZK+Fw9LH2xYBnDdEb
wBREhvgPb2UoTZGfp24bEiB8sedfGyUA1kC4kjjJStcSs1B9gYJCAYN1jfzrBwiObozF1S9QriHy
OecqRcOJpVFRQiDIK+6/SzYrfALlSHl8t2MykDETok4CxrNDcHHuIah5nHBSKAp6KO09tPBIqeZe
B/Eaty0EVMtXrM2ZQlgE2IHwpazsCkvYS/WZqM+eyhsQB5VyFA0/ez9QRWylio9moKF1gbjw4qJx
bCZuVtNbC636s/NpUXLbt93rb7bFMPI8DQfb9S9L4PZeS9y4G1a4VEjVTb+U7K46e+Pf7W+th0i0
6K7Dd2Rb3reoI5IDCL1gAhYiQq4E18MzmrOkX7zNsC9FqZcbLjjXVAvmCAalh29DFqjY+Pj2bgP2
54MtC5X0gSJRRSLOTmDkD8EZGHYIRJs72AF3+bHcfQruTLKf5++gB3+XLVhMfoVMMR7SHCnM9MOx
/hahg1mFK4a/L/wQoQuSC90usoFrSJghkfcFav4R1ynvaDgSrK7ekRG+Atpp/rwc5jnRajKeicI7
vi+jvJeqlhLyzvPKeS/68LRY/oxrzFHpHyn1SYNa/Y8hqjh13zK7TECKCRhJWcCWUzOecQtnPCFU
/ahWp5of9kDtFzr3mPKUTsLpbU7VGJNBDZoi1IKrjfLLMl9XEk9xtnkx1v7q9WacA3Q0foYmEU7l
ybnXF+uD0jYw95PW0d4BNZkRdu8vX+c1Ds5PtkC89KcmXd3WBdHgXztUhRQeIHWFSRwlUB8v8DfR
vNNEtdWTOv42+ZwhJMFl5td7i0kt+D/SyKDXeLB0u3TqiS+IssaVG4pBJY43IhO0Q6E670yUgR1A
vS5i6G5OEns+2ehhouwT5IsJH8sw09iwFg3/xmqqq6sDY/0hZ38eDvMFWyhyQPMLcpGGkD5uH9rc
spsWyX7DpmPNRA37bQW8e03CX1zZvHKFSHix1Emk+X+IYHAHGV9d/homNK2va7Un43YvtXX8Q5DJ
MHXWsd5jrIQ2K5MuOVinj+T1K3Vnbp4eKkm8NADhXhhl802HC6NApxUS3jQNhJcjpMKao9JIO3SV
5O7YMlTm/lMosNfZRLk47j9jPkxnLgvI6ykeTmnTKI4HlDVpeoEnv0+VCXOukuB3GoE89bcB4Jaq
VJu4it3j7/o1so5rkseYeobZtf2otb2OhbXvQKDAFsTYXsn+vfefXFUPi1hNWfiiN92jzuPKPKQF
KjHsQgnpD0fV6Sm9r0xoqEmSbhubh3pwUjfdH/AhZNjjWz+Watq+kMsQ3BGjRVkJsC5IEvcgg/80
+h2CR/UogNjBIiJiomcT37yY9jjJS1qvNS177bD+4MlUuAcuwXHX8oEB1yzIbMl6RtzPU5bc6POH
NFCRnthhOkiPsntl2STpbNkMAdvieEwpYo73A+JzwGzHnt+amNDN4qQZ+0ZiiFUfNkNF6CzXNATS
tC1LDXcEwQtZE5GTyNjjbgNyzNH3f1djddEDSaQkNP3BubUpQGYV7gNLe4V+BBnt6gh2NBa+lYXn
vclOqh4i8vyorFm0gmYkxuseANlSv3phwBrXqP56KKjwR1ELkSPEl2f33OM/km7PXJn4RdjKQ+Ki
26mU1uEdMSwoQt2/INVfA5Tz8B9bhXl4ss7HW8x7VcdlH4H4KkXB+hYgEBNfdtmw/NWk7+rhXUoy
tYbKfY8j5h+nTvQDJCw+voc1mDlVe2RvKKQnrpszgXmV1nW1uboBDQial72w8VYI0tDj/xjIAgNe
hqgA0Uo0pgfff9TQFFSuB1UpVdBsUr41zfaiawlmmsPMNnnncPPSQc9oOzyzIJrcG5D+NzR4DPoJ
sSjf78h/MzYW6Ah5YGAptcme6SthpsnecStutOvkjAtavQHqs7kaZTDccHVs0EpbLfdTNSoKq6uG
BJ64v81f+hj5QeFW/2055lsCQ9Yz2azhmd4b+Y8ZQ62QBo+HNeH2ZzEVpuWvsrgXp3egjym+R4uK
r7FGNEkCzPgjbIQ7rKFP8PwJSbX9q5m4DFmL0ihQ2tycVdINA5pUXniJS30Za2zhj422Y93uRtBA
0hVGYoYqlSj3q/GFziuUQYVN2AgmtRhuXE6xpZrjjpwVqQOSOXRDtF6zKbjZeM3uv9Z0SBIUYhgB
nbZSmcjSoVAl0joyt4LAoA2KnATCTCjejRJD/5uO/Ssl1qIWrjFjZJIFIO6gSwPAkPrRNxc+vmZY
Z2Kxq4aY3U2d4ozl5iQwL5bkOF+YaB78hv1dCJJWb8pvqjhEiLAsK4s95bZJwk/6n1doE2kJskm1
HLkxCMOn4xa2EongY0FWor2PGG8BwQC3nSE7/jq8MzLVTLAPTHSr+6S2AnWGgqHNjGsMWQdGtt6+
4U7V011DPuMkVIgDOxOGi97An2GOmVQeMTx6eqVhUjly63qgrSdETpgb2vGwj2cw0AcXSUQ5RzD7
TZUkwQes/CGyUzccfT+FJ3GoVup+iROKg1maHtkbILoii+fOepFJAzdraula+wAfOq/Jl8zRkcE1
eKqR1SX6qLar82suMM5wWbAK+Ay1S0q8nJdmrywOEXfyuCW+YCDNDkRYfzC7ha7nQBb9R6eTbNMQ
AXV2WUqRzzPcRabqyMKC1Kr/sksX3VcsEoU3TZAOHGdqSlgH6nMLNdhDWpsY9zrlZ6nWvc2Uyq6V
V5x33qVV83oLHqPjdimi2hWdgZx4ZeSgmtz+kgVwu8pOQILwHCdxPJ5XgK4VQUub9IZdoNXriint
gDcjfppEu+yP5bTnirkLPbJ0ZJhf2mqu1RZ/hJCF0Sfg4PMh2/8UQVbtE5iHJcbzd1KZXqIgAcGz
8NpCW7MZNBG6obhSkUXr+O6CnqRdxJk62WBQhqZysSZjChmbgwS6TqbsLZrA0qgHEDMIWHRJHhQP
efGR/28wDrp4tkLzBJwC3t8D7yM1J47h0IX7lofb3+AE6lTDZA4/YDqvfm72NMhywQYcsHncqsyo
ofcX6/E6635K01no1QLG30n7qxxja3clI9rFWva6IPxBisFe/ZrMGD+1TgpnPL82AlgFUb2KH00O
WnXAoFjr3T9seUv6W+GtELd5d0y9zipX6qPeDh3VD6FJmAmHbjTolzY44J0T4j/WOr6L+r6V1shD
DDph+k8s7cnBEknOg/uRuJw1lpYZgy+jYcUWjJTJfS4Lthgw+u5pXSts+EIpj7j4nA5nTXlswgrY
tbMPkrkzSM9YBukhHYI1OEwspZD9L1txI+fNZI99Q8Gkaq00U9hpr0c6rQdCilqoWi9lsrAjNvN+
4OOwZk1TrymwM/N3pMEneV6ekaFohDWPh8ot7EBQtFTkm6bbcUtErnhzF2slPD7Bkf/Xm/UDFe2n
Q64TWCLmazgdyeGdfN7f8v3/2Cyg5xBcBIYNH+TRReE9HECYmCLDFkshP6F53QJ7CkrqtRjBPNkf
qN+WJ6Sw2PcSpu9eFxxBqAkTRqPAM+jaYisXoufPwbRlGp1xL6cedFWl8Co9wx9NYW0Vztm4ph5o
M4inz6iFrLX+L1MjG6YtGTQgNmG2gM7v9xRZ4YH5lbG7NR7TBj9VNNbK679NfiNPEiZiegM95YWO
uOkV13weVkd5xItKW2inDGAPgZrhk9er1HIZ0xXK5urJFDXjmfu8i07HyaM7Qjdd0YaPIzeG2YZR
3h1y3Y8SE5tdGU5s/Om8POrtmU99IK5pfgSNuLzZCVyQmLR3oFDCOpQxEw7w8cW4FW4kGqczQHAN
KuBGm6NLv72us5gycapjvztFRN0y5qxhvTd0ehchQtcxDbOjdCn/YAu5X6Kc50XvsCn1f+4aopy7
yLz+SncZ/xOokvIeGHBbeg0PLEaaB+15k+KncfiQobk/AM1lVxKBazomEe0J/bxnarEnX8R55bzf
O2bjp0I7BtoVc8I1DPtswLDmsVsP0bYhDgojtrkIjZ+GubLIiaPNpCqoEhaTUL1PjlRuUtVYB9TN
BbbdFaz2BHmzszVzX+wPWj/A9KjmaaKeIiMZ5WMcpuXExwiWNmg8k1f22HPyLthUFoFV7WoUtuyK
+SGuTIpNBc2amIAeZsUcI9QF5hw8V+ZHILGwcjEWH+SNlA/wjOvCVuqYeDn02tgL2BEbmIQVkOTg
Ptca88/QihRArx7qveObDgvJkkY1fWMIpWlptVNlVjHNpQ8BaREX4DKx49bd0WEtRTvWMiZveaQy
d9YiZf9FeDuX8632KRuyYohboPVaJ7b2mbYYmxxHw9WHVJQ+tDHubwQRhIexNu2UcBLci6WyMkCJ
6LzsGyHC8Bs9wNUndA6mm5EjhxS7PY+8VGdDioCX3fligATeXeeWx9EJqN81nYZnBPsryCLpNU/C
gJvlCzHOjRZ4NDnr8ttkfKkVSTd3UoGQT/o7VvymHSH0Zu/HoYaW7HOsXEKNgl8DKdfipvOCXhbw
+iIxO+7appPxHoO5gq2YeKNJp3KFGSVWfRphHE2j/D9WdXmpw1PPYjARkYjxIzsf7wap7LKr6tY7
yi0TUil6vZjqwpVFR4f9T20vjyyYW3eCz5eE35EjjFiWEONeZm4CKvYpivngmgQ9ApsH/LWwapSC
Do8fvLy3IAzyy34wjEbFCS+33HIMrM7DXBsJQQWldnvuZIzRNck5kA//kRWVOyrMtUjunX6ThHa+
u3AMAbj43fQdNCtj/mYbpn+dznDFiaODrzI6v7qOflLz+ssCt281yI6oHPDkS3D6HwBXFLWfujB5
zOa7YlxT6U4CTdZn9NrIphBRECRvpeDu+r/Pq/pMWsrjHyW9uHVtjVSqE71BopKmHJCyTvFsTLBW
CqM8eZx7fWfBrSf/Gi3FioFyLEPIgxY/LfxRIaZfXascXZfhMIimMPXFNwrXFqEKXsPuuIXRThLp
Slt9IJ1GSM3+U8S/KRNXAJKcHzlIP2P+7a3ecXEHe493ZW9bnoeupmh50h/3z2Gfal0i/isUOi+W
bQxqnPglkv0lRvIFI1s8/SaGdftPn5ab8c/uaqfBfO7Aq7Pz5000TKaN7z5ipq5OVSSL176rygpX
YnbwV4XLzfgh+5xfuaZ0Etn44hyPGGJvKTNQK4W4rbd8+/FjhuSxqkBO4ZyPlrvI3SaoLszevZV4
7DIaTiG5D+QOuzDjHoF6nVYBhDYlxSBOx141Jd9fZMCzCx6Eyz/h5p+3jqTYDKae+ujSsFpeE6F0
8PkRhnhrcf2oADiWRzNZ2Tqj68tIv41Oepbu/aN4bt2hs17YIS1KU2OyhxtTtm0w7i7+1U6lq0PJ
oZnHYZP3fkOTalbRxxkNreFrcU/MaeFnLdN/k8B+fNrhWwFqTbSX5k9/Vcs2lVhh/uI0SQmKuT2h
HoV5HkH+iTWh6nL0ai62kcf9u7EwZlIqM+TVPHhvT4A5l1onu0CYX0U3FNoptcwStwUaC3pAR4bl
2T1ueCNDREO/0cF7TbCpiGGb6mDV9qAthBLIYIA0uARUCHu7kGr3O49kNbrZz/6CEkojY2PvdTVg
mEJdRL3cMZODep/up8PHPXZpFJ+lYrNcCob5uHCbk+RTmIsk6/SbwnRQ8sBRsiI/SVjONHXe0SlX
wUtgh2hK21HJfHJzCAEGtdoOspXPdfZuk/kGJ/yflVQwDaiySp6znpR6e2xoTUtqOAzqok2J/mWi
f+pTd165cupo80yXHIxxYxO6oTypZV92dAM3LTtZao084yPpNGKYvEzvqYx3VYwNYBgwYbgCLPFR
3xyOZ5DgVC/lx8DJJly6EtpNUZ3l8tsooxwPju9sBamM7kVmDGSVxR1diAiHABlA1BcQTx053tt5
Cxv+sjCO/BrAYCzZcC2uZh3T1mccyCzmjXotGdejJs26LeMHmYdabxbn24ajo7TgjKbVEHlr2sxk
qdBJY3GepwvoT7UrhmnfY/JNm0RQ+Z5Z9+uPM6B3mc+1F/leiFfcaEs/ttItr8oJWuqtMBy9qLIy
mFOb5Ge32pLe7pXTCU2ubr7aYop3zLaeD7j7VkyRkJOIk/a1A7B/GrZ7Rsgy/qADMK4CukcGaSNJ
gEyMJgK+oz0FsuzZmSfWf0F81QfeGejrvq+eBLdTGt8aLsTCgc60sJCOcjIidxMzT1uedOwaegra
cn9i8NHDtjm0KgkZdoqwV8ByjfwGDIwRYu32z+tAZgh9yYegTrEV/S/bkThJaZteCke/784lCdyf
Iz0w+5MQS+WdTWRtrX7+DUAzIjT9gXw8yj5Nh/L1XmrhJsKf3SS903PoXUytMMLm8jd+MeJ0bQ9P
FjLIU+DXq7mcVek4KHS4BUFl7ivfY65acShugrpM01aRtKDHSkBssy4u5IxG9NUP9nzNjDqtOyT5
FJnACdTDf4i7MGAYgt0ht+bFoYqsgPb4XcBsm9F+KshwPZ/MOoA8sKZxujA2Wb8UZsS0F2z6189a
gtoR34/Ttsysn7FIogcMJIJLUr2qdBl+vqB2skUONSoubjSYJK8kMkSuci6tmDh/d9CL7dCLENcB
5223il6sqYFndFatGAA7WaYR/9XuyStih/AinC+3XtylplHEHa3OCKdZeZHiC1t1PiZj+K9lXDou
MgZknxdj5ruAlKfYmLjMx5EXXjWemIGFSj7EYxPV4qPYkHsagOjeKSu7bbzmFSDesfXSKUWw59J6
uZcpDI/sxaot4lGUU9HIB+mmE9xLMcgsJatHGjB1mpeZ8awZwwjbkzabLxQLaT4WIJsf470z/8gH
jVsr58m7tBbrqPFsf5yHAq2GwL8dFVTkWrx++H8SVRrXaOg3ZcNuEhaGlvWjHwPFPtJIEoUR3W9N
14lcMtQ3v7oqgiCl25Fx2q1PMMjxAWOttGMXITvh0HWP6gnMhaDkLiwEHQ4YUcqhJb8vibjQNwCL
Qkc1lfgAu2sXKGRjk1nZ6RU17XZB0D8OdmyyR1QIugFbK6Qs5YF6W3JsiqrXM835IdHVZ7jdgfj7
vy44mf2dFk2hbpHyPr6ndJXKg0NP4yE/S5jZIsr95mgv+rMWdV4cc85PltAavhKM2RLuHgxRxAU1
xrMQ5jJY4cqo8p9TgnqUMFAcYIULsyFIXd5KLZlyIJKAQpHiV7ReZTmI+xMp8H1DIIB5Qyh7bSfT
HaEa7eRUnOrRS68Rmdqfz0+9sSkiCrmItbCgnt+xdHidKe7WpN+JCPBtoIv7ChCpAtxoiqxaC5Ve
GDre5KAvfHJKEkVI22vt7HNAJEgqO1cAG58z/FthEe9In3JCFFjt986r9sSePIWoaR72Zq3Y1oy/
+LhwrTX2LweIqItBGOHxRbHVzo60LNEGxjRXOlCdSzmZbzgo7Cp/d+xnLFnIzzGgk+Pb0Ayo+Onl
V4WjIYrxreV81RXrgIVmPmI0lsD4iS+7QOm6AzDLpSL+lxdv8W7S0jqMp/LE3WgJi3DCQK7rp3iR
JieYp1X7eYpt82YUxbncw666DAq/sadmsBMFQzUi6e6nwIxCu3RgP8wMLlPM+r3Fmtk2QVo38Jrs
c+glBK627s1KJdiPSDALGNRCuuPp/DRBWg/ATxEeCHCzq/Lsqn5q7H1x/Xo93atGxwK684gRBgCA
WhEjpGIWWcdpC4xxOkYsoHff2D5TqTkBp8tkyKDnwvG/UPHX4FRdQSzRKFMR/5GafY7afLHEHC0B
0xdN8244yL9nQdA+S4GS4oPI5Lf92uLB6MroNou6MjjpnOoKckE5hD6EkId/PdRCj3qCzV3RG/OD
OrBKk6FC4SgB2EUBNVu8uR8fswCkDsidTUKZRor7XvxQIHuw4c1BDaQWR7lKi1YWiQkzJAeoSBZX
KeN9hFK+kscpvvb8DknWyK0eD+Qy0qsdakpJ0cWJX+etLjMBJo1sUMzP2LfGJA27S7dw4MJVLXDQ
mgtP04eHlV/TFJdeCFHcNuGhzrZXJhZy6GkQamltocH48XhacEzMidd8D1nH+NwiX/rXkfvg99Bn
Cd+gPRZfjDNegfgDtpXtosquep/0vMToy1J8VmKEfQILBUTyNSSE2Z3PopNvEl/wg94C8k87jG/d
pOypQhGTTtwsX2bCr3E7XhZOKCMpsNu9gtMQ0jngXYzEjHGUE8V5qeOhXzQEXghjGbhsJAEZmQIw
kabiuPeTonDxuOySiY0YxH+W/WZvZQW4k4dPBm9TenhTU+52FR2cF0q5Q3cH+qYvvYqLrjS3SExZ
01ipgPYPJ7gJfPGXbsymhyNMg7Ax7eEVLxC6uw9TopqkM5+bRTh5DlCcvgeDf1G3eZWL3V6ridt1
usV6OOexZD4iA0AXWFoNtF06s53jc3SzTpSu0P/fmQ6sDb5zNj1WXJfWSyICtLZ3Fq8bccOS6Jru
t2nUGr3V2VivrZ7Yn6ZFkV12psj+5U7D6EYhb7kD3PLHmbqCid1ok9yGzKwsiBEjCSqjQsiFLayT
t1Fibsy12iKT4p0F/oHtYvFGt0ceBj9yjvPtOhT6kzytwxkpcWii5iHoC6AFPcNvUGRZDKDDVv7Y
8+Rn4Gq6rEhBrQpvsA6llsJTVdbNk4KTFyJn7lVUFHWxTuq6/T4sMr04BgMlslGHx0f+JIIbqaKl
JuaFr441TYfkd1J3RMDGzrYXmfDtfuBaL/bQgGnBF3lySPAE/JwAtqnFJuVlS3tl9JUl/yUYuIxY
dvnQc3v1sEE6H3pOA3lL4nqQENXR1ImOydnA+y5pYn1ZtwjV59sN+7n2uevSgpVKYeXkC7YpYcr0
lHPMCR8Oh6LHccPQv8xoo1MpI1kbZdy02eHgPhGjA0kJlC6GZmSuauzRHCH4K8fpt6hdFEKBO+Vg
9+2ptZeqS9R1LwtRA3L4/skMXgEOh2CN4Ik3Nj30aBuueuHTMBsPrRL96Hegp7YQ/iNzF3UrSV7q
9FgkTk65ZEHXZj1JDwA4nn7r85Vl/r6qYvW6S3djobu0IgkwIx5nhSbbHMHUNbuFwhOj5IlhmyP+
2WU94pW+Q5iwdAoeQS7oCoKco/6esmBqe2NziPtGaA1Vd3T6RJeh43ojYARroTtTvduW1Sa1ypyx
FkuTDDK1ODiQLCFOYDcQhRU89S7kBWPwGECyxYpKKF2g/O2obPa3SGEHJ7oGZHOKVeR31xx1WNga
k2eFRg25bgoLnEexXgYd4JxZ1/fEwWIXzObrMj7hv3wYOgouBLe/nfw/EW8G3BlxUUUhD5JmUL11
LlR0xvU48ArlfmYzL3d0ftTXnp6y3dUfWKBevOB0+A49nU3aR6lYl4VsqCyix/eC5pi3Jz+784N/
kX8SGsmBXZbhjAhJUm7UqH4bt2mopTsIYKPJ9mfO2dzQrH5qG68yk4nh1yz61oTcBwf7tr+Ayt2f
S7zOdZ2Z2W+hMaUs8lJJi4XInSfh7Sf07dyPEYXavRAy0Wtm39dNDrP7tDoDe2hgDxWRQ0uD9F9a
yEyjvPdyQGGw3GQo9DDXE64BSXd7U9qbSctWRPc5zL1bH0AM5m+uXso9KHQIykLCG1YIz3E3ZOMo
tDNmzqVQO40sPd0KqDvVDylCEO1sP7vBDeDhflfNsEwOLKrULnDvA2OdN0O2DN0RNEi39xkv4iCP
H0Uawh32RM7KwjuZZu6NSPTqdlcQg29tcHPVMe27SdC5GSFigrBF2QzAm7k2qVAt5BUFf2uSNKsJ
Fo/05LhHbM8ucLZjFAqyn8BXiLMViuMtG8WGy3KnTg3CRixrQ8NRgRemeyeYy6gt+XLhtkR5EMpR
eRYdul49kVoyELEPjGWFRHtau1RevawL7YlN05bt4kQ6AZ4zmzxniypZ+IwNF5H+x03lTAQaoWbF
oZQUiGR41VeptT98D7RzcII9xBd1qvFqvXTC8rzW9rCqJAdVOXX25aeTqoYtfLzgK3wnWYkaGYRe
zF6PPx+nk3GZh3RKxrTyUEsikhhrPI1OJqCeKlA1fjXnLOar6fRWUD9pW7ZG3o7+7yllh0eU/NzZ
CAT2r/VH+Lx8Orks908ersLO/GtoPPiYFsMT1hWlmu/PRDU126R4A9+tNLF3io7eQI+1KuwFKEpT
EuNx111MPItDLeLpeaT2RJKm3eOJXN7agPlg0LV3zO8rHzBnYpWXyMYlFpIq/yhge0HQ1N99zoRC
EtdhrxtGoszdzsj8R+2XiwzGtkbwCnMVj3Oxiy1ivfLQLdYAKgvRxfbdMq/Xj89/Apoz/txMNfJ6
+YgitYBss4i3xIWYZPtzVTpMrbd7yxG5uu6w0FGVQXwq09Or0KKFVusg62d6DRxs5qQifC9keS7I
Y9XYapO45WS+NQ3S4y2g+uHPpULHWIr1Ds8q3GkP/lkjV3kIOIRwKN22a7dXR8PCgot0uMFSp8y7
l4ZWxHZzUJY5Zm4BO31HOnDV8CqrzJriYT2sWU/zehV1NownvRky9SprrcQTvw9+f2cb7EcjeAai
hItcqmlvqP7TGHJqgU3bcjmTqQZJyJUgGuK6xPCN4grkQLtsHpggT7dN4Glc88MFozpj1+xPKrTD
nA6id328gQiYI1oa0rd8B3IASDcSZte1wL0vuhkOVwfr+8hIC7ETvjqlpDpGEa0hkeAjdu5GT2o8
1fES+slFlbDxfVETEZPrLPTXUH8yxFHaGkWnJ7h6uHymi33iOO9kEzc603gabdVBeB9Ryi5sFwAA
qpx8Qma5ZwANPBBrXiX3N0N1X1/r9ANuPKCjz5uaJdLshFrAk57XETNKhqGcH6ezKj4yRE4LAqkZ
kUp6ShUrvkvBn8MpyDLrgowF1H7sTC7hNDnSxwMNaUd0jwajYfkqXUjDZRFyPsvF+OHLFEOkn6ki
njBi8+4l8LDa75YX4Gc39WnKKkyHnPEXd45rs61uTLpRpg1b0dI8Ovrj48R13oe1M3CZ8EWR4kYI
KFBe1e3tNlHqc/81O4jqAdW5n/yWIkd2Axo2Wy4JGocB3+Tamrh23IO9JIocLdFfb8BSj6hAejYJ
pelsxNgYYqENaHFXERGZ52aL6JU/RuMbffJycP6/YSX5ObMmZi4VuJxV4A+IjYD5cJrgU2OTwpck
E9ACC7UgjGjOcgTVF8GcZnedYDftF66WkuYzaWBPSBIHAbVJqCz4VimYMDHaPanwSD6Fy5zDb/8l
f2XYxFfQkiO3DdVhpPRCkWbcLIITss6fwRwLriLyMO8zBqYA5xawVFDQSq3XxCveglyMpMnflrMh
kch52vJzwTCb1kR2jMssD/B4gwy7q3PvsCXrWsKMgVMm+X5qUqrRgg/0ZpfY8OuEnJ5xKGseQ+cI
ctH9PeHpGOYtAUn5Ps1AZpzXh4vgeYwM2ueU+3Fmr7DYUZDSv1/zD4dzGHJCM6g9WelCOihUqDiN
n3UIwfnE49xCe9CQ6TfewJZYIVQzLFTWa9Y6YU+3HAHJvwt1TXvR4IReSObgQk5kq+1Gga7VcwJF
LC2fiB3ISCdbq6rIiXol2AzvQN1bWxPrFNy4YUdTe+Fg0J9tYAwI1+v0cP4aBK+1hMsK+Ve64nsT
xeq9u1lnwBO6bk8UujBw582wz+GE9P0Jg1Ivz/L52k/WktmBn2vjj3ZsCAwETfZKsGJnhO57B1YK
vKjdjvqRTOC4GA6Qa3FogCSKp/I18Vm9oupESsoby9Umh5IGlmuDCamZdN+w/MCbA3GtdTQYEPYE
qDqtXPo8hEtc9Nb5XH24X7KTkSxTANXUCqPzSmMqygRvKuHy/QVBi49tTAGu2qDjvOGUBQD3n75A
tsLKdBwREiri8uyl1CgBR6iSpZ/yB+1iV5ZQ8OKBIWqfu+kYZU1zCvuYmm4rCC3JGxuCCG3cUG/h
Qteoe82hQ2VBzKg6PBWDgyZzgJzae2E+5DVjTCWhWumoo+2yULtvTZ/cZih8gMmSJtRFvFfG0LxP
ZFrj8jK9WA11y8VVbsjf+oBdfJ5xkm9rPNamgQoLlw/oxJ75z5a7JMnk592luoQ4yJ+3yxEYaY8j
Qvex/YRQ6EOgxk7mcQRCLRrbxBNr+Tw0i5Wrw6TkQ2Pk1oZxPsZNSFhFcJtaq8Sa45HvBpj/47Ny
XjECluaCepAuHJgvAz1Byd5mrDAdBFKmKCS74UjABeQBS2g9uHhpNWLbpmp5TofNVd2+4eaog6zX
q/EKrPPsaEF7Ujm5PBwxi1CbxpuvW2Kusd13eUPMI6UGenO9LxVsAYXlRD0srvA4qarxdN91uoA2
IpfZBXcJs2R9wgTjXg0nvVFNKUdsoJsLGYK9DeWdPkwP/oKuMb+zKmmpwYjMpOyTj7xxB0gLBDa8
EvUM6KUY1FEQlkWsIdwpucjv4u/9t+HdqHeGXhdq2ij58lF6HhddEuuQTZEvJk0Md5hmjD6tkxUg
mCSqvg3OKt+KYWstrU+812bcUCQJsFymGrLiOJzMdmc9m3HaPYerbDRuua7ZxD4pO4NLgYoAYOvR
+N12ecorB046wQ4Py/A1rTVLRW7tmlNo5B1K/Q+Lcc0HuneJXQaQJQTeNgoF+LHZNxhFwXNM6yur
n4lxCr6MR/lORWiBkmR80LFe16AnoGBfYnSoCEeFK6A9mr5NIxdvwczCggjITf9GYVn2BdlYlXq7
HXpSDGOwI2/vQf2WXYNRhYPoD4revGDRC8Bb9fzLom0Oy0WHu1nSixWPwXsxyi1IOiXV6zx1Zmru
3WLGfdiHRMEQfmA5vRKG4P/UyZeUsF5eYnSPMN0MPEaquH8qtPtVzLwET6pHMyA2dvnlx6BOekw1
E1Yg53vcmimgK8LauW4x+52HdeaE5Oa2RmNd/vQ3YoRE6Pf6PQek4oEgjKzFCxnAzhzl9HXvGDym
Ax226vIL6i4fawoTpsj9gCM1HWGNjZc8lDH4hRzr/AHgYujPz/fTF3M4r1/WPa29lRWRcb8jzmFj
OfeB9iSgWDBw0sP4s/yxwS3QYP0PtPGMc10ij6p+9NcF6pUkf0UFCbveaBH5vLkz73Y/+csN/fe5
oGbrhFi0R6+Hb08ftgxLVv2T11Eq01vv9NVp7Vre0unmuRd+KhHY2FzhAHsoGW6Wex1cUqiAo6f0
c+dw2R7igwd7SOut6DIkdUQV/ktkfgfiW+2wgiuXDHq/irvZmFqtjijPSYrRCuGHZ7Q26Dr1Fb/h
ApbIUxEqVqdANPILVyUJzGx9sZXO+1g94m2XC8ulzkZ187EBMNGXaGA/BVD7aUn6KC6vdBrt2iFG
Zb1jlZQxv/QfqRWgksKtKbW/UEAAwvyJyiZ/iumANEnPr9l34/UjXSZvUhJz2ijx2EL2mv9iHeNs
/c5PsDc9A1rXWnnXb2IhAQxFhXfZecSMeEPuLmHhLhzZp9XoLppLgY9xOJnv0ThEWAq3msJonY69
7GBi89T9qUjp7u7poYFzgX8hGGd2ZTnAu/pQDgcxt3zC494sMX+tSny2DoYQRyBcsc8rJdX0gK6Y
lwXOAk5448bTyJvOA09UK/GhzL18bXvJJqwBL0a9O7eQrgQ/vfkELnQREVKdfNG0V9/cF4rbyHIL
tSU4NMZ4z+xkoS5OQy62KsOp1M2rv9fL0kNtBB+01mS6aqjKNSYpZjuCjYXvqwRwYjPGL8GRdIkj
GzH1SY58H9tB5CDmPHPcF1k91fGDhWn24NytfAS5n/DgLx+zZHiaYjz7I5p5YaYPC++elym6lOWc
LJf6LcNu7OEaEb60jQI9vGNy/cONF2kjEELz7LFJdmTtz6J121spcFwxbUbtiJUvT07elnvBxQUH
x4Ctt9CPBQUz92EUPboRtaXBZS81MlRtuDTfZdUpvPFh7SGOExrTAlTOVpZ5HcyIwu7X70YIlTCY
deoix+i8xPsn9k+Eg1vHx5YV/GZCEcBGwIjUWgWGKdK/WubKqgA5KhsHqaFL6AFv1e2jEEMm0/3T
ttKrPa3+anH/WqER1Qjm93Caa4sA5KUv+8hmnfew6LAlzTkNC7gPHWUUcrMpCEXg/vLK58HXJgfe
OpXDqp2pbKc0AwDgS0K9TuOVgeJZ0FYz74R/xQ+6FTYNfDvi0C8yX0xhbbVKDCp7f4oydWi3QTh8
9EyKJFCagEqzgcxSWD3/gs5Z10i45IbA7MmWia+W6nr5aw/88QfinxVmXDQ4cew/bczG6FwuMK6B
CJ5zO/LJE3IvoQvhGGtBvTjh0wCbDl/I8+m3yW6baQAJSK0mY8KU8y5b4Riwq4ugtJ4daVwFhhyR
7+LJ1tnKKwOpg+UEgYgCs0WaslEpQcJ/RQN38GKLg3A3ZcJTdMWptRtNd350C0THZm53ojsRLYnk
pY3aSx0a9Tq1dI9FJhB99kSO7ifLlihnfKh+ecqsTSdBX8Mt0LSBa9Vy6VoElMynNTuZ+TfWuBCi
8zqDyyubzWqO0802zRUddkWbL6RM0brLS/QJdM0OuGB3bd9E8E0i4wdQpNuwUbTgmVqSfJ0+roRy
HDAnMs1WY67FRbY3inrwGguOSuu7/2ByO8KHSdNWZUIU+6VVktSYotEINyCUsXaoPO+XmoNRbZ0x
EA197laSU+S5ayrc6dFkl/01OHdIDI4Lv+3M/E6cWE0yztXGOWVE4GiQFhRxR7/8Bjt1Q7i8QE2z
fe9F2g/hFwjnPtpUcUzEPsvRyaZ9kkRz+4O0gK8gRmoYHxZhzFVVOVMwX60QUUb6LDjofCUsdVH7
LC8I4ev6Qln823Q803OckEl+Gr4rmhwy3AcpOEbKkRGmiWaLv3C73O3QwM0z1pATqSAWUgcIdG+N
FuDeyTl9bgM1gc2bbltHJfrHByVbeBso0+bzMkxeyfWahB5CZ5ozhTz3XiUh9lz3dKCjrGZ6QQ8h
qc9K0j1XSeWWDLGwSqgKUu8U++j01Sm5efe4MdwaVUW7N63a+cCltDVdci8I+0KVy5Ag2uSzaV1i
212d7RQ3w5eSE0ZSqF6hzNW8hHBmBbqhzKMo3fGW4q8WskmVeyIL13iCtgftRoY1d2o2k5iRroDm
FGVxv7t2ftvOxHhdY297D2y3e17x0XC69Y2Q5BPqDScYGx7DdMH1q9F/6yR69tcE6naGt3fx8bh9
33mmqvYbpTdA0/z6iQAheOE8L0uHCOM8JAJATUPKmOaaaMks6FS9FfxiEkw+Z3H8gxWTf2+n1mwK
iMiY2pnm7xN4iBS6AvWecu6ebQlhPbc7bK3+TDR+bNllFwaWHI4sncx4+PK6ZQH4cs8khITvtMNk
j80TSwcAdjlTdofbgLTfdCCD6LPayzpE9X1cIDNJ29NSNjnuM/DwXqcZOuc1Z9wFiYiufjzbmmlT
S58M/CbOPGx1jxLLL3XceEzu9V10nXUztp0cJxb44tYDrI9UIwn88QapuEx4VG8+y4Zxq/rLjewc
zamsh3WUV2Y1y3YxgjO3e1y1FtcDHUCZtgJU86DjaG8Mk6rA6gcoVVCYWaIuUhzRxCKAQGCKO2/4
j6VerPp930pQGUuSILPNlk4loRIRO2VGBfhPSh/HUcFru0uO5lf8Wc1br/8CsJf+IvWjx3rHwVBx
gvEfS0eIsGHbbGjV1rLQ5gUTjZUHFr63TB6tNcYmIMQw33pH9KjN/5p7/rwHQg6UZhU8EwYuUWkU
YB6MEmfxySOhm802vqkzgETPvFylEZOjcFslJv9LxETtO325k1dUelwxI68Nc2B0GzCoaPs1Njvf
bQWMTIQbgCQ43bU0QftHej5a9zjTRkklmRtb86DSDNoHrssnr6U6a/w809Dw+wIHPM7osti1G88k
N50ECFwBNJ0IDV8f9dZp1dWvL4SIL1lIpR9f923x2uxRstwk+McQdBQ1V8Rip1M14IW/SJ7Gd4vB
t7C2RjNx0S1R14+aRxSP2GWaaxEBu+V+WJvzei5ak3mIpl0Os6GdQ5NBhTvjf3SMJuzzJyTfQ2V/
XlRJ/bbDE2tr++qYgVLV64nL/+OHubeGIwDBZCSSNqeyYgl4C0gY05oZbvNmxLkOOZHif4K2mFy4
hm3T09UDuqvtykPWPEeisiW/X7xvjvdv8fHCqaBJeSGnWoYFak56v1C8K5jdvvcU/XxxtIIg8sZK
u6xX6HK0aUbtBk2xFYhXDxbzahE3nHwEIzU02QFd5tnGKnYUJ+VT0v0z7TpOApLa4nW+AjWDhsCI
lN9Nucf0QS9Zp7z47dcer2+4dVA3TDkA3RpCB1CQh4GoxQTOJmCXMno0j5bkmW88JY0xeaGcTDsf
V8euCUtR21A7xlSjCninx8FXhKi4jgRd70gnj0QFXhEoF++FBTwQP2pNa5Zdze3OcDhX0BU//QaN
75jpXTJ/y8fML1ky7xTIlNqTwH74zrcll5zsFzQ+dKDk6LIJceDwRs0tzXlg+T4q6cClfqKj8MVP
i+xRDmS3D87WRbM2WxOtmkoxgTVt0XoDXogqKUVL1CWPPNVqR968BMJSwX0CCkE6TzNK/2yMNZji
dyzP9t4i44Ss8IF9bKfzUlizyrr/gXT/382y9TESo3qirEgp2S9KSAhmmxz3tftGrBlVfeyDJHpR
6hnwVoV+eLszcnpfIY5AJUITcB1cnonvOyA6ZjkHV5yLGhQIjCX+HArznIEuTZJLkt6pP44iAVtp
7XQ0FMixKuLFgj8rD6ghaTW+132UFcHQaOnVEvuGkds6FA+YnIILCppBXALdmK1pFzO6IePJBga0
HAcLd5NeGy3zdYGUOHTIeLPPzim3jyITgnk+zoExTKDdFft3onx2OzguAW4HA63iGoYk0mXa2TXw
QDMAMKO2ON582y0FVxKO1smr9ZGf/MfiJxwyvZbB/qDniNVxM5DVfZT5d2SfvAe+WixOykkeWqaS
JpWFwN0XKjPGz3PA2+tCSMO2S+EPvtP1lYt2kPZjI5hDRxo81xQIslyPg3CU3UmTVhyLGHmqH200
e3hs8z6QzaZpSfqt0mzHPEVDHsCrAvhRKnIXpL/+jMue/RCX591pSYUpthiouskerkj+mH5pN7+S
iSbUg4yZ1lFvSO3COV0rvFnvZoybMomhHjfJk+beTs0ACj3E2+TpBLDgpqXleBzvX+T9pEC6MKCr
z9R2H5+zs2r/SQJy1egEmfwEj6rdNCh4Y9wevAyrow5f6KYtxTtBUuErV27q6jfagt3SFS3LOSVX
JmnURpBqdw0qISF/6KzmK2kUfU5IRaqWNSQRudkZJGEOTOQALpxvrf8JpPr/OtUNbA/LOmPYoxHl
y9N+00aBwCInba7HGWyS4/ZxSVjZoSbJ/aGHWZVuObCEh7IzGCeW1Z2I6AZnxKGuz0KVO4+nlKEr
KDj/8aUioyLrMj2jI9gJ5KtU1g0MA+wKTv+Epuyaicab+CmFjNqQpwWEW4iaQ7Iny9kHB50z71cX
//zD5J/xhWwLYSn/fwDQQfkj0b7+8iv0Tjshgu+GCSGxP4uCI00EOfMtrNstdWOnZZdv3zNhAeHv
ejr7Zb0+0QWuhSV2tvHdMHXMMZw0F9tsp/62r+66hXQ3JbIFkV2ZwjDQ89GMcLqcdw1qBk4Vo7l8
16w6GBjltwCrT3R9vq9VK8NuBJHAgSmvP6INfF/KHX/oap1vVxRx8TFykxZS1yiJWZcbmwdlbvMj
T79Hlm03DbLXDFI2L2XAsq6Vvp4+miml/QqtPvAHW7TPfAWnhetWUkyk4pk7XPq6UZEE5zU4JIRE
4c1m6QcRcMRQAvUmEbzWDyttAn4MERcwNOGCDCzy19sUM4/wRAIJIJ2vqBAniroxIB8rc0t6qsQk
ET59sufQ6CjSJFW3x72fc6BF6MCgy6fp5kU9omGgIirtv3SOTdI/oThx5JTm0abXiK4a5JF+Vw2k
UV6J3xeGGYPH+kycoEdAuJmVb56W2pBKaG8xRaH+pUUvSG0DHWfc+mGjruHUizhyordQssTdgQnY
Se8Vm/PifJcXeZubRF2AU3zCVPYrjdaYSG9rysPV/2pixEnFLfrRAqVF2P8toPmuRvUrLGiCb7Dv
uJuxq9LA72PIbn75BlF45M4wVflEW52E0HDS67N+Id9Pj0cnIW3lS6dzA0iOj9SLSqkPJ+a1cLd9
F3lcJU7h3U6wCEHJepqYv/ubGQQC/77kNcIJzISRxZ/q/zVtEa9NiFo0fDsLs6HKQiQ492q5RWmw
P25uL1UvHZ0g3800ZpIEC8OMtBzKkhUNylrmC4SZSMs0fE5LAsacMzJgqM1H870ClXuu2XBnRI79
ZUVvi4KtiVkXrgYGIEjFkgCvW2Flr7zwVi+Qu/yysgCqk0g9AzD6PNzk0VZ/fERKaUskCqUIbIJo
Wlg25/br1tiJkq8t6nNSZUrsdJ+SGmH1y22GXJRrs+zzBJ1doiUxRzo5zyXG2X3dIUQceMCVvviw
oWl1fWlre0syr1rfN7vnneccMzrXgUILzkqY8TLS/AIsLcl/Hp/pUwOgHhSyk+0rhZnPoxpSRpms
PD1FvpKlYks7KxpoXN7mqkeHAjK/3Rh4Yeaw5CrtPPntiK8URe8PM2mleQLHwElXhCexU/US4nA7
Qv1uuw0ca8c1UwSBskoiRKqVvidvIUC3a2ojQCLCBjKScd9aymOmqJ9UOZYTlJCFpobkBBpsZRa8
/M8S26kXQcE3p2zZVdD+78deKwDEtromSNqnpJN2gg/YjEG0QTgt/tmuA0+M82W1vaduWmKEXLtR
NP46Xdq8DMjDeFpvFRJNJWkZOtHWHifZKayAJZoKo1k55ykLAbaD4CZVr9Ywmuawp6pdnT6hEqXe
ASoSykojKQpbKCBLGo6kTj9WaA2pTUG2I3jzXPldEwvVXRk8dIGZKWQmxjXQpprCHO9BJ9eBtTBt
6vm0mU2b3e8db4MwM217AjTTxFN7mu8gah+o6HYw7mUsiCuz+KbtY7ch1//4oIWKB2VhcwCdJl2l
SpgR9oqX4vm+Eu8dArzKcYtghRbdGA9Du7yA8NDY2X5gQ1bpe0fux/FkEvNtHm+eXrIGzVgraeDL
rH65N4W/m9I1W/hqCTn8OJ9d70BIAfsXSqii1lKgtV9uVwNwXbDuZjj81wt9ynEpTHos0R+D+HKc
2Uh5I7fYR3AXqAXTpulNuzVZxm+Ap1CtHAeD4HuOz/FUM21EX7kipH683Iwm7St2DazUImZZEjPZ
KXuaRaXQeQhnPAYVYA50i2IhdFCDq0moXUPwWX2c2rxv+UQ1EtaMPCMJdUTC94P6zTqsCAc3pQxe
ARx2ocqBw/TrRWVprNFOGCDpuMJmISyV+dJ4V3mfv/P2vQtYKatHiYYqPMl1+dVN5nmc+rUrZl2P
biPdSOlbgBqS0YgdeoqG1Z/R2dcpYRbhnOoHOE8T0hspSDzNB7wmMfbWIpXhBCAfI4jdgSpJiBCN
2W836lJmTfdTX9sT2pmQicjdwggWNxuPfpCvmg9aWyQPdIatkS3X+00TuOsFb/hSNJVc8f38LDmq
SrjvhVDRkv/aRzAMPbIt9G89JXgN8cl3nOWS1KlXCg/f1dWpC4sMNaX78RqNSjocHX7GlKJOhnGQ
/nJ1ZBdIUXNtilH5DGalAkc5c7FwqGJFAiwr4fOIIMq3Jiq2/RdMiBMLzDVPjowYKMkCwfvWBHRb
I8ZYvdrsKmZcdXPWXyBnBC0t9z/ONdCYakWW27tNhYqlnyFKYlNIkaHVxBRu6aYXS5MuVQ10hdMl
b/nVlWIv3ZnaaDFvYifklC0eVSJdwWYKxS17+YE6e/IH9YOFczYSbNvM11bLFNjCgynK7OrxxCIp
oj1+CcejUl48BUIdnWKvmyqMrhl8S4Mny2gRw8NZ41qyZ+N69Mi3UzEdZ7q3VSgqUVIwXSW0CLU7
gzSWhIH9NCqaMVhV+8cH4AZ8xnsXStUXil+TA5DZEJabewLKMkMfvD9XAdWQnYO1/u8K+FmQ7g0V
RmoXjXGr/g+iSpzqyjYL58ExgMqdyYV56A5SsIhyUmWS2mFXA3XGr/ztI3DXIww5Siy9hdcS4/sr
ih1fdwVkFo1nnKqLfGO2CXLAaMV1SH0YXEE3Q9snSIFazny//fVO8YsI7wgFJeWpknM5KBlopoNG
88mqfAsxt4NqrayUIEgb2ZAQw89as9voKT5ewcB738YgukXOhx/uTJguhC0WXIyMCbx5gutI5MIy
ZMw1T26LQMPb3NaS8kGBOqT0TCaNH7q4ykb+QZ2GgCNf6So4LfED/VXpTAGzODB05Gy1DQsWHo/C
U6CDwwNbZ32DvBQOQ8lStxbso8Q1SfpQhJ1H5IIuOQ3rx9XS17zb7J5w7Ffru4E2c9QW2hyoyhkL
iEJq8yayctxeu+2ssvBBlH1kp1m4sq4h4ICKdMnZar5Fa9T9c6RqgKvW/ZmKBlzm/bxX9GsEgV+8
t5zzq+IFlQyU/I1SBBtGZ3YBcC55bAcL2/jSnazSyvKodpaJYtjdeIo9UFR734Y97Bp74aZru2ES
vEa7/UPdwHuIsFaDcSezJkdSvXg+EVPfzvhpu5xWLZWnoXmLYugKEagpIgnfUgZXJmtOwZvse834
tuPX896diE5w8xCOzyXsnRwPtEDI1KZtjkDuQ97Wqs8hEpj/lw1Udw8ES5FpNzpNJQIn4Q296gXq
7oKD/732F08LlLVajmuHeEfUE5j161qyb09MTLbS/gURAG04Tmp2WxIwPFkB7xWPCOzm33aaH/ov
i5l3T7EFL+iR4zvh1aYyO+KBNMVptBTuaZip6ai32JGUggOe6n8KzEwK7BoVFnFo89hxulHra/eC
U3GCA4hoUEMojgFy3KViGZY1RWBz0eLSzdRB4tIj1/fe9xJmVTJEWxRnE00+cAyHeIuTsyw8ezSZ
pWaufsF9nyY3GpQmCIrj9Pg6OBgbgleN/1vee50N1p9qW4sY4hX+DDT3ByRIG7QrW5Oobzprn5Xd
AVfjj8tpzVn6BLLEroxVcj2hXyPOAgCplCqDdj5FzB5B1ckXQ/0pxGiWStURfuVm1DSnNMimqW3j
kgGkzNsBqRUtMqA+Vib8/VhM+m7pg625X209CTylNVaNBuEiM6jRzaq2YLGTieDIzuSzWJRPZvDU
Gdi3xs6PK7nj6gPXH2hlFzUcS2xk0Q7wjExuLrnX9fg46ijUhJUxX890ZOZ7PGKN7AEmbCegpqN3
yMdhXZZj/bO4JodzN/iFbPbe8xpSUH4VydI9zhN+xP5eZoGYhlziXVQTAHbTZ9QDKa/b3ng/jqJX
MRErQMG/TQmo46VvPNqwggEqizVHsN4/4XZUk2fnQHhrlgWyAtE+8u7HFtqd28OjIvYEyOuQOrlw
tEuL5Ga+F4zPRKljXEWiXxIyGsrOgk946at3+b/htoV0RyeMogO6bgy+z0XFyNPWqEToAgxGqUpB
NsyhOySvhpLVbKo9MGLjiEe6X98BSDXi+uc4YJPncx/50LYVizekrfwQj339b2eq43l8wMe+ntPt
5Usm/Lwrvn6lVV6cXv2m5kIIBc8/MF06Rp0XBN8KH5/fON+wku1JkNGsToDo2FfuwKLXt3gofJRz
68PSQbjXLeix6pw3v9wTq0y8IsMXbFbtkJhQtegAsT0MGpzQVygmYbeN6nciWn9lGRLW3dC+IWPZ
h7VBtwP+2BCq5bZ3YvFuzNHdvFQ0BQqayH0mBuS6cVQMYImTith67bTgGpUHslgcZE4qV7H3DbqG
SwYcmU+eP4W2V7lLXcIKh2nAiEHYxjPdHajKJR5cfvdfeiuxBq5oSwGcznSiaK64im82tFU0YmF9
k+U4wRV/Tz1u2Z09CoE3PYued1AQpVhL3Uy6cY2zqtRR/6UV2V3jAwzTMRjfmHZkkuoOmOUAvBS4
M83CpC0Kug3IUKDXaSudHFRolVIhhHsMLDjz9A3ne2HJanxKAmCTghkpOXt4PoLIB5wXV4oURqTU
JnijLA7kx2e+X/MiOnyLLqhdk/TRhSf/cGM65xn+ire/UyFpg++ZXufNZTmE8X4r/b+PTATs/tAI
lrjqEs7ReZpS7GbDJu4fbjVO6Q5xXBRFLSxW5aGxnq5+zE+cAxqXMLLokBFcFpFk/hUrPUUqEDnH
1EW6duEUx+fuJ3pTYlPq0PWxQL2CoJjkO9QaQtpXs3FVaEtDSg8hpr/NZrmQMz78FRaapZDC5AAp
GD9L6QtORWRMjA8dXVjoehyqUFleQtYN5kV+UuQOhHrPj7JwrL0o+mqSWCrs5gjBm4Szmr/HKW0g
HnqAd9wolgRs0UQU4bbJPZ88zxmxuloRMmxX+dKdY/CCfL4C/63+pGkp3KNZ/NGBvke9gxQuSmd8
VlbQIW4ZNkqov3r9XolrZrljz2AUfwSYz0nkdWEU7NEY5mWQjJXMQM4tbX0IK7yGz7q7jZl3AU02
K95fQ9zXI9w21/Jg9ZEqgKYF8lqRcj9DQ4ly/vGJ5uXZOCxCg5mMLpJuqkCxXZ+qfOORW4siv1ug
as1tswnRpZYqmw8/A28bvs5SHZ7F3fdIgqp0440POa8lZUJK95fX42pV8MThUz2g9vWyw319qYG6
sLmHRE+gLus1Uok3sQwFNR8AVus5BwtlVr2JSzhYqWwfT/kXepAI72fu8fAN1g1lpPvyHM53uRIy
6u06IAjqlgi9SWdBVvU3I5XjPmhgIVWaL2UQFKAkCp9i90oZQGPmxKt9mDLf+GWE54bAEqd9TPC5
8qB7ct/swb+BL2io48NI6i9VCP4bMG9SarBJd+m8HJ8k+OFfe34cqHXAt3GrquJbAwPkpO6gGplW
PSw3PMCUiyppiofkQ4qvdSYh1qhOpt5+Ln6R0oAvKuVUlqRHOPXpZP+JkmU78E3aZNQWrltwU3cG
5JomiTU5nTZeD/n//URRP1LTeWm3Nlv1WwS9A7RQOofnVqA0OcKvOaT7KfhgfVr6A+A/wlQ2oEob
2uM6cMG1QVFoM/bji4VLF/bfU8PwKJzqaSaWsrYcPLHCgGqEmPyh21oe+z6lgw11WPLuAabkV62j
CXRzt7KV7RzCP7zGUeZvaVRgN1ae4AG4WJ4q5WBSHcctEZX74E0qnhyR2aWF5KhCyIIvbpOpRi3M
cWANEa/pkSnSqPccx63vQf/hPBUuyVAn5kqS3gBYDYaPsP7rBrr/3iUoTp32eqvyD5BJQF6EZ8Pz
o7ilQ4cETrltqxovIeHuIa8Tb0y5D69PQYmPaydqykxxNxv9hWZuOoyM0u9sPBZ+s8sPeplvi4af
xeyGC2OKn93eouH7VKGsgVI0Uy1bYhdRsUIsnBXBDPHWWDtvUBUO+0qMAeeLT1zPqbCmPFjEm7bJ
yKaAcbCcPwX59s/8DMJpQTHst8pcRQLVqL9HTx3038fl29PwfVszlC3EPF1RVlODb0KilLwbMyD8
MKozc3mxVpr+cXopgjoILvOB8prtl9IJgxSh4cnFKtxTPmjTXjXdjHjbPBhGVmHo341KYiu/NSeH
kTiD/JyXqDFe7oE4R8WxEXQz44Rjl7LrJMtjea4CROZgxh7AZrPeEGlL9l9Qs9EweiL6YME7S0kv
yfBtR4qqXNcQ9cviycIgNEzCcbNF+N/8elrQi97dRyp2tLlYcaia4Cz7kykrQAK98Aa3GBoPq6Hz
qJa8YHUjJxYTfhlV+6PJ4rjjCKF5az2bqK27rNxbuCady6IjizmgaE92PXbLrkmVbtI4noSGXn5m
VqxM6CpBIwcKDBE+pmHd/mS9JLHa/UPQTCTk76fnoEK4F/J5SUJyZS1moyBRAU2i7/bxVrhqxBYx
MLAZjKZqJnWlg8hyZ8GzjwedeDlMqiVCBjbXIj+jSMi2gyu8JlizsXGnC6ru317tjlpBxTvpyf1l
vfS/Xo8AGLmT6kCBq5sPZdk8QQpnE/b2woUk/LwOuiPOYkMUCuW0V2XUCLc5hkCp9Njbsfb3IpSH
qKdLKhxcmciCm+6I69T/6K8GxoUMZ0mpfpnPEP/fg8xVo23Ba6zz2QbLtwbpl28T7UaSZt1nOnpL
SwTMdQm3ijIOuA/7RRrLASaTbW5cfwUjIB2A7OrR3xYgo9daHKGBd9ZH5BVt1T18rifE2U0PxsQ/
J66x99Tf4TEQPOHbUJcDN9dEyy+SLs+PgMSt0g8rH3W4TJiL2BGhAgtSmDXOUSa61oXHdNyrkRv4
81C31gvk08r7Z8qWvnbGjO0n2V5MnX2/f2yHy4UQ6x9gKa5Q6toajXAKQFS5zrGhhqnsVa8wKS42
oZES3HATGpaT4ISz029olkSiWXCGqY6IYfxgP61DJvhZf2Wf03TqMgXdlreNfdTCCFJxQIhlBCGL
vqgBUHX6iNY+IsmW7JLnTTze6TbtpyxzY2DFiZX3NOVsDOHU4XxklQy1Xe4CO1sSdnnUaAi8+2iN
XYceMg6JRwGtZkJXoJRy+sxvpx2LVk63eEJDMPZUh/dCEgbbynaqUkTqwswD8UXWm5YrVdsVULz7
nfcEGMza/M9YT3NMBUpQzRv4z/vJkf7wKeukODx3phdXz+2q8rwL4jJzZorXMe/lTQh+h5ywFGos
OD8bGpVvE5E4/zRhCNtV+EMxAUz7tzyuQ0h5HWxB5lrPw+uBKkBb/xm5uOUKkYYLKvHn4Ei19egX
4IhBz8P4KbSliZ0lKumDI8Zhh4HW+OOL3qUjFre5vuMlde3ItW6egLByEjgqNLDyeAyFp6SN7QY3
KNdbQ8L7m2jOj3+xCBhiArO0fzwXDHgBEqK27DivpGgGUaGA3gYk+mTAj8NoHDAl8RlshSjEHobK
lSvTyjFPYuJ5Wfbp4cXJXGkdHL/aTlhLUabBgp41IvD4piGP9Rort4hMfk0+DL9cW9Bwpt+iMvjs
rdXca3wTihvP3gJ1NECNFQjmR8cU0poGs8zbOvc0x56eX4RInd64J/0vkq3J+yENu9U78NF2aQu2
xLTHXnYRzCD8x+6kkdWVkfE0agJsnCkABpy5SiKsHx2KiG6ZqpNZqFZ3prBwJo+CyrTIBxDuDOab
KDaD905zbOb3ubHhN4QknYOAkjCYTIUl3c1xfjuLXGY76HAXPHXoUnyPLwrynFCdWUGSsxlIp9p0
bhSgHkVI4ceOMk89KdmBx2mpWMWiVJYH2gxqKasFUCzogFYN0gWRvoco4wBIpyg8C7Z6av8kShLh
eB8mJbCqny+k6xmwGML9bXllTePMnbUCrw1ghXD8WvfTuFf1U2LoKS/S9lDze0USu0pFepUYexbE
mn5YotqIOjhVc+jz/xMNPwzlUJpAJk4LvAx+QBFxA+u9JqvRf7aFyaVWWLT5TSyJJvHenfftLQdR
pXgTZ8BUDcH48JrTXHZavQ9fpgWBtg60yUHuGPT7s6bx5iUWupUXt7tVhGgRBD8QCEkIjNzCDUbL
GvKEWcgeN3jKIm30qGTPCFMz2fYJRImUf6xPZxlyIZJNxPtvZtkE1fND6dCa2ut3zJAr+j+O5JMZ
21Ha1HNJU4UJKX4NfAk7KoZ2hloBXf7KQpqsE+N5uKrJrmCir+iEi9jkbXwNu7OZIgi0JxDQqUrY
qNFbRBf0Bzh8RQQzHd4tL7wMy5FunXilG5fE7u/EDISgW8V5lj7Vunn8MZsbWfRspV7L5T4fbDXe
JDU9Q/o5p07mZ1SgFebda9L/K5UD0CZiL5Cdf3WV9hXVAvanXwxnpn5jOcVISYHohxGPJ9tOqY6q
zwkAu9y3miu2nc+jkd3uQUedMhU02RW0LvRB8cT0Q737Wj/0yn0b9h8DWerAKUwCNZkze3jqd4j4
KWfgsk4++36KHMuy24yd6zpRpRiZRhLbyvFemOnV1ThGdTEpWM2NdsLvjY3hZQjf8MIGJnXI5fHg
lQbzKvr/05MsY54GfKseF09cgVPy0vnwUT906uuoSvxXZ5sgZGuI/IypbXmEcjRLH/s9fBQiV3Tx
FqI88tWIHkpdZe5yCUqEMm8ILz7+/pe2toMykH3HebX8VD7IDnayNvaMTMZ4t6rLh/oMEbEjUb5V
CDkT+vu6iKdt3HwjTGtn/KqaIqhvENTn/+VqEHXEMc0qd6uUp10H6qjdVL3YNpVujGkaG1zsJDkB
ZODsHPvrVGGKws87ySnhae4Jwzi5DqRtj0GMEBgmRJKdPKu9CLvbXkBJeetCo62x50+jLJcXiHom
qZM2WO/Y0hGUYnPh8wGUuHJfibQptoG4uYQWZMOR5wns8M8fvvKd/UjUXoh3XyY2P9rOwZIXOqJ1
kCg1oVQIk/ZTrhEDfLlE8czRarnlsC5CE3rZ1id5fWMExRoDC9wxTKENu5kd5Vy2BKyMBHUweoaZ
Iwx7nO6f7eMjL+bf0k3mvCxgsbUtilWfoASJibNY2d43cLsnViVAHdGjoMbSJ8SRgjGv0PfEOHEV
yFJdIiIsKYyXm7/nAp1pSHFoUIREm2J5BgJ5o3OycTyKAl2pSY7A9tbw523PzhLs3BJA5bzfpn/E
kXa4rK3JvkNwfQWuFu9UzVBafqX5tCj1RZhcq1EBuJlp9E6lWvH+RF3S7qsxvaZ1C4IwFRaax2HD
IUaZNcl8dExCGPu4UuQsdmcCWI1gZC0VFl5+RKG25qRHyajNJmrnCokHwTaBavG95aW7+AmCjTaH
XlvqzUvj3uzUOdiTfFA+D1eCUDphab8dMWLmhr9hNqScF3UhGc5wL5wmMPP0JH11Al9inWXOnAww
apHx4FwN3Gmb3m7YYVSiCgyLbVhHvMNzo4FoOgFItvQ59/IeaithMulgEaDu0PcNeHiEbBiZ29gB
gXmwJVbkr3cJ+N9cf+mEBMJeH9DHF+BzBve7l465E29NV4AbhYTiD5SjbWU353V4vKQ8HWc9Ot7C
zTrlGAz2HqPM+FMQk+2qwvlwbmaAN6risEkoPUOtu4pOCQis7GtWSYcfXJdy4w/MNLaS43bku5wN
cMqy06qGZiEUiHoM7cyLmTNAUk/TBzmR7ShVELZUfSZ0g0DTNtMEkx53KeXV7IqYA/DKH5BliAHb
RW331Qi3Dhvj2/C3TWdYfm1vl9NkpssLw9AwQN9P3Mux8DqdWsvxKKrlD/eR3fHIhkTdLK5Z5pV1
Jg5hXLy/8d50P4dBGJqzx6JeLqIRqvVD3md1FRvVfpT7qt88QU2n0bcOhZCuhxQY+rVuXZ9McGTH
3PSxC8EGVHuIf/ty+A+KG+j6NIwgyMXANBzlFvsJp7WVwOkuyKwYWAKFzLjaeREwLYbiT4DaVCIi
b2Suc0rd9AQw7RDK5II5l2o9mgLt4O7VAodQbRRmwae4yN0G5bsskOg4XH4nw0h0vlxuoZBQFK1d
RUgrT1ZF+dEtMHP9KG2+rD7E4AqCAjlzN5NHzszXqIv9E3Kykar0Rhp0hiLsd/8y2DYocF7wDMc9
j8tli9/6mYpcWR2205medWYCj0aOMbMhxTpwqSWbPVYd+W0vB9SeZPKV0+1SR56B6I6z4flGAQ/l
b2ilWxg+JY4HJSl/Si0JHbuZHWpn+EwbbZLFC6p2IQ4/pKsoy8utJJuF0pLccdazQVqqbcjGeEk+
56CTrKfy5WmTh3q/HwVqg8dpd8v3q+b3Pq6MjSVVVESv3OOJZsRm/jImMYTeb6ny5V0aw7KnNwcV
M8uKj7s8MVWhhGsexZnMNUYp3l/Kni7brONsOPNdjxXowd878s925p2/MRBN14wkR+PkE1D6kpBY
8zX8pV1W8TjF97Tr6Mb2ifHPGzY68MIk2lDOQMGkrzqx55KDGVmJkiVDG20YiS8YyJFxjG9PDe+M
hdQMeM+E9dplTW3e0yz2+yPiVsmMZ4tuYpKlWW6fR/AuKMfZWlg3pymwaK0oiXEfYdw/FGDPHKMh
NLeqirI2bbb4Y9jX7Znf//msKjEW6Gs4RAUcQ+nFZT6Gi0RDQGQ8r7vPqEfGyXxH03tAhg2LRN2x
tbUqJ0uxEZpDpQEFdDjcvnka2pj3GvHcsbDIWVK59AxM8wswAkF80LhD8e2nssQZ0EEEizpsOwsx
0xLuKO7TdNEf0bs/DOoSGg13Vy0BGaTUEbc+hPUJXlr1Ek3MoX9rPVXTvLlgoGKY932wKaz6achN
Km6FrZ6NpqKd2pGJcM8s1oXwKdOgXesQ0Gspy0o7muEPyDqYvAblk29prSZ8v9Afklj1rqFtfBz5
uLqITAIcyzeVTYMjP3j/NbFOX5xepUt9ZyepPqbf5rHnwuIgf/vV/ZHLAsV5vGXNIOnA4FQeKhYt
vCdsB0pBAnsnQEnojUp8G0Fdq90B+96EmH3hFKrhbMOzRWwMZEizRm+Ov70HN1JB9nw8GgobFGQc
8jv2XNtOJZy5nwz3mS1JBf6TgkwOf/668r7GOrIWkIplppRSM2f1+zwYZjH3sN/aduV4IUGkjeDh
h3+vo+jpGYcyR2GrCJDqrxE/GSlm/9rnljgzHqN3o0nS9V8SxhnzucdXm2vUmbhU0psFHVYh5/Az
JgH0Kh/vMM9jpm9cFYBnsoBCjwzh9PNm0NdlNRq/bM2NMKUPPwAgicb2wRmEzwRee7accshHtgLM
LsEX3O3l2JQyeNK06zmkUF+09z/9Ui/d+LpVSfDaQiiwWWnHTg9XYq2sJDm+oHGjQltiySVFOU9U
nFqmBf3pTHPwqvZrsHk+eJP35Z1UB+PVU4BADr6eKQ3Km45Xwv+edJWNdSVeIJqd9ISLEa3PTrls
HSgl1Nh1+d2yyFtTtT4JTDIFmHKmQMFpcIhbaje3niFuG3KrnicKc2WG4cXnmDh0ABVFJX5RjKNc
8J8tHBlESwxT/7s+HUETRoOJfVwiK8ZmCdkCXU9KnuQL2PeDnAfdRKA7y20rgx9BqUfzzsvxR/a4
TPv30qGEFysCVwag+rKii/N/7SjijbkzOawJWjEzKPqiXWv5WanSKprJWQk5UykvDAwN41yAjnO1
6C/k7cSomOJNlc7wpWwIss7L1VWfZ7q3dUxeD9fcksOU4s+ITWUmEiv6VRUNpSv9IQV9wR9FPeUR
FT+BC4mUEIW+XWgbqbGyihbgCvfJd8ro4C3Wo8opfDCN/Dw8Ibz5yB8YhoaAziapDE6xlsCz8YhM
khIuRdbbXW3fnm/ZYeZP/eSpwRz5Bf+5mk9//OKQZe0ftYbh4Ys8qrYg+Kacq3B5RbzchVKiqTYR
I4jOGqgTRJoCCfmaWq9TwaCZMPhQ8O9KcTF8ypeyy3AJbA5eNBWnjLBGoofrlHv249VdtGMi6uMu
xm9rfTjRE8Mgz8kvmIubpVWxaEPE3XI0l7QdHS1ktkqzlQcxjbiDvJoNaLc5cJWiGj+m9eAQHnMV
zPI5yYMiJ3ka4NEhPvw7zsNDOmalEC3MJ59BrIyhLS/mXxqGx3YhsRFb8DgbyD+WosuSAYtFuQ43
t3tLM97zGjY5/Ujgsn80s/LVCaUxOhNoYTGlQPAQqBg9SzPGQhQkXmEt+3pBcz2FlankXOPtJeS/
57dX+v2I8JNKvUusgLoy3u2Ut4wtHTDweqjZ8PyfNIhLQu5wQpVior1Xy68JBcWeY6TGNIcUNPF1
tLaqSgTit/aOUxfn2czb3POenLUgQkKi/I7T4VABOqXR+wwBIEuZbQ103JUHpJNH2f5foOydVAuE
cHk+CxNkx6KnFdkrLlek/DwDdLTiwP1PAT5OWNASvRLj+Rpyeb0Ub4V+iXa4ViQ+t6EQAh4LhQQ7
KX8d0U7ZAzrqFT1Fds4xrFk7yjdCQdVQv122uzt64HIJkz7hdiUezf2h5g1RwkZc96DcIWBSsPy+
M3/7eu2ZsgQmPguQLPZ6nu6hAN9Bi3lmweuneNSFoU2s55vqvH5sQ0KKB+q48RPs4B6laukgqjoV
No+ELJoEkscip5H2TAUUfDUm6ecgsRNurvHxiwY1VoU6ISMQXBQ94P232voHjqGeAXVnj2wFXv2R
Bv9txL8jlqny0j8cYV9+G/ty8vdiMqhTlhc24N0YiB1uOKK+cRiaa5pSc1t9jYYbCZJQ+a4RTkyL
+I8MO3RrBPjnT17Glfk8CmG0FPINtkELQufJni8pAHj4v1GCe3hhi437R3eK0nnx3VgBLZ3CEfXN
7o9vGmPidgyHAhGvB/U9laBNUBby+7OZXTtt2S9TvsRcDz5vEneCgYgUU/drWjk/e3A6Sr3gRuYw
7mIbvGhm8vVgMcZOae/nn1cw3MXHT/lYYx6+b/9MNf1bvO9LsodzTKzGMFJ9v1xAEtgPOIkgh2l+
7bKdCGsERxskUYYuY0jj9gHUNEoGZK/HYQfhqr1W0GZurb9ruPlFH90kzHFi89cnZ/7R3PZcV0qj
vyQd2+9fLVy/VNGrO6P365X8ANYc4/d9D+czYA4AafS9berYQPLlzTZLa4jdGjklBnDt/OQ0pYxv
kqLMNih0A1t0TtUDfmeOzQwZg1UYgV4fYQ/BQhmtICRduR3qJYhcu/hDXfsX8LG/i3joZhLOglYV
nP41szXf9WoDrUwpHeBXltJ0UBzD1MKUFQf2aClyPPUnp78CRvx9GRIWWmPms5Pn+0KyOIhhLP1q
a9VY3Lspwxelu05v64NGyz3C19kMNsm87XQDa/0S4CLPfcXGQoXftRo8cBh1TV45x0jYfbBFO79Q
WveMCtziLvIwBNVY5sz/7vhsqgtNeWveoZlec/2ya4oQ7TELDuecr+L73frDb+/P7M5w9f00hFtA
rwkYUsj3hW23LAFj7ORcvXhuHCWnedKaA+snv4VEHbhg1ooqLfdEW1pgEppjUC6ZHZqZRU5QYEES
Z5r3KvfaxlGRNtJ5gtH5Ycrm1Z0f2HT9VqVQh8RGAj+6UquGV1dmcViO9VucBpq+IReD5Em9M3lp
gt29NEAJ1aL6UDXaNMpU632xlPVh1hmoibE1TFM1008tXVfEmPbTSYNS5s+bj+1O4ZLbk24+q5bu
YyCBVtOxPE2fdjPpmXYX6vbvdu7AOYbICBL3TXaqLvicWN3mY6pQSYGy+TfhGXlnnuOnGNAEWGXq
mlY0+ZH5T9QqH33HN+9g2Ng8uptuIrushNKf6hVup8EuA1j1EY3jzJAYUXl1tM1qA4xGfG2iaph1
++/+tXwfHPzKwBjonWyTb7fCmji34YXfB0UX8bdBzCBgaQmrKkOKn2akZCAUiIjo/PyFO0nLELDe
HlMDB0TXYD7mX5lCFrP8b/tidl2aoVNlaX5pEz8754KyjAJix/iV1o1ic382RCuxBBHKfiwrAzuv
8yPW5sEij5YyVYl+QdVBkQSwgHo77v7Ed7rfLPdHcJWorfsHNnKG3fX9Ydx1DLxrdidc8Tjyx3zQ
5dsOyH3RwLVgrPTzN/FKrw/PGcY3I8OnexFXzzzKLWDqNq8GOXRLK+0HIRe7P26x0tTUaUl+wrYK
2Qds8kY3fXR7QhBjP/u8XIw3Q72bkJvmBQ5iqZpYSi0bfV/l3VeiyTHfI8NWrVtV5nY9u75r7kfl
qk1o+3IqU4QN+eNobz7pnIqLLNlR9qs6rkjKdWZlKATJqeBVLirKXx81sINRG3tR0NYZRfqoJ5Uj
/UcNdgmoSVJVu1Wwuw5g3/y0V3BO2N2Rw0tPNQAcZ/hGen/wKojyV4dR03LBfZcgVmYtmHo4jX3i
ju9g36tBHsCGcovs3MSPWcGD5/XDyhAq1kuUtY1jZggbbLGuIpbuL9EI6t+hlDhJRbziEKK+PSTk
a7PQYWSXfaDaR3xHYMonMcFva4gPg9vn92rt+yy524AVz5j9m66LSM0TlQ8KMiK+lY9S9e2M45xx
QMRNcpVlGRsVgNuZdM/Zbbl+DCvpRm9B/IrxcRA+7fs/4wV1Mavk5kvdZOJD0Puu/DR3d3mUqnye
r6Mf8rLhMj764gRJUn+oFCY4w6oPfPrtmDS4fhVQzOwK3S/2TPqN7nnBRRfVr+ZfBZYLxInOheoM
RWKtf+VqJ9Cg1y5INTSqAh1/aD480Xew0ladWp3Zs6Q72rClul18WLUehNTa6QwuSfLH4Fs9bG2R
9g5Y/a37JlFvr0Kzf0VcRgaih9mCxt7lsQspH8SSDgzOM7ODnj59qrqIcTgEdVLCZw/CAvkpQvSD
1xKWCTKqO23ALln3rpqGtYJVnsXTBQWuKgmi7aBT0AXRRfp7n25c8R+KG59S9qbpvY3qe2vWOf19
W72NeEL0LOnVRYbYd31CEZbqHmZpS917lau8u7if2TW6gMuFZU6eYdlJ5znAXpPZvGJhVtIGwoVP
CpUPU59frLmlgspdcGBknpNr5NKmFBEZjle0Gnexhdqyo9TAIM8oojobfUJ9G5/pav89hkgOTlDM
Vg3BMt2i7+qwgy9M2D7iW+ZXvs6UcLuODeFbu4C+LnjPdo687dOJnzL+GGfFE061y111EKj0QGMx
eLR2vnzaKKWNTgM1nvg5KyvOkaZBMYs7WEmxzD1hLHMk6KU1sxItIKe5EUJukqKGQTU3xyt7aeDn
lCmeHU07ukmH6G56eL+768h/1fq2r2eWwELHk2ryVpHz+n8KXpAgJ/lMxcU6QyhufesyJ1+Q49No
3EjxHndGV4NSMn6zbmvxUqGWVSmQBN/5HvrGFecPC32lnourCaCrHZBoF4r8ABhoboeY6uHLVh4V
1l79whiipEi2BTPU2IAqOZ5BSy3QA+RZCzouaA7ESQ1OF+Jxqr1o9aOWV70wPruQmFnWz3+ugWaY
a2exPGk60m6LD4urwknimbpwgBk3QWRb+Ii9f6B3QcFwcNQQNKhnscC0Tyk3kU1C83AWaXnfMBHq
lwz4fsp2FAGoTrq48d4kfWQex7ZenKhfk03A5SJwfbNQF4mHrfDyvrMZsb1a6PjkNryGCyhrDSZH
oTHcji/vXc3AguQkDF1Cg7XPNlXCQb8k6t67vnIj9qmagTQkG+vsQaZetFAokyr10Bv7uxf0SzoE
aszev+XyLOW51izNNCJcu0pWJ62XecbAbgbi46hFKYwyQ4zBypFfVO8z8HGogwLp7hAHL3RwxVSP
gRNIoSjuK8M7Z4laGclQUgyNS6PDb+LQdvr/SbX4MFKCemlAYLuTRGBGOIv1eUNL2QOLID7TO8pV
4lpboVH8eZdsjr8oqAs7R/hd7doj91Q2a/Rn4p4w4lU8pkKFAJnayHt4epA3Tge6/J7ovKrAh6vM
9rLKoqim13PPjMSF24nkKdtzNWrzv1JtfAfj7icWhQTYWPG080ITgAwnxbBYkR7PslihFWZMd7iB
0uMFVv+yzMCZUP2uJwILgzjLhiVtG8Anc2gPoe6ANPIfQEgo2fabQdRB3a4s38fDaJBNR1X5S239
Cs8aEluWyHNpB4jqmA2r+0wE++Mwy7medyUav43LyIcRp5PIRSqsVAtoA9+t8leICXoGiTaEd8Vn
GN9RiVGS+d0cUvQkEleftOkoibo4qJEX0oX6SWo1HC9Bjiv+GwKC5TSychzZCgHtd9cixwwNqwPU
0xm27zD0/YmADqspWL95oOKJAKSPDTQJKBMyZDBsUxZ5Uw2jCowpLzjqQQb8KXXzDFSSoRaJifRm
84+OwmMsTQgzynY6TfAdwyvkxd7eGZJ5PLbWEzo8G8+YJ7tSoF+fdk5Q6yl1l2DH5txJORbJJbzY
DwUWJeXPWgnS7/qf8ZgBtnxd0YrpNvOGHCLRthKCmOuFLad/qRorUEp3eNEbAeMvDdOuxSYk75pJ
16PLmMo0uo9tSlFDKtSWR1POz9WQ6cMMpwEAYtkHOA6k+9P6OlQuYCVSMzQOL3spjgpBOWq/wf/W
psU1EUbvx5kwGPEJJxOhSIvdbNnLqUhOuOUzEPfMi4J6u8LOjODEkaQeGyi4n7tK0JJr0XqU1du1
73wkuxl7NtvQ1B7oERxLljEgf7oQV9in8BlDSJFZs+0VPBethM8G6mMCW+teGMgk6qAa89ijLmeV
fyV7y7rtdFqJsAJkHNAMiAWdoi7KtLFI1i6FxNSnoH7MOSODxk4rBasEWbAgRY1NPZ/YuZr3gWpp
CbYdsz+gMclW83Cc7rveWyZcL5/DtPWE9IfjRoBkvZy9kt1DURltot/YQ35VeJ0jEDEkId5hTkxh
V0JTAnnviOs5ZlEajpZr0rMpTWB4v0nEMT7w6bCs5wQHSUAECkHYw3olLT8F+9GOdGkpF83k0rya
uNGj8u6XWtoZ/b/NoMgv8RX9F/X+PuFRArjbQalMGe/T0OrM//e/YbEX4fPoGeTpe7/40k3yLgGe
BTiHCK5ZMO8N0KF7wRxEggNdJ3bgKNIkifZbM8ETlMdnCQQNZm7Lh0zvbRjCFt8HSDS/eMn7KI3g
8zFS1ZxdkxI9BSyvwWrcLaJCS1kii/VcA8Ued53pg6hplMV5tY4eFnJxwJ3rThGpbyIWU2dLqgc/
PVWSt9O7a49p2nq4Yrh6BYYO6df3L8vdjF+TED4YpG/26ZzAtSGAiORcz1aoqF2pOrxnv7rUZXnE
C6XlziTffNq9OJgFOmbeRDOeSKJmZXEcA9uWx6PtpFiX2ZXrmjJk4nZpFe8GJP3SfYkcIQD2nf/o
O8zBSXOQZbr7ZkQvlditNoXIOAKM7dvdUJL9ni0UIoAyetviqjE8LzM/mg71TbdI9mcM3g5Ig/NG
ct1PSVozLlrz7KS4e05PvXQ9r3Ouk4Vcisgmaaz7RrjVxXoFFk4Q5PQZkSOATF9OqFHT36Ulfdh3
UbJan0GLkl/dcnpu4WkSMVuPIhtkg2UzG85GFKv9+LL0WKtaY0rR5q+mbHMer066gVDcRFM9CONM
007rjIDFMYGZLPJ8CCDD8uH7LlonyUA6fAuNXm/7sJQzRIqj7NEnH5DdBmDfTy8xky5T1Yp7U9cZ
5iz00ouhDbuAZ93KENUtfuVKw2ePwjv6AJDD2CDhdHhqoXaLHcv6CQfyeo3lXHJ46j7fPZ8gHj6f
UbkzHxR4WkNSRBvA7YNee6U+cvWRgBJYR+qttIt50MrmPzTu9AziFE4iXgkh1xgbEzrbPnnQYX5N
VQD1zTAUxN80ZsCHav6QU++DFTljj7Cldm/UcmxpFC9kY+0UKOFaWNOUnBmOfrfYIgu7LidygbNL
xj3zoN3/WnCntbpiHcgCoBfb9IdQ3cz/ShP5qzqvSQtMqcu7MSc2FrHv/uMemgJaPoQY2sGUUZfp
bCxq037S26woai/Q+VtPGYZd9ugloPc+9dG0iMOTSrDcWlfSKOj/89DmCT7WENQJNntChTt8IJAn
ZnRbpRYh4q7YJwo5xe5FFOHvEpcHVyMNCtL6h4Hei1V5UqrJtFbOZsvhe59SpDdQ2wI6J59zudrZ
USB7bavkv4cA6P4YOOAgKjn08jmAUdC1SCBO3H48o+3JPm3tnUUrYqjc0Wky5Q4pH2nvpGg9iKhq
yyCr46apyIKydnJe4H4b65K7xYni0SGefDz12rqkctHJ80J8SnObOJg4RMUwG8bXB+fzDYle6saM
R+UyOqhbFywSG3rAaXpFOTTzZqkGMWfuecW9eb+6UQm9Ilhq/Y+Qrx57gPujDg9y2lqlTnEB3FHP
j4aD1F+BpRBFHKx25nWDnmf9/t95pvWtcOzYcAuK1Qj8Kbh/JdBeELat+U0LjBbEWBe8A4w+doiU
KvDerFhSuyfoJaZi/sXoUBgK8EtLrDpFJFMtPRgr+1yO+TvKN9vPjFxCxYthMGPO1XF6y7MQY3UF
Jf2LRJl8cnAYUW+sLdpsx/8DBzojoEU2yBo3YbbciUKGMf+C55CPIWd82HDvJLRKarPW2wwWAP61
yn7820Tk2f5Ona/QjM/i4Uk4wZ4By71SPn6VJNf20aIRcx3YrPv/QP+5xP78KeePAGsLlBIHn7Em
ghSiGr0kQHP7gC25HDvwuQh4Pjl6tW0vaQpaNnU1rs6HfxK7ws6gHO+NVNfwaqe0RMUbpBsQioBD
XUO84bBDr8aD/z/CBnUnw07/HxeZCSQpHz/t65B85zC6Zu+/ds4W1f9DQEIqq0AciRLwFLt6AkTr
ukvpXpSZ/DHnDpIJo44JHvJJxswA5aAO5Rpmi8WDN9TbV2+ENvuB4U3v2Bmy99ecrhKuW/38C+eJ
xiiuv8LeHfz83yOa54wtd5ilqT9Trz50RKuMOGE0F7jEgJ6LanoY6zWwrhxWbS9qj9xOim+X3f6/
A2dxfm0B31ZNxNAEmyXMOMq5cKSDyZu2dmJjMkgcdcvg3DIvwEvRoOUtUf+ibP+PFk8dB3Amlrd0
4fINfxtdFo1mg+IjLGWLnYrd0AYYegqSp1Sv1pXeqi4Q/rLN1pbxM6JvGSGEwJE1/5J877pUK/V4
r06T8aVt4E9u0OSFIgGiAia0UiRm39YEzC8kDlBYwy6snTPVxhCm0jeeTixOS1nmM9LAJlilzaYo
9xBqZz54S6MzBqksMT+iKneEVmpfDsvVe68xAlg3Wle8FO6PumQX37d4J+FaVkwSYuPjbqdTgwQu
Zuj1ko2ZbPedBFBLy8nmNR4rrtUgQFIgvU3lVWu2DjyxMaVQ+CASAYHk19U/VKOTcr+PvMTdVcqA
vXso8mexY5e6gUFYfYE0BpcBm//XPa68+YrTFjLh6ZqWa+Ps3QH8jt6zFYDsSIDs35NOqwylE3NV
mKrgUMrtOdLXW1EubOVRua5lM9SeuCPZp0M05dwybs/F6B6m0oGspqTqvQLO1VPrRgjuPn/gwi8o
cJWxtSHo4mbnmCHh5uKo6nXOLxjAbh63lyg6O9+YRvN1zygf08noqMo2u4EVn2MmRx/DCULDgNwS
9CxFb4pKG0qYP/IT7Q1UOzLgM5LeWZhjDTfSTuNs4XIGLicNfyDj+VwRCz+oGJTBdp8xV6ug1bpO
ZxUo4FFYcwJfDsRHv9sU/he6fsOss2ivWy0Oj0WGh3JC+SD5WVltA0G1m0XfZ1FgkEWqode6rtPJ
BzfWNLGg5T/S77AboxyBKCpDvgHjWsFYP/ZhgZ+8G6v/nZPSvgjCy7obDvj1frQ8OaufAE6uWMH6
1kpJqpYDSNqeJNZ3vN1NaxkD/aE8vDumVLdOo/4RExyN/YWvRXgcVTtvoGQg1j8VORfTrHSF71ZC
deBsXCQxBVwACWBZqs5YN1N7zz0OHAlZa4/bYF8BFWBSsYWYPWe5iONlF2Rn5qqkSEuEdY98bbJw
ZxRb45MhPKY/3CQ5ZnIJE6tm5SVKNEWVDqRNJpruLzb012Ubs0Znx1gPMCwellreKfgQA+NheliY
qrACcaU8kjANscsbRqJFtwgYBx8dDJdt/8HKm46IiRCH3wR+JmqTKLdflexQyyg5wl12hHz1iOSh
sv15ZlfCk47OoPc7ucXjNnxXghNAKDaoAgwAesIXTf//R3efESpwi2pYPGL6Wfs8g4XtC7q+Pyrn
6/o3srJ5yysA5Eth1yb5rfPHTP5/VYDxQ53Mp6wLypDiXIjE0uFe+P7yFLPO3PQHyN4FXAkmtCQv
i5X00PWxBICTIIBiYkMXqvCp7FoJnEhV2Yma4XgivoMbc9QMuBPuTZSmuEPnMYZISxLciXMWPZBG
L7uoQN1LFT/iahsXk5WrvvmBUOe+ZqdxvJKuvcs3yO3CbhhNyeqY88evsPfOIADi5ADt6q2pneJo
6EDUKA/pgkTHeJ3RVCO6wYYqy/G6WjM7zGL9LBy/ON1txH6a3Cua1j8sxijMIhJcbv/fGiDAQB2K
Nbml5lJHa0/fp/RKAzbkEYFk9EcwcCZsz/hVNFTSmFJguBygVZ8cDFj+ixkKx+QxAiKRz+GEzrKp
TseSjoFFQF64KdfcPDuCqDTftVnfHvDui3rHTZtS8Ehq2/XWNaHdz5FAoBq3TepaBs22pLApgIEH
eKTEU2/1iEOku4gPIFP4zkW0sqREa4bBfjRlzx8u0eDmI3M4SKFe98EgMa0d8e/7Gt6HH+9gCIwB
8xzy6BzJEvyuZeo45I6PbdBpJOKYncGUY03XtolPhxr12qtfXaqGUmI4M5XhlczZvESVM+KV5UeC
Mlil1LGAzChcWY7rgbGRAk/CMVFZ0zZXTqLH/iZgiEBemDvWIDD9OZr/W0WXNfFMVa7za9HRfiaE
YbKK8MnSm+eyhmxRE4dqtMEfh6vKmss4T7+yZojJXxF8zxoqyJ4Zh5RO0W14sJPGLHSjAOCT1XsV
8piQZ6MW2FczI2SChKg4PsMyWUPLJ4cj7sWKjgK/uIRNvEKnWqJBQ3QRUHUFDp3lqAor6aFHqPDJ
sDM2ZARwii432fwhCooyzAqnmJRLPc/lxx+dD/dAjHD69pSpu2wdVUGdE6OOub0Ugeww/CFsAj8Y
uJWiCQHSDCdAbpoYlXLmAygQXSZIJtqlvdYMdz8xhKkXXGMypMRrLT80eXNilvPvmkWQgyuHr9Of
hkNeE8ltQNO3a9wIKAU4gZYsGAyIpwuGSf2mDcpKA9UQjEy0pbXPWGttAn54cZ0wiukq55AHkOIO
2Z/TlmjieL4gbIBPSB5g2ruFm1p8p2k4H/IphJ6Vfapb3IxeDoV2/wHZFqqJJ6RJE1rCZ3fo5q7P
CLqigD1U1nimktKnGJDOt2zi/Aut1wf1/ul1L4h1Y5UKTxpkIX+aCd4J6FEe8vzD138+aOlPSfhP
LMwqQDKyryNpKmJV3RvGqVk5Gik6qb9EgPUmL3gbKyYi4UdKC2radhqmAXWip2yKosaIdc/OvXCb
lJLoejQ91impVg0YhyYb65K1xY3MvrssOS7HUtJUfxAU5Hgcsbgb3LG7aGqbm/Jyg022+iMhQI4p
EE4wb+Jr7utYW2ZrY4KrKMDjRTtBdPWm9hVrrglMl8fbm7wTW3iYLbCrLL8MaCJavAAkSvQQaVkh
IjuKg7Rgdpj081yqlKFH5cViopUjB6C/1sWqgAEBxLz/WGdjAlOV8ZbFL6iQzSK9tsYVEiDt32CR
qwimh5whqWX3R1/n7YWUK+Js9XyDIGQRATmDHj9WJccOHSqapL/pWySXq0TTa+Bl0snHcRQHS/ko
dzD4YnekY09/YW5DLIkzcl3TOuIOBYMiYhwH4muKTqsFxNUjFQVrRnuqApe1dV9Zhaxm3tDLlRFp
Y17kw+ribMJL7/0PfbyOgyJ/NPMi9yZpFAwTN9NUO218yy+SqE1VH0jA14HklIiuQ/OFObsyPUbL
kE7JLUraojt264gB46U1EWZIjhgI7zvSAHGewe579V41048DEdlKyufZV7gECCo8JJiAzCZIk6Zt
JV5BUUp98IgB/muZ8tgKY+HtWjzKGX97TGtecJnu/DfzwcxUdFqFkRj/75cRuyLf+aa5HW0dLa77
J8TwiT38EKvecCX8Srp/b2chO1azCdSDycqYZUhJ1FvbyC/zOGdXuAvonuUE2ngJf3Jnlz+UgJXJ
KTCWSrDBj5fV4B3VzUp6f9otOttiAM40WHTgQPa3lr1ZcpE4ShImYqrk+Qf7SJv9F4VRK3GjnTrH
AkZ2/t7JSHl0Lrd0XKUzcyfSuNvYofbPLRUhINm7h+KRfpsiYkyuGhvveyPTR1CD7X5yOP2+kQDm
EAYuCP2W3pUEMmWXtkjRvX6Nt6LgZpBGcWpAFgMULSJbvVsiJFTBEyyNldN8oby78ErDyfheuQ1x
Jhp2tkZg1fuJAmeBpk0rwWwUBTthbaNVSb6ew23ZrMjWf5hFnqul0ryDZB2hwiLQ7rCd0CPPIcxq
y0eNAshlOu/LX37+dLS/1uKIOj8lc1TQLHeLhFWLrLVrjijTqYZBxwtXHs6skaeyh2nAGIRxCP6d
Wa77XAoznHflxl7CBeVE7tuYhiRHyOoXcYqfiOXfyCopmYuLP3HBXiEcbFu2eKhZet/nKDSniVe2
ctfhCqMH8VI9fx3Mr9LUHLwKY0DOIWOUzUfmQsf0buqN+Te+TKFwcAwusYLVpXT1tMTIcIEWQ31q
k6bFlA5jQTjyVSrF4+LLSJyhMHPTVOBUyQxJ4fyCyqD4U6Phbl8ZyQkyd4IuYOdmXNMVvDwj2HKF
4ULcIRjEwRnvE1oRQwb8lvTYTFgsMhnumxUf0EGcGmM3HOGtaGI7Hh2kohMRRyz/hhxmSg46EzAI
mPIEJBoebmVGOph1JrqCCnrZFSDyyP8rzlxIwB124XpU+/j34x5c+WzqS6j86zr2wX7g9avCSXBB
ZeXs2Z9OGDZrUsOvjhrY4C2GIgVsKE5odh2tLil/303d557BfgmfJeyk9y+IcArr9W3dd1gy51F9
fvaKAK9PJm2+TY8O0Useno/lwXGK/2wa6BRHQKU1MfGnMD2xJouzRwpZAjsXPrrx+HVeVTaYEg/6
wlTFU0Z7qMwjbIbA5wmgGYLbnRroX9j3sudEqLkghEVHmEpiCBH+DMVyDrcVPLvkCrL4ZaPiZNbY
ooUCSyZK9xs6+3l7Sq3kuE6kk8Mwgko1DpCF6ZMH8ZgBr6Az1UAqNdzRhA4i5INjK51gjEqu594s
SOB8pHrPtjp0PJc2sLgOJ01DSuY1H4TU4AFYNvyk+JzMsw4gC+sd/+wOE7p0y3U0x0UjCFt63YSA
tVhCqSzkBvT7635VQ0PK+i0aFYc/Fx13qPizBjsX3MG7HHYOAwRoGfNorFiG7HJX2KpXhoDAKwz1
NrSbhIB8bzYrWPncKDoFEnkrmAbrj91p0h+oSSfl0W1KPFpGDhklJTqV/8vzk7cquOZQ/cRvVMr4
MkxeB5c5ReBLRQ4t33E/wh5LfvqtQjTYAwNaAQV5DU2tmvPJbPxM4GIw+0sIgRlzMzvXxMH+8mAn
wZblZviWeaBPTJqK5lhGcBTZc6kLQme/UsDCaAcw0Kv7KskGKHNZlOKgpmjnT1V1qugHUqx2Im9I
8LfGpqFysdTqOCC7gVt9t1Ksni0av4ALeR+gAU5/9y3GBPgTNwNr79rmiv8JqZ0OhYQcOVzKR9he
4nYlhqu6jAJYFQB5Wlb/q1EvrgIO9dE04BS14B6pfHt5r62RzTWOVI7Vm7jBBcvmB7y2JJn687w3
pLt7EmAHUiHk75pZmxahENJYNfTwEuN2qf+EPjkfrkMeePDZq5hbqJu7oYiGcnXvjxp02/b3xZGZ
Ts12/GTRdEJ6f5zWZnTmthZcU0JLicLynnIfPoWIL63rQlHPZkdg8hOetPXwEJyjgObYUMtA4vhc
fkgtIFWXH5EXlBWv4d+A2hS0Br0g6R9I6YOZbvUsH3gbKn086cqeyUXSy40xLkL36xsaFh+E+SpC
mxyKB3CHqJ/CcAjPuf5rztRj23Sfu0zeJD791pgNrJPmjxw8vUfRvxqWt4yDGKUkUSJ383oNKUYG
dIg3DnK3WGDwdwyMit9vPjEZkfa8FaO5t0juVDH7nM7oJYIVV6sZjRH7zlHYoMh8jOaAh1d8l7Lv
zLlo3IuydIM8NAEXnXB8LaKsB1BYxzV8wUReV4M6fAnTvFvwPXrCUykgxSiEi6t+xGTT1w1Lmbti
A1Jx/EEu96/5tUav2I6lKKvjLjs20I7Toj8jmbtsTP4++brUhM9fMCnd6+jFc+/lhHWSpJZW0jW1
v0z+jwCd6an6QliTaz6sZuUnKabtVn+LTKsLfavqlZbnrKsxd2dS0r7g9Y56SuugJxutnugn1KIr
sf2Y7LdwMHgWQtkjRnWXpVX2ULpOtoVxOc8RvsUIEbxFFVIDOe45LctvkYo1wilAL0bWDc4q/TDF
G5aJ2o+t+wVAuUJBe881P+2LvRNXXlxxPGMbH0ODuP2IQV+Ry9IWiL0zaWQfT9zzwf+XRIpq8qzS
+ZqXmbZGRuB4OjK6KpOotNDmYLcyRElvIbVpT+JPRbgDyfbhgMv51ozZ3MVtR5L6kmrG9d6UOkuU
TPZJi9PNX8cF3GxxOOCa1cVjMEG3ID3k4XH7HWE8Pfv0HWHGEbXmLqTUSQwq29oC7WyhL6HRy6Fd
XWmEl0jikgEUcxwy9Uk1/IBFWv1PX+69LxILQwez9ivRvzYuXbGjA6d920tHODotezurbVaTYYe7
CPxzYl5N0DLk35WEDmxLVpDZHQETImztVrdYsaDrr/chZAvksb2FYZqggqc5MciUPeOTlSqDGaKj
TMVvqRSDX8NhRTOn/6WEPobJouo/YCvRSLOSPUouz/uCBRSZrbUwtjMLhUTW50XKCCSTHLkzOu3d
Z9fgLUTczamP6CDszrFx+KNj1ArhdVP7kp3ntNR5oBiSOLw8gSjbdiNfDcqU84pT8aIH5pUt2UGl
mTZ3Ue38aNK4zvgx05glNSvLN/R87fJcXMgAxZW/XtyjD7CxrHZgfOGxlBHBlUCcGytBNT/bO/bL
JDnQ+l+5gWjU7xcDTtuQwOOfNTyWAWmAorbVywvC6qgkHfFAN9kl9crHwYbFj/q2RmSGoIJ0d+n7
MShWbfE8ChUhf1zlWRM9tA9SbBgM/JmqU1TjFre0jRwrMDyrhVb4px7cGPAgDR9EMMnlZlvF1bN9
rJcKaJIeOrUmy52I3/TBxrwB3ds8KYIk23S2EOgzMM4Yhv43LlwKk51szrcFq2yrnu2TSHRAO2vB
AaGm3Ss8B959XeTssWLe6zk48Fl15Iyt9NIxGcGXegO8jhVpab5nvfpIHd+/izXbMGXcNzkxWpQN
4cVt1c28d4akDsl+lWrsCQTbfhOOgPbeVzjRJvg60ebgsFl6karfsnZIF5KhZQ2zFy3iJNi0VyZi
7X8wBzuAgPUJ7U8oKiUUr1CGx/CqYvwzZkZ5p2o3whRrCzerCenm5Lb7laOhd8bZogfCCtdmUVlO
+qXaaKoyc/ybKd0+Xor5Mludndwmr2G+ygPVwLfeDhwGiBFLf9QJHygPsL1LqK8gfvDHBeheo+oG
dNlK/S70vjXeYo2xtz1u9eWD4UB0hM9ryjONLAZPooCb3braaPhEKpeYZzKdDNFYCTP8zrBeCVo8
tM7S1QcqIjQYDnhfb0QI1/I1DGYkWaNiG+BAQd2vG/AGnzj+aI23sN/OGHdkUDPKHWLZeLh3ySpo
2ytjiKtH5LaKernsARewHtMuFE3eGY8AIbTf+AZvq9SnKYxIGg4xBDGAMApluP7ZJBomAVukU4bH
W7PfNRoRbybTe7VzCTulVLbyB2lrAMhRybFqZbVWfA/yzBFXffS5S3RuJSfFbASLnO7UPLdQUV5N
DdtGZIgePIMyIr4TQ70NQAhSIkB6VfRmn/82U7/0gMfOFx1eMbHUEKvLZ/AWuH7uDAZS18lEYS1j
FVWHTWUF1ODvyCodtLDtRC31gVasSoCjGzB+N5Lyh6x5L3+7sLanzzRiBnWgb7NhFXK6TyclZofN
vuEFHN6Mc2qBSdCssoYX0OWAdPZ+HnY0Z+mzMMR4gXHSxW8YCud1+fW7UsHe+HcxOIhaYuOTLB8Y
Mfftv3baHKWWAlce2i24nkDIGEIf3MRGxdy14ZEeqIlvyf+9ZCZYusVnLN9k37EULQaRuKN4cyZT
U0dZvsHCAaBFDYMEa1eYRnrBuUmwEigYu/UPPTOvWaNbohzBCdyrHDxfY08KdnrPGdaoQcqNuEzK
fCct5N2NJeE8dI1MrWVGNHCcSh+A6Cd+AakgGdj9Q9FPsSojfgziYUi5MP57NgbeNZeTwqziN/lR
MikklqnXv93vUrTdO6tHOe9SloYLJxrbBaiThc+hAegBDANo5pz/2N5XAQK3IgO5NXo3uYTCJWl4
7o+EVJxADl1lavQL5ombERBsdZ3JclwF9x3cPhOxPMi/Rn/peTR6qHLdADzH3RNM+ma8JbfHYfeb
nFlgsf841Ew3acpY7UT9pkj0wguMrAbX2HZINy00TPcGlg78b+OuRY8tYVuRP6yQgT9ATyldjsXW
g9ivh7au0XMC5qqLbmmfbqtTaP3SApj21VhW+cBDpSIUgWnDu+Mlz76qNGArym7ZK8O+dpBEmbHw
bzJQ7P6fdgPcLcjdI87ESxZ/kFmm3BwdnKj8CQ==
`protect end_protected

