

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XHE3IrNUR0rAgOSs7TaneZOCem+xKOaVUndAgQMQ6fiqQ7sNz2l5jVXfMEx0J1E5drsp/vFpyBfK
us9s0XKVnQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iNP9Rj01ArmVzHoVSW7lElSGoWnbQe/FKLklfFiFiJRRgWHkBTgJfwNby6KYAgA4XLe1eWz88cQS
FukoZ18JES1Zuf+KwL8zwISn6iD7iixfZNEwpWFYjyj8XUfUUjAVZiCjZg8f5vwPfWs79Kh7gZBj
vgDcYNXjxLehTwCVO1I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nmobDEi1pust/app0GNcoN+V8y2mMEri09/oF7dQ5ZiEiG2p7rMxs0iS5vx/JpQ6fiI0X0AJUPZb
worjx3dSanWZxlmpvUQW1C+LK9h5RA4c6zjOdaM5qZ/K+NCauMad2OY8ZgcddQsrreoTh1nJ2DWa
TaZPLvv5pf3U+x90B55qP2fEPiqbYkbzpATAH9u4NTH7sLWgjc2AhgaoW5eC8oXtXFv8D/e6aVTG
z+0zADy8vVe9/EfQm/dJ7Jg0DqAR5qYWGcVn7yVF+tPiL3kEf6FJZBjo3JgKIu+qAthsglm8Cx+j
2KVIa2CX5Gw0SJbZkMW71N8rkZU8FopYgshYqg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sQodddsOwbYSlSsSDMNCYLeaJ51uv4v/ftdtzRqygsJNUO74ZhxTo7+viqM/zY+gFJjqy+vyVh6/
lpYCCvOfPW9ohlsyigMit+d9OfUAHtHOnSwar6P7DvEbD+534I8OBinFHuDcHnDIFirvT7RdkfNd
uCfMWv1oGIMacpnu8DitSYvvt8DCB+bHlF3ijp/IC+P6O1hD15eQnQpsDwpKg6nnVcZHA+6NbT95
rwOncIqFR4E+wPstj6ayfvxsin9AXJ/L3hE0nmxedSpKDKOwBjtiGDED3rRIS/N2OZSt7dsYgyAa
MHSfsznlBT9CuauHVihH/u5MN1losnUyYm2/QA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PcTPY1NzlVv/1miCbWVLH41v6m5uRKf5NQUVNklgE08sx21KGWF+V/ICQGqfMvIC5eom8kSFM2HQ
dFf8l+zO8zFaHEcwmOu/VP5gnGydh7qelqNx+0jPz05q2jp495ez4dMFlOZ8sQGQEzx0VockI9xn
YjRJ00trguEtLmc6trk=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lmC9ahCx71j1/ZSeKA8Rkt1tIlMKGNu+RHHj5Xtwh0bt4FfcPDS17km8+8ppXi7OUTyBXSIFrdK0
NooakhmRZCmMYOTdKwnxgk20HqIlahm9Iu+bxjgvH97W6T5jJcYvFslglttPbZrvLoRpnSfUfQT6
o0EtaHvsEFdvL9+ScRUKPku8EqkOu2Bw/VZKo9IMnl0FoU5KXba9O59tKh2rkrbNw5L2gwOiI4hj
K6KuGhkZNMCIC23+bh94VLvhhAbeZ4zYdMXlsjm/BFrp9rW2/KEFj1X0Rlmh/dk5PzuDb5p8oOdz
YKZejj1J0rHlMYssmi6qnwXn/kI09IersaxdRw==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
anbwWs0l97JVYhigoT6et3H8TOlASkW/Y/8eTKUdRC9TcUSfTU88XxtY8yyw1fQpzUYR2pxNi2ri
ijWnRd5cdXyd57zrFR97a5gvOC1uBQO+VwZqLcjkcD+uCBspFim6ZUmqCQtPaJptG7SMYEatmSeu
5AOckCi1UQBo3bcklZM89hRwua0b9rPBtFacTvBkGGMEj+3Kb+3nEBjrhaIJyprIebvMvsj2unDq
NZN5AyhAJSQgoJgaiptXgMjTKV1UKRQ+AUYG3Il2upp7ugSL5p+QJ/8P9M8v4jzmg6XOd+GGtyl5
iWC6yFcF9Yjeui98q9M6xYivbpBmKndva6F27A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SEfonlyNG8YAcVnPx91iCPk8borIGPaWiJLZAjQ4ei/rFpUclmCrmdDaAEKl2C6egNjlAS0+sjPS
Y+zDUbgB1zmvlc/tdhSobfHENw4E7nVpOiO3LpH0RNW+vE5gVHIgH14HjipI+MnMpA0WPM1yKTc6
9vNke9I8uopfYKPwA83sQD58OW6+jvJsOUI+g8qfuRMbZKYy/Y+NS2tS4ypXR8KfAWW6gdUxjrnw
P6T3WgTbG/zxJarG4sORWn96Yc1NAiD44AkpnonzeL86+briHkw7CsuzAVLHENNjRtcIeC4zYXDr
LMlHg9gcMiK++n43ZX6hfeV9cJnsZRPwcJdMvA==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lo9lKufC+4lUbxCisEYQ3GipTP95COa6tmahcp8LSG8DdAWaHT60LT7lpmYwIBAutlJSIqVJnIHn
qUrADSaI85BggWmFFPiBJ9l8F429HJ2/9X1wD1vQmQTxvt/NBuo22uXQ/9tVB5jGm66HwdD7M91B
vQ/PxfdS7joZd4HlMEsJLq/DbvxI8yuhcPiR9juvFHiU66JL+blx5ETQSQ7BUFQg9UthtE/ZNgFO
J3eLiChOF77wzbPzU9J9Ypvm/Py5gy7KUuzfP0RlH7s+PK7XKwdoCXUWxfvIJ8LKfFQP+lp1RpWV
4tEypdUV2MqqFIbhXuNGlk4AdOtkcO7Vh1IvXw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125888)
`protect data_block
z/MQZOOlLCWC03vE/cTRRDFAt3CuA9ZFbZcL/sQMZbGZ7EtwXrZVgZRkPEYgWT8WIYEIgIDbHWa4
2efCzuO0MPJTAv0VV5kFX86qMb41EEhOt+V+geTqZCIjPq/SgfOTAZclpnTUV3ua3Ktm4akA2iFn
VU3XUXEgs99GsyilwpY5lkpUlv31x3N6Toqt0MLrkcBiDGuHWXJeGVS0kdcPmOL0/4LunzAdZ7w9
efNB5W1oHF01ylmYOYnC9KaDVmSxYjZcpUyT1XKqhrR+THN9N4J4JX4zD4duYmDg942rZyEZk1J9
F41K7ut/zD+Kzn1J1BbqYVxzxgpTwAzPtDie+n3H3b9vwOvfLGu85VNOxcpOZkUYtf9vbwTbm62d
VlbyTir+sVxqM5s0gcss28QQRxX3vzBIqLFulqfRggVdgGYTvKke0NJOpfjcf/i1IGsmeW1DT2Sd
ZnB/7Rxndkf+i5KFrYrsedZ2YMyT4xDz07sgHNVJGKsq3CTj8O2Oov6yz+f9vp/HS5jJJzkzol12
b1ubsMXVla0Xzhk1jN/FAIa8S8RRg2DJVH+pbuELd2FFpAwoPpm5RtwszdgrFi8oSD5JZyoFDM3g
Z6EAouRlhns7edmrDP5LLdlEHIEpGjTDo6SnL4XLixmCnJt1hK4vjVts7sMcOWkgSw87SLD7XMGr
AAiocB9CdAxAQHLBTa6N+X/is/EJzNV5eOZdYVqJ8ZXSGsgHtlgpr102Lb/yjfrhlxNOwevlDkeg
epmuw5UEl18h5I+MXv2mLH+DpTFV2Y3Ar9smbyGodjyS9Nf9+OpuY5n45bjtQcSXQ8+ax9AqSlr7
RQiF0e/5ThMSHmQAqvFvoistj3moFFs39b4DF1kR6tsdlcjVS1JV/2mrbgzBQ7swxMAnwbUd8EM+
/E0MtcPoL/0FqwFGV1CGzHuARZ4wfMYXNBi5+MEFMaM7bvUw+0b+T0TcIck2xV458ZMY9PqA69Cu
R767KNKdpyBRT3I3ngfQIS0hGQCf1ES59XkuNT9nqb8pgcCiPvwerNkVmI9keCX+dEfagUAcYBx8
/PztNdvSdzrkrws8t4s5Je0Zt7cndayoauOa6ERxu3183MPRe7SjEZytB4hNsmRo09juOY9xrMpS
WFtPpSNP2grfSHVcKMI13CKYCDNFzEX21V4UAHsAk6kcFmZxwMIuoTMJGSqHz6p3T81HTCzmz1ud
sOn9NMC+zKHBGkiJLsmvkU5lebmy8QljD9pBvv0SP8GA9qV2eza8gVKkSghuo90OKcy5Y+4Q0SR/
8WTGrhP0I4Nx+ldp25Q45jVDb1S9ILBsXQeq5OyenpgZBAJnQPLOjcu4NBUo8dvNZSibPDB83UDL
sIB94W9+8f/Ao3whvl5GFYSSUO2XXUhqf4RJ1q2uZVc3l49ftjPGToErwzoSHLP9zcetNBAlVkpA
YBFN9eDKJOz30X5Ou/Mwk4gcAxPHdzxSG3IzW9gbohQnw/eN+IZQmDpR9nFfgPIrWEdv1lSAq04B
FMDcoND1VFj1qlCruJOhPbczYjLdoiYPKXVIYmTx5j+K11hWECfhmiW+KYbWb+xsXgnWrhL8q/4r
9nGbFYIm7+ZwkUtiJ07jwW0j9dx3blPPAf72fTC7QynMoGaIp1y+V44SenW72Dcy9naUGMP8Yi8M
bobhWziSAV2/PtpPYHSYtoHoqp0z/EIuU4ym2bC378BAmZ4HibS6n3RONgY4ZpX9x5NyZ1Zv8hs/
z9smyz9DUonDgUwWlavh8OtQ7EciFx3+A2bGSRZHGm/orVsVJ2B34UQnocvddIhvLjw9qcPD1AUI
yStDtnRj7Goo7QqKk+cVe3N8KTDBbRE7YxE3kS237SHIojQFJAr/iDNWbBnOL6uHID8oCmxSfu9H
LvTDPepIPtnHAv1RnQY/yKQ39rpP4dIJK/QaZOREYduPA/tFPviK9l+3fMwCKL0pdw0lttSGe6OW
1Hq+Wy9OItaEprmC9CmPFfuhZyw84yoFefBTiambyQGFPCJEpYc2t6STIf0PZ8Vu4VC4GU1jmJTh
u/o1QIKAIB49GldVyBOSuDPoiwpzAKzlYNBei1a0E+AUOz7PRGOI/o8jBEB307L1GJ9guvd/K2u4
XfUBlkJoSmEgE5adZ7VOrlW3n3NvmiKjjmSr4ff/m1QNigrnOSC8EyBpV/hc72qUYUdFmZgllaI5
PY4+aGHdSlY5dw64lh2ersrDgMtXC97eudv2P9L6jbEEGTPZYmo24aojV//CB9gMOzBgijREK8CT
Z/E3NX+a/dwcucyxbKZDuum5Mn5VQCQguXLCk5O86zGLpbeEqc5DMmbN5gTRTt2a7smPzLHkReJf
7q8Dp0vqBt8uR7A1YeCZ4fhDDQPT3uZSqSBzgvQB1ro6WE/ctaA0dtuECRTjXufxM0GHESYKvb3o
CQz1WHg8CMaaANaLfJ7H8puY/Mn+xhtMKVQ27nH0fj8LGDV9j/oHXQY75CvnaOIfQQsgH+BeFzl6
4qkDLhOkuFAxJeqERTB+F7+vtRLgXsIkrx/5qYlmpydw5OFDR7SqC0PFoewLsw0zeBTgVZjXm1iy
MOp2reVyiXLDUlpEMHwsgFqu74gzh908daghTrwmvjbit57IW4Nf964nVfgSV8Hu26xBE9SeYHqC
qgvy26gM18bHZcwz5qU6pZGQBkhxKuqppyoABgsplwF4SEJK/IsbxsdWi1dunfN25Qj+H1TRoDjG
6INNRKWwXdU9d6Z4H241UaMxf8gD639VoU5GUBR23a+QUSL420B/XFfg9JxzurwrwsulvkOLKfNV
OxgoXLZJStW/uh9ptqfWmCib5ZSLaWTXyPj1OEyf3ORrw6IN9IH98LBDR8OX3/QdxkMDcHzQHlvf
DOfpkBBt53U2x+5w81xrS0uB6Jo6wwZMLf3boEnlygGv4qMko1Rmrk7wu9nYnwHbegSlwmKzVysL
nMg4LopbMoe8x/YZZFeezQPmeQJCq46MKAG2DyxwPpPWJS31dt4tLmtLHcu0gU9bPaTJl+fSFGF9
7A8zLK49LvJ6gHwcudkYdRPPiFW2wbLhrwqXUQYV0SnNXW1+ATRl+I38x9ND3vLAZvv9wm6Wynvj
vnvZtGsIL/JO6g08xUdlHUGD0FW3VYo5AHoqV9kU4jFvRYziot8e0NYTOCj1cQms89XSgyHCcGG3
qcfGo1kaJgD0aM8wQRBOnFajtXga0njx6PPJXskEcNEcg5k8ioUWXn18mfPuf+eSNMRhVJ/iD84s
NRi8kPz5BWxfZxN8AfjLigPg6VpiAC+NSIbqzq2JdGYtDkceU+mUz1LSpQJAzdc0t8mJH100dmPs
/3fjnAoHUOA7nUiJwbRtsO1zEL4zlJyqvT8wePByCxSJSKn/cseMfDEuY9bhXAKm+RYBlp9C71dY
ms2ZWTBwRMoStLRR8ahZjCplsRD2bnJKknkziDFxM5AXz5H+wDKaV/Y+4mcGJP0i3bW+G2ZFhdgu
4kk9B+c/avzxGf/n0WAOoOY6AzqAkyFeQIhdlKj7qqVgs7DsbskPuECLO+5iwKHFlFYhS8lT5UVk
hlpYZ/Eb007JYqadMtKRXeAN+pjwzS55HZzoIEZtjn0JNWdZTIdnshNN8OcGnf1GcyceUhlQOXt3
chw6aBHBcSrvtYJmJ2OFSJ9f6cCZ2YU5SRUvv51X45rJGXORTFZUodcMjuYl/0ekmIVNulVYpjF7
sMlHeqzIsy/aHf4cgWF8nB72X/KyUzw+u5Pa/ye3w1Bt6I9DAsQr/E8gR85SnwGefC47WMc/a3ni
BW0hcOjdDy7226hhbTLtPx6/sLospEseoAbEf/47BQ3YA/8c9+aiiSu5I/FpjFAMOwDWHyXc2fPn
Rxl9HeIJQfyuzgDl2gXlrSvAAr/qIsQ/ew06J+ELrjgA2B2z/rkAQeRIizeNeXsqdtWHB8EGZNxo
CU4NLoVmBuSJb981njNpHcDiItZrucQe8OMPedvo3HR/I2P06Bch7xEtTJ8K+yngqDzm758J3xxK
6a64ASr3JOCGcJfbWfn95ZPsmWQlvV/bixaCkiSwZfzUzCYdkdBIBoZI/UXewK8TkkoZJTVs5t8r
yRZEQsaiTic2zILuW+EM6GWhQJYw3uim8XX59ObG8kTpyL/TQMrtRPVMU/1iQ14rKDCy58eFiJni
3YoI0h7f/Aa3fuI35GX0T65AUn/yMhcs4n6UZ2Hr2fMmtEDpgt/M2f7WjdLTCenPtzXuCpRgafzZ
RG+4uy7WBCrKTGGxGFKetTqzGnY0uFUrkP9F8SVSLSdKYoSTXbqKiSMeH/6DS+920UceOlaLUqmT
rdREzk2ODpw3OVvj7GN2z+yRjz+9ROUi5hCoGoJm8AaUbWeM7PAC7UgOM81vP94sZ9qNZf6kruMN
2NcwagA587VdJKN6AsAzoGYHnoqbxHmOHpNpgFpIOOAeLfegoNldLEYBRIKWT8pSmWYkoSTjbNGK
eQcSFx1e576qjmD2gDtUdQ6n0AIarFwCSpVLW0UF+tpzJ1Prk4GXGeapX7gSB1bpgwKgSamVp9Ci
7FNKv/rNY1zw4VhL3Ct4pv168KusaY7lutW/qXvd1iPZNK1UTVl6AWOLVD0PFnBs6PgM7286CTTt
+YjyTmO0B6hlUoQvr0VyyK3/FlxcL1/Yq6szhJh8htw6wQUCBpUkiTMKjiRLX0hvlSdOe9oL3Hoh
fu9nTEgLJulg8nZj4JhE1wXz5OyGCRndYdIRRrxt9dopmv624LhFpzUfiSWccp4jREZsaFCY3SqA
ClrSf2kcDMkIOzU9VyZ/q8jawn2VWaHE0763euqPVH3F2isYCYM4Gkbq0HlpXm9HyxxhRz2qf3nt
RwmIHdYx9FYa68gom8zFz+cbsH707D6NianM006ruqLIbyHEOs//C/WNqIK4/i0Wm8HnkqJbvdvp
JEYDZ8VsYZHiU2fU69tCCS3uuULV+cs4IGYYenhBmILQ63CUtQ7vEIwYoTk3aep7xuDdLJ5JckEo
T8uxD3fjGeuf3tQInfb9OlwaHfSx4B8V3v69oobjDO5t6vYYZrfhR68co+1yAzaY3vfA5rEfqfXp
dUnZO1IlTfppoLu/lzPb26j2h31a3VsZ3OkG/mrDYJejtcnmC9DWeor2ygRXFz4EIFPscBN1EpYu
fOGAz3axd+SaD5I9ARY8FY/qhluhx8QJetTKK00IH+wB27Cr9UbGMBj+Nkk9CWP+ekvNX6CDNS77
LRZPRYHPNlHeBdI7yL10xW2Iy/Nt8fSIpUSgE//VNRsEmyD3f+Es0aFN1HlkEg2wzCXblQPjiYUT
oRUHmzVcsxlbCiQ2ZUVsEInWtta3LpXdzQ1Myo1wiyz3lWilKppwrkj9QXU4abqdLvVUZHR7D08Z
THGZT/mQYDvv6OWCN7PK1xnaRItZCAS70lX/umsLxtkGZ46IYc8TzP1NHdk+nYWjiYrNaxPznkjD
rys1ZFMenP/XDjSW6QtIuDbAVkAarsWNUL9iFERvPMf9SBDt6+hXmrCrKIr+Y+3TBZ1NclEFBYau
ANacms32NYuRjAMaNso5uxqCIlp13+RetZhyL9rUDSO7f+qVw6BdWgQJb8OOI8DJ6EeJuz0N9Uir
+O8Jk/9GEYoydeLGYpo+0ht5uA6jQAOEXtgFGpjZ/NJFRgTblzWXhWp1CqCESKmh7cY0w4wcO/gS
qmG4XHPOeezxvWBra8R/7KcA6/1+VwCf8HCpR0ZagdjDlh8GiRQ89/O2/hYJ+W4bF+MrWlc/h/cH
fSn7vTHBxurFXS/QQqHkpj6zB8W+QwJ9aQyJEoaURFqS4eOo5B2dYezHf1RbBeu1d20+3U1Kruwe
VCgSWAbodV9U1g2pC3oRILjoGOaAlkwj1KvE1o7Gu1Nwf7t8GSjd+1hJylXvlDZ5ZAq5Rqc7q4fR
oKHab1u2WzLgf0WnuEzFlW4+mPu6144UUxCPmZSftWQzLuXJWjg4tldF2OojoulIEKraljcph1UL
CrUo9wXC7rSwz5aZkpGAsG+m6gCY8vLyrYXTle9qbhwgIAajOp8DpxedHFZzddZwGDg2uQf9chDR
6ofuEPbQA+x4P5uq72CX4W7eEY5ASDRVVejXKS4WNNSiNMj/wP4EogEY+UMl6b1R2yQs//elgNSL
Fq3hf1hyHgTlnA+9Bye0S9ws9fbR+sK3pTzY7RkqbkXXuBK76nKbkD9iClPtg3zF5Mj7GgKHjvI1
UnYRElkCJj/diH8O/zLZW/k5JbgM79wNXfuR4dFKLMu1hhA6lJ44ZvQVxspQprSvOpyROicWQSBi
9gpiNXA/YCUaHQueasUNdqJlv1Z3czy8bkOts8VxvFlDarQUuJdXFR+i1GIsfDpzP/po3/Fv0zbd
3umU8QDlvFAUhYuo1taDLtpB3c/vmJTtpRSb0VMcwSEm8crjFkIyItFTrPw8beFSutwa/rnx58Nu
/5CGjHNyss2Y5h3WHlf/9Eb7sM8Hv433gY8Sn98Fujy5NMQ3lgy8vdfmZAvbtVJFwfgBQ+5im/lQ
d5BgNMMe5h9kYdK5IFVPf7fr+7JD+cz0gsWVyajPHUenxERa2kndsk3xGZpn9ZjiusWFl1JRTDMd
bjZIi4ALDp2gzfMw6rkJCd71a3H3zZT5mvnpl/8r4bo9AmYvlxZnJncVcKRMDWAL73uK+mWKOUd9
jfS3s+qsKVYilB1WyoJksTfZmR9Ek9KS8/PSwIOwAR2WZKTGRykgWEallYlaogCUlWJVIcBzKQtQ
07R+LIBaVaNk95WaWlNCAjSY9vRLwZy5oCw3C6JlhN04y2iqCBoT5BKrhNBcS6tzSvrKBoQMUM+R
qJB4mK1H6TWE76uCZU6CjMN4dhcR+JFL/rRgDWMX9M4xrVlX9ZoEfuFa8o3mZlW0zCRR6nG7QADr
5aE8UnLo2LtuYfysmfAMlSWreLUjdOZ9RmgG+fidTem0qQcM2cHjdR1DaMnz25dnxgGJYi5yjbjN
Oz2aUdhtFj6yq7fwGkWBk/xc+ERJsfQA0cS96fNjIa4PysJHn+Ko9watqMRn3/HzZE+02W3zg2hx
9xsSRxNvo3dkOtbuS8bBVp+CxBHotdGUPD6seAwRhTXJfhRQDN/hq78+g0rp27zFngj5VmA98RKM
Ymr4xL9wGiVf7qmvan9FoXc/cutxb4Jmw/SdnoYuFZgUrsRLUAKLOmpW4EDZfkMwv/2u9+HGBS1v
4wBJg480QaT5cFxNttbKI+MdTNmIL4uIKWdiW88RTQny764DsMtBnQXLkrr3sBu18XXNbVFvt4D6
MDuHQdq8L8SEY5xMse93+9iK/fpVrELwJKTUJaYoynQcrbvki43yxTY6WmO+TQaZXIgon6slHfv6
pWLzMWl2NCAv+eLHKCEeoffdqhEwajc8/jhVwM/RTuXJZkCyb+Bbvr9ZVK2oWAZUDj0Rbqyusqyu
jUnnBu4Jaof1hjvL1GnlxapcyORVtzDxB5TZCBz0UMt70qtqqRLSw5aiMlO7ms5WYi1BNh/IDWdv
DaWLKjQl/c+B44VcbdcEa6p0+7DV1iVwFU0I3HWh3fgVwz0AU3z/PZPtYfgnMgDWtF8psnso81Rz
ac2Z9VFWewp226EkWJ7FvpLWGBsZ7gPCP3c2RO/IrvL80I2EQibGwCi4fW6awfUOaraoYjtlXO0d
H3OhxkVFb97wbvZJ8W/jKgfqYiUioN+GcJyjy1eg/ortyi2swd77ADOzgNtlWmus1/vVtOkrq07N
HyVGAlpWDoX2a5O7bwDGBw6v1HTdqOmopSxAGNMu8XW7vq+VYxGtQIX4qV5xDaPjsiS0Eb0V1PQS
ME/NUMMNR1RaWVilnCaWL3Dpnv4XSgNiFR3lLycJ+nWJ2H0vXN041oWxx1sazzRJxfi8BKtiyohD
w9NIKB7U5g3dPcFHojUDz3hmksSaOFLI8XE3+vrlUmG1YSL2Agxv7vjVYu2YcBa/WF6U0HxVQ4ex
09rtTb//6MwgtryywWZFuxEyOiRime8dkwArrZX6Ihaaf0BLO87+wXLXWy+dcahoneZRHbOxEhhJ
a9Aq/Tf2ZXZtS7eWRzsceMPYBbDYSlBpx3ZE+JSDk8yAv55UT8ApjT+DAqMKrEgtU/Z8Disppd/r
dx0NlYEmUoVrHdIOC3w1G1fwfnmF75swFMVvRwL++mvbb0eZhta1scCOTpvLEBcXOBqBJkHln1Ep
qBpdUnkw8k9fidvodRkLZKqFamlV9L1aJPke543g8717ytwXiVTEJVwRH6nzbzmHYcA+ooo9mMbA
HYLN7US7r6FJVMRhXIPrbcpf1ZYRTKqX5B0WjKzAYHPVTXAoDEiIjvjCq0KaKB5+bI2SzeESMPDg
I4VJagxMTT2t0Fqf0nPNTATNgAAghjwTZVY+agLaJFISwyE+dKHQnKXpfUVVk1vJv09/bhbq01rv
vUgJ8coueIQ6S88WGNnGEbCgT6rwhjFw++45CrRCdo3QapG9/rLbm9TnpSC6gym+YMuXlPm0N+67
OpjvmV0rluxBekhuZY23TjNyiOk27k6IQYtp5Xeb75/DPCSQMy4/SXKo8OnT+b3mivdsgHLqyoAc
Bvt/H0tkKtxxquvN+fh7WbOez27tEBOBb9dlZEze2ynUIpzRUZlf03OIiosR8Mnp8dPmI+cozmDc
Hasbjpgre7hxaHKE5Obvy5t6Ur99CxbbdCva0AmCXi+JgmDLCZ/dZ6vCwT4D+UciQj0o1nNwZWIq
QAbsrEEbhmLKvwr0il6gbgYvlU6f4Ir3Gk21LpgkpfF1SsGpF6CGjmR/V9qxyqOYMSbLtFmXII7K
+zJBfoexj/1buRNxNopp3SICyhw1MkANTYdPhMN8+Sk4w8QypKqxeoHfm6DVU3KPk2YPYf4FvmYz
YVHrPDmaNyQUh+EJpLEisTyb8Sfnr1brslvRFNA9y5wsGuxwQYeFUWvBjDbhzW6uMyufHwqmvZ6i
dDrw9XdkppoReV3P8Yjl8Cbnzyug7fxv5sstOwBFDwJvZOWxJS+HoV4JtnrOuIJTYdBuqqFAJnO5
cGKf5DoJwIh3FE8RFoBFEljIUHwsmMjES81usLjcUjITbt/03rj5Qt7wp95Do6OlgUqLcM08WI3Q
xkjJOlpSOT/Bxm+5dOXaaKKiTMvWB+PNOvqwzJbmxUNMSA2IhTKIqJUTLg/rmq1fUrsdpTAlxYrY
h/r6ams76eCzaoQdjVX0cFYleDl5jCiq06lRO4kv88gj9/Zxrhg2+70sPuNRpMVbrO5wNeFwsi22
J6+vOy8Fku9NOkJPTpvqguqdv7B2DNQK99mrP3HJ+572thzvNRbXn1iYrZQTXeC3MBCn37GXhJ0U
gs6ItANJB0wuHqgLenVmY3p1sDEO+Wao93RK8I8L3ydaWqwHpntJaLppWFUfCYAxxYoJT0wfCJ8g
zOj2+nVJwiQtCiPzcIa1EpWaSOykCQMQttTfWBAUl05vn2C613Eo3xPoa/k0ipUmuah6IeinHu7/
CSfzd9NQQpajECadv2Ug2f88KTobGxYmgSltYGMRTf4SZzsJ3aFyjDfrQVXKCNMZkDp6pDBVMfyu
Zdm0k+MdiN+gRYSCURr2ZWqZOfyA6Mb0WF5cG/cQAjy1freP/H7JcEl6U0rWw2eenQtlHBcG8s3M
45Gv14aRZVoTXcF+kVdrj9+wATvnkIbspGwotX396Ltkl5Eo3upUkD5Wf985GqCzwRhuzAxZe4GD
EnZYTph+bDvc5G4924qhnvZH3tIwmtRzOLzjtz7VqdZNp9P/DpFJMm+VsD12PgQspwZmMeD8d5np
qwdgTrj3VCWM3jwvu6CUyU5pevPUE+9Jqw37rlMpyHo38rTjfQFvkPuE8GWzJlPJu1C7lIWNc5KG
2W5EghRMYNtXwwaWNKmJQhjRWbOQRvZLSE21es1Wrw9yjgSt2Fbix+iD+FljWt1AzkJ5Qz7mWuS4
dQI8J6jeXKAs3KpLVa3Wlz/QabAnHflK8HCwyRxyNDB3RdFqDWlJ4WX54G7gom87l7aOXiz2+OUt
5mVB1RWGIQOmuQEVruEvdwk1/BBGOVqtQoCJfSgPmYgooInqginrPxygxKry52ERoC5+dvltlXRB
gvPRvv/lQqZ0Drg96ih8Wo3tbdJanVse/qk8eVy9ImH4tgKcXEmJcX4DKdGgmvn37n9k8kFqnWYg
KnAMfCuQaGXAh77mSJtvO9LAgE1dyd8NPa7wjcZL6AupwiJFq1lm/p49u+8zCURJMbqxWW+m2Y7f
FCL+f9mJagVS0wpVVxWbeSOAp26bItp7mF43th2LYxSXbc05BzWwnbdfwufUtwNSgpGernd9HmuK
8WPYFq0mF7hZDGneKozDb/N+akwLnY83fnlfr0u5sIG/hWma7sreBBu0GDPM2wT10yW+gky6KjzG
cRDLnGy2K7gGKBhtCWSekX1UnoaeEd3JCX2dtuEVuRpi28kzRCv9geR+AxFgYHUamRYRBkXuZwrI
L+X5gcZag/d63m2sLxJHn30BTrej5OQPTKbLPfH0/rad7do4vKYuVV9c9AUhFSQ+WeEO5/aIDfTM
ZCQ9FqJnujRtfxjlXDz9ekYRcuO4o4q0r/oDFpMol4ysrg5D8Z8BapoU7a7OW1kczjwqRwQXkHXA
JtdNK++L6k4xhjQYN5qYgi3Z6KPbAuI/mJXANTD7D4Zmd2hPaVYGg9jHvTHHXnqs5EN1Bb4TaHqh
LwCwBGPkrontxCh2763RehEkWhyB2Ti0rsxbdEeHhb1JFJGbHBQlYmP6LBGl7DN+V1gLWg/tBu81
oLoYHPK21J3nkqf004mIGATg1jx1LKiAkjfcxye2sHw7ab5Or8l3BQnW+yaQ9C2kwRS4D9YBxOrp
utjST6Ux8stEKvov/H//s633heRc193EDCUnPkFOXjdWbn0al9fRtrETtdHb4c9HhbL1Kb8O50hb
5NQ1D/b54ATlituYdzXXyCLchQ+GcyhPN+OHAK6KH/tpggVwpOhVT2jfYaw9fBOMvO5JlrKYuCcq
JNC/nMpkeKaZDX4iZSGvP0vgM9DMSjjMnk6IJuEsM7OEw4O7pRbmwmtnh2+m9fjihrdocKvS9k+j
CorDlVabC9HIOSayFJM5t2FKibaGkln3JRSfD2ziV1gmsnucH5la+c81NyH5d6f6vh1htEJyVa2B
jiYsbuh73wvIZ3+vmG8mv3E/xZByWCQ+2hF1zwOn5eup5Sa4CjJGuiB5K1bzB74Ur4RHAEDZG4Z2
0guUUeDH7aFavKsUN0vVFh76RY7yOi+5EUjI7fX/ICU52N+L9O19jpZ7vCspiAcHditurziGj9eP
HBfSgu6tsFlua2UYlfgCraQpAuFlO6qvruDGG+kVqCkK0fQnZHNJEDwzxyYW9CkDZ/fyYApTJRxo
lVZwSn+0A8N9KPfnU4q1r+apTMZYhcQrihkVaiV85kZDoKNvVmbduCeXkAaX0VAQk5cpIIpiAfc4
DeRp20pHPfvYdk1L9MOmAm4tWr3zZLyGOOWgF3NKRoGWYBmzAE/eoAxj0Uqi5Uq4LdTWnvGTK5Wb
gUci5CK0xKVd4Y2L0lD4EHRwiYoqLq4Jf+W4WB+QPoHZ6GL5eYRst9wKGgkpSdyt8IIxH1tx12mu
kw+bIR8oGjLhwGR46IYRXelUhsmcB3YzfEkEervl7VHu7xHlHQE8bVS21D/FC1CNfl6J20rmIzt7
RmIABmVnfgiHvZX9sSGXMuqRry797P2u45UzBVcn/FV518ukTRhHZ5dml2u5usqTSa98PLhhVMPe
XNNBY8UIDfUKb6mIHDR4qdVrVldAp2PIrpvLNSzWlusu3eAUBydxLe4fzK760qbC4u6ksIi3mZNQ
Cq7J18S5ECtDkKXrq1rEoaOyqPk1m7QAJGazJahCcLKxrczpcX5wIg/+8qcS4cGOvGGHkFeAUqam
d21ZZ8CmSgNocbaU07hQxItoOs6dsBO5m7XRWl8ZvkaNZs20iIhh4Yr6VydB7WiOA2qJIGg5eBAO
YnyvAqB0cQS8pb3MF3qmMvSzt+yQWSMMPJ2iumrBeey2Lf7/OU7GPGuQ07ghp018QqKZGirmoZWh
EG2z+2dD0uVcN9prFb5RfdNARWn7utviCBPc+MBj8yjCu30Zx25i2BCCImi8iHyZzZlN0rdmBCnE
/YgjOK3E+vi+8qv69PxEdmBFxz7VbOfg6PSxDIq1zEaP/i96vfSapOblgFd13EApBJNih91xsuKh
owGZKaWwJY5Vp0n3L8youjPuxF1MHxOQmTW7onu0TLv5R8BsQEUwGWmkiQvg74/Aaxs5mn1y0oEu
qvhZqgxOKw82dykxIHNGHb0GqCjbdWopEMux6vZ2rhf2EqyI2g0Sw4igWB/foJl6gu9h6zjfyj+J
EamCaBvs44+yc8xze3gkQWV1RHUmLvoVPP1wbydPaFNt1t480FxypiOJ0SQ3wNTYNaFIkioAeskF
lLe6CtUaa7y2a7vOORjW05QFeH/TWsarB9HlMEUrOxcGZfKSFmGRFm8B4aH2BS64PZxtyEGvnrfC
L+pSutNzqwkBLTTazbwLJyVdXotq07OwnTA3dO0LD//YVIQ7qoLNmA0ZApiAGOtTYoefb6UySkQg
DvOFY38vM1jvQRhcJMcemX7goUS43EdHKDui+ujELC9/6VCI2tfWI9ivyHhhYBn2hVjm8uH9liOs
viWWEiISV3ByvN3ejuhfmU4LFBKdkZ4oNxs8LKw31gqehdcgzMHIvTu0uL31FHYaYwwrLpBZQwMv
TjeCdIq8jcVL4+oZrDwwc6pNpWKsLNXSql58DZHnWsE2hxPzxkL3JLoXoC1xOLuQUpD3ByD/tfKA
r7vNejzg5l94gKLrqQ+veCp8VvUFe5momx7D101gnhhguO5gMueWJqNCLjQr2sxYn93Zi3xyGpQZ
klhoPaq4QXGBmBDd1zCGWLJkc8epIGSS7Vr+GOE46MYxwqrwmLyZ9YqlvoIVXvuNiIYj5bKRR+bl
4eF808gvPRYDmK0FlMDC/sfantKK7+KjslZ4/+8eEorTVyfTXbQoslZx8hAV2TacBiioUOvbCMA7
SJOw8oaYfDWJPWgCiRxjhCj8J8Xp107w9ChIXDG8yxqoT0tPVhn3+Z6knT3DENcqLMhTcmVJsui6
hCmic/dd6P+3pt1xaU6YXui/jqGxeVdOvYaIYCf/M+EAU9Q8aeEJUmHM/EiiQYOv91yGANiakgn4
OfZL1GI8mLK8Vvlb6HIQxBFG5dFLXSkFVzi7C33OQqjM4hlW9eQ2miegu90VGX3oO3DNreCv1wQn
DH+tt2gpdYHMErKcbuNPojFXa6jyLrvLIWRW9D4+SMJXMBUXuR8Ptond3+BfvEdH6wJ0Wo4IlvHC
I81eZS7NepcrWJifaTq4XBlWCNmlGqfBxD5y2Zu2yLhGAP4ZmQyqrCNURLdyb9Sq+CHov5oZ/WAk
8YltZQX7jGekTpj81+evLSuNOgtvoZN69BwWqlTTRsCElJkAnnXLTcDU7p+8GXnU+jCgJZZ1WvBQ
E1aSV2YE34PESj7piqqOZ8aOUW3cNnIAifFCm1N9Eaq0llx7VM9GrOtRvAEm5eFtcgzLZ4I02I+a
fOMePWNXS3OheNKVMBblK9mt9hkBXWpiNQEI7OVlfz6+PQ5xb5+ScvT4hxbgQtdioQ90Se+dnnmP
okgZu9t8h0pej32dEbWsUdbC3JfXdDXKrp+KS3fv5hrO/X9Pjswgat4U8DfV3afnFbzck+a8iCvM
Rwbr3OhWataNsEuwWiLj0DHfOG2Jqkxhbo2jSsyHj48U8m4w/sS4o6LNwohjoWzMRhYS8Aauoiaf
YSyn93GOUxU7oqcedkChbReW99p2fyJUERyzGTawkCg8l3QetoyYsCIRlQuzGv9WCAzCnHS5cnja
94l2HPc9MdY5uCEQmAQ13bNZtUmrsQIeaj6xDNRIjNaw2FYOqe6xStIdQoqy0guALQx/4E97J//R
g/Rwr7BjzcGwBQgUKX2kJdHs4rS90xsgn0wochgWAYp0a9r/y1sB+7jFUYpukUjZzYyp8yOHMhkn
7WYSgivhzW61H6FBRsAg905y85k4qqrhWbopT/k0APRl+ikp/SmZaeteIME8AvRsmGwVCzJE+zYR
G0nyP5ZnEAC2pGNo1lWsjOZbscG5tcamrYXUiFM8PCXMLI5YwdDDWMDbJs9X5h6S97b2SaUc3lG2
PR4BIQ8y2xKTCKBs/LX3HMd1lUfqVy5cCYKq/13PlXIt3VroNdF6cScs6btfYfTtTUI+q/GTtiqp
bToQBHwvpOHmCoc6qFDUJGnhk+9/YqM/AkmiKBKD+88Uk0OJMmQ1kIHRUyl+/Pka0McbPH08nbK+
kDKKbhH5N59TeW6WegiHOlr/inBLuW/OYSMgwQaNk9v9FpQX3dEpvUt6c7Bf5CfRLSYHtEFZM4mc
UD7gd3lK9JCp+I6iTtKgvz9qcdLAj+zgK6alotm1S6gRl3pKAbDKp1dyZR2oCaztmsO7g7r3LS83
cq/sFhF/DBgekm32J73jh0R4r7ty61V4se4KiXRlwiBDNIP7Wgat4vLjALiYQfqSYAa16LuA3Pa0
CIV6YsNl4h6AFUx6746nlNKq4ft1MiCInheA4XpPQivUC7WVLmpqye0l5G/BBQdaHDr4CDCQOWJK
ymAPlji3k0pgmI2ilkmGOd+pY5t3KM8INizRMJzPl0XbOiQ0wj1lJRK2owFas+I5wY2uirRKG17X
bWSiA5+Vl/xNVH2prGIkYVUO4rhxerPjx+EbO2jq/CbCx+koKXbw6iYkGTCXabp88mG/0zUpbSnR
D2LAbrZHuB0aUk7n1ZYUI8ARjmPayR6HY+/PkcKLJnHBxWb6+hnlxMqkc9n+eVlTYDt6lT5tKD3G
DNIe371yyJ04Adc4sVygrPuKsMUOhtweQrTAoi4rG22r3tXK+3Vq7QRASMk8gDWGMfREDKFkuMlp
hBCgHoNNzUZa9/vgDi0GTgOwjUQAoItbwMKtDXkEZzSzUTUxSnqKRwrbJjw5aoEdzWXkFllWCc8Q
Lzcz22WzhkBRiap1B2sPRVbylHmZGIUAZlNYBCiGsWnEeJp1QxTlRMB90KU8cZKRbzafNVSoRUEU
NnVaQSsC/WFV5H1/wGUSgS5RIkJXGRiHYtgr03IXKHVEhZNahLr4vM3Qs4F9NoHBuexnfawidsf1
zeGAHIXLayEYCTWugFjcQqlDTCxjrirFZbQBUfeP7IXJw7fAZbx5mXYI/Mp1O7fIMscGZUhzKSmU
/ZOm46BdZSKWOczdo5t5Uhx4Kjx6Vy8pLpFXQT6acP3hF7m2m3FSQoCALMut/knIG4X4gThPg1d4
uZHDvbLll80cYQUK7A+eoOM6Phc5kUyFYy/MNhS03L4jTmYF3AvdjjFbLiKLQf06Ux8sxWXpzLnV
lDAb5tybRogAT1VAH/1F1Go8iMljDJeom2O3rY+Nac2cfBx6kVE+UoFJQeG1sdwE+BuPYdwzeLWP
GtqnCn9F5YfHc9ldjtbQxyof0CAGpRgm6QVHiRdQ98hqDbJDfx9cxl4Hzi5IedpP3tIC+GsDfKkT
ouxuUwlw21/J7BwCdFRpTQp27G7xmicxhtAEb3NrqyQCKR3JNFzZG/jlhIkxEOjeyJtynleJrOJr
501TFnec+5Pouo8AsKSq68bScQ9sKWtKaw3vPc/Rac2ohAYPIZWKpxA3NgpuafArSaOrbtHMdr1L
pbI29gz4Mxc3j5ptLcD+RVLqLthm5DsO5paUcQBb6EeS1S9YVf8QM4pXzUy6EwBIcyvvSpFwzqgb
UFNwgnn8dKSgBwdjRl6O6Evl3VG0TPUCNXLGtEBx7KGs9m+Wd6JR1DKeTHJ4c1JkPpJqlHAg+wEq
wfm6FGfjPhuz45f7VTAdukaG+vKLryXKc0jMvi5StEnfImSQzVMR/UDn8c+qf5DYXgbFnuAtQeUS
VH++eYL9N92bjog9eXb6GTUGizHHy7EcnRU5p+dyHstGfZbkayBC1vC9EQGsuaPuyFg+FBRS8dzg
nW4Ks2pVKz1Vzx0aap6XTBJPUVhGB1jciT2BlnocERMxOX5yhEeHgtkuCTdZw8plrkt9FOPUkESc
ihsIY5WJP+B0b1DEMrmV3InkdexXnJfQ7Owaltn+Xm151HZIBxHwckldwwQDkW1EjzAW3rGV1Kca
poAmmlr2PgxBrzgmSFHidrwRX2JK178yj+tUIPS8T0nPzoIaocH2Auvr3XiMleEISVuzfzdn6md7
ywyYTsJpsBSWYmxJ2b0YgzZNQuUMNLxWi8a9VjMv1D/nlkInCua1LjNvs+xr8/1BKyd40+aRugji
J4/rJBpAcx97bdn6di6yNIIEiMQS2iGcoGqzvANValTtQKZt+b+QOciOQ3R09w5fVaQnKIlUUzZa
UXZFdVx5xKws3VeNFGyX0btJNmwxrPprR5LyqUZ51dcw074cSjvAfPVofQBCCFERugiWooB83aMo
Gy4AZZ59JEgYAn7D2Iw22YhS8m9t/ojk6CRjkEBrCcGeU72vxiCyIpZRj6cyI/OLnCUpGsFgLP97
qvsRY5Js6QMhm5JMMoPbWNG7cuX2x2/dSFYaujrCnoXZw1aP7K72dR7+nkVg2t0HQdQS2VJesR8E
46+5AS64k4ptMg0whPYAOcQZu3Ujnlz9EiyKG2JKyudI6nZTRre4rcb/mjmJYZCDNUm2RdJTRT8J
jF8QGSk2DkJyAEb8ZFrjWY8VHpTXKj79QQjIy4lDm9EDVhr/ZMsdZGk/O3T6l0GfnkXRK5xjswBy
2kGXhVTRuTiZe3F7E+CTS/3wARZFdSxwqI71tXh+yiROP23Gqz/yJuZD2cEwMj//dN03RSHU+k0H
2SW4hfV0DcPTstTziC392LB67lOLE5fqpnPBMHJRPsyZyUZpYh52Zijztgwz8wroXPdW2HSKgfkw
u0O3RY9PTmFLglz1LkXxRzMl+ZEAYZwCHneyXQE967/rk847BmekCIV/jZ0dQa5EMI9W+LRJ24BH
HcwHTjOW6SHLzUaslXAUkLi6Rgkkr74AUjmNE7xQLkbNllKHgPGDXCnWvjJ6D/sMW2fPb5aoe2dc
upNmKi5b0MNi0zEnATTLBhYI0mDMqJokX4ftaEb9lK8vKFsbZnzAIgnPggTkTs2UHLw+kBLUzUzA
K2y+jdJetTkIO3f9QjFgaoQq8BbcaKo9kOuPv6ihLJaOSIcpC3JGb8ldGXr7GJkoSKU4BSEZaqI+
5CRcmF+PxmZQCZ3p/I3KM/poz9scZmYNeGACSHoZAE8jSJaQdi68+F2YenUVy5L9Rfb9XgG1c+MP
584b2x1agMZOP0oYSLHBndUf0mg2Mhtk0GlT/rL6zxR36BLLgdeJ+A5dG1tUL3nZ1gMlSmGdJrI7
oC8pR6sUjR+kwLWJEFen4+DXcfF5YhGe/UIeikMqPJHQRodV6LRoVsWQKU0WYjXyzljCEnF3Iw7N
X2r+7E/giBHnIkyYf0SxYxh3HrCSlsCLdci/4IrapDg+zelfbKO93RKVO67ey9vVzZcSKetyKu9N
uN9bZaScnNhG74941xRDLPdOFSkw3BJaVR8CZ0NjmTv4fQXJCWEPS3c3V4wVl/0w1r4jpOYGmLGt
rt09887sIUBHvLHbHrmfSzFfBQhSwYj1bt1WaRbDLSAXIQasNc2x8+6DgPNKQ2xFOiruvC31ZxZM
g8h9AtlVw0jIINyjnuMQfcVHfQ0XGIbbZSfZkALrAIitJKE0GjA5IjvK07HmxxfHYyTiSojDCvi5
G2DJP4r3BVCdEAdBQXUOqk11c1vqMH+LQosKuy1vCGV285SI84ul2VlUtBLALYrFoX3+4CB3XStM
8QQdRwTSisSp3Y+wTeJE2VgHtS9pkjn81kg66Fm38SIWrDJtCa2HLVmKDhINEfS3V/EQy5WFDHLn
0GJ9XIHJQe05/VvfYK8Go04CIrcw66UgUPCBwcFqsTQ2X2/L7++MjfbJM812Sjz9nPKM/tF9rJsF
ojio8x0c1Vj3qsJXVZR5C+GyOhKXkrYBD60nUdwkgrwKvR1MW7vyBrTBb3QmZHfBpq5wuawTyIWD
a29T/N30CT7Mp/rJ/PysUYNH81KlMN22q1KijEnOkYV+AOOfq3vEwT7jyM6epn5+ladGTf+UlJwm
AFmxHzzKHEadHNiKMo97kcXk7oYDEwDQYOZcDSId3jL3vbfPwjdMImvbAFGpY8zH2HXki6kLfr7J
gu8I5TZoq1JHM+Ew6/3TpbCv3HLdUKu5dMNgoKfhq5Wrj8T9OfEuZslP4uh6ztbl4qTycbQbmHFT
cpc+ahIouLM837gHlXctq1+AksymF84SEZ6NKz+kmrVYU3PcaASBBG8CxnsomPGrK4481lUJKUPH
dobKi2bXd6xQYig5NX9lAoRiWcFGrK5lWb6m6yXfiqrlPGp8Y3oO1zOisCQyHT32qUmEti8DrLKK
3FIYy7B+Nkp4FctaYT8lrY1urWW/CfI1lcZtroWsJ6m+SbkcBb7S9z3EwSDj+FdCKEtfM9B9Ccc1
ItYWi5WlweQdSq2EsAor1BLmplUnhGr9h0/4YMgS+1sqOsjmRLjEKgI29POnQh8MJ79atx/gn93O
hIwLlIS1qtErRszMdI5hLx9/Jpgt8p8kBSYehDc3hNhDeHbPFaI4TCCKrCInzU6KvKEV+FcOOgAj
364smb2RrJNYcEInMie5o+59e2szT1mKdTO8GadT703MvCW37enfMmY1ktdQyPaV677ZMSMocuvq
b3cR4ccDa+CT7dvpPQ1KQR19v7WQDrnFY4EUJek+hwdoIQ8bvKvClVT6Ls1WNuF8Hi0yDTUI9gSA
7WITu77WkUTDJxeE/Dx8EmYAHKUQuqyjEMTTKngBlaPVn4pl7L40mYpkBI3Gvgt9V8cMx/YnhX3A
0j/eZ1LI7r7f6k7S3SrJJd0D0nEJdXgWgRvquczbwMnhrQd8bvyiX8J7xaN5wRLeo1jJ7NpKxkeB
kjVQgv4CYcVzo1VkjeHmRsp+mnQJw3o3UnTp85n/ewgd5RhSpNUGtclxzzBL75L2eFQmwFbqTpET
2ipM+1V2aehHiHmxCZnN24iBJPegIQvbMTTN6IyO8tSSOerSkFvcP4ifKNIIHSQmdqUVLdi3MpXt
PgSjGcqeh850ttv9E7rmYOo3pjiRdlVxevJrAcaZtxf5xcBEfw+pXiX8QLueYnztGstRPxRNJoDo
ieh86eUedDQKJbgZzKe1KhzggDZ9F3bQP8QQJouIG11k+8ex1LyUdAy2LHD4nYXesx0RladUO3fm
acRjrWf+fqqNZXLPMTL0H0bKXVhJOtGe3//7YFej424HCeSiD+n329iwJEj/mwc1hZINiSbYI5bi
p4L8WUrH91PdCjyV1+CwShuZpPY0zwiItetzclVFqc6ZKC2rZgtSBfMQzgkhY3b21pdU3TxbmqhC
nDiYSyEgAiOw5DqpXyt52IHLWTQFgFatyrqkd5ta1MUSe3Lf3DEQp6RSGR+DcykFVVhNixvxIV+T
FxzKt5wPW1YWwalJegUeyKltkDU4ikOt02KCZCWW0Fl6W1fZSxLzgxXwV5OVP637J9odVttJJyA3
ZPBqGkH5AjB+J20/HveQ5vle3j+PQgk3pT5RVnVcqfSKgXqZbFiTcXowZ7s1wS6hBLCmPIJhZ15U
ymUl4s9QfD5vNVqFqM6iSKtX4NN4Jd1SxWwhj2IW1kxvZbb6LcsvVpWNU6WTdU6d3qSJNhNZ/zja
TrkX2HJZbxl2u0IcPj6/grQnPFErH2DJQJaVYQsF5/LJUXvtZMwUUUaRz04zJcu6TaUEQ1b0qGSp
MzIOALHoIAqO3DkkOVUPdAuQs6WNQxEqgSkRtBtDz1bOddQ5XELhJpqtPUO+ef6R/yXIj64ygrL4
S29ws6F7i/0i80EA4F7WZXp+SXWYh5TNso1QaANXGjcfOLphmT3Zpva42Nnm7q6jRwC54jU5p1cQ
HM94yo/hpCMlnOe4JFXmKyXp7H03pJyFsREdwAmoVnKjX0FjifyMg/Sx3U9WZT68e5+l5yMtbpUe
65tHUYTdEN2pr1mNP1UKrq5B3Q5BUjPu5vmffKIB/eKbMA6ySiHX0em5xJPSlrTJjZC8qiu8u2tQ
UNOoYVbuWa6ARONqEPPON1FC5hrFXkJlbQ4+icogbOUTaYtpkwPZKO/7A/ZljiVZkJMjpXLTu74E
1SrDVxhUSw23ZRZwzIb1jMcF55OGDpGU/oGMSXCIeX/k5pSA9jP645eKjE+hwUe3KH0O5ffn9AB9
cpeb0sTthwUC5TCLFn1wywTuwXYZB/9TjKLfZNFjL9fbBWyMUWR+hEBuxUoTscRjn7F4+kQ3r7nU
Hh9psSHYa1b+MbnEamcJ302ApKHnpv+qMtwsS58N582DQ6BsrC6BYNJJ+hccmaboqxWmdYvOVO/q
79yj0f9ZsyXkQsZLyDqsjui/MQPjsJyTEtIP0/GF1uMoBIO5/V9hWr8+DDtB09aqqinU9jhOqk/Z
S71+d0HPVztsAtjQNNMct5hg5TuxV3Apkno9xGNTlPDCVtd6axQmuDyoNQ06sHT1UQj0JsWal7Mb
XQ7g8Yb8ZTaUxWUQyEOND4oY9DN3dG3lyiibdCHPRLQ55gxlLGWIELBfjsnC2xlrnGFIjBqYxd9u
5p5ga36DGxGA7+h9P8CoL5/R+NGZrLRYzTBrqYV1WUUuJo0A0RUeHMNbVtVBp5R2iS1W8MXjWuVo
npCvY8gxqRdRGSeDbrWk2d8kXUI5PBu3EwFaeDrcjESpD9t1Zcy31nOa07jU0Cx2yMJ++otQVZdv
c9aYIoiAcjz/qGyt6eC2q7wYhY/EQLYToWTLUgQgTdFteKDj10/jV/IyzEe2IXmZSRiQ2ZPjs39U
HuqjnKzR5VB74qMHjlobjYPSzOHZFO5+Oi/qUJX+9LSL+GrikGE47xcvhwYCs3DPbMdSgCd6GIXd
XuRnpyWi/ErYYLmY3gGZFe98bIMaa241nf12202/JDINQ0iE1y5kNWvUFBQHIkhCR29ioeRI1mYp
fztO37+1OwF0tmjmMpInHT/Y/TUbt3PRuI+/JKGZVXuricSUq9I7+LiUJ4yeWmt9stGb1mv39J+l
3fdijez+wUnYXtqCTQ4EDeDkEsSzB8ezDABAOZBmF0+sOXnjANnLF59atvYXP8YruzKQh7l778vg
qFRLQnWJYgmIsjsXyWqfOzEyl+Q8fARWkp+CBae8tb17tRbgHZVFuXbmZZcLgMI/QDIlg7A/xh2s
XVgVqJJS5skaEZQaHABY7Zz02t644EN5I7pCfFbQ03sRA4gtsJQpxTjVBYT39F0FMB5cvDfkrvln
IcTkMh8PX4sVxVogjWFAQ0RxwsjuQJAvbtS7B5Lwm9Q8G+/Lz+it5J6r6ztKOmExyqLrICVCudV6
hURLkOUdkhkUsO1svkWr7/+EKAfOgEy7zEwHaB5UWnVIEORuN93M3ZGM/eZvzYnLXD3PeoxThed2
gLRhJ+Qqd7/cjQDtVJvGgQVvJcVdppqdf7fbfRh+sEQKt2vP/YesRVCc6XHnIXaE6hyOMhC9nLHW
EGO6XmHEU49nkdTAKDlMy2ZAJd+nU4EGCU/kXxWkICRLlbu8z8XjDjg2A4uUy/BMZyYHr/ZaW73M
u2Ju+FbgSHn1S0iCkqOHiZI7lWNaw/5C6IlR/203RMGmNBJ+uGyHbBddpgouYUcmpXSNEJRjoIxR
VdUfbiafzdgy9bJ/x1GDixi36iA+XFThxrEpCp0hdFfvcGRK7XTzgKdccZtgqYmjw7BCqPuovA17
4yrlZ03gXgLn4MGAMvhp81GCod2Xu30NyFZorh82CPtbR3z3CiA8zJKIwSLYLs2QC0IgjJXaB2mw
3LbvUOGHhLi0/V/rXOOXLG0YQRp/p0zHlGbEelOgkHaJpeiLweplCjvDUOEwPzy6se4hjIM2jTNx
xR8DvqVMuLtiFSgrhZJQh4EDhtR8x/kYCpImwcCGHCuIpvJlKyo84OxLSEPBE+gYVIDaktP36wzs
fuG9N/8pJYPERM+b7/KQ8tSZ9RJZAML1jFbnmmPvS1N95bz9OwXuTEU7xJ4ySPLBXb33oXSlirzD
teFZ0RDCfAp1kK3BOWKE61SOKcGsbX3RNQlZUhu9PBelM343MXsq3twAzfNYssI4avDLSZTUnznM
6Mb9GBYeBa74Ht19tixnIpctPziK70XMCVqtEuFAWDJUPoFIsCUYuqVqc4Yoydfv3BnPV3E8QD4q
o/U5M1pIvNFAs5kxwVr4033meNKGuwAxpLbmlF0a98jj0zJ/Tl0zV60TKcyYk6/SGQaZ7TLwSqJw
0eemgzBg5htHaPCHgJ1nd/RzK+k/dUt9+zp6jXfD9gU5VyL8jw2wyVMOx7ZZzkk7vCy+OwCAuCGs
exJPiOv1XuhyoYQQlkkm5WSZ4HVKJjGL9STXKHZhZYfa119iq9Z3Swcxbd49X5n1WqyQBu+bL/OV
QSLjqei03ijR71usK46vV2489EkPEnVGJKQAzj/w+PMI+Ei2m2Ky82og+WsHvNk+lA9aew+re8ag
E7u5NPFP/1PiM9GGZpsDJuudnWdw0zgqTrH9h2yHidhv75KyH5pen4b6PCJZBvyZefEZhXMdmyZh
jAEvBQZICExjijRM0wboOq41oY2Oq2PvZVHx3pXxz9O/PjBUYnwWkKiB1hFQXQSEGm/71xpNS1Gp
o1bwJ7UkiFyod9zFk6OQtRlFsbMY0ivvSkWgboKicrCJkJz5mTc2E9gTyjF6ggW5EFZAdM7mTQ5V
h4PiK29inghLz3+nc9+fCCHbVSTudZn1Xpxg2TfrjjTtM+evwQtP6VaZm7vy9Aw6PjvqlpC71Iir
0XgyrVtKXrVw5DorcIDgGmaXVfQaF895+JbZ5E1R4jlP5v61Kn2HoP3HG0+dLcYcNjCpBGlozpDb
BFsOPf2jp0mUjW6Il1lvEbofmkTGzN/oOas/wUV3WFHWqO5iUBOcQl/Tv9ZCGKy5mS6XNd3BNLT8
I1cfOkwD/cNOJoCN6hoWalooI7nRfX3zWKuPne8s98jDAC0HNeXoxl/ocrv6a+hgfN3LrBnM0L1h
Vf1p8wtem8GSUilciZCgHXpP3IeGzaHPBYmG9UYbnvu8KCnGjyFy2XnyKDWyiFDhMsNL/VhfEpGa
csWsVhbL69DNeVtorsx5JRv+pamaF1xcE60piIS8Wm/vcWjUHMoljFx1jROj0MQvS3KuT4f2zo3L
pKUJXHwBuBMNowq9u2hHh2bZuY/si9vh/Ur3n8C4fHhnLDwbB3bo0rzkDYV6LDcyMjCn/igiQEh9
PTDUmhHYlcTJPuToW/7ekBquz6mKoDKepRP/rBnLZlP51aWNtO3jCZJLQ4Ldar6TLHT3veRoA/Hf
b1kVB3pJ0KXxbmb89FSFhktb888DqEU326+SAKQFux7LcuJPBoC7M1j3opMzmbGggRBfmJwy8XEN
Y0FgTIzJ1Pek/mZZw5TCAOpBZCnwAPKHQ93MKiTU23TLIzh3ZtkhKCx2lzgOsOtYgIK9KdisY2ZO
eMNzduNwQmYBuUBEbRN3kl4v805up5nFVljcQGqWgCsIx+Xdw/TIs1KO2Yh0G5DoDWAMuVh7Lhuh
aYKh1/HYLz96uBlUK1qlVqmwVMusT+oM+tA/cVysuxb0K+TFb+I9Kj/8pi1G0jKvEjRuAnsAC34/
supllTY7a+A7Z0n9hVu6/3D2jFQWs6TGdZjJ1q/iQzTrc+Zq2xDFwCZWaBU0NfImkulFTXLqCnV3
dzPBnJneqg5rywax7NqyKKuSWn7prDdix/wrobKAiV534uEJ9wmTuTW72xSQaAANU/C9D/nxgxQF
Z5kamQX8zLsMp5tqI7CL8rvezpZb9OxiLCF964jrT9SypPPCki1teMJXXNPSo7X3ek37DOmRZ7WE
CjRRQ/HPuUL6agpgCbIetJqFEU0nKzx6eV3o2anHU3srdRmmAfccy9CU5LTM/RTOz9rGSFOgJKNQ
2qvuWBqiL54fWAIPfyIvx0yFVmMCpjxwgxM4tPpp4UBw9rVBzoPYvHefi85jgrNfik9LXG09DGym
ltE4aavtQ7czyzy8gKUPw+R4MtSzkMwBczeliw01+KSi5jr+dCs2dSYNOQCg18Csb0WREPiObSkU
AUcB4viThNe6Y1Kqf4XFyBhGxuuF01zZJAJf6hgqr4x7UqOBHaaeynZ7XYS0LQ0Sl7BW7TQ57bmq
SMCvZ6KSXGvozjzm3rpk+DWCv4TkQxOBa5hbBrWd5zzXWhUEIS3AvZ/O6uVbVJN2A5/xh8Xn/hj4
U78dxaYQctO2VH3hrTvxmqE4GyLjBW71s2I5OL8Et1sn9t9s3L03btYB9YhzwCdKFpmUBE2keCSD
iOumOlifjSy1M6koTpnoVfcqSCpf4z5r0GwymoXR0r4rM7ws7TfKOG8q/USUmz1ZP7Q/4lj+ZLCs
K/YUqPFqPk4fBWOD9kPNnoCsOJP0v7Xt1fZZTLBI/av2cys5u+e78npoR36IrW6KOTtQRwXPUKPP
5Ja0CMoMEU+8FZIf9DawzuXQe/g3Ku1H+qpyuCmaPGm7j3MNvjbwf96wIFq4Jk8kN5i4ahNZBsH0
jsIedNfBB4sIQKGsd4VyNSh9p2qhtxMku+yPqCrZdcRWnhgoS/kD+cyNPWC1xqAyUNdp9mTP0Fbx
kY6fYrs8QEDrbzf1hFppb2tuoeyypsDte9fQMnOB5I/xMGWnssNA/QSCMUBvddW15Prp5OFHhWVS
olaUrsnMI0Efs4ZB/k2CJI9W1rKNZRzLL1NXpzfvV91wvVAGFGe8vauZp6Q+eql3bcsMJT71YrMr
4jiyZXEgjzUWs74kp6B2QFgiFd7MfZRBr42X/6w/MfBFtgd/aWAkf9LWKWYai0Fx/lML9kUHOGm8
lz6A6hOOG6P09HcOsqrv3nEpH9uMdvYth2YO/oNkrWj9X9KGuLFioUwEQEBWhrnL/s1WCWi52goE
OZDWnSojEc6Xh6k7lMMzZhG7QqVx5SN9GfirAsYXfDylKzrBsF3J1jYsu+F0nVeqZcYVPwaVif4W
EFkDFmiJ7P4dHG9Nv13PTsRtj6EtCnFoiwO2GK41pnZHoeGpXj8jVwlzu8A8/lLsFwyjfuS+Zvnf
5BBl9sufmZwh9CCv4rjfbjajWoazN7zf007Mt9SDjoYjJyVfS1Q2D7T8fGf+IsHqM6af2qQ/Cjzo
eEHnCplzjC5hO07vyMxN9fzIxTjo34kxAeVAiNzTX1wTsiLk4HZKlqhgs+gEW4+IJioMcSYD1S5y
XLE58PxdXjwpXzlSC1qFuCAI4vN5bNr5Blt/vwOYRgh5bdn9bCJkU4s98q9gjY4NMZzUJVh+7TF2
lso0CTpfxUE3ch5hi6ybYKXmZSLtx8M7CNisFc0PxTl48fCiZUD1alVTMAQ4FAucmwZ9P3hoiJLB
t3quMi+2ebXYk27ksIHQhGafH85Piu3w5l1gbzDEtUiX/da53ZSkH8X7tiQpmRARaGUWz3pgJUsg
aTROdnzqbSLXT2/59G1EWZKxuA71yWYdvU6p/5Uamz/PAk/KH7pJ0AObMQC37Vkbejb9vfW7SThG
0o/Va4Retn2zX5RdAiVy4CMsRXhGDTBBr5NZoZLazLBtuk+/EmOZg0ME2HcIQTFnAcA0AGvkE2s6
Z7bzsML+q1EI23c3UEbSRAwnKEt/aXP8R3bqw/btlG4IdsL0xZMutjpVCP+G41IiEz+063I2+52O
bscLc5ELE0SMEP4PXHWRLigQXT1b0AiiWXyZ3IiTJD1jYkmYVDoYfCZanQAHKWibadD2QQC05ubO
MoaFjT+p6wv8MUkWXluZf+yXW1pgMnYOcUI6IpBQU1OTZlohbHxPbiSBOIJlPiiKCLQFbiRVeXga
AP6J9E6Mva/hOmkMl2TM2eGN6/M0Ofoc6Rm/G47j8EOH5OQnHs9y2kR3AR+zJ8bxmdwyBYgHcAux
3AvcxIy9RymWMl2U+7I1WAAyU0R0WD0sp+upF/fNQSEXxVYAeiiRcuuGJ1gL5hjxDIUyBxlvlh2D
bm9QTWPXeJZgQra0qfEPOhj4cmNiwydnluG3Z2/3XiQbFoSO4G59ydvTVD2JEBkkkW7IGSnYaOBB
VCo/DZoWAgWR0TlAFqTv7anYj/njkJa30XKNwyVBySEDJvarmbOvJo7PUsjpRS1Xq/WZX4r7I26S
7odZqmDOrMKpnuHbuDi2q6ZcoB30BqATDkv/Xz2XxhYCLrlfk8p2ille5VrEX3JVu3OWcFlv8k/9
d8ASuNfStNzCuVmG406F1Ry59UPT5u7bkzFHHyeOlAzaVqMGWYh76n7PyHKqc07zsKLDAFEgH+Sa
v/B+UHiHlxma8hLJd/zCQfi2vfV//BhJQTM5UZrMpibBhv4HU0C/IMpPKwUtRvO969HEbUIgCjlK
FO0ncU01FKYauM7WucJPjReWgY5zWz3UHpbphA3FHAFPCSrzvIgtxUbVJO6SDAKHau2UjnvvLAb3
Cji7DDzjyYejawXFErII55SLSkILmEHr40HaSUHqfJfZ+rStu1BQfxeIWP6PvBftHgBCRj7IN2Ua
i3tVC94a26oo2ysimlwWagCp6pVC3fUxVCBbkSFm4Nkl0nR6x4f0BwekJZPBFVeqaJ/H5w/l/fpa
WfAyuNl5bqaQLm2aZXHDrzukd3L9/4Ra/taWhc5KlBNdf9X6HhhUuUjfhXoATnsP0sqDj/c/188T
Yb96lT+zMvr7woWK22hUarx3casiL4c6j8SJkWH69RORB9cPN9bs4EpiztnrReDdtvAKrSVvld5Y
mvmCmgqF+oPEdL9pTQ9kOi6zjTzXx5phlIbnkd9DQZ3gZI5BmZnPoZdmquNO1Ho5PME4kKEQH9v0
Dx5aaMvYYOf9uilJpGfrorPK6fq1z7SeSzFjnWpqVCc7i5aEPMCKL1749aIPeIIy3+jdh4ML26k/
w1+zToxsWFdeHbILNwN8JZpYWykkNtPhHyqCuM6nTXc9zw6r3qwznIPhhm8edgAYrHEOrI6VkjmX
fvm+AEvVKjQWMMn1NNXO1AGKfm8Bt17dVz7ORjvjW+RJjbhVbzBOQkmZMD9MrdYbx6YdiPFh9f7x
qsuD9c1+rlOcgE24QBxgvHX1xJCygq825M0t+zsfps32s8H6rJv30xBwPq+rM+azRDFlks+tS1iD
yHCwduZ/BDPpWtLLy4+zidaXFlLd5r8kKnjNcVdPaR2nvh81mp34vADiATyMQQ7AvfpG4iL5wdon
kg/L7GOpPXr0dikWS8DyCq0BZX7g3N+ULUs4UTZyFdXHIxTUFXdKQfXHvSOVaCgsT/RPqqG+llqr
riOM3dMcvcRjW3rFdnXsW5JOkqnyfjMdJtcOOaMd0+Ig0zzx5syKiBnR8FGgcB3z/OFnn6QUiQUR
o9qP1Pw/VWjDXzTNtgT6JfGIBsq2bn/n1NYCZWgUcWvHbJg9TO6WCktrD5ljnCfif7W5X0x5GHKC
3PGVKONLF1t/o+Xm8/DAoTViFEoggFKvs0MjDZgIjGmhFI5thMoUBSlUIGvLAXMQOKiQXY9lkzZh
Yp5zjNqVByx9L30rs7YaVLeNfNqmKJP57Gar7G4uXkJgEG5gVD4o9KkZkNJvewuUNU2+Nu+G01I4
yVsngRk5s6svYqxa1HtrH/NFUbalVHlBdQxUTdYnUNR7I/tuwfzqY7BqxSqauBKkVDKH2n4nX36O
BTgXTflTntSVeNPd0B4qDqWVtMr4VnLsA3qPxgoYfU9KBrPK8Giz6Y5iIxULHCAmCDW+x4mhmPvu
XbIN9XdzsdAOBpBrB/y4ogjAcU95nUGwLanDPYFDdVRxpz9UQtXAGwR4nQm3hpbtqJ50oevpe/s8
dhOaRX0qsbsN2Ke9KwoKDDJp4bhgJnKY9iaHxy50y0qu0EGIjaPKZ3VAICIK+jG2D2FiZ8CdzsLo
5CuEeibyK8ruDJa28EPPW965k8ZjAZD/rGm7+tbmrcp+lfIxvzLXeR/ShslMUXW1Cx5ZzJGqUJ8A
nNOQCsiyrdJBFfBKq0zdTQMv0iRriSkyV+hjfcnZTtaS/8JFQBgEQAMf6nZIWA8p5QSbYnqZFno+
EWdafV9rXJMLTWmJ5dZTUcxU3CAS3gZcxPK1/IZrUMQQbCfXSQTQjD5CnqXiw5TAverG2JvBF/E9
JnnlRo4pY3vf7iksoVRxPdqumKM1MFRlAgcRbruD59RVljZQQjgJwdcBURjccZRbcaqie0IaNNhW
dsxh455Ads8lm5SDYB1ITuiqERuWVpU5XelZdPtZFNSxMHVv00MJLOknPcQM75Gu4QLxvweCxDZm
TGn+NBpOG5Xp+zEc2SuA9jpRto0avUXiUVxXlzAmf/fj9M3rfFmEcfjzImxwUw2oiAXJ76dBb0dJ
hT4K5VuaPV2e10fhdbZHtCwbxJXWtSHtPinBP7mD2ANwvKrbdZScQrsxR3zdNRQsncVmrLwgJTJS
7d1D+Q6MLq/XaVz/9O8t+D697wERdworha6IhgyMQAigxi5wrmA+7Zvt6D39kY4DM0dRtPkuVEUu
EE1LiQkDbqzegunym2EyFjnM0V9awyWaiS4kHixLz00mJ+dbmT9XrHDUqt7uhSU44w+UUB4sABL6
xrEIoXOQynkEWo0L3BKoL6HhEmDWQJbSFIIVwqDl3Y4a1xk0ioqD9vo+LqWhmgY2fAvS4hNLfBU3
FxwEqTUiQznIIgVgMYfufulZW6nwBrql5UYKBtdcuKO9SNlQ87N/eiqhJy3jPvthLrYXu/VZhLKM
N6tpazIiFmNTE83hXhTXu7qUG3J7oPGUrcqPh1pJW02GCtR2koMqE6F3pWkohgS/qsrqWgJIWE/o
j7tBsG0seAKPwKKYamqjFPIMSJdqu1M1l/Y10jWc0q2tKEtH4LWFjBcsjr4ohv0522ZiaYMrFYDg
tr/HqpVEXRXGmKsTKYbCdv4gBTyjXH+TseYA64FZYKbtfweXDYyMePnA9WYJd6kBBQdrvI3EAoPV
ENCFIUj8Y6Tu45YmuDgQgp6UebLxGlMsi5Yhxdb7GvsPR/dZP6bxNu0KMW2p4P4siigWd5WRRF3P
LdNM/EMcHKuzhk7rQfy32FEdgGGv0jMLMLgGiQQ/dQlUz4WJ4muhFG5wKzHQey2fVvjNV0w1PZKP
6iHo2a3WC7fI2igY23JCkKHExzuKyqHgjBr6UOdt/kNSjjUIppsXBiMudWj0ke3h/P+hzhWHRXQ4
JN7p5EZxQrzGV8jNKuyeH31+2fsOCUzg4OzVDP/TGc7WsJ8BbiU1NVDtc7jPTKVsqf6Qv1yVlXI0
vtkKzcnhf8LAjssVRssO2Sbxn6TGxUshN/dEjZV5XZO3mgtqVDxa4YEKzD2rO8A5vuyliWWaicuk
oAvjPyCg/pMLpTR1gB2VVTLeruZ/vEBDGQbKbWWB9KpYjr7B2v1UMAV//6Iq72e3zu+tzR9wF1CS
aEquo1Xo09hZDjFZV7RZt9pJAUDF2mJ7jsdLOkxKXs0M6XNg6kr2iXQMWK8TFY60iDHGsE1wY1Jy
KGiwaCgj1Mrp7znFU+ZvTL5lI6ywGlWq6kUjRh0tweDF3CMmBWxDmDU5y1RWKutANa6pTvZVa4LY
0/9Thngg9rc4JSSmEV6X0C3+wU0LX/NfrmzJY2LLphFP17uVeb09TOuyAWU+LiidIQQEYOJ9PnY0
hFVO/ZNPuweldsSPntbwhlG/tm9mChGdRtiBAu4S2Mm05ans/Pj8Jk8NBPqpUSXfbTwdSZIWsYIr
q9SYGPNnZGjK2aDIOwhSWurskZvbA3BHmOebBqxNiZN0W0mfM90TLyzFYnbtK1sEvZ0NosQRwjeq
d2OnVC9EDC8CcTfE1IbSCjyLLn07XZEGl0Xn0SMRBbcT9iActdxkK8xq+fDgmkN1bmXH+rxRIt+0
0QAGylO+iehFUeTmLdQSKeRY33DPcPcMa77r1OmSdDDXoZUrZXoUu3dhwVFjUuPupo2xa9NQLvy+
/dcVsBfLfDstMf2NUfEXqjhK7Yk9qNHdh4KT1Dy5OAi9S1mirlVZbtupuFGPg66WD64N9x5IMg3p
9ukk+rTwrzx2egKw/tuJm95yyYzAna+9zY5FABPMoOe6Fc2sfWbbGfGBjdrs2lgbUqaG5nn3Xg6C
Ccs4fhlEkYzNsCuO+QysRjwyHXbuTQnzrGHwYEr57VmGC9SewtgYF54gQ7YMNzPIZ7lYPrEHgJmD
b/2a1wg1wqFstulz39W2jAQRzhP9GXU6j4izVXy714S5egt6M/egX1kNeJaP7vDVL1W0eGY9wTZb
rklEgKNG61VlVmvdvBKSk7n8sr12UzeOOW6u1vmJaqSDKzO+hOp4m1I79H/H2Ydff65g6yc6Xz8Z
AyD9bngAkNq3jCAmjfMwW9OItksqWFZqyK0UTF6nTdRdMO8OIdTseq9X/PsZlj32U6VWhCPz5/Uo
idIePkbmp4rH6TjzkFxWH3MV4CRTTdo4DdZzyxjYB3V43Q8/3aF4/IHNuco8swIi412uA+2epGW6
tJhEMalF22a7RsQW2gxWlqkAFmUOvjsNlUHJr2DSg4M8MfofuILRG/EwQYUStekTK5b3cszGzg9F
YWohJ5V3T3D6SXMhXeiAxhC8mqFVFBveOISHQLg+HNfvros6KNsWzpv8XIrcRVavgddqV1R/gVBl
AjTri/sPluMnqTqNaVCzhv+egf//HaCEAnm6UZyq+vU47lLX94bQH9IkVysejLyTS+2h+hpqImE9
YZqYJgKeicyhaXVVs7HoYFTsqr11S+Qpv0GgmrYI+wT7oRX/WEoBmf7G+QnUlDDAsndecd2bde9h
uPeXCdt5sea/7j4HrUAyQ44D4ctYRzK+VzLumPoxPefXI6UliYHDUgA81UemBvIfzQuc5DVo3aRB
LSy/4hwOHfNDgLXH1hU6/WG46aCASOAPm9OqIZmhQhc2CmLgrURZJ8S2y+qCeRaBwE4xm0MEHTB0
w1F4QMfxRLTaQZmNo9co39sXFvWtGVpl12T24Kt46qR2NtT9wXZO0AIrgsmBOwBfIusdcrt+6chB
FTVwjv9ti/rc3adzd3zWod8ZYGNm6AC/zHEiKEUFSk4NvO4Cs5D507kZ9n6KrOrG9Zuc+K37BRAQ
mIIsvlQvtdYMeOoPe5ZKOZumBYlD9EM+8/E1nSoSlpZHCyip/VtWgZqB6X/nOWQQfLCvECRg1Dcn
3jDadM8DhrSNM98lsrhHGfhjIEwLk7hNaGlzqiRVEde82BLqBzEVruQGEPgyVhHN72W/mkP9F7EG
X2530SevBLsvl+j9n9dN5lW3vVx4QGb7pyX6MlRkfyKZRPC9WILckaRT/V4nc9SVsc5vzr6cCTDN
/VVUDS+jgZan3a/Q8sOgsuSFrT6nx82j/a2vWPcN6IxC4fOV1YfTzhA7a3eXdvoWVYpCNmbJAc1h
sGOmhksRy2Yz0z27dx404nmCDXaY3NBvvlbsojKObx8ojbAMpyk2y5DAjL0Z0qd1tDL3misrKsKc
K4Flskj91JAxNca8LyfryiEjAvN5+xue1CmXc00JZNt1vOrNsFpU4JeH6g+1IRcPsLx17vLCKjYO
qzu5UESo2uAqMOJW8LCxpuBWELkls52czjcC+uGBj0pwv+iBRNcvdRv/8FUCGc1t2dOZnrTyw7A+
HRo2ZhpJ7xhNjL0vMS30UdjWVqONHkROg2235m+0Hn9EPlmIJbI0OpVT7U8dgn4hRzqCHSRvMXO6
5Wg5ytWUKjVPV+WLGhLg6lZJOcvBzLbqVN3tVswSRJvccsVB0RBApp/JPmxMuTVhWv9jej4MZeSk
+2BbCtAAfYUCuPGZ6M1eMZfx4Y0TT3Dh58KV3fXiUGCIvWZP+tTpyV8tsbV9nlN/bM3qvwUHPnPX
/rlN/lRa8rzLTplg1578V7v8UgH1rrhot6TAeFJQ1on6qoIBnq0tBFgkGOvim4TBQwR9cUgLhpzo
kYRFmtfUSGpwqbRZ1pzMqEP6rKVIfI9ZSBNoYBeZGtJBoTKM/bjPB8etGV0bKGw4tSOVKtmZA0b+
IEWkzP94yOLaCYxor9XVJKBWNp/62xurBHbX4v/cHuY0dg2Q3ZDfXB8jiat3fCZ4HV0xH6aXklP6
9IUTszznV2JTtVlQtF4RURjXQ9Vd8jKd5vutYULbxYDKdxOi31ePYhSSxGOCI4//BTeGUAk+KBnW
2FWiGH8yOqdUPyCU1Vbe00IuZHQ6BeOV2NIHA1AGmhWuYk6x7KkI9hqQBaLwlR0ogRLgKVGM306r
pjPakQg93QxT317+UBhQiZiho8wKI+34/Zus49BPrLbYRtw/5W2+lUiJ25y0BqMQeHUIc8GFz4If
hxi/svUJngxVqXq6NwLpXfysG/a8EdgZ1mLJly/k1ebmjArt5tP+xxhGAunOO1dXyI2+CvvJYlKz
enZMOBdxTo4ZyImbmr1cTHPxc2i+vL8A4ZFdZDPLKW8iqN3WL2G/1La/S9cVnba3mDtIRmc+2+3Q
McGRPG65v/hZOiuFT3WQsfCXJZ6Lzo8dcbLqqbBeLhGSkcrrmH4kBs7LD1w5D6A+hShRGgZPnH6A
wOt402cQjZTeOGDadmjW5EsUv0mb8C0MrDuYKfRObDAa/ZQ7pUagIWDR3BauZxezTQL/npKQO5CJ
qE2QhL9jkW6BieNPby6Scza0PTfkITtiKT3DpJhvqsThVicOSoy9+GUglPGP7xZJFURFSfrhQ0cr
+V8GERIe+PQDPkhA6cDHq+3OJVEwVJMxbxE2ninMEkpw3Kuy3z/nfyxVk8S1O6vx2zW8oLcCE8DH
HvfcyJWPPIyIxuK2R7hac2dduVJuO95rbtQyUX3+3K/ygpMsy5VvPImw++du6ugsXwkYz4fcKP1l
3tuhGrPqzRmuLBk5cONFhSJdsTu8+5++u9iLS+KmPe8CDWhz7BBwiVaocrimj76F8qr7fncrMhr1
mNw4ku/p6Xs7/HNy8Vpv7Q3GBqDSX08MGhUZws7NlC5vXuhkHUCRfqbbdezytecM58Et/z5Bhn4D
RCQXnAdOdrVOby0Ms5v6xa0PA74BCjbKQvDhnjFKk1WoQNmK+7AXmKhrpnmz5FYLFFKTfd45hnn4
expXAUSRzYL28a1IIDvPBq4MAGIJxL2DnMHg+TrxMonOZ7fbwY3Y2EWKzrUfvBjQtZvyV2f/k2wO
f21uQZBOpPfIjj8kXesKY0zH0eT6Nroe0jI1sN78qPfbWO9sOYwxJlBesbbmdVmiLlCXHpvg8ZXr
oES8lUif1imGm6UCe87wSS1IEOc/KaFXrXJ4VwtoB5VkUavwJCpU7y3UR1ssMMKl0/aKS4Qr6Qxu
DSt7pLRXNb2xuuHeWEInc7BfTNTPC/dcDU3N6BgRLO//qL3Rr3pLhlYpdoaCYI3ItELARz18Lc6K
kJORF/gJBxZsQWLxmx02xHQdkYp0DX5D9y3pzbF/7rxv8Yjtj+hHOxdKeJ7LTavqAJa+2/FrRdHa
ZYqQcoNLmrr5h9747oom1LeHVS0Kx/oTxgr/cIPUIsXsiszvDg1j28hIehFEq0MpEYhc1LtmVsG/
NOrBmLuGbgbn0z4zid5GSPh4/j8JEQXt2aJOB8h7uaDlLDWhsm4idD/5ycVt/O8LoLST/IDeRb0h
8NibRFpqYhE0kRurI2qXhVb+qVLPrOfrVV3LygJeWMortRrbHhRS8ntxoduyKanpq2togVuF48nu
hIIKFilWf86vt2X0pyX/dsOlA6KummOkX4eL1KM46MWkKEryJOD5mEaSboMX0SS/JE25mE0Nx7ea
Efrv24rUzomWKtW2QlGH7dUdLPDbslJsdRSW9JviG3fJe9jNuokafMIL5k2Fg5RE9d5Fc/PQJCQP
hWi9txdcrJiADdSfek47sHejYUntJ/2Jq9wg9P51I5SCZsyAJtM836jmSavtY+zxNAdC5pQuGDz3
uu+iUp3DnoAAX3PvrFr31mRfYuoqIojcgOONC8UgkghmT3ITlUKx6PVc5D07hAl4ViD5x3nf307t
cQ/5z8xl0BFoBFuDtk1HeXw2Q7rhI8jDbYIoW+GvLr9fgoQbpBNMbRCNAuTcKVGcOpY/YEQjkVqv
JX1REicB7yZfVod7j6rXbqVR2ZozhxcyjfXEr0TF3I0Ou5uHJzXA/ymKnIZN71S1Mh/ZIvRrqbC4
oVNvKC8L/J1wf1LKSJ6vmzEy65Av9AXTO7upjUMmzWC+eRDVGxaXxYIP+TY/qrmQS5H55oDDjxmb
yaA+pBXDuQk7nTuZ+cLNhiosU0H9rVXRzqFxHX1kdbrQeVMy/Gfyd5K+lHRDp+aZYS1xg6ykOnfx
6Hrq81Zm8VyKQY90LzHwJyhAhEU7g2pPvLqAt5RCe2cU8IdiduiOC28HoS8INuGmob7eZRjWrEpy
pMPikQmMin6+8TxnQBkx/s75HV2JuEsu72VrcrIt7BVfM3/X8dH4PzIIORk0KCsacKfCVb7/0i2b
6OAvJRGwDPYAN8Qr0bUJLI8tc3NuCTcwLh4dwoursY7K25LOrgyUMH79DWbsn1+EXTeUCCs+N+hT
k5+XRRj5Ws2JCAS2v2mvccNKXIH8f1I/aQq8fn+G6UEKxdpTXbEwzsb1uiyguJ/Ztha4oKOFvsPa
XhghStCMfEtGjCjRFHOKqHIjtCAUabHDmGjLEiqSnbM/Er7xJ+KdqaYZJt7iNRypTM0Yw9NxURTD
lp6eNSW0X1c8C/nmD5tMrsiq5zFvTF9iLYB/aFWKVW2xtLGv8Q3tYuLfGOJKdI8OgwG51BIXONy3
Hdhn1LXW8+S28tGtO+KymhaZ+CXiOip3ynf3qsUI0bshP/NAU0m5WckS9rWFz1SmR+yIJqszAm+9
ii78Djy/ZjT6iNcIczNYPajU1lujVLQKaa8+ExYzYvjWxsAdgZR4OHJ5OXUz0RWb2mrYyNAma/A9
LdnPOfFkam0gTRcaeUR9+yeJRQy8jygJuZyYnbI8bSCZ8AFDimQIxoW20mncDsKUMKPbiHx51s5z
Depgh6GDFEQ3izXwRduFrW84GtYBnaCeDjqg4GQEWZB5f0MNMIo9yFWfLyRBEFVB7u9UHaB9x5Jn
ofKe9YFh8DJAapMvUsF8mwt+GvH6/TwhDJ9FIF/ucSSu3wqlULoVCdVkR1uqbcIr5sVf8HsvRL04
RYoqzQlWieRAvwTCtoLgh+HPkjByC9IU3iw1DH8tECi546g7IV43bhtC0/WUNrm8bzWm1yh1zsqf
jFrdc4z+dvdho/pxQ5bzuMT7rOoAbfJDr4809BvD3MlHHHp696I2yJTLXq+BktJh9h29AfcM5mvd
ve+MPVTnIBCsc950WdLzpEB3g62nDWGoEtj2X4NWfxgDPDgZSNiIyHhpF8bdjrdJPsVuZBVS5uYe
rDrmonUosQ7mdlSN+or3BBGoUWfY3qSvHCU8dtSJRxs4qEoEDTL3SLXRanjSHS9MYf8cqKYrAPVp
Jx0BUbWjHxHyQffDsi04KgfURV8x7B0GRi+RZfhO7wYIpd39CGzuCl0Uf5kDXXtn7RiLmoc2wN2M
O8Lqr4PUIgAzhPEwsKgVcV9AUsh5ibgQV3sJwmSglrDtyiobURsYrEhGdur4WnxiPV8ADiOjbBFB
KCyN/G2gWihD/K0WgddI7lChzPG1oXTRcvWvqaYkNeNf3l9pipnhyJWuMp/IfJqaPPZ0OV0Kl+NC
lnx5KqTgtuYn/g8ZeKth4nzBt7K9oTOROschbVm31mgYSAExKUmm/cNPCTbT7boBhztPNAi44GM9
1cA4xtVoLtkI1i2NJIdSBzQhtd00EUY0BU342abvXpkWy5+eO+9RsQm6yFmH7eAHvZaUv3b2X/SL
6/9bg2PlmLKXtDqpPeycoE4z/gP07FyXG5IAWowuGzzjJ9yKJANgKVvXY1z2rIwT0g94eNcyzfZp
QQDc6zHiNyfq2I8F2ge3S3Zzzbhkrt6yAkXsbyKWrtNxWXYvN3RjcsZ2JrnkUJ2gHU+8cFoCysM5
23IiWKDvYl8qQk7Spb1r410ou0m1k+L/JZ/jOf0fpnLn7znw0jdJBMjVPaOBKVj6fFKr0+fFcwBl
K8v/SZjuGL0qHlHKEkAANV970d1vSHy4cO/1z8vvwW9O3Ecw3VTNzARcOa+rUPio0sdOQSyqEQRT
MVtTS1P/CHHXQaln1Jc6uyBXeiA44CSpBhNGjBtauM7t4zRtlx/xOvEjuFtwSn8cYc2whpmU0C2G
atmRruyUhRjy8WrePSuuFeEuS8N80WheKKQUikqAKSRUGy73oRvkmLqZg5M1dQY00udXdPTDY3DW
lknAv25myxGHGv8uCR7ApZhQW1nbQANnHNrZtW57jr3UxuehKwwgZH3HrlirVOJUN5iUFWHw8GdU
NYAHMattqFTMu6v6yETL/2BV+2+8zZpNFpkGg8dWnCHwGTgw7/orzVeUyn146bKIn5BSEN/jhL12
k0RSYQ2YwkiLH+DujUS0pE+l1L7BYOwXOo8LSnNmqo9fhkKP+HdUiKveFz/uQMH1nSPcQNr+fRC2
S05AKRJcu6NE4EI5KgGQ/7Mb1HoJamMFsbW71mqHVMdsjUqprh7LuEHCKv35hSxTcU+qD2ooR/ch
rs7L4xz03TkaaBjST/wyMJiw5SVffSKJ7l6lgfXbzFRRFAnfYtDmo6Vx3KrOlKOwvD/zK68VFk4O
glHsf8SYgBE/APuhO4vsvODULCwKTRkKW3agL3xX+9hpIt6TzcD6bLwfw5gmHZ0bFQCqaIMnRgvn
DEoCBOaxGONNJ5coDQ3sV6/iU/jQHXqaMgYAOfLDdywu3EeP6BNYOpbqwTmSTjW7ZnwLJmpFTD6j
vpukoilTZdhk4qIjp7z5Rqi3kvctp9TJ1XPQ1UPUCZMSSLlaBIwIq/z+MKRwQsOdBMHwjxPP2SUw
woF1YqEtdn+Sr5MhzqA2ybwYtays2V8bkpjEm6l3NUSPa2PtDMR6yg2wlJgeVLY8vYKg3+vuF3JC
H9+NmVtpNwDSMsZl3qSihQkXEgpRpxbS3B5smiIZuppoCIPqssTtcNUqtdUA61UfG6PGTDdZnSx3
GNcUxzUdhRjHpWVb60PTNkWc3DiuuQ45UM5VEGldkgOF4CwwSvgK+6cLHtp0FQok8qiO9XE1SWhJ
WPLHCqJGkBhTSeoT7gNf/oHhBqH/1wYV/LJfSf25HNkeMIF2MUjKW5pMMH6dlCBkcas/T2fouRpR
aORaMI44S81fdcIV491/QB9QJ/DPzLjSyOUOpAXxMWYCw1xNRCIBpg2uZQKXaRUg2loACn3GFX7D
N8Kv38lsadx8iRJysbB7qD8o73WpXTEgPvqI+DiKn4TKJwE5EUtGW0CynUDGDofC78QO36ygLP+B
+9QF2PSLlOh3L7hN662L5LhubiqiEsflabaE+poFrTsfok8cRjXqE4wy2zqfsi3PhaP3s3HWEODY
qEsEfg0BOe6wByDFeTLJJx7MauYvoMR1GvAxBqyiMix/5vvFryEvQH5ujU4YvRcIkroehqYalmmO
KO+1aF45xbFHlWVOS75SgZYJH3VCAdY+yoMKXzrEGPof8Z7/xXU0l/FCLGRi2+frCDoOZYl+/IFZ
4D9E4EIx6fSRtmaKfPbzP5xWhffjx3bqnuoBqzwHqp6ZCL/KctJ0ls6glqr0k0MkD75F/5mpriZ+
sX3JVqj/LSGhCQIjQWLXfrvApQHxsHjZzQ+TiheSNl4gGDIqBoXAf8MioB+gBUBxkCmmToxHe3ze
c8dyX59efpho+RIvRglHWwxKeNep1omkDFpx4hr8gCc4eU/ckryUm5np5BD936QgVaYV8FHbwDVU
vLb7eRimxbo/1fkE7T2XwSVnhbjrnmL8BoXhMhs/D02gWmBOLcPWm9V7qa4mxoB/MLHS2p66UGp4
88pyMJMR4XdkB8rCfVRuhTBczk75a7OrPp+DrXNUo4QxboE9i1fjwoXD/qTi0oQxxYc53Efyu6NB
x2rGRfQSF/7vjbSvxKeKCyTvi3llxcr73FJdj3sSXU5m3IcoB5vOC/RgYhp3iw3UDyEksYQ1IFy5
jnl0cpGXtjnOy6Dx5o2ff1EpFjeHesEwV0nteguMiA/p4yWxtkhWVyP8GNRcjCzaPEOxWOHb/Tmo
dgPvL7B6GE1+iQNFURpPKT5Wcku41OGzKGWFWeOQFsiB638nPhfSzp7qYKaVm8eu9pCov0Y/99ko
C93RtsG8T43OeXye/mJgzL4su5BwfrkLWYeCAO+f4N44u+ceoTI7j72KwXFoTeIQUEpcevi6e1pU
FUtPRclUt0yW0T3df4dUDyXdocv5JTweMd/maT5PFWIeU6HMi7tfrQ4Qg0aZH4ptWSvnvc3qPwxh
XrVYcAt7Fk/ywFPjIxgycEN/1JD+oL3IcLKrK0MeR60GXCCT1tccv72DbZALQ9a96osAPf5x1Xwg
Sv11NhKopSEt5AQH+p2/OShS3Q0damKnbo2e6osu7vU9Zk3ayaTVRwX5u67Gi0lC4j/tGMWAqPQs
cyoJ7TBbiFNCRybiK98SUnS25YWI60YwI9937Ez70jTMIthbvyNPO2DjCbdbAW8IzN++FqfAGwLp
Z/KghfgOssNeC8GRm2r7CQ1U9H+9n26J6/bypCcAc007P6ww5en4zPTNxDaIP//7R9UroP6Yjp1P
42HLkQBr/Tq/aBGXdvtAjCiO4qyMMqZ5DnVPwB31ze7V1wnDPKrDZAKFNWLw2v6eOnmitxvnxfGa
DWLDrIkXhvU9ZUkYkH8+mGd0fXwz7jnfYfO2D6hCtf78kJA4Ubmi5laN0yPXG4jRwgPsktUDvqJQ
5E6z166M/nEAHFE/lvUiTRdOBRDOa29qBT3kBK+3KDlufEbjBMKZRgr4vyOp6/Ojy6km0W+lxWFM
0MFslpt/tFMk+Ji80DdjVCQoDFmh9FWnbGCGOl0J7jpBupIepVdE86+Z66doo/84yhkar2e6u0k8
XXLnKCuSnAhCToGw190/Ao1U/hK/JQs9qqdYTYBDDjzMmFKwqO9IsyJtbUbKM6MwsLu5PHeFm1Og
zclDwq87vppwPPUpvOuadjFypiezuTd5K8m5+TItKKPyQJlM5qYtr5WRzPBHsBrTI3qqnxB0PS2t
bZRnc0cKDx/2/qenSy3LWplxT7uDwUVAORobBCyNUB7P6LUnvqpjwz5mZUoYqo1ieK2XJAhbp1EW
ecqWMVld+RYpy2zH2jSE95iZH3EBZnJs9aAPqs3zptsjVjWRWNPsMNN/Hxeg+anm/0WuOfgoCnM/
9bXmU4Rsx1VxAlHfT+ebTPvfawohXylkdApdPdVwbD+bH1N//bf9EgR8aLJ1rSrxuaCUXrX+gG/S
VrbI1/1RgIJxHM/HNa03qYqZOhgZw4/BB4aYGjRd+TmuUiWsuKs1RU3rgeO5moqEhi5jUlO+Z2I9
STc7Rw4xMf7eEqhAqA5U4xbfbW++CxGedkx+PzFTE/wAs7O/2NbbstR6YTkKxlvkgc+IZvfGUAIs
JCUs6untbCDBPe6Ef36Fco1X7MyAXB6n5SkTWoI+GCEFyUlOsGtyfR7fGmeBJfo2jWDEdEdPqBiT
HXpDj1XGYCEDKXd7no1FL1vTnuKR79JaJP5CB+kCsLQxV1hIWV0phb0QGJEwVdEtfobLZsaV0SOj
fcnC9yMAC1eErPcs7qf+zGwvZjQEGgh6T6mfXESJ3TKteoKKCGf3XEd7e5k/6kocKuZXjN8IQcJl
Z3M+P5ltFNs54KfoqihJOS3oxK7ncjYDuNgnoPd5P1ElVyUBiFgGAp1pcCmlPXB0wLkBZRE/PJC4
dqqh+t9Juwwy43aA2/531WGcRLy4NqU0PtZnoa5qCxoHKjQ2lIva4YVlSRVq1vX2ITbNUgjm7lJr
KrYq4tEyJvGd7FIGRHU4IsspifuBZxC8dFjUMOlGrh22I0TWPW4zGskDTadnP8NZ5b8GqrGlgvpO
WasdQNYVL16Ni+DhZlvylVn/dabqhZ19QSEKU6Fmv3NUtX06HV0J5ngu0T0UuvTqbxUzhR49JHDb
CUoe7M/rUWEKxgqzgrifU/uJaekEKrsQ/jrFEg5eifBtoulLh1DN4SMSfJw017EAV/YXF/F7vzMK
16cI4437sRecg1H2YGfUADOK1SfWDszJk20ILeC/GlmKWH++dw9PC7SCTW+SnBo2DxlFJ2EEkPvS
c4P1JUWvc4dGDJnUjX13TPG0gDAfF03wk0xqcZIcr6HOdy5nOi4ModxohVVrHgoxcSYnOe0UWN+r
iw8SlYs7y7OmapYbXSGn7aOKfV+FDLInIS+xPJrjhpuETuCX/q/Ynp2iBeh598RlxuwDI1yQUsbp
thpzYK8bksnzOv5z0whO1Tb5X3hlO8WouRfrU/C3sa0pJMHXmqJA4pBa/06TFb47xYZuB+lHR9LD
fmi8vAYRadEUNVMqnv3X7C/EdImVV3ZHwbHs3ENBnu2P6zSDufmna86nJTdy/9rm4omB6qB6mN6R
rvXP8V6vkP4vf+KrtO9Jn0RxbQb4jvql8sfpPDlKN4vqh5s8tsWeYk/1a/+h19DrZFdVqb0KIKgW
mTdLOfZ7KOXIUmuZTs5zv87eyths5yycXfcb22tKWp1MAka5m1mDovbhWB6NVOiuoyMCaDQOmZfO
4p3LTfdhzoN/WGBZvnuq2c/xOxQSBY98uUEvTSM2RLzCdXbS5WT0raPEyingoOyA+WiNZ8oXi3dB
1P8FgHpAYpng+XxteSryY6tasFxHtOkk19uqGJ1RQ+AxwLA3678vi2I3iN/soQiVBwz2QIHpkTY5
7Ccnc1rCIEFNhJMxbXzfIP97wi76p+/C1aurESEaf8dQ1fsRvkbUnsl8al16578I19TeR4ZdxY1Q
usc1jQ7lSyf2EANrI1UYMa+EAOSNz6urHXN3nEP6wuXoWBbQe/T7xh5P5GbuRsDQ4zGpBimAiROc
i+SdQ3MNUhJ3o4aBOa6AqAW6fjmAyqLJIy570TP4aC9Ldm5n9cd6uao1OpYCtyHz5Ar+WU2s/9ny
XLZudq7YRqzolrXrQ5AbrH5wqiZDYXVmXbzqgT1Zh9OFJ+eFP8JAOmGqG2pzIP6y4OxdTAOlNlWQ
WhZxNQINAnH6mNhInbBtGy/Biqt0tWPRN8FgrU60FUGE7N59NgXs5Xk9LpznOMJ9CMdxu/Eb0jgS
743Dwuva32TmkqNmphhfDkLpBrPDHjhL1GGj7CcTU5qHZ3dHncvsrFB8OY0Q3SOlm4pG8yUgJRFm
MrAqzFyZq3tBKZexZdE3z2bOfHne8lFzIp0MkRThAWV+ElAmbau1AJSDuKgmJ6Q7UVCnemeMzboL
i48ZFxHaOK7NsMtVBWVXmnN4iebnEoFZqvYdy2phl02NuoH1qiIkSTTTwgq0/vynW91eOIJSxhJJ
d7S5eQztxzDIHzH+I/DlqGok+TRqUT7yTmlBaixUqrZJTY0uE6IEQ7epVsOYuCWL5FCAYzoSwrCp
TMOITj8Tqn04oI/4Gpa3xGqHWW+0ywFzliNAaWou4p3GN0WKHT+xt/qde4MTOyanzqAt4SayluRn
QB0bi68nJ6Lu+zX2fzwuooqDSvdrrSDrQxwU70pMTB+JA2zXJS4w+WUAiySRYTJ9d2vJkYbrZU/7
GRww9NRmGzyjQ2P9GCgK4dvIETZwCoHtxbOjqA7ckJDs+zwyqI7ub7jX6vfTs9YarhCj+tSWJGAH
RDq2iAhekSHIg3mv/jHAuQDZL5d4A02OB4scMbtNRWDSXzGWj5nxttMOo9VjDGS7yey4lSIL+UWM
rwObDDGU/V1uE4uJlKfTa2sWSR0+Ff3cSPNh7iGPSFBa547Tzu+x3s/aksbhY1+ZPpfL99zcA4/I
tBleSzjQKky9DOQJ8td/MJ/YPDDLw5munLAed4cuJCv4kbOpwzNPle7inFH2CUEbAqo5ChBklbdY
NoF9bw2PC1v14gkaiG4GfS4J/ZIeg3IXKHcEKwg2IvXt3m1poCHksXeSBWAsHM28p6PSR08jGfov
plvLElR5xtWi9rSxM2rsh6tQOyYCoUZ5e7i5yKd7Qm0d773n6xHh5T+6c2L9DV8JwRYu2MsVqZlJ
SWk2lm+Jo2g0Eq6Bjfu73lKfN5W4fKRwey5GbijNpkO6EbywTV4g0Oynk/7XhTur/InoGPAci6Wd
HkHMNk1uYGt5c4Y4GRdTTomf2SNjRh3ccGOgJrzQCxVOISGmOid6wU3bzqjwLefxuH7n/zP6tx0O
rFxZqmL7wPrs3PuQrdcI18zSxqUS4vqnGf1aIl4Pgeii66DTmFNIc6Vx9Y6kOZ1yx1d9U9iLKrUu
l5y/JB9BOtpJ4lUZZlbVuqNcBBKOOlwMB9Jj6ZIWyYUNoVKlXS61cNpovvUKpW4oSkK7P43hwbvX
NB9ERMEjMi/Bl5oo6I9NGo6AwogTG1wpZ4YU08UXgQeHBKGLqSGT0N1vgd2QAqHkhl0FI+V2/LAF
/XbvOUJqorLtJvoFjGRyJ5MH7D3U10seMh24ub/3jHveAfcT6gyNqGw7D+IXJ/eytsEdF3grADea
klWUGCPqwqUE3PGkDhl2jkSFUo+CoZnssfWTRG3wCywkqviXKfTtOFIjvpFRbzENrxxb/ADc29Po
Ff58CeUvIZl7jzjkggFnPi3js8+eecrsIXzfXICXE1KwHvsMXPagYW1BZjPBvDHYQEdJAW7oaaIB
wsyW4yWlsSF157ZPhKZQi8muw4iK15PDQnHb/7WVJ40HBQ6GSN9Mzr/kyTuKmqmUiEE6cc+Eogt+
pjZ0cf+fWKe0K24Wi/WvN2QqKkqAs+iFsmL6CcYK8rGurNTlefUxNCwiLG5c91wv7wo5FNF4yqDc
25Sve12ty5wkR28nMzX0dp6b9EhmCGUsW7gRAMob0vM7JU01REWykej7c27VLFWi4GbUcjFdCbRX
AMIlZaLQzsTwJ5aPvmwnujdNEvHIZTRtotbwRqmccVSCR1aJeSg0TgoY5RIPiy/mixSKtGUzd5wo
ekHEy9cTxNlzoK2qaWM3nwsEmh8O/oAFTxFxOnUyIh68LfJaLj/nZJPKiBIegOsPKLrvVNt4Ne8G
0721MDgvMFAQqXQCGlOpTnrj/LKI0kHblP8yycLT6fQVmzvWWzlmjfMYbb748ISzkhqYjga7jYAn
EOP2bntBdP8DXBqQhJm16A0Ye9MGr9RdkrVjUlBk+lMLgdma7AjyArvjC3YY28a/V7eeQCxW5K7W
CGnUhsotYq7xvtbLhS7Wmr/1g0+pF1ak+9VVF6+MEvZTEbpSzb1lq5U/0S/c9c7Xvht11cBMzfV0
Wi2QDoBJUWQtUNchLPEsput3M5Omgi3iZoO5zm+Qx1bSDiord/lEHBqZPH0C4ytztBf/4gvKTryM
Vy9exv+bfsaZYUPkJRkha9k2LiyHfTQ/uB5E7GdLBS7BgprBYJFP8MwSPC3KimO+p4RaJYQES3Vc
ewl/6A0kg3ojINdNL1mxc3uqyO7ayqvA6z5A+siYDYSHetnlhjguTS32iOqnA3ym0d5gTksZa5QA
x8Fvp4FTJ4tD3cJIoZkBqkKndo20HL8giEPJJ8ZSN7VBWJ8qXW9jWOV6XLc2DxqmpNsIReM2EHj4
j7TsozWR8IqCZe6yoTM5jMWUWf3aRIdT7HSBuujOwUEqjxUyoggvajQSKPYU5K/qkh2WxNhXifjl
f41DBmGYs6BjJ3tvl/qre+cG2i8Y4QJfe9LFvK70/qLozB4W9oAH0HoMPeuEVCbXONZlvELMhVBZ
DIeQDzdvYa0gc21s+7fY+KCzGi3CpzNJmvC6I7/J3spYUjsi0ZT7lZusA69ljM5Fg77vLMW+stPm
HcymVkjP8f3lNV1k/+23qWBE9VRmLGN+HmW9yXc4F0pJdcV5VcA+vfrpD7ypnTcs9j5Df/HrlpSd
2IRrEMAt+WR9Nc6sbsPQn6yrsWF8LSZDZh4Ab3yW8Acwn1cXe5e7toKItp0QH9VbsKIZ//S4z2AI
Ue8TO7BAzHc8Kxbk9nvCGEnKJMjSIyP5yyLQEaF35LjG7XpCWeJYwZSqVPr5oxmA/Y9T12DN+VLv
Yes8OXIeOrEWNIFtx+cnJk2NQ+2mvrkOSdzvsWE8dluGMg4CfTVZFfART0f31PQqT7Fj41ZPdCkV
8/vR7tC5vegnu6O87aBP+zLwjYYXzRCaJmWTtNrf6D1iOiwtoAA/1O3UP4h4HBLfJEHmyPn3PKd+
qGU0XYPQ2FbtX3pzoHSTDbMAJ+67OtHlSpDS7PPi4THh2/R8IU9p9km94geQM0zI9MxntebzAeK4
Lg8GXLpagSeCizRHV95tgVfStAeYrA6mxbZSrBsJW6gwAYFWket59xmiDX8x/AXTm4Q3/Q74mZYd
V2U10Be+TyOmXLyTaNlf0NgRMImeQQFTo/ceAKD3+D8sNYjQyA8ZnbEeqEtcxI02dnCf+fZjGUPg
e1jFhejFyi/Y4FR131VXMM2fcAH1j7s3raMVlO5HIZl/l3JqlhcTyQq1MFmz3a2l84EixZn472fv
uBtQQt45PaI7tgVHrIeq94ZmO34KCyzxTn61PUpWUHV22HLUAfQLFKcc+TnjKwphK4q1kbx/Vbxw
mHjm7qdrKxp233x+I31dv+Q/dDtcXDIkqnU6i+7CafoLOB9q+ez03B2m18lTGCFEB74Ottf5yoq6
m5lBRpAQ97tCPDB+X8IRClAchPIdQ+nYmb0yOUQdai24kfQLn79uChhyLAsacrHpSGvWoUfueYv/
FxilYbzyGVeEiKX440aMEL+CWBgLsUZ8DhZMuvHrx2uZYC0fSY/taSvqA9hW2c/FQXEL0TVhRLf9
NhYnfmMbVfCX9C2btfhtqi54LAyKanMdj7nwstixiBOidYj7KUCs1oryQxMAJEHkfL7f2fQvG6fg
ucAQQm0+wp4PHxTfvKiOzIs7EHUAVQjLjCxhUxsch4vGGQeKYJ7QkgJTRSX2xCfEnB1Lj9JY8KPX
+MkMAlxlrTLPdbzFm2Rz84ZG8m7ekEHzQGL67D9Fg1ftkBWEH28sF6maj/oRQnxEBDIScDZLFijg
icUskPMNpM1/3k9XPlKqIoCcEp+0nXaRjHB+lqhwxOk9V8F8Ve0b8l27qA+koSeJoy8t7EbTO0DF
1ia4+wKE/ayJi/0fr50jhnJqhWJ2u+b6SYCgthdswE0GPVNFcNoggooQYTx0/6MZ0D7JAxom5O34
KxipuHQ0TrGcWqEUzQGrG/+PRGlLqSlLOA2oQ8iTN3mr9nq9Rfl2yw9lPq/4SRBG0SIIzEcc2Mb+
kdH9rhoQ0aoMmZTzHPtcCXQ0tFzOzceWzRcl1l1htoenaEGXVmf3p/QkoCeOUAzy0ci8hSuRwX3v
zH2ET/Vb9ZFGX+jd4+PAw1kqPIgzbr71esPvO/bezsBoynUBSzMMLW6qdxV6fFwGJ+hInuDTS9+3
h76sqynzzBG8suMJlsFUZE9MDpuc/+9ra8GKgRHy5vjvY6iLoWITO9nmFtQwXVJjcJwXf2OOD9zX
2bdZwf90i5Fb44K/TO81bmz4Xzn6qZJAZCyN4ETrqh6APbJhXyNUu4MlkVT0iliOL90ES4R4SkxL
tKtJHBzjPSvqGMqP5FaJmSPf4JaG4JmBLtXI4Ya4OmTNsn49VyjgV60CR0wLAbpYFMImKFF5h7DR
nddJin9QCB5HfNjkxEuqIqVBRk08GTgfOhBBdf/pACg4DAk2UMQD5XGH4ZTx6S+tuhXsxZUQkojj
BEjMQSsPwmWv23S2XG2e1ME4w2q+A94EzajMObeVsocXepxLTWl9ygSuJRzwkhpTGVSV9J+ykK56
uBVjO77TOr/keI9EBV2/L1mmMbr8OCUKN7nLwYn/qaetct5PE15RJGSpwDqfJ69JFT+cjwgiea3h
LEA316wGU92+OFvkiH+kNfXj6s1rf7fTGURFbwwGkvzzOp/YgpPbJpc2ugTnOCOtyoATYIupJkYE
0i6BNQkZMOdTs6e8mRCqutjWlqFXdyEyHy7OSJFmjoUwZ13gDL2+TLoyw2+LDi25UCmYNbM/RVrC
unSPQnnKslP+Z+Xh5ohyz/UkMhjfk26L47N9WR1FsN4I5NFfnT66HNDqB1G5pIT9yTT8pzhUOrZb
hQ7XwIPGlxvgpdoC1r3bqzT8V1sIJasMhLxIm7egzlIOSaKWMUjFzqSwBt/nesvaiGA5G/KPjI6Y
PTeo6KRF1xMS+VbvArK6nF7tJ3xmEiAvpiUTHFpBqREn3QXHfAiyyA0WYU27WlK2jetxo4hzV2vR
GqUypD5xJLIZdDX82GDZG1XVN8gd4o2WJp0W2d7rpoUP+6PdQqdeQYZNmI4fJZndKgUEuJBgFV5m
dy+aKY/pPa8ETI5iNWt3F9i5lWm5fKZWGrnb2EBDzyVE3RUyyYTvP8ZhX21stgpIgr+znAoufDQ9
ooWy1TXhZJDEiV1hRGsdGpF1RyTeLBMyOMgCUupT7Nu3OCx+RFQzjr0/vbzog0BKGCBOc4mjLsnP
ZcNa/fUyQ65VOaQKG5cABKsmS3OQ0I5j/P4I10dhtHqx2c9tfu3EkX3952iHekmzcPi+RxDUG7st
70tAwZGrb2n3Sfgcalt1JORMqbbhnziQXRAWjSicG8KnEWW2RGngFIaZw+eofBeFpdq4G2xT1Nsy
gcJ0Djn0yMPuk9vd++HUXzGfKySbXoC9WMdw/4ZwizxN145ohRilu54FndaUnCF3phpa0gYitNsh
JqNSeusfysYSBMF6pekiFkUL1qPGwZ7rMvLNUM9i5bidOFEb3KYYJAuTo00nYARaPNjPbq8H4VQT
RW5vBmY5HfrexcNE671yY8YdNuiXYurjveBtx8qzceyXvO1KhLBXEL8KNvDICeLHC/QqC2KsmswE
peNiCGjM3ULAQUUyyWrjgIdbFEDR5me+WojfqcRG+AxgkNkocQsN5OlGFpG2iUGqhrmPjn9LjEH4
CMw3MbuSVrVBuzuQQa6MqF0WodPhBINB7eedGN2/r0XnS4CoxIR9XKGt47txfl3AWkINij6LxTOH
vnvdYPQSFDo814wvA5L/WBiZESFvVhidXdyhUN4SUkGRT0+GpDoAa9HER6zbBEpafy+ZYNErhr+6
smhWxiekKmWxegr2Lbns6VaQtNXIyMPF6e3kZ/r0h0O+SOseLeL7GXSL0HjsDO0gZPvLTvc/Kwfb
RKwboMELSy/DtrfcolT2eK/WJ5pUIhSyNGsHL0QN7Ws5Mt+X9n47/skLw47dhjrI6CcUZfs0/rR4
78/kRutP8I+Fo6Qz8L9CC7BCKSPUOk/zf8opngFNoCTVszWKA4YXAbyPB1+65cutblb4mSpzmydz
/ZFo9zwm1pHxv0hgN0f6hO7ewG5qfnO5sTADeJPg57KkLg2VT0w3h3IZtp4sHSjE7y0kS79keLoi
Hb/o+1zrqyHNRMUFDkIZHr3hWjQYMuyJ0CJGdnTsIShkCuSOAieVcMkgUY0eVJaR4Blqu3o+VS5B
pRyqgAwd2G7onw+jwksILX5S+p/TF9WZxwxlPwbaUsDPQ4wYsVHI2mGt+F3dhjvxa2/nPCKC2326
MpWI7Hp2eglc0OWyVVK/a5DZQ8rJSVvBi73DmoipV+0/rw+4PsXm2qj6xeFrKXljZEGf6L83lTJy
R+30O1SOBLr+ahrEr+RsIlQIDluAOw7B9vFGce8uXn0brarPfU7KOknwYlYV49gyyHaoibiwcnDa
/SquHr18GzLgCGqzlHc2SxyjaNfYMDdCKAU5Fj7XjTLaTcsawbeKiKMo8brCTQr5R1D5jxNrIEiG
v+yll2HeHmgqUvnab0OJyjoys9psFAvJ7E+NC0eQZVNRNLyp4eJ9EHUkSTbxNwNByhJrdAkHi9Ve
UKWuX8rULKMlgP0u4evqtJZPwvYKO30yA2f+uwpbLMEI2jnP26yPBWDqNQh8NOHToURlE7mpuip/
n4D93R/Be+Uu/ipa4NAbbnU775k9qMsSd2JGXezI9gIh4Kzm+3cfszh5vXe4nvtEAeKPXNXcDU5R
bR8r6wLkxlWifAnoqxik546nEqGHHDNm9w6o8VGsJqYC03D8X++jtML4qiioh3QxbbWV5GyXh+k7
TEy4Qd2uS3kLdXlj8eW+cFkEcFTRB8TQkfC8YEC8AtJPeKj8dgFSKAIlSsPl+99LGfsHeJHtZoGL
6HCALeLdO+KC+JXkbHs7/s3BVGpFMRkyBULstfbGQOiSE+bRYV6f3in06tLQUYwLzkMKLVU/2hPe
EANB50It8vawstr7xek4xAvo92OyxMKWFcVWDywPwBYwzEp8PEyNozNFRCq6+kAOn/9N4MtEsuPL
8PmKZk5J0lNyA1BP4CvjU1YjZWGwyIN8qPWGPOMyGWKuFOeG5P8pGBZKH26ZMbftfoGSYi2bM9uT
HcWvNaNvG4ipPxF/PZrX+gG0akjJon2rmP94/E8XU/7161JT8SbcYH1fI6LGHfsl77Cc18uT0iDw
YJoiNXd6a6pkk/3T2k/4J6gjjoW1y8iE89y0yt5elW79ptsS97okPXr/W3Qnmh91EMl00Sxng8gO
uyAzUqzG8IRXOn+w9TcYCYWjzZP5Vu0/Gc2kgoBtOmQLB8no7XI6q0fKOPz0/r4OniWdJS41xQQB
2JoLeneALz8zh/vL17Ba+A/9fyesx4jeBIe6y/Ynxh7oH6rXFMYSJnFUQxL80/BfbqVbnczODc1G
9J24q/jcBfaJU7UNuFlTbxQ7NGStWiUn3Hdoi/QM68tFCUwwPh/JrF9rqEeD6UUSxkJ1sR/9624X
TzC1kgbdWBq9zUQZc8FwhEkRFrLcqGKrbBw5GZ1T/f1ZqB32nIhcHU7gQeW7Lt3AcIrEcZaIXeBU
W0Nx4XQuidNFzClvO+WF0sAWz+wqk+ZuPd3b05wYN8tTTK3LGKHkRaG4TSNTyDtEEAbGLfFGIelo
o9Ea0mwc/DRVzHeG67+ysuJtvuGqIqSIchWRHfQhLC0pKS4Ld9kd2wgvZG6xvjiV/5m8E96Aqnzf
mdE7vFdQq+l2p/5AF3CbcA1pqW/J++crnrh/vEuOysplkMLBIsplSMhoYm1j7XExrMQgIFROkCD0
CgWQLcdW/c/8mTZXh2ND5D/1sCjyBLa2QQyzQgfaQ8urvK+UPlNVAaxG1altao3m844yq/ssnP1N
yLan6EEbvRRU1kcGHNMcEg7LxYlm6G8/tXWlWxdi8iL6jtMD/blYgR2hLOUfN8Qq2LsT5fK4JdQJ
44zHBwz3I9iy5eyqa4kFy7ofxKz55sy6mZoB8Zmbz0CanAfKw7x8qDtpGsokBdiMDyElU4zMmMPp
fCZr6Sl5tHSLDyJKOYft8yjG8M4ewdih1fI6NcxiXUYpaNX2km00W6oLWdfq/T76DclqJtySffiI
kmU4fh2inXpLKRfad6/hBr2pEk1nxOw4iA8Go/spnswbcuCCsNAAXQbpaQ+wUTDRMUFnQIagwkog
6vMu0uZ04s8UykCJWMJgrV4iVIpCl0gYf5yy0YKQPVyLb4VX34ffwzDPsO0A6962CAxGZqpu7dRy
rXcnLTECdHgCOwzC2Hgz27PK/VMFlfHJvvCubJbwkWasAoIm6ejwQa+4viKtRBcuedGrquMMeYAp
Q9holCEEz4+K8wOIg5Ca9A16K75UNFFR1Qj5aCX6siKZ3b5VXDWYnUun6ozkAd5AcJgRplV7y+iM
anCP55PJhEoNkxd4X0ZmoqmRqnEv+1WLZWKOzeYIZjnLr1oBuzshrDFVragDqkFIQXLwOvjtsNK3
qS9rhLISIZtZhVTiZJY/Zqb7aXaGEslOOWW6ZywbxsHWCXPmV3lrg1T2R/vWQkNRPKTIxjPbcDRd
ziesbgi1CU0u9xyNV/aoNWXwfVRp6+iE7lwJiP3LoeUXfZZ+nw1eUJqDTTgoQVqfvWgiT/i2iDL2
qRZxyIOEDYnT5PVnh96m+j9hR6qUTbH/ylnZ37hZ30fOzjVPxrLaAP0DgwB53AEZs87qrOUB651K
e/U76AmmDTvUwEh2j9bbpMk+hucNXIUr4jY36oFGFRW9vJRS/LVW7IzcO2kMO34wZ7+DqJYk5m69
7kbllWfBeYu+rJEJZlIFV3NOkrAqyE6/QPzNaFNfhNJ+g5TH8Bft20aclOD21tVQ4nqaO0sm/H/7
EAt6ICMmTmnvuOcVm4MdddEZ04HsJ29m9aAS2Q7S2pxuQetRMVGze4Mv2DmKDExP99kavczAjBMo
UNyqEA+iXS2zIpB37/JYP6LeRHp0HzxsVVDfZu56QuTbbz3dMB2i5HblhoqH0wy0YQp5aqJohC8T
LWKLAjI56utcPrTE776mrWV842TK04TTdPS15Q1Lr1vpcUiDDtuxzKxKJlG4TvTW9IEbmH8B1MkL
zNKzfkmHjT0oqNCM/Bxl9JaxJSmNwFhW0pq7+fx7rPsOlmzOAB+2RIm512KeZSUW33i1hq9DocJj
OJRpRhQVXyF1gYWA/NPhs7aemQtRQW+mU/rH4IlFYji+Ey3DtQwWmEO+1tvUY+hOgH27RZLRaOKX
9UtkoZgxRw6jtXTd0qKdM2oBir1Q8FS3a+FjJlNBHduexW7t4+aaPD/DuSHEbFTILu0Rpy7eO3Ql
hxthYHgtLuzYpulanmgIlJwaZ5h975BjgL1AOnp2KuGDMn+CHE7VMB/uW8BoKEMvb4fsMz4LEb0c
X/3l/xGsDjLXSra61aJWCtEQdnQJ0NTr8/HZlblGjqhyYahCBTBZ5xSJDkSD3l5BWZaGIfI3gsuU
d2jlGyxbhLGK51pXXGs8bH+A3e7RhHnEMqHjwfHte+BGnfQ1YreMkMrUzFNR1vCgSiUyZgeZhoU/
AFxPQZYpR3fDtsCPWOdl6cxA8G0H9CNYTOqV9hMP+ZQ1r24ilwqkbAWa0kWDmQsUHJ5kR5nwIhjn
kvymU7B/PiF7CDGfSlLokWV75yl+Z/iN3YAB3mg8VdRbyyo4qU/DcQjMWdIqOSDG7DZqcmDwwEq0
qptwLcDIGXMymc6WpgFbbqECRE6f+raW9HUXsOQ3SPStQ3ReC3S7q5ILFtvg2udZ94pDdJk10Nhe
aYJHVeA7BeoG1JmgIqg3tPw5e459adc+QNfFb5xSKS6zn9ja0nGmmOxLrIMU65TMoOgssELyrvUp
M3e5LhYwcutg2n7JdYhk7INimSEdPMZzvviIb3c39ozKbuF99fmyiSAB9HaNNu/EQ2qyfW21SySl
3F4knPSxeTvBCot3t8oXqeKJv0tRViHG0EnzBiUdoFvVd8aTrnqmC9TNPyTWP5rMJzFyv8LhGDNW
n79aOHyUhyT6WlspN5LLYF3aHTPTsWdIMH6XyhIi4TbxwxkZGentmuLVOPGxB9r4Q16E1Dk9Lb8f
1Bt/os7dGHXdQAfeZKTKZ4P1nSVDQ3oLi5mxzW7MKP+W2I+h1GCzygsGMvGqlVhf8cg9v1sWEaFR
ehrssNiOPjnS1mu0QempKt9TyeHHH3VkqivPrsriqh9yAi8sJ9R2qNjGkjfTXW5Z1KHncDUmEDLx
14Lnb0cfxo4smJFqNgyJb08OXe3mhjmr1DLpkSFBd9dZmsoSwYDOAW74aTTUIbupGBUCKAs01Zq/
XsN1xUvZqNKd7+Pp7M0HbPTXJaVQpAofLmU/QFD3aaoA4s30i2MGk2Lz1pbbOeAr/Oc3R3arzsd+
Yiwk79lwdOHGGCPmVpeV8ZDEVhL5JuG941PXp99Qg7Mal+vNSnEXRyoj7hByDRlg9CinbsQ/AC5I
Tf5kej6ltHifqpFQrGDWhGZ6dIV1gJfffraPjAUYIn4rSXeIVjDIYU0wmo36z3c87yOeqLhg8BfZ
LMzmE+P7p5JzKGvrQLXmBddDp1hXI/mGZ6eZmwA82L2RQ41iuvtmk1kuBq+jekX/zfuxf5eKRCd3
clRwfdnqyTso3JTQOA4YxWnxQH4DRLme4iin/IK9dU4kt6JXW74XEz86H7dR+3CWbSam+qXqYXD1
SuXDa5B4cjSCtzsenhj13y9/969FzAWXa+sP/e5z4RCZTb0JZkfE+RNzz9hf/khd8RdzsH4y/Ktx
6oIz9n3x6EY10EhN1gBNok/6TRKGjRk5iOAMOoijwhpeg1OheRFMOhF1iv1r3mPOWa/MXrIErdHd
uk6qpZOMZEHPZeuhO8qblXW5s/6skP5SS5UEsBbDnE+4tFJUfOvOeAMwo5aEQ0FqLnnOYVkD7xIq
nbbq8k3grZJimxtUCsTvGC5MdnBoZbJzEjoebhPx+Eb6X1pHP4oPdeBuiJT42fwgynihT6gky7xE
oRVsVCFZvupxDkl9oOr0iipmV1rMRF2o89rMl2LuUyVkTkkO3aVA1As6++sTHBxdHDx/RYEzHXjM
w3hGvN31eUtdS3LQikzyRxWGrXJYuzdWpOnHEwZdPGCFWM7eG0VvMfP1910aOrTbFVmhhRFH5Hf+
UpAckNNaB+OqrMUooztgLj02SVY7TCE3gQRcHoOcacAXHJhlc83A0UqhhY9KAXWJ+D47SN9IfO73
2diivQEoV8OquZ5K1NRyIu9O0QES+rrM38rsNZvS5SfjTQuLmlnKf99F22l0yQsN7t8PFPcAloMv
ktivBdw2XlDAkfRvKHv/xvtb5osnnJqptYgKaDMfi/NVbMjf/xU0Sp+Vo57EmAuqXWgqnP6VNJXZ
fIoUhqmfHSV2u89V6n5XmV/mI5ezxTkd0lwAimxj31s53RAXNbCr70LvIh+1QFN4NoS+ljXP61F3
1X0o/OKzK6yGLhK3I+jrwfACQXefG16q9X6+OXowe9gB+Wp+UjXqC2Ig3/PHu9n9bNnZsZZ1cA2d
QpBQGK3bF7VvFtyU2WHmNG8D0TV7H1sI8KRYAAV6T6EcO+uEe3mdviixDKPGd2melZgkGUIN1Z6n
/zWD3/rxEiFJ0lILXcfvbnX0YRAy8FdEu6xn0bK6f0x0uPUTEc3F/DT9G6D2prYiT9n2Qd7y+4E0
STRhFIt44BAIPjE+ClOLsA0O7FtcXkPTxz1ZfsXAStAAHeTUSXWaynICPlqamMpcZT2fhmh1ST3I
bMnZo8KFdnvPXb2zZMMdSiz+18assBOmIdyGrGETG5VhNQ3wHndRo+qkIV5b0u0E0gByQ5sZkP+W
HE2TKTjJoS47nmTlviJSWFWidXRSgAqQh5RUdw3oQLkwu0WrzFyutPYKIDgpHWQly9MpULtE1A/C
4wt4o40qlWaIhYpPfFJUelNa6sVj7cPkvtiFD1GyVUITJi0X1bapqPqpTPRw2B3jN3aW99eGfyUc
daGZk7sIGNqTtXSIxBp0t0rHaQwAztCMEBVpOaGV7wuDMGXsMot7qMiODd65kupnwK273GWWkNsn
O5IQXFUi3H+8vUnyYYjeClpLjMqTIHS/ftDY1+bgHEir/Qyw9lSBDHq2+mMh0bcjIbUes0ymtphk
z2Cvx4HFhSkiVJ2ST8dmR8EQ/+5asXEhFBMhpLKlo353StAgCIsuHtQHlnYnLQXSKPKbiYCnZAVR
bMoHj/1nIevZfDXCdF1DpaDc0GdgExA/VxJWJP0/SON5go/chNR/zAGPDdD4aVm7AYRrv4cgN425
tYC3WSNGCGh6GP1E9le6lXMt0hu6ivs+NdpvU6JCkUPzZl14ArVtuSpBfMtOXCUu1bcJ9kz6UIr1
k9QOY7+/MyEHV9/lOgE7ASkZochn48UjNdxQC52/4eeJkaYvojIUr2WV9KMM0YbLvmAt/na2tYK3
LyaCPrY47nwPkUN4xnAGFbmvR5uwWyru4LQqx2dv4hWQvIzNFS1xyJTDzDBAiAAu+n+cyChOhOfA
r1rdXfaUOB2f3UPTRVmMypD0w16qBBJwcUHLTaVYF7a3DC/cLxHNkqyDyD3m3F8/DVwU1sz50tj9
khFOJdKVNOlaKN2ZbMWMGW0v7qjjaOxxrL1jJVcElO8h1T8I+cCapsy0WgJKwesYaz5mY1fdzINj
esDGTXwAJ4kAqOrE/30TPaY3otun/g6t/xtt1nOiCqv9iryMq4HZwS5tD9C6p1myUfHXD/P0F2Vc
eyFgaAeH7cbYUWPux9pOJcB47ipZH+znqbo2ekT8F8vEXXTaLB7eC9hZvNE3OWqLY6ZrySKvj0Oh
mK/UOlYmCxQkONtmnFQoPyDCS9TDQBqFPZx9p87nHVgqOUT3OTISGlhTqAUv7sfmehnBq+67qO5m
dWs5beiQKT/oSBrDD+Yx69LluvjhnGfif8sMzJtsUJwpfe284PY/XBZBXFRztwFQTkt2fPET7JVL
IEbWRjRDfj2fYwq2Jx0R5plHv9fI6xfWmMonndeINRRI90pZkh4Y4ex1ZAW6S4pXOVe0zwnbVG5V
rWcth/+EoPt4rP4+kJmyOPjvfJ6YND8naBqR3lJpc5oaianEx4pZMu5i+jNIdKGNMShk4Ja50Hv0
gLYKz8Sd7qI7sNLTPw3CCtXvTfwL4+weK+H7o9owB9ME2L/YdsKjm2S0v/dtLpYTL11wYf7HcHNf
/YC4Axxv9cbf6flLVU3oI07yGHT0RWsBYjo1Pc8s/oZWbpXZLaKMMkOlzB8tWpseqaHWQSpTrt85
e5ucLLd/DGqDAXVb+kzd+cwO/Jw9A4e7XK1JQv3wOGZG2kP0im9ADnAosseGCf4DFk8dFZO04NEi
5LZZ9ENLRlS4Bmyxbm3MOS86OnajwObGJxBoMkDPEK5/W4PlVBtIJH5MpaC8l9iupFqqskscBopt
EsHnWvRiLoa4iRmoEKcWFkvJayAPq1sFygcqvmxO50M4K+PA4fwLYMgQlDvaEL7fRbizDImXrsY/
XhTLd5ztPc9JGOTM0zys1r3GkC+24tDK3mwFKpo0K3BDxFxbZ7ftbeR+C7FVKMqZSUiE4jhxLE+l
lGIZUMVSyaso+cztFRHync4D1NJsIIwcSUmmWWtg+Lamd+/Glh1su6Btw2G9OOQ+uwo8jbleZl3E
soRfX/4ioQAgPMegmawIJMMYSdDRx17WjOQhnrcI1qQ2PSreGmb6ckKbuf9yGAf13COVRkryxKVb
pTV6NBDvbeMdP7ZZqpgOB+WTcxKqood3z3Yl9M8vKe7rngLG1cw3T8NUVCbVsQDeTfCfrUAWnKfS
+ZvxbR6gE/PPXCnRfQ1XWklXjbYy93qybQo/CvOFyrSzWJgflN4/o1Ert3TczVtbJh8ftEIiFDYM
hfjrPpgmFc2qICXh9bLAjfDcjYoyopFxomNB6qFdQdVOtFgiWAruseKV/fHi89mVl/4OzqdLn7p8
apUPspqGvBSe+3MApkinln0rszDBcDot2/hgoPVnCdaA8UhZnXZkxswnXY1BIn7YaHzObsJALErf
DkCVXlfCAQVePsH1qWIYD5YYJRvAiu6AON1W7W7OpSiGSbV49uuv75c05LsENpP3Eq3ZPbFMWCst
H7TFoQXshceNJm0LtRqFWx3xjVKo+K0Qywm/22RBi1iFU9SiUZjfok1CLjPsBiROWfisPcrFFuzM
lSZUuG8vuwEpbZVDf5gaiYBh4SDO/zJNzqXcTMCkp37F44INrxIoQnG7bCfaQjTRKdXzV/QwdTTL
p+v/+4sQFpBn9VDH0PTKDwEqXCnv41OSMOW1kD60vfEkDltACa5ixMb7tKT2Qa1xMY89oEws0SPG
7eI76rZcqu0pkRw01/bz/9xSX74I5wXGQKzXUBSZmEi5VWjhAJrcjwjQHEBlT+JGxBCXVn4lMUQ+
IlSov/J6I2NN0Mv0AX/iXBcd25b+8ZvGZOSZEuVsxU7tKGMqsWY3cQTw+/s3b8WOkldOWqhGECee
iah9Wliyo/WQ1vCB6Iq+GFpetKsvB7sS/eTo2zcAaEFptGdttS+D9YFm0KkRnwTAycgvQrbxqKVb
Zl0d5i+Co5UVNUeK7TyVP6I0+pmQCfdPm+KzIN6YZLHAqcB6FHKWyS2sZXjAQ5iIvLRSd1picRve
Q5xyUGt9dqDCgdYQD8F//7wQxG2m/MQmyEtrlVOeCnbj/ZXp2RdQee3rZhxfsw2V1+tDRJudYP/R
O33QRkkDz8tt68mRJ+QCNGIKEQx9CJrwQUg2ebqtd19d3eaoGf2yoUfm7LtxFHAcS5P4F4ceAM+F
BVSLGX7oNJPnaCfHm5mQvmyZi4PPei5yEqZ9bDPp8myNt0qeGhOqSpawLG0nz4UmHRRsxq5QVSRx
fwg/6QDJifIjPBLigLZccNUnX1QBNEEkbytGEhU30lphHQZjAYGFrhE2flrQDR3GiibS4Mm+uZIM
2DMrJG2TkBPt/F+CVl+ySOVNMaDixh0qiE7pkUQRPwNE3HnlEjRM5GWzVTIB7AQG+aJdcrGXnQ6g
zuXdxyOJFPZkuu46eXDXOlTGskV7g8tVqPKYUMjVbza2oHBMm/bQncIyMb24KcPJg8D+EErqbDCv
e6kY13YSsg2iI3WQzNwnraMOrYXmpqqxgTZZyM3aOz+ti75Oph9ltqZaZ0TXNqwIByqw9LMdz45w
uod6RKJcy1PB2q6qYgamYzLxz9Zs+GcesTvBvXbTathiSicjnK/BPkB8UOqkrBRN0NDAfdyd7Sy6
Z+OxVjW63q75rzrLfYhptSvx8ZSvY+AjKx6+6Vf2WhoBpd8hGGeptrzftg0lUU6IME7nFejPSOQc
MOHuJ5yNvLkwBfz+t2ppKTpzUeYKvbegfQaza1sp2+MhWnSAzD4hG5pLWVVHGxS7c7oos/YLXqaP
g/inXceMGQlGr8Rgd6FVnpNtysNylBOBtsX6Xj0RZrfst4+xnh7dSF2R5T5Ri5hsi2mtOj035YAW
0GgazC06RhKfBOPpLvw3HgTo9quBU6NLtAC7Er75uws8IhwMEzo14UPB2ExUtK4J3VHg8/Mq1WfI
+TF+dXm0HgAvGYOcj6uKj2wNcRiJsn8at9n2p+i/RctXfgJruZeL9ylpFekT/aQ4++TsJKlbt9Hg
Rpx3ng9oXCIVJPP104hTEXAACs0Q/BMHsccH56VafAW61rgX3PCMyU3Pd1FpSSw00yrv8CTLAzza
BiM9Ek2w+8CEntmxHXKrFhhHrv0DtIbZyRtdm0JrHO2lsw03aFzjHT4v0WbRH6jlELrVQNiDHvDF
ylcyuKuQDKtaDFa2BuotUlkNWaIOzKCilbIdFgNYFdJ5VG1XjJwVbK0cBmnfJBwkP+FkkeSIRcVL
wkS1xnTbRrGteZHAYf7oOh0pAqg6qf0z4268vxYc8RrXK2hvqwOYk6rp2qPpiBdyvbXH3a3Zk4Yb
6OZpR7B2g2RymsFLRPVKkrPIWVdmaGk2+axqTa4NmP9oqRq5pbDlG/twCEtv6ysZFXXQZ7cc8r+c
OIM/rAst/Barl5dVH7ba4bcVWM5NLn0qCUai798kszOWAo5uFQdFXRrYJXXUI7gRS6oWctMYgzVi
44aSy6JVI+BJ3nwfpHVgAr5bgsTVqvosFpJL1ZSNKOc2CWOzGvnD4tlpUfouEAQ0yVb+hchLSpIk
CM7RPotXqYVuCyaYzdp5QPVpwDxbNKg+5RvEHSS9H0aSyUZ/tSoTK6POcP23IQjiByNrGG2mis8O
eyL9/jWS/V0Dnqz2Y4IjBbxDvMMnuHPfs40lSpXRfp5dVWt6jr7PMF4u/gDZRSOdCWw0YgDDylhR
ObHkNJ7Rbzl5cDFfk6poh1xDY3vTJCEn+2DBt76C5s75Pbw2RNhirOlPZnD9f/WqPQdZAiLkBfb1
zSJ0D9PSVAGWtZumiq/FYBfo4VNAidNzVaiSrh458i/ao/Y3gK/TpavOBP8UBi0nB54bGoDrm97w
vQROrzAGeHXP1nEXfGD3LgRzZtYTAJZrTD2skYI79FpRaej0UYZ0RcqZ+/JkIB+Dir0xBW1Jm731
HkyYv8um9nULeG7ydY/EeEsAHK2Qwvp6Xa3TW/scuI6UnOVxMXn57haAtpMJ13pprJXcJ/qRcP4V
lRcTdaV6tgk/gaRL3iXF/hDMyEt8uvJwnrHptiz0lFn9IVJoH9q7OJ8b3G2xVrXYpzURW8dgpWrB
nB3JYSad1ks1/nayHPFMyKl9BZy7STtXPkcLoG7KCn+Se2q9FBckPfl7zb6Wt7d4umajCbT0KHAq
k//nezknnAPhVyBPnWfpkIKcbpcV6LmhUfAT18J20iogaRvzXtER4ywW4zdapZEfq6FrkQ1KrSvR
bi+MlB/nwQsr1xx+E4bWTFHO2bMPhNRHSTf+bj9f1XHWU5IV0du88OluN4Bs0noTx4phP5lVUgin
5j6ubGQCkRReqx3lDpUBj4Hc3JuFxoFA1FWmQSXDiRN288UzUZ4eQkyOVGIgXtzrUa1wfQQNZWQL
sxpRUnIOpG76bQlpiy95Ljpi0V5PxxTPByJWCUKkciWGEfpXTFhxDcq2J3/4F+aGKFj7i9kmkjny
jXZEBv5w7b1WWI56H2SvzjijOGoaBFg4Xf5RZzuljA5Uj1+av1Uxf6yINp+zz3r2sK9l7Ivwgvtd
CCRC1okQBZS1OESjECP1Qxdf8a0vVV0LCaFgKn2Anz0/3wLu1r3/OW9zi6V+d01zsZ3UpoA+V4ZN
AEwewROBuxoekF41gQNmUL/US5ZegoRoPv+pixBPgUopmd9JL92ryn/y6o2TDxRz9wSBmN1Jsvkh
2uj0DgfaWjQIff91hPc9CfI4wt0m2O2IwmONyNb5UKU3gbq9h/EFbVHFTv6JSocTnSDN3Khcpb9b
5GCKt/gIh14cOIfk50cnONBnFBxG6lCp3cOrL9WI/vlC2kVlYdYBU369YIgWvbF/JbyNAS4EDcg/
2UIC8fgXNI7bpYW1knyT/SLhj+U4lQ1ZIhQe7S4UOC9mOSsnNJoA0JEqyM4yrR4QePcp0jFJb1sr
/PNfSG3/ru+xus0lxy3Bg7nbSxWSqpHkDMAVxEXqkaBj+DBQRTzMBs0zN/AMjuCPGUHfU+EW7o7g
68USkWKfXDFtyh0KOnlOwPSQXa+Jj9xa05D5J6DKZZNwISapn+3ea3NVBJlzrQUfS6DIAF4BH2Dv
znQuTgkr0K9rBTHted8G68Xnm4SFgmZ8gSyH2Znsz2UzYumQIN5g5wsyZUgF0nIwlLOf712eGn9q
UQ7pLcCVktX10EmZFe9C8GZZwc3eNJCovdRZmG1M9OGGG+aD9Fxzvjs0HsecG3Z8H+Keos5ub+zN
Eo1MpXFfEGJ+QiIm/sWz8ReIEdkKzhCfsBtuKP2EKFySQEfzzWhsESxVw5tjf4SRDF/46EFjLZQs
YMRZ/qAh67113sMVuM55rbdYlHyB42KBLsWl/xGE/yltSiL3qDv+I07DPIht0dLzN07d3VKTxulL
6P8dkAdl+UAUves06gpVTvBiVt5oPKBr37vVWQikAATh7zi7MvEPB5m/Bt6ZQh2VNL2Wu6eowyXb
epbo0MyIxdXisN+hAnR4OSNrQAHTU61aZldn+7F2PJuxazwcByNtaNOAKYp0+z9WBSuftdnuK/5T
xZBEJ6IcwGyITzTlxVnfBmGvMFIkfQJbJLfJm07tmRUeUJ+85zhsUyR/3U1aNRnJdZOnuX73Ng5j
w485rnHsC9CZ5PpDzkmjOvp11n+1DSJJM2L9dFY41vcOKW7chOLBnnfnu5ZaWz3/f7zx2fUhMtXL
ELB2NhbU5k+5rwwPq3cY6M93mF6LuHoJZ9RSnfX1rGGaSV5NjiyM5nvM+sQqVuKmUwIUJFcSLn1p
2lNAgx0S0KEC/hlyPQqn5pMspqa8q8KNZgqc84qS97kI8yozLJojupaPJRT1kcuNjFxJ+gxOHW2x
45l5yI6rV4gRs82mgyv9wZihKcyGnBk+9CHOXZVheAAUivyUIz4LPNJVtIRgffZDDnBc5HJZx1Nu
dxpB/B8NFH8Kd6qy/0/1pOuG6H/wvFtPw1z/kSIqCMAqND5u52xjLk1nj10vPSdKJV7dM85pkagB
+H650FPFlenmzWMVpKxkZRvoK3UlHKjIwd1nC05lkeH11QKSEfaxP63IvgBsgduPNMHZlhR+Kyhx
6hiiuW6MK2/v1uhDyYCS7216E3lHmn5qfCfZb79eqhfNgSvMS3cTnH1OgdhLpiMIvTGPqi+7owDL
k5f5Cg8ou2+F36+NwNKg/YTzNMWk5YeNQa9gq2GaY3Aa8Gh357VMSS2JzviXeyttEq92nd5TlhXp
IXWcGB7SzcQbNrKTajim9A7AZ8z2N4fEczhA6Ir+/17sIu763KVGutUfi93OBJWdsB7Uy2CbW/Dl
vmC3c00W3Xg6e6RcZ/MA0ynK4otgAod5qeeDbFoOYpg9B/wJkk3+CNLrkVZ/lx0Flq/fvmkyvsxy
7lPRIRrAK6QrMRUEyyhVycTfuqOm0si66QEx3NQZktTOgzJh03ezHJ4o/+B3lxmh3QgITRfCPuVL
8oo9IhDoOb0XXF/j0xMw3OJX5npiYlfCvxTW8T1ugXUSVXjMlKINOHrTyVl+2832FjPEbFie3ZaY
FQ14Vl5jCK1SK2a3K+L/14hcsJeZ7ifQNMJGcBITsapm8qsVDomlfY4SwPxzjb00FY3qWaGPVhop
znd4shVzJ9z0nvn2BZYmpGbZAwFc2pFripGnjo3JYK3bh7bbfO2U+M/FeepFSIMgmE/HOAtqtKOY
ea9IpRlsOS36yjP6wOCRaDXV9mYcQsuYHQmJvQ+sEGGs1Frk/uDCPkAckfOp7gzoxROX7+G3j5z6
5jtpCik2BYk1uhd+Xyb/wLb7guUDYPl8QWwWEq5xRBI7gTqb/6MlTSWxK/VO9+0OICT5urW1sd4X
s/BGvNM1xHq8ZUIzi7SvHQWfNV2A0mxhL6HArFl13Ch8eP5fGRl/TCASo6OGb3CrAPxvwsemi8Np
vzuuu4QGFpRRB8+wr/dCpC79mO4G3nG639YJrKOhOUqiAT8ZlUN/U15ig47l1fE5KpZCo60QtjvW
O+6UEJYwI+Itkauxms3Gjm23EAKxNhvh3xOhRf/Fb0zDSHiMLBXW25zQ9IZgGviZtOY59oUevPj8
E8iNilKvAVnlhZBMNgPzUmKY8vXSLaDa8WxiqbIPTehEfefoaG2eBqXkOwi95BGZ8TrRq4x1phOc
QH/ok3aMYJd276XnfMzZGD+3wjjAEYBFkUH4+uNyNgAFQdwPxB2RB4ZWqAQY0i6NYVZpqlUi0Woj
QLs3y0362cQ8jOhn8XvVygp8Hts1NgyqggqWDL0F3r5Qjq+MMa5K0LNwtNP3zYCHiiTTsYFTEMBJ
Qv4Zaz2eqwrQ32W5R3cOgOkqIKaKmpGquFlg91AFabMGPKMciQ8Re1Zys8YLJ97529JkqRBCNg6b
sFHiR4FApsq+H8Zhk/TMSkTMjEOMd8KIFP3z6pv2yQ7GZIMR9oVxxEoYb5lMuK8JLWpBdEDEXeyY
fJrzg6Hhkrzk8U7xuaFMcpCpj1rV4HyCswoFixCrbfwLeYisoUD5hkwZyeUocaJHdO1CvXdobVKC
ZKm/kXkbJQ8k+08Laeh2iVMHJEsT685Us4LcqfvUig2rt7swWI10eEv4LueJE+x12ipTUq+asZj6
VhHh0hsoJjrc4aHXMvstCkCwKlGWdKWXqd1tkxObhV9FiV4IqOS9TgqOsuCs1HvHYk3WWUvU25xt
2BvxhsNLIfBUxKIB0IfZUOaschH1Af9hQgWxyGfGI+6HZLaErz2iVCNdCsP8KdXdTreOkpXeGtGG
SGe3l9sch2A0ZXCADF2yuLfKUsPSyb4mouT8wORgK9g7+TzIrKsAuIms/nnimK4yA+5RUKV2IZuC
vfkZ934mpfuvVLqDmFxjIypYjj4o7uDfT8TcoOQ8mM/ad2ZGO40bSGAifSa2Ib5kROYTyFw+fls9
llJ3RqKPuOx0BkZWDUYpvH5NQmhvifT+qSMJmj+bq0ssRhGGRLBG9NUCpOM1Q9fcrwspMzbX40lC
e7sBIUUD3oeQDkAjdOJxDdT7y55QX3YdxMxXSvkwW3H+4jTvKxrJUyzuRfvIE3230QubOUKpgrO/
dIHuO85iHf/XljprHKbNM5ciUgtitSQ4Z6ompnzMlKtAyrjGqLsliJuHBoS4ijAUHNNAn3UNPe7D
axAeFes9FFMY7XeE0JmV6QoB45qRr6HO5YMKvBtb4RWxa5OwAHlIcl585pyJ9Xyw88hPJZbcZrVv
UhX+8yBilvicT5abd5b9y4XhTn3p5jWOhTvLKg9F1UmCgdfxPDre6mMBwqj1rqGmh3i192GaQ8zl
2JWTixCd8fHpPiENsf0zHYK3hw5SqjWTcdqWUxhv0GtBPFKxzSFOuCm+ec225jNG/k/+GJoLuaUB
lfZzUs73KsK+R+YIkxV7185YhvviT8oAiiGTK5O5xYNfJxaEEwPBQPqsjARagAPNb3mYVHQbNK4G
6heDYqmj/F1amsG9/Mfvqr5sFVy/+d59MZENR8x1YhmWCtlD6wIZvqlufHJyhWDKAGaO4wVzKeHa
9ZbnKtgfYsQiMzsVC1cdbCLW+MVcEzNFBI7U7JkRf8ptLN+DFiQpKNCxRVazqsbXJfZapwnL4m1g
oX6Hc0fgE5ojBFzUmYoO9ofcDdn0oGkW3WPIwmpvKaWymdEjcNIl2UYEuRzri8ZhkFTFYnj9VMpN
VbAk/E0uEnUt1/WozadI8YMtjSKgwI0Xqlxaf95UsGEkRHKt2/z67Sf4I4eWngJMdpyu159Nph0w
lLnI7t9KAIpWatvo3ILrNZ7d9/pJcRIxtCQGtkKH+IYzZBNAipdCHdQK196bOsItIVsZh+qQmKHk
dYV7OejjifReCbavqVq7axLteRE9IQ8LTmxVyD0Zjnr44OHTt666EbOrONb8s6tP01bRUtPib3ew
ccCByL5nMYluW43V9KSQ5xD5SJ4IKUwVnEW9GHLpMOBOJrmWkVYsskFWkRhIBl4PK33BEPuES53F
rn/porc1zncMdNptgqlEBtL+HQtmK8phkcbwVu7zRi8kmBL7Nb5bfzODxQsbmnRIaBSp3hPseIwP
2h06dcwPWTnQH87v3yet/EizU9ifUujNR3ZZQmRycBrDMRxp4IwLqu5R4LeK0Qb79gwA1WLvg58z
F+UpcGzuXiXHJgOB1ghyLznRVpD7yvCwocuWjpTOS9yYm6MPbiSPoSgFg4dH7bK2/sH6iC8nQ0Fc
F/lhB0thrv+irAIMxli4eKZ//vZwJ1yxpcSpycHiSTONFvmsAt1lWVqCeLYv/dSAJOR1r90CEgV0
kTqlFlRH9JPjevm6kEDfxSrE/suBeIqA/KWqTVN+qmJJ2VTNj2eF/Kd4LkeQB8XrruK25KVd3Ut8
M/7QOcovmfTtFvvthgOj8Q20pcukl25U7Wt5+XrOHH153PxPwnF6f/6SvSX2EbesPg8G2/VEaoTR
KfK7LEgv7vOlP3FYrTN3gEqUR2GfjnAo9Hp08iqp3inXFgKu4fv7Ac5c+tOEifZ+AmOM6Fd3FRUF
1QTu+CCFNaZKAyxS95BWwXq39zYMwUloVK31m7bNj84aaS1FmAr/1SkewVjxN0BQ1z9Z7fumW6Wj
FXY06jBofTpYZB6rVzk+M7YMHvfyTPVxloP8sEEsaX2138douA8u6tijVMCSu0+DHFK2ieHEEfrk
RLTMtX/cIck9jBZhqr/gQwCmRU8xd0ecZKchQycD5n9XwxH9EI8vhBelZQvC+ADaoB8VR/TLDLD6
grAmn+anQ5CgK2k8EuNUTsyfhsc5wnRMPslY73WZJb7kBfm/awjS/wNhTFbKdZeUNrRi2Gr7g31u
n2dYtr5Dq/a74JofixZmhlVKbqpT5ometyjLIoLE/TNnZiBuv4JojA/A/OiotXQECcVPo7ETk07H
OgZ6D1mdyrwuk8sc1hPZPRtPcfr63aDMVNpXC55Tn2C6kBE21tz1M+LkoUzKDL9/tDkgBs/ccItc
N+lk88MFram3sRb7CRbQYPXIqZLGop97IsutMwqxO2jhoSpDCbZSwSQQIsGMH+DiPAyGDPuo7NX8
o0wWg+q8XIpwY+JkOijDA7MlS1jwV7fe1YUx9nIqVc68OKRtDN+ZddoyQ2wwW79tOnEZeB1CeUBV
rpqRxEll/ggci+9xVr4Rh8PCiEJaxHbEhlFR8NILB99Q4MOJaHy6nZ3GQKWSd/OVHw35Ma2JK1Mh
dcticEem/s/R2ViF8R/T+qxm4S6GWtq+5tpVGeT1tiK+yQGSLE/kNtnyl0sisxJFlZEuvDhd9ZdV
7R0zKNcqgT4/yxw8OWAc/ZSia/XmZ2SoZb5evpf52e8yZieDOEYHeSXI1+2F+EodLipPXzyiO6/1
HepdibkNftz4r9b8sbA7Z+AKi6kc1yBBN6DUElqgBmk837LDfVE5DXOjzAtyG7NO7VLmmRXM18ze
KE+TYndPfxXjjc/zwdL5gmmPi6diJDpRrwHHJq+YtKGPpFQWOIUKUhKjLVuEb4mXl1brWp4hzXdG
/Cp+0XHdQ65jXt1Lf4UJ6mBvFhqfcsgZpBz46RgJsQXzVvtjN+zMA7o7rzGMISzaaMF/XmXjY2c8
gyMqv+ShO2xBEtbuN+cZYrDgAkgFEw6NI+TuyVEgt7+hSTuOBdn2TDUB71Ssl37OWwomoRSZtYAU
Ev+0lPgqw9Ye3P9uTcUugbAtUdOzGJP/D4WNx79HFr/QC6U8Nobp+iCD+60xSFZnnWfp5oF2QQhD
zOUR1OlRjzt49YBerxs18WKKPZmhaniH8dAz6JofSCMylfA2fJTyzNvjlZeJ+dFs9ruH7RDD7+QE
551FYoHRr9p1CgyWheB10PfYE3iSAdK0H03xuUAXc47UmyEiraq78TL+uT79b5Vqevtcj6mscdIN
lon82/1Qh4bzhKi6LgU/tMBkOm9zMzRHnweOdZrSqBYuHbXB4yTS6ZSFnO874+MMa0WdaG5pJDN2
mXZ16Fa/mCsXLnGdFWsi6rCPz5FX4qM8xcQRdGgLwLtT7medb/zIFxj0KIfB/eHIQGQFsnPreHS4
UYUitMMEhHxnLM+0xn/Q6dHaljYiNgrbTN7Y8YR0wPTGrhsBZBKwYLiVecv1hvJTBccNSBWShIki
Y234XQURUrK0102i/krb04RQul1huMbIjvwysorAbrmXhjRW3I4EYYSN1EEIjQSz4bXR1lH6GTDp
JNjLtUQMCus1QOHr5iyK6sQDRA+7FtVFQ+EqcxGQ60Y1tBsizSFWGWywpFp+pIilRp/DhUcFede8
/Z2eBhs7nIcNhqnj3LZyTusXgDNyRfD0ErW+c1Enxpx1qL6grAbUQUZCVf6ZjQkS5nkb/qxLTXTx
xwEF2Wouj8Q8sf/99jkEEF+JoWrk62D7icaubBV6VfB2J4z1Bnhytjdga9xjjJyCQjx0GaH7ghHj
RcY/CzD4Op6XE43ncVd/7P89+8TfB6STrUE9RW0epbDnck8sKUsuNoGIIylXfydMk8CwnEKgCmJO
eOQI4NcMJdgei3Xy+2sm+1DeWzMHj1jdNgIH0EuyYVh+gefcwWyrVfYBhq07bkPQEnmQH/QUnyfx
pIJkX49lB+r6WidlifsJ2qa7uldmXGa8N/9LesP0rYAdo4sF9jJwmfXkRY683p9/oPRP/3DMjxNk
7w3fKobrFzs7mkPansSg+pxN8rVfqHzKZ19mny8CdSZaqlFtDNKWaQZ6kgu0bpPASxzhIGu09Sia
coZOSyHPZIpTYOwfYj4IFkcJjGrv77pJpxqiJyfJ7Myj+NU//a9EtPZRUvdJqTZ8BELVztcEXtwW
+EvHLLCcvfsP3YiT6USG81pF2PG9tzqeFCEnO2HoIDaXNrFXFjeDJ7yaUGoMcTx7xRr7HpIM+/CR
HkEzZ5gShKY8nvD6ib3KBG/MvckApTn7FE0bWPqkfwb3Pj6M055GUjsq2Fy8rbXN3E10NuD2Zep2
6vFVx/6uWPmWGEppRV6vBewujAeyLHboxlo8GkrGYvz39JQtYok8qrUtmCbpiPJZ3XPZRggQuHBz
CWx4leo5Wo0jmKgl48ABH8SCSl/6bOP4WsSzimEZ/n91hv1ZxJSdvqwWiaIwmsnGWRhWr2mclar5
1rGHRl+bwAC3RRBAKE9PJ0Orj7Mdm3ZUFvS61CLNJ4ftp4db8GXy/ztMrS9XqXw+K+Xxo7n9PBo5
YuLuFtrFM8Orqyp80SmX0fiCZbVX9oo9l3xO44n00trZST/+RyYzZWrfiQ5M8E8sjuMi37RRDWv8
fXw7JHVoTib2cjBGn027r2kqLxUsJc0bN5ssMy5EywHMkCxU2qRZyq5x7TT5xd81MYGqf2viFsa1
I70s3slp3Y7NHuG5eXg3ciK58paVZZj3PhJkjMkTw9RlNyinSFS3emPbYdtPw/CbsbgO+uHvWT5q
HrwBA+/YnlUF0/Oh/NM8fXS23R8DSj4Eqo/0H/77ai5EykqEqOzmCO5xS7w/B5Z+PGuqtAZz05a8
JDc7QrnFp1JZi+kPhFF2rKooHRntSGCne5KbhNFLr/ypWhmABxEQk3n1Y8bjoz0gdOR9Sg/l/Dms
JM3dff1X1wL2oRvCtPjxwmWT9TePVbOhMgy3jBkn57qQZU76ofAZUGqpPjWI9NS6dcvj6LaRbVUv
RTlSVIzPqjwryD+Q4ZRF+53y9rO77rJ7tXqQfxUKBjwvzAc6riIl9pRJePSj658D7HOgeLtxFri6
frYqrAWd3NK0zqe6VaAvdUXXeNJltXenVwLDkJ4hXOFjqi1+EN193p55zotldKeNLEvweNFyjTEO
wCPpwfJnakd0TIoFM6LhsoKV9cf5v/QuiUj9yGUw0AU4zVnrWqD0mrW8/OMnLKWDqv+0Ml4+hEx/
h63JwiICMir3Bn+TEC0ptiIkn+lF7X7Z0HcKWr4btosRrD3KItYZG/9lXyux+FeT1j/8rzYOxnwj
kFzU0C9XptcWPqBuaQnSY6e6Z6A1Va8SlulqQ+9zZgyNO4qzRRl/2aZbxUMMSqgSIv+e9OBmFX7b
K3NaEJlc4DPj83comhrxk+WgTJBSnp+ewpTLY1yRQvu9lkPA3G7sSg+4p9Gxck6SlAVWSjA1SBcp
BKVlJ2wgJo2LHOJl82gfuawQaIHGa4jCuu9f9GKTZskkGp78qnx67nJnQefDugAgtGGTctg1quFo
J9XE+jQCMX7ZaLhw+TNKYhQc565LlCuixSyM2wlaOpet0ncdsYrM1OnqEWxZzFh+GMxFk0ZWzBZO
NgEiLxklt8wKlX5rpt+c/SbEQW+y7AxGjpKxhKgz25exgjTzbxMWGnjMiFJdGfzthjYnt710hAtm
dbkzaubx8KETSWRzCD2lFDsvwBhGNU0ZJgOiVaMxHcQx899i7hbgW+eRTOixp8GodcxHzO0p6h1Z
pWHZN2Yk9PIcQre+pFijZGwg5bgeH4lQniJ9p8Drh4YJQvBHIsLa0/j2wTu84vy5wTrgcrz9EdAT
XOn/12bcxck+5yPDkFa2oGxY93N/ssMexUdAGZNv/M+P+OKQCXp2r4zd1R/x6NpEclmtLnjLmtKU
sj8QICLmfPCSU4EUO2uOy0/CrKnh8Fs1oXRD/FUOYq8bH7UsuEGFBxTA1XLdntPp/Wz1F7Ergo6z
jyfZi183tC4Futg4IyQynbi8yjlfCmEmXaJu2RzSFxe+AsYLLVtqL8oq/qA46wv+qhW+2pS8yAjo
+ImD6abzp55qqiXlw9wTWz/u9ODbFQP3fpZXBE1T2PCnemXjuBg2nVBf9zKPQPzf9mh66iYnSvQ7
H9hUe/n5EqJceKd8r3WXTI7hgwDNnvY1WOHhk287GZqi4HGXeqNuyJNDwQp6md/T2rETO+Yf8o2r
Aaj935l8VK4oMCmaluhRU/EuFDUx7/MXdsZL4xqePpy2HNBlYAE2kwDcXDmnAQvEIV5F1w9WSJZi
6HIIr84L2sQPI/jKY/ykONnlGBmKIeRsXE/r1JxHAuS3L974K+x0VHbyivMW2+7B12ADTSCA0U1Y
U6bDTOVUdRWQ8THgrarUBYeXP+WlBf6TE4TCKb4r5s+RkJeYxJ8zq6tVNlOmgAs/UUObdQqNHkMT
UHbFHSXjYTir1rkSU7Ksv0EeFSRjg6ZxYRv9v0ZEPEy0tYm4dY9KW8PiN+Zwa4q+Tukvu6TP2G7/
k6p2BzKNNeSQjpc9QjjjAKdKODSugW4Bp9U70iPhC7RUpygRQSPf36Va+rF9PwiMCAt2uH7Lo5B2
8zmvS/LnQvf5aOpmZBzDClYYWWdOuo2iEhpqA0RPqqPZYAd1+8Mbidy3MS+kXPOJcML34QZUfl+m
+gRY0VmCfOC2kZaJug9XQjj3TNqYTB6nsu37K0BomfcEH53/zqe2wd1x6qst3ukv/OvbHlK/s3FF
uMoOhUzBw5A9ar7vSMe5ncrJeDsiFufoRYH4g8wJ+lNavD/esQN6fCqmY3oJK2o5TpxEkpt+QZcb
2AItRw0SdWC+YB0GsLqd80WLnQYHXR0BCatoCVrpn8f/unQI88FpmJnRvJ20m0E2Vdwk/7e+Xkdp
o5GxIkK/fdAcBq7yn+Fv/lszUig4JmIWpriLRkA8C8la1IeeLYSO2A3SlkwQz++hu6l/30r36izU
QfLdGbG2bXRT8vKMy5k04/s71YH8dX5ElUeqI/W/p49PJxWTjDP85xR6A4s3vL/dx4++LBgiXtaI
dIpd0+V/xaOA3n4lrKk/U9oARPBE/V70fQIb8PLCu2+4aLSMVIiMqqJ/0OyGk4JZk27WKe5M2Ukh
X5VdBbg1+OhGmn64clhPnvEGZUXal7HkrIXrgKkWo5qpeDBOutd6Pm3TJt3xuJ69CD6sojHNmh/S
PNsoiPMuHy2sQEELw/4g5LyU46BuR+xicN+1fTL4q8tZyNYY+xWRx68S54/0EuMgn8RX1zAvWhnW
6twDrd0IGkM29o2XKRkxOXCo0A5jwQ3YHjnzbXz1/wY9vQgRUMz3o2u6fT+/p8XBL+f+qIDc0Aw0
6qoo2lxledYpafSG2jswLIVxt06FNeFjdx12uc++xqKMhQKTVxoUc4NmwSN6kIybsLOcXtpC+2zK
Sh212elMCmeFrhxIYb4rFfYwNIX9WlikqdR2AlEtzSHXj6NI5z4TBLzu9hpQ7qatzQAjW9fXsUWp
+nzMaxTB9bPvtRxDK8SYaVAVA0Baq5OytS6OVabgLVvuf0OuuU632sOlh62Ca4ZU1kFPAud+xgrR
XHsqWzYP8ggbkqmYuJtqOioyYcI4qBb8LLDy0VVo35hSPqqRcGb/kagHGuIBL77q0S9s9lgbQ8xJ
6kGH7ef8aOqMN20otdi5rmviUwVGnw4pri1zXr8zFIR9F15h8nq9cJuEXO6IzNYARhfDK/PIXrMJ
YaqRnhkO989G/UUkI6gTcoRSY3NqTytGvPJy7My6Q7vH+TX7cP2n3jB9VnE+pk7EvAG1pyumv8of
ssEDe2btdVPyXvDA2GHBEyex0Uw73XGcpWqf/WjDEs7ExVR1/yPjvl3lU2bRUyvMr8gmxO3qqzBw
BUzF7TiGoPPmme+5e5sGTpLLcUvy7WZ7fHF58rd38h95c3Sx5/1NFG6/sHfdh/49TGDMrSC4UQXm
W6aKrdEMb/US/H/uScVyV50tqsqW21ufO129UARn8tKGXXaOk/jajZK2QtGcEWSGw2a7RuLPb/tZ
AKNjCuy07Xjhoi8ftubrujWSoPqavBBGRyD8X3U8lPJAS7RtxkG6W57ODh5uz+aVEMe45n9qH+HJ
qkrMg1LyrqHL7boWk53eZPsEHWY/Q8qOq80r2KgEDnPQaDzbsVTudNiix+k1hOJLb9uMrLNNLyFQ
Q6V3ntnMXdnLev7QnfJunK8XAo47yvLjARooWYdJ15cjSiFR0H2fFEhgk2uIYkPcLsTDe29zvaxq
2w4bJ7j8+QnBIDa/D0yY2V6kqz6ToscsVzDw6YhKwET8C56lAGIoP45O9L0RQoaPTBjj1FWwaCCe
RDwb8NQU7vfnBZtczDpatmNHnRlgQAB/7GAJciURy3crlc5cIRaKCazKW5AcMulYEQIG2S1bDvNS
8PDO9Ld7njqBwwg2CP5ctl3YhpNvvL9Lu64xHQk14jhqI1CYTFo9WqOolwG01ABRYi13e8scQ5qM
4Xw0SHMg4MWshRw8Vvp3YKFRGtkuYoSEzu0tvYAaqBltLX/gaAQJHo0xBglN71K9ZCKxuAiAW7Ji
t2EL3CwTHWRHRT/9MWbpre3N8wopP5xGBQlxmem1K8oxc59yLsdmuamlM0YxXBHQNbj/hgp6hGx9
8AdGhRQiiSIKvYFuEaS0hSnOVezR1yABIuQqJwS1IpHccn5bzSMtno40PfVUE/MbfyDGt9BYbPyv
XiK0OPqXxrvnl3x2CR+N7jgettHxpplQQ19sPtwULjZE2Uzazc/kb4NFgiDtRAgOL4V0DAOR//fw
8ZCoPBTxc1I97zszCXlTWMOsnurHtJT9948YkE3I1/+J2dJMjDvUc4xu3NNNQvQ882bl43xSmqBH
PKUozLkgvYtvShWm+fu0k8mN7uO5KPlYoPuf5Uu7UGubUE5UjOd0+WMZElc61og6PIc2ezjdbcg8
woQpOwVGNm3IF/IMXJpVjkET9xoqpQYi0UBwcczHfkKRddlZz26bymaNqlwL1k9Q14ktCNJCm74h
Ra/4ivp8gdDSgpZMgg46yHt5a69o2OyQl6MImoOndNUz0+Q6M/Ldwdl7YogWW4AcWVtgXUZNk6Pj
qOTHN7bJM5Lb0GebS0rgW+N7qHHzY546X5sgw6jOLquY61mG00kxydsx47fJahXgsBR37uUjZ0WO
vi1nlzrPbVhcCnehN6MKt0D0W5k90YMCWzpBD93fbxRyhep2YzbrdFxdpyONxi0s9ugB1ywB+6in
bEM27Gz0Q2TS3EWuXijwDKHGSTgqZiasgo0LbWeUSEOnKtfWfe1Ph/7067SZP0sdOZrjWI+VnzYW
i9I49KX1xGfxelw9hsBJZBl5mih3FLRrqgucdpII6L+OhEZU43jgsc46Qxi1Aa4N1pypTu/YgMmq
I4qB2QfhSc+oj+nXAiC3MPGp65OLcC4mo2RjxJHdnwqOw2HORy9EU7PYtHG8dTgoZ+Qu2AfNoBzQ
67xbcHLQdqfyK41NsWSqcNs5PqKMBS0Z7043Hy7anguZPyFQe/Dsn/FrJwkUr5gFu7+XuTwl/8WM
HBQY43sX9qihoKpzyscnZpqJH/HYx3kYT7JHy9P5lRc1wiBsB/AA3XCdq0HY9SYWaMVaIfDTtuTY
HwCl1gBu3OC0HkXnbs/pYclr/KmrBwwaGTDf31NPWpJZEFLpWKv8S5d+qN+RxJPyTaNMTSqV6RYA
GrrEQkp75/P+UxRAlyeijsv/dolZ3AzvKCeqCS+JEDRPfsFwn6aES1PaRrSu8uAjch77NXhRKko8
ytZovKgnI3bVW/hYbPsdUiCMM8ymqDXc6Vb6HkxKNY+ycPkwL98O7t+DN+Eb5m7Q+kQUkccPqaQX
JPrMfn5003DA7uvtKcZrW4htDV11IeXf609CjJKQ4QQKsiFnZjA+Yj+S3LJWe5pZkhrvynV/Mmyq
hEnnvPeznjAQ8YtotVFNVtU9ipjgRrN9ujhJXz7qpiDdG5nyJnJzFjWeGXE0OqAZ5tJfArz8lhKk
WKWsa9MljcTw4hrkoNKcCKBrcdojRCdd9vEA7we6MmuleGFDGRYoEioaLgRvDUTe+lbWdX3mr1l8
Vlds+tFvyIWwQiOnLUNFPilsMqGEf2MDapDFTfDA9AtEwKRm+C/LsvEGtbsAtcJXpvi1I3ZVWOA7
2lbmEaE4tD7uYlH0kCKXz2ojkoHkm1DwyFhwYODAqAxDhybBEVOuRR3mEBuEKZt+/vi4fBLfhyFk
vnNdjxNPAGsytkrhplOtlpahf8tvolwuRAPt0xvZQPLH2tAwtFbUnxEEfMfCACjwSBbSfFAa1wkB
dwX8nFxD8a2/Y8iU1ErLVA8vjqu5uWu+l1gkGkCIEIeNbOpN94Wg+XVKRUIlOpyxyZqy6Jxte+SB
9RTTnA7F0dLThQjaLZ7ivKzZ64pq+60R04Nob+bvx9S2pBv3QY2I1Zkdm/tQ7Wky5E3aLuP6mzG3
M//zyjVvWF0Ubhgu9X0x/oOdMaV5817Uv7UywEr2eRte7ujrNHrVHMxmPWl0zK8ZCv1TzclJiBMh
sPrfvLmvqeHfx0xfPtOYhUmNOBVw/ThqFOSEWoOhPDNoeOAdvn5JhVkXgrHceenM4aK5C8RthE+h
epZObtm/rU6ffRELOOhJPU2ANLFTewRg3iwpBu4IB4PIDueYZmWz3/8Y9eFliTIQLIUi8SQk3Lfa
/Y8DzyurYxOrLiFeI36vPR1xKbs9gFn+f/6uPMivcDyT/ay3WAgFmF09FBqsB7nVny/Kev3/vKQv
ZP4ky+q1pja3SLLdXSb/cIhg1/ebDjyOEWsjJ1npz9mtnLalmRZLkxvTn+jCCDplMSkq+GKO6SWt
eoS68Ntxmpkzt0781PACduKkNZKim44j4WSPPWb/CvYol1hi/zrGTYH6pIHtLFF6gOBaj1yHdywG
kyIafTxd2TNdMbR3whgY5+QlhunA8UfD/2PAsXyqLc+W0qOrJzuEug7ZBDDb7oEPKxWzYOqeZHGV
pYX3Bx6GefEcTCUK9qQw1nUpO/D7Q+H4xYKgGph0u4nqQpZozkw4Yr1NZAnha0u1flADkl35ZHHk
PFrVVDw9fnOZv3Vkho2Lqak0Evnq/2qL3KjIlUP0fQKmmwLYeKH8ilnveK7+uA9l/d5zYpMBpEHf
jyYnZxwOWyNBVDanrCyG132WTp/rolGte300JOQZ91dgEW7usrCy9QqXBLnn1GaCeoW3pHd3uvzS
xSODba5BNf14DZwVjFFQvsZRh1ylrRzBnTkKU+DbSr+SzncjA2rwdPKJupoBtPUox2vnzoEHz2Sv
2vXlEJalHhu8bdaFqOU0xhWQ+WIvZl7x92Dc1DXbYMBl2Jx18i+YPQN12L0awn0EtBhIkVebwchW
9dhS+7tlP99pLW0yidbPg3rnt2gg2C58vTGsYhF1b1O5JyrpkVh15on+nTvXpM1vj5yjruhtrAbz
IYvM6Dd+NVI91w9Rr8W3NF8t+ZBPwISg/ffmHFIg9DxAo0YwbqF6iz1T+FkBDXupCS5fvWXR/Fcu
h50Q8mINEH0Q9gt+Us+rpaOBAdlVYrqNuhOxfdeZonqfMHSoIho9B3iRGf9YRiP3ktkQC4/7N6Um
M0atGgTWPqdFDhyhSf0FxdsMuVhXpRhXQ9AAk3Cte5ezkEst9VIXjdzslDByiXKV+SEGC3Cas4ga
o3muSOyj2JYOJfhNEim9C+Md5BGD87HGxz/ScQQ4cloViSHU4hsXuF2bx9eVVV0NH3wtquHj4AGZ
+ABJXI+TnZtBq1PVaM3IWLWaRfA/oIdwn7Wo2PM03B+RTJlBclBY4AKG3TiWujURcqJwB0okaU7O
L2NZq75DIKAvqHvC1dE269DyiChaJXy8qmMQ+AcVLAi8TjYrMd2QBDE+LTj4SpRDupRmhusqKBId
dXmq1ZGMCYZHOUeUgL0zQvyWzFwYH0nZ4ImGNx8Fzk7glzBEIdANiWUGGd99Fq56iWy8poGaThAG
KSYx5gLARvcxQfKRYa03DixIHGvm0LDtp7RXK2x3E4ao3ilE9wPTkLLlDhj25qOtCcP7CLujnBEz
zaCYyPREkQKTxOK/MSVH/BxZxmevMSsTmonhHCrayJ/6TEZ6MNrfdmf6vj7rRzssFyZnRUOPp1dI
sBBtOPfXBduvEBVc0+jfgCSzyWMchyIkh3LOOkewkMbp+YNamuD6ViC7K58htHpjdmcoBizwcJ5W
uo/jsgg7OITpptBXxNOapH437N1yyNWmqC60Pb3ZjQKzpWidwXd/VqtMRQ7DB5SAUljbTj+920pG
OYcWJ3Duqom3F/9bnUQeVHZ1OXY5dc+fycpIZR3hNlJ405lhOM4U2pU47e2Ioi5inuQUVn0Y18Sd
LtoR24nOTgjAU0YfMMfGvihgtpLDDoOlnF10qsJ5zzeN139k7KTUy2KDGqXPISl1RnNTkjs+CjMc
h7ayXS50J8FSyCv6ZWb7nQlE3EO9d3J15KRnS9oqcPlZDEuykS9HPGCc2pEpX/KhH0t6hRaqxEtP
wzQgQNHMgsffCLTYxhJOYeZGfWSz28I26zUEhXVlSfKPrqMLVT21iDITV6Umb+24MXryzGBgOJKj
vnTH+cLT5pIOuIBNnf08edLa+DbXxX/9FFVJPJeW2YinbRwjm7IPwg/XF/2GxuN3X5jY98KZ+02A
Nrl6mkq7FXMBYdwWJy8JV0oV78lvsIOVaUDFC91RcXO4tbALOdUueNyjr7K9OKo9iu1s35NRcKeN
hRjjwJUs9PErQk2qm6RJGNzmnH7MY/IuMpJJ6/cGqtGqqmSeVGG+k39mnuStTQmyfROkzgWArRxW
qoeivopULB2i4N8w4yK/GzP6t36q4s36NxLQs6O6+8k+uHFpS3F8FyryDL8gg9ler+9t0ZRifahV
8hd/p3cBpW/aBcSdK9/P67//yuJy1+NoAEU3nIjuZDmC3Vbsp4m902Et1zGPUpNpqPwDcHnQdYYh
tY+tXeb1LlzQov5O8CQnmoPfMESLukytkBL9Q1AB0Ojjb4AUqxR1KU2/8/T8NaNrd9VuUEBxkRkH
luc91EA3Zf93URdFbEBBzvu4HJdikg7rdPd3Itq6WXRw7f4ML0InIBOGlGSmbVF7mZY4tKR5D66Y
V7fKGdYLUXxXWaqwsAsHgMyKjQ6STt3nCxhbU7tau/FdL4McEDSSR+LJMgmv57oxZGnZK+9hMtwo
noyNNIgkF0vVRf7nf57H7be0gSRzQteigoaweXXq+C0BowXsfH06uNzm3rsFm2OIvENeBVqc2ATm
mdbkjxJUE6N4eqTEc+zGR7AzUYCP5UQYap9LKk3bX7n8MrxAHnD6eX79KyfoUwQ44L60TR4I4NKW
dql1Te38aCLfgYaNLJvVMWw+QpA8D80KTzs7jHFlU8es8bWjlgIPNWm1YVWFU1ctBlvAoT7xgnb4
Tsp7sfoHvrblux40v6vjtT+BmsHY+Ni/53vixp1MCHSl2Z1ann1UDveJXXfFBLNXkRvS4n4VD7DN
0GLxv4UWOnftr7Fgdc/FfH+JS92om1KQyRSiYjoFUDHV/eoP1fPqzQA6YUOdFvzcCQgcyqIrri+c
D77pUhWse39UfKTupa40eNFZcRM/26iqDJTGU7obPtgcRqAQwJsCzYf/01DgNA/9IJbOjWEaFylY
pv0h8LHCruH64/SFTc8uilBPoEWRwi8MH3E485bGPMeq2mJwQPKkrQIeb61JF5EmUXX18mZHPfnt
C2yTXxYxsDutpJRKWV9egHoD7U+a+P9XJQ3NaeGYffg6IhIU8B642Y5iZOxY3vNlkCFqkwA8Kluk
91lL8n+3D9u6uzQ/5YE989GYvwkAP5kJ7A9GpDiAr3rnoJWdGrGo5+kpu4Ktpw5QWy8Ej0YZJ6HL
z45WOdo5/AEruPdimasTUzcI6KvyEG1dX1w7QgvhhxeWnS+XMaTq+htVUYhQUtBpRjYZoBGAezE1
djl054SW2QxkbJ5pDD+E8Y7zK9eImXPMv3p0DliB7npcA00ynbRw2Qp1V/fb52hknIhpgtMlLUfQ
JtJQ8cvaJvvP9zcOeYlEN4IXlKni8cJX79SjarNrIJ3ZI588hv8uDRSMU7JEJTPAbGb+D1Bb5y23
yCtVQaBxSWQ02vfO2G3hVew5mT0JTP84XEPBBK3tH+gChJT+pSUjh5Y3BenqMwAAK3vG5GFEr14u
gZzViUQbZwHLB/qmjBH6A5nldDZletAcCy/r+h0LC+paknFxrt+etXGbUQi1GJm9BlIUP+K8rKMB
sxwzon4eYFSrUQBHMo3S+YlxzkzhzhZIHr19IRH6aA9QGiiXKMMksMZDACyVV3LNMryj51qnJUQf
55Iw/D13sOHc91eaL/0CpEjgXc+0ZEpmtsC3LOodhXdwbv5olfFRDJ6Ni5THMzoK+LQHN5qJ0a1t
waFKo4O9fbfE+GwECa8n1UdfbVBbEklK9uAnzB5iwOlDyH/8ML3BLsgCHi7d+PjJ6nYNlUHPzV+O
wd2zSzjhrxIKybBthYXgIz+MRN+wbiWhPomoB0EA8+UGt9Oig0xCRhLr76b4FkYqbN4fYQKqi4WT
ZFnQwTw1D0Lsm+6A45i0G9jhVaGslfMvaWJM0lCsIpncHtndCjJyFh9/SUi+kXorOO0lsnSrCw2Y
+RK50ikPY2vfeVyK2wYqRLdvn8GRyJk7lPnU4W53JhApZF9b1LyGBsKh8LCRCIj84aX4ubQqBpi9
lgpgZjvBBVwsX5kDaHxO4HqymOJCZ9M0626E/gGnhUR62otryIGsvfiTR1voaIiPLzwejczbHaNW
b80iEVInPf4OYNL0IYQm0cU2XK1rcgHLeIAm5dMLITaS4p9f6obD4Y9do5Wd3me8qsqDWn0UN8oH
jw0JVOqvi3Q7zabKxRWPEDSlDKOHEkHXBf4PlsReRwFB7000MYgf1o/bMJR2wvHryMFzi0wxjk8u
UQC5Q1yOY1YOlbppwMOJfh/+VXJ64AQwp+SOzpRiSSikDusjPKZmTJBwCt58V8bPG05lf+10IQCW
nlhoWvKDGYpuY23J8hZSqSiI4UwaFtHhdRHDdFzLg5NUURXeJweSmIPkTfKwS1vukgA3uT+3a/wQ
dCMEzN4eLZNPw63mRK8j44q//ZJ2LGIjmfHewflU4h7WqCGxMKzwGf8dhBUnOfmoDt3IrkLS4xJB
YqahyaFGVwm1I70MW4BxDRTmFwzZP5oQbnMTNW7+RGAnObvyt7OFE+K+vktFTufw5fw8LAylOEoc
cfOCF4tzTjpWuRd+etmF2vuxfh6yJpts99iGW34WhggjwCecSnMpaPnm3QpdU152JjRJNiWrZtLy
pBn8xXEKWoFWDiQjhJDP0BGGhya4Ask5CdVvvGQ/YjWUwFVyzhIIpQIvcbN2qI6NoQTS7n9/wBHr
rHNSN5lWBkCpxbl48GRMEkZJeBVEJ2RSZxZ1Z1cUCpoz8vVvtayQSwOzhggVOOt1VJXk+GUIELvg
ayx8Z4/BO9ipbpPpNbVN/T8NwacV6U9x55SqJ1Svur89mYpURxa/ordmx+Qzz4x7Mo8OHujmsoQ3
awiAiKdjZDZ06+aSrwYQuFyvio3aRZFcxYbFWDpDEkuJLTy9gj0mRZowIHQpTyjVEqk1g/3XmYsr
fE2ROYMMRHSSIBwL0GSFUqSvnPCtZydDZcFi18z/q9GwEZqI+5xzY/X17djrsoOCuGT0K6JRJvBi
63/OlmyU1/gZbBsmz7zkIzMUl1P+AzAtZp6sDRuQXbSBkewqbBB69rDcus+xJWDALA2qxL6y3Gq+
J/jUyRrhpJXO2781AdMu3NtoqTI+zAiimX2iMQK7l39szhG05qG3+3T9TOTAReZsYE2AEdAUOOU8
Dy5i/yMnoD/JDVIHNSdpLZtn030TTKpOiZ5DaavCaYrgMip3IMUlQRf4ZWj2tyxfguAk59qrq16t
fbsUZLKquDV/yGJoKusGYFQmSPz+co0yRj4dMvdUMImLAc2TgZcNd0pokM4aWz1IeFPuzwi3qK97
ozIDbivY9PB7E6mrHN7mbvdYeE86PjhRB3XZCKwKGCLUfLXAd7TP8/WnmML+nvyl4oQbWCjdau2Y
iSzpEtKJkXcmtIuTBVmTa3BBRle3wToVffwlR7Qzwr2PNP0x6lhn+QxMI7KONxtpWJyzWXrhroUA
xreyv+KNvstvzrBzvFR11Ml4W5mLL7m8vxNMc41g+TlVGhEZVvieeQwKilw2gy591ac3FKj71x5U
VYIM5+2vrATOcJGF0ibo/Ql9gTUxWISGJoT8r/WedLb0TYLL5gfFaFrGKWMuBwGdNZdY7gUFUFFA
senyG3HHdRYzPa5FXkCvaYZQdqkkQvAs4V5YIhWPzgfaXkU7aGjxAwSbqZFr0lUhWSjmYS2rcV3Q
GdUm4AMKbEXovEhMJMnNs6OeGYz7z2I7BD5BUwmZ5MPPzk16j7MahCy15kQEYj28fleaW4hfpj8m
RruoybD616/gktDRHGYCUNDKKehNQqDN9177AN7FvblZ5rLmA+NNz66VT8vPEvuvK03BO1iCb14c
1vh/+9bWia8wt5K/2thbacB88iji7Y5/pLyegp/8CW4VQ+6TH59AVb7lPKr3m8FMBsks3XnDN90d
Dh6RtGCPfyXourlSbi+bp3LdOrYO+vp1re0l6xxsTNRjz5bqR2TukxnU/PIV7fVuf/Rkq7glfJBe
PzDEFvf7S7PWjTu4U+XidcZpQmfKM6W9GsmObesTyDjuiy0a3U6mmXZGkRRlN7PAsqpvtTM4m11K
Ia8kYYxvZL2ikkFriQM7Emd3U8riZ7TrLbtcbkB/oLssv6NWHveSDPX9zrRS7fmbSJ87zLktKJXv
8tR9rl3LJGtavX92ZOH2/lYsLa8P0qyBL/MEyJoGpvveYkeDZdDOCMRMAgeN9CwLVFWB/hFqh8Fx
PGeBC/QXHad5qFF64+gqmGqomqo0nQdcpmKsh5ta4GqyRrsNz8kvRddGccxFCtWKnBDjzfXMr+w2
DPkEhX69LjmUwkh6IE+TfjFNgi3iKrJYyNb4iw3KDMFhkuUkSQnYhKq1RL3eTtWwc1s/nSKoSlTH
MGS5Q/FNYf/OdHJX7i39UHrjb4eXi15IvgD78k5inj7MWP9vIKc6hSn0loDU3nMbELmUq7Tgp7sK
XTkV+qYhwLJJ67BwDP0NksDiB1pfcbYiAif9natYun51pAionEhZW59Ek6r9KRv72jIrBdUhwrOS
hFORJ/n8sIUWTbNG4lSshfwmxsP+wETq6HDP+KnPzP2KCzB0h8VOW4N2xFtky8gEjTlK9L8ADLBV
8t07HUJFFtqt6lw4fGgltE6cP3EAe6DRIY80D9lLUy5EmfZ3Xe2T5jSW1uOn3AYK52uPrGRC5Kx/
NkMiE6jNco461L1eGr1Lbp9LQhHxHOimVnkkMX9MRkDvfcofoFLSNvIPVOr+TRteRn2uJLbPduOq
Big74YZBv7Jd1nsXbnGqLgDXbB5/brGGJ5bAJbPhay4ZBmkw6LBHBn03bbzRyvVNSnHjbKOvan/g
sURpQ340GBBULGJDxDhTfdSHN2cwjiUzVSfs2S6LkItW4xGh8J4WJt/ZpWZmk/zWC/+xExuGhxLb
LlOaqD1ujkpf8hGU3dwiFambqJLYeBNHBzWss4b6+VQFDGCnhItrPbT0ts24IgEfsoSGZoHSPkhJ
YwP2kCclIO3bLped4sEAIVEJTirRMYJI4AnGLMt6ukKvhI/yMZaV/d6W6/vm/S1t0mjPNxa3HVR3
ZJgw30h5ztISXjQv5fg36uYf7xF+aFK6ANWZnrXh+PDmhBbnLJbKGwQhXD+e/xRWjcRhQDShYYcF
xD/qsufouO/PKfK4XCQyWi1xfgA/oQwD2BcUzZ43cHccQS3adYmAnxamlSaLZSrfAwkcYDmxVoL1
BKrTfWsiatSsuOHgmnFjW5uEq9KdGw1D46AdYMyEjvMUPtTn8V4swieqLe+ssOhAeRMumTKYq67i
37cV8yFjfdP6d70kBdUz96o8mght82GMvdCAJwyG1JCi339JHGn1aNHzF/s6op8KfJaV3XA1PoGq
9sMTxXy5TaI2b0EjpV+V4sRhsBnCjDH0KrUqHB8zcczBA/iAuDJjYu0FJ5CUDdADCBYU4fH100Br
r7F4Gq86N/Xrj+hDDkMEC7BcSSuG8t3RUxTw2zT1KA3MOfAfPSxje21uOjcQ+QyuhxuBLzujbibl
vxuTCfzeyz6zMmMzimZjZnov+u9YlQA/WkeVpUINxobo8R3u+ncmzUJfbyaU/lroDUDsFLWk/UuC
JQ/yHKckGq4/et8YaFHgZ6tT3lWz0ynPX6T/wytowMZ2c7FUgKCVvfLuGHo5xK3SKrEYaZP7mLSv
09lQy5R4evVf1S1sZUWXzjxyBev2l8CBSwFx5raUkyaemxw26+MhQ77rWHVaGmpjz/3oUlg7X+FK
z9xNKiEIugPkQdtsX7pG+1tsMiVAkZZCv9ewL4n3QsqJeUIDdXoNFez9tbgVsd5CGSCK2B+sKrA/
IfBMUZdfLy1f0PCCUf89FxWBTfIx+oW6T/Jftm7FTwxT2nidvWdWUpC9HBrPgy0kq5OLXzBt8U1j
9WLeP0iR7yLgyXMxkDK6YPaxYyi+pP+S0gNyKORs06jfnBFOjQmzZL1xPKfdfOjs7lv5aymWcVdI
qrYGMC8ExS+3SMTNCRvoXvvI+vOr2luJjU9AU9yq6Mz8Kw0QUXlMpjRXVZ1AyuaSUUZJjAnSY9AV
EDbQIiL2JONzm95lWrJhXKZjmXGgGfdjU58Amh+IZjz+xeeFaxT+gFn4ocSNGtB3kH25AF58LrgI
bIAcw2JhKqxafpEUhWqZHX5Bd7qDZM29lIYuP+uXlxQ60PFfBV7iubAgJyer0KwIvAlROm3L5DeI
/1edqF5h2hA77/C18xhmDRpdhYLMLe/73WkoQU+0OwkRpZqJcr/41eNK2Beio7cC/qjnNR9LDs45
lqE5vdXlMPgjX79PFVzRexdOe+jjZ5jKsZ9OcCRxT8MrWXllmo5WBblC8r1Ye53gK0pPCEDDaxd4
bGi+zbT2MryUgffz2r+/psmJKNaJ0WBLns9//Xaxhb3gxSzMVVIwuKdjHnu1RhJi2ZM/A2kWtB7H
lAZST50dsyWXRBegok4vCq1JCvH6jXDptdzuUxyNJcmttioQO847pSPCuEudt7+fZ6Y1LW07nW4u
viARFNPImUmnyT8YL982+4bgt1oJ59hhV2vbeOBpLiziqbQsrkDLDLQHxaNyvM8D2Re4lzVgQyS+
SWWpCrM1EUsJMnixvwiyX++LWQ7KdHwXMS2tjLSVL596ik3ryDb8vTPS4CSZR4xodIpXPHqNb3/Z
MfuzTOmOddx61R/qsmzWHNvufVvOaKtUbhQY+WUGB/b1akDQ8O9dDQBGMgaojsuXa0hJ2syCnAuE
VrjXJCuudhE3Bz5AFuXWuTjv09ksmLJgH7Daw1L1mQlWF9Pv/x4tNGUN1Uyh1xB+zrb19Xt00R1o
zKdhpNUcrzAasOC4wRNUan31Y6YMTdFeNt+Y77EeMSUVdpMBpGTR3a+6tQn95YMNs1XxR9ffFhmL
juPYHR0HMY+6gAE+iSZ1k7FbA8JbzJMpc3eYWHPKyL7JyvvVG4s1i8HcbRldb0bUMjtNdFLt1/EY
1pLw4ec8xBXPG8Dh2GY2YfJBSX7sy4SiWv1jjT+mG9VTfly6CFvsHNEBVCypuRRLeu1/codDMLrb
iqcR0n0sRi5aUXZRMte0ZKALWkpDbiOmq10aPLEUPm/NhW40S/Pt39JPYfZq/hiCCg6HxddH0hMo
OkzPrmZ3OJ/Yz41CJAQpgdlH9jvHZw5Ame0FZEbf9kSguzB6CnQHQQ167ua6a+QW/27D4d57garn
sxQegULyt8oVuq4FmzxCgmEPUeown0dpR6CjH+9C7OE1xe/gc4BSg/n/MBMfyWci1mIm4wRvZFd6
6QrWCDxkAxFh3hw5wD20d3XHQGeLsggRR/5pj6iP5vP28MDG5DxsOHt208CcaDYw9r1GoZTxmoqW
OY9cVU/7C+pn73jWGpIivVYeGxfIgC6OWTNSA+2qC6CZim6Vs+hFXu+IEle6c/NqXwgzJP6OfG9s
KhQ4lBVnzVEWrSg2F3bAX9rbhkslA4WxRMLFQBgBOwNedRsdC+9dN1PvX5jAHb4HJr3WpGgR/H34
bsYrAmpeswF7OBnT2gNr9DvDfXL+nhqUlUIYQJDTFs/OeEGYksvVUKdvNkiGWnFJiN4seZjS9wN3
MDRTDeFmYdt0n/+BIbcP9KNFA8KY0u6JxLCFy7p4einFQe3wGe5FPUbhtMRcPjbZJXgiOwxUSKLX
fywX/VtUTZu43rBM9OpJPeE61SSbIIRcH2xtQA+kpUHHGItNFMpbP7UAXlZ6C/6Tm+1wXB38TFj6
QI76tzNnVqqY8N/P2B97FLBVeybrmTUYz2p4WKGlK+ZsF/qqOzKgBFS2Vje+DubgfwyVAn18cW0y
U0m2oN7wDB1LL6RZe76WWJTTiYpobHbdBax2RM38yOtcJTP0GQZJwVxzO1GlcosNeDFCEzTGnyf+
CmJHhMmiLvp8CU7tfxf45Qxc+ULbmJLeERRF3x4myB2KIhMc2dIYfpmd3+9LKOiiJWKnVh9GnZ5P
vf4MrwptgvgOO8972c7L+p7eRjmEHafH75lWQs5sd0QVJuzadFHlru3mjW/IYLQOpjtrJJ2HIF0Y
NcEYcFaaJCE8YEgVv9WFbBgBXXJFcBtkqWOgeOo4CvK6tXFw0/zuB6lEplgE4CU/hlNhJ2qsaK8/
iXPoc/qL9VzK3FBsetFzg9eO7mZENqD2rw1oAILMn1rR097aX10Vh9+qMA982s2xOEq4A7a63JQL
8kS+chi6jKMebayZRWAJ0/41gvZHMQS7Wzhr44UChroyabh0a76qb9ePaqjV8y43yo0Xa4SuTr59
Q5zTbUQbDu7bXHSNGBhEryPWnRryqk5EGZXk5T0vC3r6h928Rvj6iY42mqA3yljrkvOL7uIHwbiH
NttDdNildYpHdpYhapViRG3pVAt1b0z7/WtSXcf4NGO53E8uqy6EmCNU16Awh79iChmQgQV4rdoy
GCjjzVg2mqzHrXkJ0QJ+nodCsL5zAHHyI8ATGPOBLhNDhCxY0lr4xfyoz5xTbarM4UvFVMWd4zMR
ec7KmU/Nel3anqswJ1Nfj+0rh+d7mH4FTUo+YLHP28IxTGT55GPkATYX6hIKFTnNcx3mlVd3zePX
xTnA6HghUGb+jcKf2k34yG7RlHLPNQg9eJ/YN91+3MD1fR5mtRCeYy7tAwFRCJ1kJibIqV+wXyCD
Z+3VnPVz0La9WtViU10NLtmi8QJohW6P7EbcUK5EZu9tUKay62bzDQiSY/2KTt8AlpPLzgF5JJRW
uZiRKevJTjDyPxvZpqry1Y/0s2AXIabMHyM2pIqdzni9r1iFGj+0UmvhhdI2KRVL9T2mYR3CVSlI
7UGdnUj++Pzoq4jQRvZvOVnDFo7ryVP7O6DLs/2HmMlrnVDFDfzknBkWffIJRJtuWt09HrRd6qQV
m+BK69+bzEtry5jPptJY/7mRX6cOQdTsLPoicSSxk4p86cnVWUj4ws8YFz+9d1Q7TFvXzT9AGpte
GciwWEq4w8wqtYvN+txxbfsGpjE7UD+Tj+w57O6ZglvfhQY7JDfYLuNG7QiKBWvO7DIM1AWIGE+8
bc1idONY2ScZM+s9Oxw08xn9eMOUQqfaaml4XW9D6ThWu/G/tZSn8u79ab/NNxXW/GR99751D/NP
3spGVINkUo8JrvF47cRlv1fpdeXrit+HVrnM7MUCtEWi1XK4QZAbAD8FgMONMLuOmbMx2l+zDxzF
xanB+CePdETTrI27xsFp0pRjYAngb4YtbYHp1OGdZ+t3DcUf3sozd+FvGHF32qQaAFZPS/hXJbc9
BtqSYF02Jinkfz3X5z2+kFsFlga0gUM6aPEzjSqsObgdkDHLr7o39TkeH0TI0fdFzi+DYdnndRgF
N/XgG1IUDuBMYSY6l6fpbFmlJTUVygLFV+pl7JMPIcs06jHedTvvETjGQthBLEKWnBwtn9l0oKAU
8Yzfw9y9HCcjLbs/p4XEoZZPeaGYjqoKjXdFjCGTJX+147DU2Cco1zewRmYD9cj7C97ig6MAIanB
q9CIpg/8Bw+bW+YN50kDs9q3Deg9ib8dL9OwuTqL40STesM1ohjAc/cUqZWU9/cV6vol9GZfNAlJ
z7G41sx2gKTFO/GPgKlpEB4B7UtWFwYnXfKK94xbQrQt6g1+T3Ikf3FCTU4P2BbgY19YtUGo4QRa
+vP4lnecCHy9YLwRKojKMqUzMuS5teBzyOIP3UNXlM6hrYxPTfJlOhjNLJUbfj4RnDPfIGib6OAX
yb1l3SWd8oIOI028EGEARvKaajWQGEYpeJRnAJso2n5p8FRW/hUKlvq9fcKVS4m3IlI6JCQs79xv
WHcrPL/SjyYpHUh1aKJzYTYBGoNhe7iEodj2MrGWCz0EQC30kH/GDR1ixB4lYst2ov5SsXn+sO8S
Y8LkTCkqshC2HVILCP9SFn77skfB7x9vxyA4768jgEaupRCPg3GggfdoPmTHZxGa9X3xxCpJ1lps
UWSL7Ev+87Nj7xxSnmREh12UYcNB+FoQuvTFLbWMzBW7NKJEMvvwvofv20RkgO4c50Rb9ZJnxn8C
pzRjAJbnBqMSFVOhtaaf5J0mvE4BQCk2dhoKYpyCbsG4iqRoRAwRNZL0HWjhcJ3bQb75vbwoLppM
dq9dekgKL74kXwR/v6lLtj/8L/QPHjzp4k6oZEk9laDEZo03tgUeCnhv0BcJlMzlId2+rjRRzrQU
QGJ7zgfmTHfjsxbcfycxNkEU7GfvPIGFNhLfD05wqqk/q3sDu8usytQYjaoQUG/zshjlGfxVjliZ
PGbxtLqgeaE9sXZr2qrjMoTdtloKWRvsZY9Js3a9pD3Z4DKGk+Lz3E7SF6Gog3rVPjAVJjifW1Ap
ZxOzShBPrJL6NI/Dr/ptS43Ha7fUfJUS+vTyk9e9jqeDbG2A2BC54shVSuMTZ1HEk0tUiWB8CQXF
Krth5PStssJ6V9qZnSEudqlApDmNqUuUrnIP1m4Q8VULYpt/6V9xSMGtvLPAO/kHPyzc5VvX2EG2
HIILuiF9JKqAnGdhOxTP56UE6O0uvYwSf9kYjh+Mrx5m/YBgylguKCD7uwZUY0HU1/g6EUh0DZmx
AjMXvooA2ucGIz31s8+ANBSxQvp0NMcL02Aqj4JHNbDrwJ6SrXDdru7qt9lVK4MP3eDIBAkN9Zdj
LHfFKPLIaOHpMdwtTzpAPF8r6tgP2a7kkP9y3XZ0Lk0Kj1I5O+bCfpsucIwjLFKmYzXWwBUIt6Mt
wuW+Ax8MaZcQWylZGe6IvcDaJD+6mJyUvpRA6gAcdR7B3mU+hGLUQJe5hgYhqqxTxzPJGkaDidKb
BrfHmoLloac+GKIQB8uSQZURAUPc60LLK2nRLuR8htxZWz6NvnqWxLyok8VAwTvSk7O3hGTZT0YR
xLI6PkkJBJQFkmWU1ggwjVYD1XyrPadly0VDZeVIc0j/mysJfriDEsZd0K8EV5P5mxF3BG6K2pte
CSK2JW3lr/h/7wKMrgHusjUlsiSMxzFjskWyY6tYrLX2MOSnEX1H6bviIaB81YlKJzJ0jv1Y2781
DIyZftYZnu7qpQhCEfD4yBLmsnTJ8utC+8jU+SDKRXJHgfXeq5kfh0/BmnkYRGBDhGQnpgtaT0jW
2W845sJLD22qfwFpz94t/BMUiX5at0Zh6g189J+86OuanklhXBIjwZreYPC4r6HRTM7Hst9rcNki
Me8Ma96+9wPD+mM93geLPezYwAxdizRpoBLKRrFZs6fj98t8uYHoTOVzTltRZPoA/eQW52BxVe99
ch0NsChjiz+GWI9ozXxXMZByxX/ACUNHxSIMufwzsFvTBae1Oby2ZWCWxhGQAxxwLO0CWfyYaVYp
MzbH6QjACPbu9JeUZMQcDgUkuP+7I+dwNniUDP+yKzFu6GVihXJU3x7ZDfkghBQxvoLx5vl3/2dU
ie9+UIvQc7W+vZY/gn69Sm0gZdmjZTqUZ8yCsLevDfboFOMSduDMamDjh/nKbCgFLgn9aII2QosE
bWUKrP0NsSfVHNuEVgq8zFIu9P9ICi/bXijOBjD4slb+5yZQtXAANxuJyDpTX5hoxZTFxfUs0kyt
z/pmCpAKDs8A8VhQ/hu5lj/Sm8nMy2p1f5LeLOHnO3eT5fdE0MHKjd6A0mVgQBFxLGCJPEqmsmzO
6fijc5qVrqdyGG2BfAE6G8cB5N8hyLC+65TN0tiEU1ZZ1YAsyz92j3yntlxxHl0gWp6nACCSSWmW
6rYRN2nuDpG+bxg2OXixOIENur/nrSyBVqNlBOPsMEwNOhSu/KJEqZZna5d+35Dm+Nl0Z9Zi8VgR
/lhaKMPUOE7mr2px+kbFBB8UgxWpUCeLhZ/cpD3tGkkesLC4lROU46gbu+2vPLh5mmW/2lQF1Od5
Whi3+DNmEOBKQxnNVGEyNTlG3dwUAacfKGWSMkWFgiDreRab+da259huV6+7vohnr8xeXaUeuwrE
wiXgguzhKYcYCVnthUxNRqayWW02c7a69xKvNuJIojVE5ZM4sBW0aCVmrWZ+JxrN36iYNlNuRGPz
LDzRrgO6tiwPzjvfw6ZijBd5JT7y50SGOgWGBo+9puTjeciR8hW4EwR31f1erqnWR0/aKJ7Fs9wa
dFxtxNa3CUBNxgaFOa0BD85m92KDrIC42XkZlneZoD46zgwGk7H4Y7HRKqs9hycPLIQYjgW40ilV
bV2la6upZ8qMor7drxae2dE8nPc+Nd4djrDBw90MxhweP18Wq4FYYqcecS/qLS/65/WtytkZcKoT
yL6Rdv+wFM5KciT6PReuDV134fb9X/szqrVzIoSg329xE2QWMiDGDjfLQaPxgT47TZqnVcZI/2FH
QrsvGdpAfaJGpt2U3i8M67bprnL6vueNKqg7wGCncFCpaK0kDKPjOOfFExT+2/ZOrhnKcUwc8UqK
ZIcNPpPMGnxZPheuINpMm7CV/GMzGydOhqmvqXPM+vxcldu3Yeajr4YTpRfMc3UzEh+T474s8SuM
QkwCB+2ALbjciZU7o22flua7iok3hoNqlYewQ7xeWRsPaAC0fDMGq6PpVPKGPxDgf5Z8nrT8ZQdw
ofQSCu+0T69w62/2u9zRniiFlVYYD8LPKBbPXZKJbo1WZ7tb1PoZNQYRG9uoMTARS7TExO4o7kJ0
D89qJ/QJsqFqOPL2/A70nEzedZv+fB591xyfdSu1z0BqmXC1RFtXqbmrOpFID3DE0ANsKJmkTalM
FOA3itejplRHooBfeIFUR9EGF7NiLHDMDwpXTNfYwz38jsze3qT7dF9j+lmd4LQz7S+2GGPn2Fez
PJSrKh8/4y1uC/K+252uQtdCecZjuNWjkF7OobOSzgoiqVsYZsbPSeGy1oka3hAAqS7EpP7cxSow
g26/2mOBoRpa5DYgPXO7Mi+K7Zhb3xB52vydvpN5/L0O16xGqDUKyWsk6vuWP2iHwLtOjHHbCK4P
9Cs6DLNZ1KYTw0RrtNpux1oSmhegIuGrw9d7Ltm8JUY8TnHK5YtNsWw/B19/dM0RJ5m7bJ2+0XDH
rdAs1zLIvMLMEr9lFkO90NrHwIB6O0TLJqu/qiiVU/Tgrb313Tbcpe+GT/Ko8JW2WRsaAFIjYsXe
dpGUwQP9sSTSU1qDYq69MhWKZrTVcucrXDmYbxw66RSHLYId4Y0kq3njdanOxI6hjVOt7C8+F5B5
7wfxdVSA4iUjsaemKbUh3pnvZc4aBqfPpJC9jyTxM6+GecHzg+mFQtVMB3iMa0Plr+2kumoWui2b
hwyGKdGYnL8PhvFfNRHY4aKlAHt4n/tZ/Y9A3OhnLJCP6yvDhxBoWD8EXeR2LV4OpIHnWCtIdcUI
2hdmGQgNXugVt8UOGrzheHAqI9xmnglgOqM603knsjUFZp626aFCH1joIIeB7wmVqUpNqrV3EtpD
6W9kbtvgVJvupWeehzjkfSJG8a7EXX643Mghd8fX+WzRIC+AE8Svr/jc4pTDSOXhtRv71o129eRG
fyO1kHcNqS+VKg51iRBKF4VSWYVCy6MP1vVyHzpV0GQaJOdn2txcE7WzzLGTw8fTrIZK34+h8LGf
GrbTlSS44tfJypY2lzBKpZMwB3dUdn3UlqSVBGVdsWfRe3C2H5/v1Tb8hZhjC4QYxxVrF8YIKPKF
H+52Wsys6f4eAQSl9ZSvdO93qdOsKr6UKevArDYkZSU9Nrf/CE6lJZjIce0aX4uNlSR+ZY2nLWGt
PERjjshcfOBDSkqV76nElfqHXw6aG5CzQgHbnqXiq4sPMAUsZqhb5lZ+zbyFVUunvxt6diNB77jV
R/XyNbvxGuY2dfSeHVWul4RgT0qahZbSGrBYbMCJ4Ebx0/yRnE/cuV3jVMbqZGDUQxTppGrm+Hi/
ra1okKOrWDVLJmZvr5W0dn0FOJxekvG25XHinpHXwMY3D1ruumLfuWFXWZD7c3w6MIkIEzQ1XuQn
wFuPJWtqU2zfTP9NMFfJSzBerRg7FmuC3T0yEvl+QeYaavnTznpmCCAiBy40YZQk/r+v2WMPqdD0
v3vgjtYHOaCbfVXIijgUhJQmbdDAEUMntbDx9Fau6G1g6XVMFVpwTrtw29ad65jnflbE6lhzHsjB
JJ6cNP7o9D2FDpobTjIY6WcLTTHDvM1Fc3239hiUKFMS2XT7z6HazHSZgtYugTEs+IlAm4SEj3k3
VqhXQCPC5Qo08MGinaawNjT0jO1Jb7zu9g8k2/DHv2UOYeZyT0ejh6ZlcrS08vaPuNy01pO7nMDM
fJlYF2DPQHQM71N67eoCYBIjFog7NDTN96tBsQ0obM6MSQz0DBV2qcxlo9yVjDoPoKFySW2LMGMY
3mw1Cu0Z7nA9D6cjYoIEcOgM5uW7bdM/AAqWtseIFvMuY6f129WP2Wb6AS9/pBEuQ9WnEuAgIuMY
mcja05m9gxXhZqEApxyf9KbGL71lFim9e+8Jgp0OyHVRLvKYoj8FhcHpdVRpqplAM0naobTz3cc9
wl8EW2KmeNPNrG30LEtujraKvYul0QC7YYwMEsSTh3A6NY07WKjpj/Ia02kYZqTFHSUU1KzO9nUn
pnPwGnYcwRFvz7P2MIRLWd8tqgiH0eOfA7sUSGLduOekiUcebB+dQaEU55qu+ci/MgNyo5km29P4
du6wVcK+2+rVe6/eltBj9Z6lgCrX4vrLoKSBNuSjJLficQfRHkbbtyZt/loerATz7+TdWlFk3jFm
VceBwuWVfabPxq4VMPEHNhRiIdSD5dPVREB5YNSVNomrv6RjITztO+ASJQQoLA3Kpl81d40HA5C3
Lbc5vmq3p+rW9kUEz6jrf3nRO++pYQpYCxbLpVwxt2lsl79e3iPyElvcI0VzueI+7blZ9nV/sZ9n
QVQGmtn8zzLB+WYXnNigTNd8/PFLSAISITr5Z7EZrK9vWxH+41lbWqMYBjjDg1z2ooXue9OEmeNd
EY5KCgHpVBT9VB1rUD8hmFju+BIwl/Qj9XpTcXYu/eXaFJoPeb55yGd4lH+de/lB02VglwP01QGK
6w2FqTW3vpPe/qA6Zt/zKMwPtPDAzpsFhwEciKOSQjmtxO8dykYAfHH/dmsDNQWWd0YmHe/OnVMP
4/m/rRicKUHowpZFtO3iAJbjZRFv4jPNF1CX9I2yxHrHzOJ2OGcmYajYWqeBySC3q/RL+hhM9Pru
rQ4fSTUgG+y8gYkXldYxh5MQf1aODMZKF0PqHRtNvxAlU9xN6KHleqkK7qQmLSbecwYqMD5YYndl
7s82ZOZO1xfNpM/NAumw78t2KWTbyMt5u4AwLSnrFWUGro5dcLMg3M/Oo56WiioyxtIZn8w0ULID
Y882vRarrsZAXqBa4SSZea9dCRGfBWe5DbW6Tz2Nqhsl9a7M2du7L34LfYNVRcvZAIzgg8NNqqrU
ig0j9bAT2CO39PAx+H5RvGikbSsteRgtfMgpbF+l1/+RD0jzeNnsEwHTT1/k/zIHoWHXrOw8MEGU
LQLxFss2L2Do3r7H6OKWFSU7SIwEwt9hq2R4+wLSp+S6FaIygV2Hfk62E1TQWOqk6Jh7sp16Wc4/
r4B6SMqINlML75m8tJTn9KjZiMyGLXeKtxNPFvqIdU3x+LeGv3W6OC5dughFYp1GvrnQ/bf6M/Xf
phbXwvBLZdegM6WZHUnq30MXm1ksh51ktyw09BlC+ZaNilKPwixoBvV6GtSLbgvsClaqTPmy1PAI
DhTQ5KCAClE3D4lyeGvRH5f48Hlvp5AUkTt398GelRAYsULlVkzYY/dR7+IdKW4Evru8nn8evQEU
Z5EZrIkkR21Jju64A9TRUD8IOt3H6PkywKw2nMdzjLiv2YyTxgY0CNd76TeuKYb8lGpgSTfgABCf
8DXThEFpfmJHu0tZfJNO8r1g7ACDwaxx289+i4+M7wNVu32ldEmCcXu7hvnmjMOqfyj2JbV9pygd
5TecY0n4DEfVH1KN6DsyKjTkvGodFvxMMc55M5qvAIMBfXFsFGFH0cvWrX5gqv0HELdMn1p4HbRw
z87e3nkIVNLBCB5xGGZHtf35BKwztMyECZpl0rkzGxsN/q8qEe2JORLsyAujRSTENL3pRYdVZaXa
jeYQzKnsWCZD/+a+Kc6i5r+J4IhWE6Tx6fz2jcQoVdGn5dgme+1xujBwUjXjm9ZUps4fdDaN8nrO
0IBAOPQrLlzjV78lCl3ldh0jXm6ieEw6rCNNVKXMs6dtRABuZxN4TV3gOd2WtPghIrp94ym/xZ4q
tRuAmSVVcH/rJv+xlWZMTYktSrHUHyvrH7GM52KDXcQ8OZE5WdMSraYigmDH6Pcv1Uq6fHf4hUH2
A5mAkoOujNAeMvo/rwIdrFWk/TSPI6XMDzfPT1WBOcdD7bWtMTb1T4RQA27WwTA+0kjIJ4JozRYo
nEBve9+Xn+9hZjPk91h6g/d+8f4dIM3sus3iEDonqnY4M/nP3LWe4N48iSVeOcvdDFpV0vNXcbaX
cxrQWKWSk6grWfHoD70JaxPrsQ22trs8QvitZar521PRCC+b/97DEBxPLogv2QOEiJlYQexfHZBA
ioX9xzJ3w3z++LjKZgxXCBEcmuVG3pEf08+R3RcVdxq1MW42mJJDegahpabo95V4ENgqHtM3qURn
EGajaAfBsYr/4P0rQo76Bb5YfxGxtI3znhtUPdhaS1C39fvWF0J1t3iLU28HA6IDeFWVcroGCxyi
TxFNRG1RnZSaYhrbD57RRrLIl3nLbrSpCctoiUZhsoC7CQsY6ii6+FHFF9yHRZjC95xlR8mznI7H
nDID1e+BkIf8XNTzxOx1NLdAVsZE6VaDK8b999AJkaUB+fQmCo9p908hMYou0yf+qkmaeZP8cxGn
CKgG5uYhO5TaVQ3X/y7WsrA6fIbmpdXDIFC0sryhI5NVCZSEx3yL4j1ipOmBAJEkWs6dHQ43VoHX
ec3El69Pv6rVL2On59cg/W4Se7MPearMskiGCVPjt1l4R0TXnIjuNyfdOaGUb1kLSQH450wKeJpm
5/Nsf8zBpJxKWs34nqf411qxM9t6b1PL00QPHRhPwlPAy565V7jy6lE1rzc1VdNFDL5Vc+f+VWMs
dQgiYshh2sjgvHDYVEZb6ctqSlJ+mh35U7u1YoQuA2VgQuKWUORULNlAh+VfYpjGGnMQzeTuoDc/
XbCue2D35c5LDur2li3ZP/6WYOCKXekeWcfg0qpQXbipW0vcyB/3hmVm1cwB91La6Yse4cvRLfjs
co/j6FDSvUGsfUstb+9qyCNtpXBhgmjOJZYwI70dW2G1ZL+yZlwaIYrZaqe93weGaBpx5oOOh3h9
Lj9MHLDtdw/exu/8Y3bFmYtow9Qw4n3S44bOQAJ6xg7osV5sqkUQ6t0Q/NWoL4Bvrl+Sycqpxd/k
i9/ve/2Gp6OlvWEekQTu3a6mkmZpROkfWVNtkYMgSVEhYqCmlhbfOIJWsSSV1l4w4suGHrekA61b
LDR/C/aaSk4+pTGhyKBKI8K1ShsrGPc0Lhadnx9fooBEmaK6xjEeGtgCxseBCvaiZaVU60to1cXM
J3H0asVgAPhMnvmszZ/WiEz8IEQwtx3DraOEbQ22qUoZ4fMvgkGqOjULzQoiwfYGW5AjpFl8AV4f
EhJCiHhovNKzw7R8uaHHkPEGwIqbOrSLLVut11/miHoDFWrkYW2bS/gtTsMkq0NGH5D57y5V4hvU
on/ww6Zs67Gn+l0K4SiNC9iYyFgz6DI8T3EC0HNxDSVkVamek0d2F9pb0e39A9jCvsmT3GFesviP
KqA73l0SaGezAbjd4jhztrBhqbPiR0akdIZOsvLAqMOgoOhRRIi1kfZsZDXZuYHRgiFzxv50+2iz
7FbrYZlvSpA1fFs+NkRg1IyS1YbQCmfIStxZyD14Sy//yk6WywacDZn9luvoVCQihcoDAEqJ52pV
4Hc4FiYIr7b3J+DR2SMkIlyB/aQFo/I+glm8UdVrPW3ea/G7vrLJlSZ4hsO/ZfvvLlCKfxQ58KF4
3QW/1vzW9dEoKcbD1xOXmXynUfgRAEYxtk51hcpcI3u2trL4FZJbT99s5m3pjAoIwLjm0abAET2Z
Z+e6l7EZSgjimt7IduY6aEMjgXKSXU6NGkFxds/o4lLDoi7q4N4woNzF7W4IwEUmS1KPsA/Xq4pP
fLhKu3GQIQwptHQesruNJLvV5GfF3tyENnIHPzdPJgrchA4PzALgowyo4w72OvDT3U4VDVooyxtk
2VEzLiAoc/CrlAaMoi7D64zIsAz53KRdLlquzBwSx4EEfbOMbV5P5O0R+MjMD9PKM5ACuRigJsxF
Knb33FgVn2mKYvIbBTb51yoPkAYKnjdJjRNPDXGHlOxgKALg9bvyXbJ09uPCSquo3Af9i0tyBLgj
1x3k3XgEtysm/vF7qBaRk+gPvNlt1ulzL+Da4gWFIu0lPyVucEl4FXoB7CrqNeU9Io4IB+/AJSYW
njiDGZPuIslO1uxFymIZOf5eFA3u86uUX4yUuS0ozFDUDxx8CzRYjt3vb7qFh0SS9hpDxsJcown9
DKpdZ6JxPgRvSpIb5GIZlxRqtVVG3+BnRcatVR1XCs/N7ZiNibhQEnAFWj5PrrlEz1u40mWsif9/
QPZ0aCoVXx9NVaxlr4FrZ1XCBFwtcSXzpfYWNXuZ5cBoDdl7N3S1e3DgKTmFWx4wXuSYOVphNzVd
fs16riYmYl4ej35y8qibq02wtxQN4jfD7g3S3wWBcKjhbPjIAxakdKJQSJsXBebIIRXJ/o/PMQBp
O+WVTPXT3wi/7iE5yqOcTGpvjR3lyx6XQA6iWUNOaLL5OLkVslRNBij316zXcAkBcMHKZ6sRVnSJ
GIlGvw1SL00AGRJdq/i6IUqmvArMfdmUythrxTWYBPKtIAsc0936yGyLz+Q8no3Ll7N/ErZnPg5M
qpgRAQ3hL/ZYfzPLVq925t42r8BTPKUa357MR8oNYT3yJmq0eNEJojXMdIU/KfJ6Xxu1+Imn0T43
3MGZw7hcXMhjILHZjuj0+y1eAKVSazUzcNrTRCazTUUvEKhiYhnYkcHiOM2NW0NMMz7OvcF0Z+Ub
LMSeHURjp5KsLayiCgouIBhT1yQcSOmWPUYYLj326o41R0iVw6VTWmEucLwF5lJU63yix7xcuz8n
i8tmHUsmpjBU+jEWpVToOmfCTlCgNOM5f3POJf1yjd1Hvhu2lsrWbc4yofQ0XwnSlPzMO9Ntuf87
N0tWUos4RN8K4ShcIviBAMIF0ttbeYf/JCcrAoAinNScAM98dgt1/WZHCDCE6maXuJsjIqT5xIN7
a4eKVV2S0QiWiwnEwiBGszum/2xYuNDwRDrrdx6IVJYm9dyVsibGNTpZysjDa50TFq2GEfYvFyw3
FPuJQhpdk1ODe7SzNfOkEfGROzF9BvlEXsDfyhilVtsjli8G0RMuxE19Qp4ZIl4o3bWZE/gwE5Op
VLb5YzyrnwoJhLvCAS3JbmaAuQht+lpNKvo3M8DneGhqQHO6gF4q1TLbqCLU7wOqDwXAvcJq3Er6
YKhzgLwI9VubdNaQJrKaDsP/oIsKIrnDK8Pgkey7yxF5BFk3aIl5eS1ViTTy/W0/NDca4spRscI0
4FCfBMoqOFvrGk+Xo07CUKlWX6Z4cEPvHtcC1HC4/n1B0rTa0d26umrQI00u0wWb4wwjqm+jF3RH
0zI9EUFhnPGYDITufV/M0aKnRS5JpjULrME+rstFoo+Ua/99iqlHvRqjZTDdrBeIxTzs26/ncWsM
Zn1NMT8s/RN5kAXAtL7+LXHVWgFU6IvbT9BiVuGhtJekJEYCf9YSD5UyxjsA/aGpka0i7hDjBTqD
urlxXlSl8OUXQqc/Kau4x2+iw5ECF0eVjCJfispuGNWHLc9EB1cIlgIuwYpVmwY7RwZAJj8m4w4w
+Gxx4ha7pJluO//TUw9ed2R7nTy04kT1QaKfCQ6fyOAmv3a4g/a4TiMbF/wehspOWjqIbeerIvBe
HgQ4unIYdVmF5NF0Hk0tCXXSxtNflrecPRAhzQIblr0Dc/Im1dJ+tcK2sBv2nE/8kmKwyeD3vSJu
Gbe5uDua8hFeU6RZYiyV/g09/96x+m8yrZHj42oyIZhjdNQjcZ+Tnx9RIRHpBwmIRhkFYd7OXx8s
+hLYiXYkeo9rT5dX//TDAr5eECZHQslNKXaA/OAgo02eoGGCl8SkOqgecnS7F4OrvhHP1o8wBifV
KdiioDg+3Oo+UEKLsEDBzOJFPIInV5627C7NHD9kAQVwbGjXC8pVNNLzUKUaqNyhcL3MXVGP/gCR
eAcXpRsfjSa/H8Yep9CMA+hgLiN5HKG5Vy1LgRDrb7ErpKPGXG571PAqQgxj6l0wBVsFBwyL/385
TUA7s9cZWzxUMz4XZhkX7ltRBn592XKSJbodIkSG9TUlRJUptsp5UbYmKDbOUM8Kp/CcRzxrgTjV
kdLuSQBSZubogWl2ET9LYfnR6TG/6GPAv1LaokGMEV+dqn2QgZHphGEf/6E/R88BP4f7O9x4jAMt
I+SFLALvtZSBQ+lg+K/MNCRu9AC6kIHcc1YV+M7tpm7V8gDHALOFGQeCVGfGsux/Bg7RTFoChoa/
AtYkWkC71Mg865lufaUirHufxRd+AgGwqdySx4hTQ4ubzpV0yGOUMzO0/fDZh35uIjUTYaaxoNGV
lduG+sgMYH8gZgS6zlGJcuJ4Qq2mTO5ysolahb3ISGKz++P6+rfbxg+pLQOipWzRveJ+TpOm4xCj
OkX4GlClWWYBn4R4PP9kfSXaNCQYF2o6Qj4DfMIDo086H50pK5l17wkTNjlByl17TqwiWiZ+sap6
E4Ng6WRF947VrC3rw4S9UXvc50k9Z6FZ/1zogEC7tJ6wYus0zU9e2n/yFjSSguwykdavgc5/huuO
eEjkDMS59iNoc9yYQJ3smD244qKFRgJTIZIpb6tQA9U8+I0tcFEV69ekg2QL9ra2/xLYE9HoY1rB
gZA8VHvP/QFXqgz5nWCUUapDcEC4G8Z5y/6KhVsBCf0pOFB5Wo4mL0FGULmYXrHh4vytG1qNhRhr
OOxVVyrigtHJvDRyZuhIz5AgKkUjBuNBBSINHotsRM6hiatwhpopR45jMQr/i/eEKXTaq69yzgk4
xCi/piYP/v/IyGR9BHAwYaNsY8V74HvxNmY3hNXbdu/jRTU6oeTXPN+JXMwyFm/DsAbAuC5c6ZN+
bmv23WcNXX5ELvs1+AeJPZuwqMJF+wzg6048jP5gXHjq8scbhG9JUsCuotl4E2sW5pfzEXVaGT+p
5iKLPNwRgLWuwQEUOaP9pQVnG5uS72foVJdhkbmjvzZMsj6+JEuXgK+41imYLB40od2iIa7lhGY/
ZnMNW7gUwYJpUeVeKP+lL2JhGVAK8vVmetWhD7AdmJmg6nuKxA2WwuGXJf3vtIjHUFqDLD0FKZZM
DOmwoi5HUS4bPN+fnkcu8uqoNolsGAaiTFBPQWUVMkwxhgpQwicF8yWV7+nN3lRgmTY23lirM9+D
HaGL/J5w5gZSaonKKnMtOErsT7t6ntmDmKiJDZtcAC7ju56wpgvtLqjDpYgbj4r07/6ymP5ir4gZ
ifCwlVS+w/h0+O2wE4QSf3TT8PO43kZntnoWNa+OEWOa8dWPkGE6WsVMRDrpX534i6ChZPb4BqG9
qskCfsLa2yKhdO9a0mzn5sLcQ86osWUGOGQ0cTiaFfNF/moDY0oGu1PqujQfRa34FFpweG+16zPS
DxjrU1fZVDAeK4dR450Wy6JOTbUOnQY+Z5PJMDEbmdnHwBxyEapo3BtIL08l2KgeW3bwIQr3FHse
npd4ND+z6yml9VYsdQYja9cNVRgH3HOPYLP3scyxzRcoZPpF4j1JIIjurdRBzssJfif2Y9fvY+cN
kx14CBRwYYynm8UDmd4cS323FG3hcmwvJoNhM8mzAW0G1kXZyQfhToALc52O+tGyTFidmWBLt+B6
jodiZW09WLAzlFXK5PMw/sVti45oPvVpQWqzCh5Nd4lRN3ChYgyfwUaf48VnTozqQGOs2R9W7tSI
6KMnseywBfx/8ti996mcOMiv1g/mygOv0pmzpS0DHy87QKOayGqs+jV8qG3K/OtSfd9SDWcBhut3
G2TzMT0x+uMHuD+dB7/XAEg31oVktiN4oiJdECY+r04jxX8w0BkR94vYCbUZiVT+wg1rF5+2QoXN
ZrOOZcpSzIFUMvDZ3mXV/b0xeuefB/1QkvB7f8VfesaiCfZmhgpnqfflUgAV0eCTDwEsK2zkJ17N
LGjld4MFi904+pqQv98R0uNAKUr67Rl5BWExSZf+IUAioKH0alQniaVqvpyzT30LZO/+CfItVxyy
1VTLAKhhpAzL/vakRbA2+JVWo45w84nSSS00B1FfQH1PZ308s+BlHtQRbxa4VLOEjGTNmPeWw4mr
ERe/3dBu00zfSvEtf1zKqdiV74aQIwAUorDYgrtQZG4cL9RM48+Tx7lTWlo1cvg3Cv9YdxUXZ7Q2
c515C2UQYwEWm+NF+MfWd/8MoMxVCB+T6PbpmYtBrpUrJtGKf7LbdB2PYeG4by0XETUdvwKRKAGh
mSl3+YVI2uFCy6YukqjhkdNPBo9p+v5pBekB64AnVKg37866UTmPnTXqhR5tFwve9k+QpyUhYqZK
taH2pbyaAaQXXzNf8FHSafLJIArq/misqaGdWJ9VaNl85jS/50T27TmGXARImvNkYxNTPX7/6p4w
YqR5MJiRLJqW7dGZt6CHlXz6qFbaG8tcQstV04zryDIXnuhJcTiBXs3ZqOk5kETlfwAkU1g2t1pt
n5KpS+Wl1Xb0x9UoRCpNC0hqiLlP8c2u3kzvc9U9nCMB/39ObF0w8z9fgmY04Yp3fwRQpN+YXLwa
S6+H3xZ2i/dMoshg4ImeCu2KvGDGQ1H26RuEmDqY0Yb4HNMqXMZO4gMJr79xuAxD828Vik6ZQxvk
ffzK1YAfR5qV+2N9o6Fc55fTPAcDx4uOH3iGWhyeVuPoHH9jFfiTDiW+qCl+ZetNxtryeDOX00nS
xBK3fFT6XgBT8rhTXL9CdOj3TCsz7BFe+1WoEq4HriD0ARRaKZ9NHdETs4fgQrsZO7DDka4Ssvrj
vHeZ6QNjNY3v+PqBtuYxkeaqZQxur0DQMqx0bfvN/rAoIUuwlb48pZ4k2Kwk5v4zPsi1tySsppo7
SyYFFuwrH519uEXPOW1WAXPjBWsW1lbDnRTu+3ZA+rFnfoasohvkZARTljxMUvw80tfsFUD8FlTA
8+cNE/jdFtDDFj/81J/1Wa1mnKiQmmxEduKKI2FY3Mj+2sUKWs0JqjJwzChB3y10zahTU70U5cKe
78tz0YgayRZYcNMIkEnkG0XbyIes9coYHHwcBOioVLZAxSBlkYBFDlHzvuqiLXY3nTYUJYA/b0n9
Rfns0OPJ84rfwQUKzzQalpDF7xSkldLscUJvbtrnYaOzOreGpW4Gi6LvJlhZJpt8nO0PdN/DDyaJ
8u/h4E9kUKfvfBbpHPMRI4j+S+vIYpiVX0nB2hicg9EoHCiyvVZz1EP2R43tjHNWIW/mgM+/6L/1
ksgixeWo3P5YEudW6LzVB3j8VKre8sWaa3moATe6dQlgEgWLBaHueBeCENEsFaDRirvWPsUk+/kd
63+rSkFpwanDPcg48DzB/swR2kcRPtRZyJyaUVEH+FbVTwOpTj9ZdmXq/aKr3tHLDtPPdEOcUbU9
PT1dIpoKXooQUvb5bx9hhKHw0XkDOLenLgFoFE04yi+i8QWHqmhQX6lUfxNBrB2aHKLj7K6M1k9x
YCvM0JH9iBjUAQ0VQJOLqluwlEurgvaV9gTVVxs+Oa5yqQnIeaVPZ2lBSB/g3igcL7YsfZ55miyF
+xW1kxcEhIcHHPVGyoNJbMyYxuK0MAkEGZyWZps2+iqpTy+hxV/x+l9joCjT2YrD0uAmh7+N1/58
Gch4Qi6yA7QT8Iq4rHlcdhI0InSimKfaL+hOWPr8/nL8MwWF0TT4PNu92EwS6A+SSTLKAb1tPJLo
y3hcEgKCOs14+ek4JBBBpFCT3azJ8eV5UM+C+aizPX59Xo80YmsK1GkhJSx9QS/qTY4R3ZUTjIbV
+CPZVMbZC+/xKwZLT8DOuqExV/ejRxcTs/pSj4Gc33B7+Y7KMWZgTwbtOZEuhGJffo9bmfAO9XHg
byoSn9b1NV9sKrJXlEXnXeLmACc9v4zdVPGPTpTwIGxfObY4J5UdXfbcIRBxySMLYPt4ezNBNXkb
Cj3UR/iwjDSGvf+VVHmafgBPh+1yUABayZHW5VI5TFpH3Mn9BoSE1Cw6O0twhRsNMWCSP13RbdyH
xVieBw5sBtCxwRJDuuB99ach7EyjoYqy2i0kXjDusrQEf+8dkzueziu2oRECwjdAUqA7MBWPI3X9
7mSG4HJg4pJ1vb+1Y6O2EdcPK3rP9lx6j3Pr21xb9ye9yOU+VWo6RPoAlxiXSS/LLxeBEQBzlsMV
1gdhYOGvF0B6IajVFEF+/sbq0ejsUFo8lXIur6kbNcTGGiqjd5NhqnBenSjWJlYdKCVc6rXJgc5+
/L1JOwI8hOaIgjQu1vvy6LvjD1CNBQEwIvYqyDqc6qPnhXg3HObJNMjA3TBaVtL5vzPU3ArWAkUp
kYp9ltHaEcSM+pIH/gnyAljjaDaJmd5NEK3EsOSoteANE4hZVTSKGu4Wz1z5B4x0ry+z7vRjDlKl
VtKKS6v5SW6lmCJNsRu/DakErxVTszg28N/WwU6Cof/TRNYDngd9EOVjKW0g3ssjl6/SF4WcNQes
uAcYo4mQmQhVmkUiovED4NGhOtknx1ye20IMAFgByFhhMnjsAT4a+JiB/VxGWxlrQqj3dTqZXoHm
uOlK7reNHtE8Bvt9kxlnrpEgaXWi7ieveNfo/NT6lSZScCRRQJdV5/SVS14Gr48BpViz2smpbDPg
UfHV73rvhJlao1r+wn/Wk2ahCjgDt0d4J1z2TEiyx3Z+BGIyWbz0yF2nd2PMl/vwtnRcY2f0l6c6
nfmR4L3B4K2oAelmoC5gqa82i5dYfFYQYsLCG/VXl3NtPFI8So+99MonHLGSPgGmw92Uyxk4tI8b
pEFb/VYKXpsWIHlwCGQ0juaNv0qmRfuDIfm+v3eAabAmicDF+A0yPZnxAhBMWZHuotum1uo8dydY
hw3aEM95h9atIo6YVgfkLFGwCLQo936hXBkns/jGtnX5a/IPcHCCq9Fgw3/2Fj/HObEArmJE97ZH
sm0HSUYBY736ix4M19G4qj18ebj/3djQsaP/ua3mlbLBgg5y5vNCdtV9HminVjtxE5g/NgSLaUnk
UT7LcCDVjVdGXgQ9V3lt+9Q/6YHniKZUBGpfhzQNgl0b+npwLqnPLnBBzTlLhEz2HeUUGO9c2vrm
Kn6Sm/i+1o6g1XiwcrjwDn/tz7mK48y9rwUBcCkHwwev2R7ck7Nq0J5SXnGNv56DtmlL6MIEqxVk
Gz8RFyYzTG9tLpLLKTZ4OiTMyUtFRcGRhEmb34jFbaGAbhBJIHziqDb739bG6ysQlHj7BSLelCJv
jtetdsydLHOuMvYW2bdchkxLzb/P9PsGhDAW0JY/YS+ZuPSXTYhKJp4Xr7oPvqmldEEBmSA2hHjb
UJKlMTT3LDDeypiW5f/S9jmMzUrR16TJfojGiyhtsRGa1pnLcP9F4pdWok7ycztkUN33PXtF2xgh
Ro1UqUFOV3PzwoTkFRzBHOpedie9XVE7lVYxClEKadDnjKu2CESLpqCmlcKUCUvETwVQBwyI9JEj
Ha+a/Ely/NcDJ3Q3ij+zjKbtGRpQ472PaZX964Q2r/mxokfvpDMvOuwlx6l4IJwvPd6GEUVTfRGG
yzKNHON/NJdtuiIwqw68498q0dT5eIZEtziT0i4tlQtY9aqwHZ6etgUpEaDhMKUTAGGRwbssByl+
o8rwtzxjAuVdQ+lBdg/Nv9PP6CnqOGo+fjAQJlUwK3MwmDpox0LgVmGPn9SIt81g3P1Egv9/nOQ0
yoU1NNkN7Bcxf5xbwGcBL240TvgFXHrJRbpxb8HyEkOJNmw1HyxvDBqU+WX6J5cmR8HMeTgCMQ8s
IDP6Wbn6F1SLVi4298gN09B0tS3aJ2Lw/JqASuOsG/zn5jBRMAf/xtGZIpj3D4rxqzEiskd79snK
F+qkVKNFFHmwvo+9pRhpoV/2LTYReauijkSaDqE0+EgAQyzWpuLkjdopMk/7v6+56SYe2TPjFlrw
E02KxLXKCpBzC1WFkWo6AOgeHyRc3h3oWWueIiUACdWkmstnL8ZTy5K0dFxFOZcBdHhnnWlO7efW
qzRp5GE2yBeusMMCQ47ieJDw0StpqMOXlt0pGI0lwypej5FzV0ZweUROXEAD6jUPH8a82EO56N3j
IkZ9WFhmsGPvgxB4Ut/cSgytVW48mBLBxMCe2YHsIWNnW+aI6HxeiLcOUCZh0b+nQmYrgdQD1UW4
okXo1KMMmewZp3bFu60jaZhcWwb7D7pnQQYlp4qA0jJGu8lDLXON2lNy9B0qMWV28Exe2s5uwOrP
g34fuTm8mXyND44Mk7UUTMHkeU/Gdgu7plZuAeAnZjxxFRtBt1IuWOMe48z0MHcsE80fRe+ooezH
gHQpyR1/qYjiSWBY+oZDuN1UJMf0+uBjpjzZHxvkNdFiJIBlKtBDeedKsCpyMwsi0uqhgLfyXa6Y
w51RK/ZhCnE+cZKjS58wvNM51fxkrtmm88XsC0wCi0kETeta8ThxNwyakJ/pQlML3RzxhGvW6tu5
oa6/2HK1VTFDotZXAAKZGFyTWlst/BEqPTtkBkB+m35HSpyzDaXFED7YEaiuLq1K+AlEELZZ5+UA
RyLsZvup6P5KCPcnvt4PhdzeP3IYFE1BwV7ueHvFv6O18nElqinuEB0Mz/FdED4PQoJPQlRqqWxv
y4P2Uw6lP7EtpOnephonQ1REXJnGYkYPjOJDctPyCxwoJIN9tNRmotcCwImmirl0mTT0mvtjH4lD
PcypPy3hb4fFrY9GcVOXeuiNRtb6Ypy7luz4HUjPkEUrXWnPYl3y9DGJ9WF0p/lPCOjqUIeMdlFr
/7KH/2VWm71ObOA7CLDFARUlnP0EqyWjInpIx+pYnrlts8Q8nAV286u/nfr94wBUAod8yQXW4Bty
8G44y9loOxDvYLOaFBcth5SNmiyDLEdj7bYXFQu2JJxyQhxTSOnVKeQ4z9j0oLFkFUOqcjhx7WPh
/do1n+hu6538YmNhaHOsH7racq9wTw0PuBb04tv0ZY78udV+UUl6qsO0cGLd4ThoOzYbdN0cJ4vr
I9o/B+qZg6nRYf+yYMmvby6R9/Yvu0K16NtISv6I8hb+bSzt09hP4FsoobyRnWjBIXP2OcUEXapa
m5eRnqNXVBU54CCILN60jKHAkja+YSlGxdkshreGSJO3v9hpyoIHkVCmIxhG0v3uAfhSySlMIAno
G6ymX4MVyt5IfzZUhOdGxabBeQybz12y3e+umttCxpzM8e9KADsQy3yTMGStSV3t2GGPjegMosB8
LYd3+d88Ti2qiHaYaBq3RR8I0GfYKOjjGuIyUzBi52f0r7z6921/ZGSBw52GafVbD9yv4ejFZaDF
dUpdKJkahT2RrGyZ6C7AGC8qo2e8GnyMOmz9R2vn/4L1Hbylqs2vIJid0S61/xJclPZ8caV9AK/c
WSPlvOtD50G00duB8r252FNviUOorkEqamkzugFmMV3Q9teDJ/95e+YZrIZ5m44coQil2H29wljC
W18A7nr0YpfiWUxZHSEkc1wQ84EtAzG1Su1ouqpB/pBuUVCZr2MJhsSAgma4a5kx1bVCIhr8zcT6
ntzh5iVTwwTxv3PZSENcnsQW7+jwhQn5ea1KaYzMrS2vCNbSC7ngb2MQk26qU/k7NnB+8kImmal1
CkpNyHEAcXqVQbln2dtqWKp7NyPMb8o0B/4cdulBYuIBIfcmL8y6ft/oMQHgQRh5IuXr8MRLIAxf
qW4RXPEBGPJiDLN54m28pyznc15h0Qavl3y2vwwzZE1oaOAon8VYT5vkTGvZKtM13SUqQfYcEg5r
TzvvopZYEHRHtNTN6jXmCtBZQWZgyjDZxyjBORS1KsgwtBjHnPtexq2/7XsOtX9WrjXCULuZ3Rzv
PkY8Xtb3cOAEv08w+zKF96D+OMsCSG508CyCXIT4bMFFisJPM9Nftozc6MTIkeuEtpPcPSOn6Br3
QF2vjmugPUrPW89jW2xKaC/4TY1iu3D//E5u2xMJ16VBT2r9NTmQlNqDogn9aq3IPi5WJsMmPHqM
nTHDXXpZifrSPOlA6ZPfd+J8dxhUIgunc0PRWQmWiPNQYy1GX9jlCPSKeSdpBA337FXkj50rS9d7
pq9fFIHDkjHvpyVehtmhvAaz/pX20OAJjgI4Lqw2dN0keazexh0ZVDsmWeLxHBBcXa2cRBU8vgkj
PnHbWFn7YWEE9w8MKG6svgieJfzFlmvx3bAGC+au4y2hRJuzy41EG2XqrJe/ZxO89eksxj/wXz3/
510kfs6AWDJoVabhHYUauMqW+DATzQi99AVt+2fp54nzBYT9OlEeOnqh/5c5THjbmCFAzSTYR9ET
VRqQW6vBDqhdre89agYJyJQmVD3IZmm4xKlDlzRd5UAkfpmQJTg+1vwvZpDlTkg/oxukAuirhthZ
9a63QrFuflssQB3ky2X1G8ABotSoXY1atdsrH9BD24icRcwdC091lnNkNRrodLokEgveOmtbvMgQ
tK7Vzi5mZcaLdETnPn4ckCfjSkqVe5cpQhFElBPOSde2zfHx7sOQdb+We3hrZhRYjhA8iL+Q88kz
dheMWJyHEh/8lHTRCFuZVOOcklvLhVUpqYOuDBPIpiQovkw1ISKhPWWzexwv/DHIZL7iYTEggP/7
CGjv69yPGOiOegIZNGuFZvsch9UhZ7sXKUE2wyuRfUrJ1Apcek+5k3qOk3gvlMzehIsVZ08Melj5
ONPZJSy2rBoDH6g4vjJbS6b8CcMBSUJf0Ssg2pUvTXinJu+0GIdNduBzF8e6KF0bm0SiIFj3/HF+
Y50N+0Qy9kJmj1o8ycWVshBAhKuT0xYyoQs70FHQ5eYyfWIL5AWNrK9z+KXf65pZ9bUY/DwnuVu2
eCJv7iyJbpZSccgUQ/53tXzU992nJPNqxRNlTZS9FO3DH++GKStSlQHlf2s5ritD+KvKhCeouV9r
cxbaw8MbZuG+KrB1w8KbGAWWrdL6p/MB6cxBnd3NVBgxDs7Gzi7DP8Hulwx/vH02+l6nAf4Y2WM5
V+/ebnAHcNy4xPcJ5NfUDpME+CHRuuUlu2hBWxbMV1JVsSqGpuZXEiaE45AWZaTEnpodn2R//hy8
8j7WD/sRO6ojzNP0BjMwy3hAGLmiZmixIW9bH15/sGrhAP8iIQ6MZ90S9ngNHRyUJo/bqpRFLW4e
cIlkgaXyMCjs/foup8K2H9tDDljmFxjpHypdc/KniidWu+5eBxP3gCGCHwuxg1NOGnRE5FEOnX0w
cWy1M18Tqj+kZTRRykd77/fFBt4bkmG6HbaXnwy2snt54AzDeUqQD2rxkK/r6JdilBNEmAKnFHxS
rS+Vpg4qcFWM39b89ivTroT7j+utDCPfg42e6ZBXZN55vF5pwdx5FgsEI7jHJqYyI4quffXIwQOd
uweNu5V+MXs7TuPNFV2eHMlhs8bO3ePIcMPrRLpwuJmJ2AvI0uxRZmKP3IpG2+GIixysGFd7f0wX
1mxDi4TvlwMC1Iiyy2HQNzNskaW9rDxvNTLhDi2Mxwc5aK/559g3K4QXBehaQMrTu+dUIoQWVIjN
MXT2LiV7l6Mc2kNUq7nF9clq8yKHVrcl87/k9pg/X5FOzDmOqnIgpIvutKQbecFcUT/GGDGerUwr
4grewUA2MbaCr7npmJGRMPYHoCnEicJSaBsvtwtB//7qaZFClUnRaCUpCru249FGj1tiIAmJTdva
i7Rf3fpFf2Blz0O82ox3zVxKZ8I6zdEj1iKqFCVp+JenhWtBrdKik5NraAn0iSrvGhdE+ymxnmqH
Ka0gaertnx0gXnEwuJIkI32Mry883SmQA5qFxHZlKGhPspaMRGlH9NbMswfR9604CnPKypZ/+E5+
tIaynSAvUlZ/MY8Abi6Cq004VcS1uxVR3ylBaMF+2UWKhyL5iYxAL8t0zhOazgEV40GD90JXDxAz
k/eRB2+16vf83KScQvcZmt3ncSATPh4I1uyudalG6kAQuONJroLqrdrY1Wklc57T6xmd1xcOPvc3
pi8bio7IdY6Cz3Nhq2rx05ZvXVlPg8wsFb1nJZx9J3hVWIJZuiM72l+PobKbmxgr+htXHGglZRR4
kUrgf77u5YjpKqBgMPcIepVwyoATLX61S7pKqV+qiEaKsAvZJWaLsiGVkSfu1GPCzhqL2cPhc9Zx
qjMzatX8eS/hIUFa5DC3+DskkkVi3Dya3hAjiaYCHkcXItKGxa+A01meJTkcO9C+k7jvuk5Ugrq1
2iT/fpkCd6Q+S7btkU57OIIO4CxVDU1LxieNGTD/oQvnRWMr1tOVJok414AxHG2hTCGxj22jD99k
h8jukFsoNITOplwCafUfHr4QYkqf+B/KGJZzjDjH+zYrJlZshDFzEHnQdcgj+nI5Mnm5wAogVFzP
EoE+JFJ42+64jxfBmAD6JndEQ4ZWKjsL0pmIzO07FdTgdVNoncRUjtXrZmQdaijVkCEmgAncoAl0
R+YdCnDTpNIIISIqriSc/ymHStQ/3BICD8lstSBIRorxjo9sLrqIhF226uV7CjyhdbU+XMTZ0sj/
ZPq4Z3qCpzscuSQ2mFlrcGv2yvR+XlpOKCVEbE5RXu2gA4Usv3ASrLHzw1pAYQRmvmQk/fu6q/0Z
l3J3jXOYL7BWn3lP8VXMjxPJ0qy2Rnx+WK2/JuxMAiiSy5CJOQPER8P1PLh4J5RohzSEmir/PKc9
JiRafCeBoUSx1aI/6SHOW03LVmWBpyo58ndvgHuCDkte8Z/zxDYrjIeAIO6ambjiHJIoKs1tJ09H
CjTswxAkUWnZrb3bXDRNaQyKeZE4DMnTrCRkEr4EdgPkJnyZRZaKdXwFW8G6tDr9X6Ojp8z0gYJo
fH1vk3OJwzDDEJ8ajAFo2FTND7BDGdDpjukPN9Sxb6OHrP1sJtor7M4DKbynE+kdhTngKeAl1kF1
YqqtY4mRwyPIpDx0vXcOyZ7ubru1HJncifVGhTVMIkHpKYb6o49veCioE+SwEfoyE7N0h1csf2e7
4tOl5HA7w3p34rvBagLRMR3pW8rkqy9659sxyWcXF+bJ9bhLUSfLUwc1W50L7nUFBujr+BGnFb7/
x6kzp08+SUaSoqoo/LE8Zcl34q6jku5JydNU6GDmsN1pJTKr6VvLZG7l1KLO5XXgg9WAe4SYNerY
KRM1krrhFP7+Z7n7DK63dQu1qVYjxbmLGpWCTx/lemJ3xak+D2zYcJsJfyBf7hMRbZKbddeffd+o
DfjsUjYeDCgUClM7VDXHkfFxxiu8VKo2uwL3mpZM9iLZid+grLB+msWDLznlmmY7aqQhGpe5CiFD
YU+Euey8jqfxD9cccMnajY2D0c2RBXxTURCytQecSG05cAgTkuLwAktJVb43IgKbjV1tL+atcgQ+
idyXaU5NW9tCOyjJ0je1feHE6WlZbcK3d4v04pQ3U9lyUDvoa90FJAuTdfNVYlL9OO1ZGbvvrSbz
uw0sh/mpA3cqpO6fvU/nx+Va2WrnjmL7lTu9PBMmSxkj6fXBs9heuEmS4uGoZO3F6BrB589kFklC
Gxzd3+yAVqIREqrXlEJYFmn0WUZDv90ZNtRWrXEauHhfbHsilZ7JEJyVRVseXUV8kqShx2tn3igU
9RjU+V+94an1XfYAINGBZGMXaBZpb0Oj1IK6q17XMnNayXRGR1yKHoAixskaMvHOCyYN1hRSZFXv
xQxA6s4MJ5YltuSJkPygoZjXFw7cCISCJcl/eAVG3uB6GRjGumdEelrNTdwwkVym166WS1jMJBPr
bDEBzgcZUZwMsm3rg9BzCEhbpK+ni+J2cZ3mSHn4eJZ7VA4NYa+ufKRUnc6CSWFUkhNuE8C02Jqt
Eu1nhiCtc6Q+h5bwl8mYnYixdTHVp6oT5iM39isuMlssTpbkqHN1UZ+El1DwBB/VMlHjD6nA3qwb
bsNUrqUJuB4Nv7mRUs1dinsQLyWJMFJaXlgBiabsMPqnyR8QI+Afa/gx8pPRCBBYPOf9khZlDQRa
9hT1JzlO4y8Hp9kLSH4Vt7EBC3tKcg+ms/05hWt9XG4Sj7+LFCBBJWUXsHRtFTfhKAahaMeJpTIK
B5oS68j4C0wUYzLhyM3itoeUtteWdXfUdMxmMhIAjfkC0X/fXEn3rqqG9kdtG3uhFGmDtFK9R+SJ
5TlYhDIwbjt+bjwmAkZf7cqqwt6xuUANMBSAhUt3fhRYvdxxOalYwJ7CuQlzisOSH4UJLEOhA7wH
jVwr2TWo42cCv+5nQeHlzjaMEb0IP4buv9Ln7P4mhKnbdO3M68GbLS5LgOEXJ4wWvpTML1koTD/3
wyb/uOuLsT2TUWw+IssufG6guOloIsR4D4EukUessIsLl3ujPMnBZogi5x4Au6YTCz88F/5bnGDn
DSwGoKoPgXZYkTj94T+kHL1+ZO7VHmEZ7YxsQL7V/iJmtT9TLbqH8BisExG2SH7tk0WS1fMXOu/5
N2Ks5hy3HDasSInb/fdr2YYBG47ssgEerEgbkaMOC7hPuHoaGVf8ih5e7++zjBe+XcMm7U678h6v
QkxPi1oZGrQ0Opo9SFfEGdtORVj04jzfvpiJYkmZM5CVdU4fKW8tNzDgU19gB6O/S9trsZrMKZuJ
6ExvyqrWdPrh+NmIYtP6iFazCv36YSr0r4IQtyHzWwEZbH5+b/mmRU4pPoN/Z/yWElTCDDUJtQGx
1dkHVCg5i/94xzdKM89BnMPBaBCRCCP4LDHgcVfXJg+U/mTGI4Pdj8XOlubqx1gsWObxvo0lP+bT
Dyp37sbCZCKMiKUm9tuJB0eb0VWTBLiFBWtZQlq+3EmhoAnpkArSzG2TN16QZSn8dGbkXqS+KQ5N
4M//q1KBstsIoYpvN3KEENKeY04+oWY9tTLdDZan+Ul3aUNCrHMJ/Dd6k1gRbonw2d+d6n3t18XO
wWxD2iP2ZURM+YhhQQWDJu4GjjWUEabreFHWc0iIpzmBP43pSnHxn9Qb5JXf3LALx3CjSgBlw2Aw
7VqrEh0k8NKRT/Gb5I1ThcqEIrEV2mxg6JRMGfuwKqEQPjae8b9beziVEsMNJIa7TczUu3DloXyJ
pfwa50rvR5VfZDvQum8jpjbrlzb8Gm7Aq1H3b2Ap8rk2sEs65gbLQTbqQQLJJ9QiHHrZocNMWD8i
1/6PyuwSxj2Eenq4YkZDKsLFIUytndGfYgoTWk7i5jL39ssbiIhTnULfV8uI6Tstr2Szxsm9tDHa
5AG3UrDGRHJmbbAyi+tcr2Fb4isXFYHDIFMG+Bh1ymIjtulIvfwUPUWXN1t5VSbkw/4bNuaGj90W
YFmD4M2jdR4TQsQLmR2hgS2AhhqsuS2mmBqLw/lLp+K4xnF4KY62r8RUsvIHnIsGWsZ/+JYx+hOB
Aekia9Tl35BCIFw9w7eJRChYwLmfHsImAKgvOitsgv9f+iMjciTTlKScgfYD787yqy2A0XmM4izJ
DPYcv8s8OJAZQXTzjy3Nl1csKGyG42NuX825TUREy3Lx5nXtOc0Aliy3pCVX6mN6Y3vhnKPppfhG
IW5t1hdHg4/v+3n+uuamAV52vBuMkxg4Hqu+w1r4IP/3NWpLqyq6/VI+nfwI434CaldtDAHqubo0
PaJh96+txxbb6Qsq0K66MI7lKjjLq5mDHPmk3ZoVaf2Ktic8A66s2FQATOk7jBBaY5BYvputazL+
c+cYINou7ulZRYePLXukcL8yB2zuWEBCrPgFDhls5SOtzL/I/mTza4sLnzZk+NH/i9Qg/2p5rV/P
sb+wD071pU+1rotmsxlAj/ja1fz2sWOIn33A24K/kqCvZ9W4QTQSiMiS5dbdGykYfrCMms5txSaY
u7R2iKXH/HbpAZp80NFIbCkgHiiWrdRu+ENmmbwztGXtnxWQll5qc1/Ee8jIyfGftXhE3dnlZK80
V6PlYe+daIo/FPi3GjW6Qhn1XX7ol9/1sY0AAOcDyow/mmc4eEw35l6b35iS4t7U4J581L33NlPX
hzfljVuI/MgU6E8FQ/i8WCaLzGLjK1j90yKmKNhvZod/gTGzQvQtPp+e5BtE1yLs+qVN6EjxE+uC
CfmhCOi3i3qrjkOn/nju/OdznaEk9g/BKQLDNfqKytnbdrgVh3U3BIT1uFJoBtBqIsWJi/lBIjox
U3LVoJZda2yWiMvbNF6UN2Q5rwSF50Xsve0PWe9C1WorhhjX2y0q3/VYx/Kzg5MTHrSsMVTnofDe
MroMAvjDysB+xUOMbzdfZLOU07xRDCunpS30RyhISeW56I5MObNsg3VI/6weAtE4TtF4S0LLN1S2
iIRNouXMaRrveZHP52FEVhLSV9mJp46Qa0EEzs3PlcUM1gr6AeJdOQoY/21lmcQOEISG2SuYS17T
qqZcTqsT53GqoS33KRTJFZQj0JyZGvAm7hBpuS3GqvzneB4c0JCbO6ftVQLExhFNafzNZ+jVcqn1
XkdWwjpps90COkKvEKUn7VnTOrONkSZ451m5hhVn76GNSgXNyIxK7PX+FLAz0zPbnqcjOsqFLbdl
9SbHtYNHehELS6OxYTu2BWLSMRgJ3gMduqDUKrYAy4U3htGBgMd/km5GdVRw2wmaHn5LOJI4dexe
1lo9q7qxpEd4jp+wa/ScDbMm+mCiyY8YMt2VqEjlG8mrCGnaus4a8lExIJSfWokm4nNS85KArZ5Y
qRW1/LbSRiA2BlAErhAUIosZtKhICgPuXgprLB6P1vVjDPKj9w95qKtRDEND9zaqkVYVU1pcWhhD
sDUk6O2mHiZe4mJByWc17CvKMI9CxgW6kkzJnTMgMomSJCi/loiX2TbFyeqN7uddhgg/gxYXZwe9
JI5W/Ibo1UCn8fDNw6XvSsSMkqjCBPM91tNKyVm9kxNwhhPIpdnq7EfGd/D7ltm7YCToF6wUUo4Q
5TWemPMtXnPvwFIcjnlaRXJKohCkuJDRi3AZOUQz63MUoVk8/Rx+5BCV0xPLSIdyku+Dp6IFfMv0
wvCDGJ5hCTuOAc/GbBHDxWBPl34jHk1BiNunWpt2EHzI7RXFRs3L0k2mS7QsJevtvceVB4MUKYxV
gHLSXQYrGfP2i+VApP8Yl/5zVdHfUvkrO1DJgFk6VQX8IsK3OEbyWmtqLBDQyUdB9A9dgDIlJNnr
rakrSrWrWtk24VF0nFKw+RiPyQAf+4NbajBaZTEnizLfjJyP3xTdiafByezaX2cAYbhiOalh7peN
tm363OshEDUD8Aa9kPWwYbFMnVZqxcJKu4w1l6JufdxywvdyKJ81tR3UVWUCIPeTmI0EnLiTkYTL
c8DAvneIIRoAGCK9Sbut+6gqRrfGlHcOl4SwYJXekqgSsUjRgtUVcbsdWQkaf9nrx8VIai8v2fCX
I7rtgpmAqpyzqc0U+pF+OF/3HQI+pg1lAXuYRFZYSDSXA++7qDAuoVmeYCJclEWeUMyZX1H6xf1x
898/5keAKuqWnLIxPI+A2me4x2+6a/EhTwEL6ifqeV/AoCmA5SFodXfol+7CMxnF1Qx6ldRUAGUj
qahrViLeQrUu5bGed5o2/YJ98IdZ4LxFevvf8pbBxSjKXiZXU1UIy4AmcHLCFi3Fx/EHzBQSvh4R
ohhz72b8TNn/PexUf+lVL6JeNmLewk6h6wkTfN102ygoR6Stldibv58KB2rlnhAvLNZlQwCzMnyX
FEU6fz5N4OU3ETl2tUmkm7raizocXy50lPL6sFN3+QswoK1Gd6yZFLuE7wbsS/wsOnQ3p1rQK0kw
hiLYSbTKip89QbEw2WWz9m/0phQIEG0FjlI7m0LbfCjonaUzP2dOu60kBmsPpPl7AeVhDPMEVpyH
akpEGREyJuIS8/jb+YxLTdrBWSsg0kOAOyW3WVjN+3h5lC2X+FfkMjGqtZc+e1P7bVgArTSAAqjt
2L1U/lgOt4LqA4P079IlKMhcHF6Mx5Zf9Slb/UVBZT2B17FcxG+0lY3W6/2faa/zFTmXpSgLucYd
CIcOI0zU46dJ0GybTLjjYLBG8QgW+G3vsW1kXemfDlKCuJzJWymAq2OwRdI7PEjrdBU/a47Sssr4
WQ91Lscxk/1DYNxqZIkZ/NNna9EYqobmhmrQPTfBDOymHRJpGqCTnlBf/ptkQGAP7sG/jFCsJbmh
eeHVar+hhx/yjKrnPmXbl6EzVeW+Agl9yvZ1Z/vrCMefrpwLwnYRdm5D80IrSX8YXEVOjiV2C8m/
/0QbfDZ1Tlfw5IGqiY+kCB/PhtrGrRmSvOi1SGBz6Z79+eh4DPcQaz2SgjzZ9gL326pSIyoNOepB
KqHQGKZGbDdEn2Ip5ylJfYdkH6uOSIGRm3eJNkvUBQRFrUYKNP3NbBLTG7Zr1SBUIA7q9C/sI7xS
2WMx0PdajjwX0WXZpHwTqS6YMOuD8WR+nZktYrcVYMkd7Cl4t50KozM3J2q8V/lJ4aFGNAQYLZSh
3vUVBi4KsFaflR633pn8hOxUWil0dW4QjL3j3W6V34N0oExU54mydyNesO5ibCQVegMgJVhuiLkL
Zn/FTVoHWRhW48bv7fbaXU380opxWAsLZ2WT5S2E4tqpwueTlTJg+5pSakQ8M03+AW/DdvpO0AyK
SKp0WZ6yORNMOdIGDOJZ3LfLUz2Vw8jLrtBsRaSSE+OX0ks4fXNtXME6sF/JTlUz3RjFMGnuhPYA
V1RVRVtfgRn9oQWfN/04LpGTZluMFzw9BZw5HWcFBuS4Yi2t04P7dacThXjQkrdSvnIW/76vVEVN
gy9UonyF6oejupIY1C4URcieDzLBFHFansQ39rTIizM8OaErAjw8yV3K6bTN9M/5uyOwcZs0wQTL
Fn5NlOkd2HKA/1NNDX1GFmn6QERtMUCxuYd9tPwUl3P6VRqP9CiTqC1XV4ITeJaM8KjoyzLathmX
AluKO/0sWpnQ6wp+3p9UKP8amUMffP9TBOE9lxj1ZM4eow6ZjXx+FEi9BJH6vFpgMzE/8ZgtD2nv
GGc4iB3XGDgWYRl7au3FZHbYf1zF7Nr3VCxWAfYEGHnmwxn59d3eLiiQGcpImwptCQVRZYMxXZMa
VhtQmFT477j2X9CxKt9vctzW5hu50bly6QnNKzPldFodr6W5LB8hGc7xi1FitNyrZiBYcZt+S+L1
t9TiMFjakNCqg7CL4IoPKIsZyD1QCuzvTwKC+PUP2Tda80pYyEi+HqPCJc9W/fUpsIO4MLHm66nE
eZad1rDWJTR/OeIfA+jdPGMmwE+qmbTkSVMuCmW8jTPjrxWq/VHaEnzp7nk8+wpZeicSioBNCWR8
4mwQpLlenR9dl3S9OS+BNsuouIrX2IwXK0YugPjMlgJehUHgDxliZIngeK8nlbwf3BXdTghgtaSp
AFMQdY7O1QXXK6LHwSuWCW9fDYR2jCjBsUlZUa0k4H10jpShgjwvnQvwO8OWEizfvJTTuuT27osb
/QndkvLm7725tT7YXhbLgt+6zsjdeK9LVsGUDmTre8aV6590L54WY2F/2FcC7AJedN1gMv06p8o6
pT/f1LgPtfQ40gbkG+cEe67ymPDpH+p/YBh5m7cqYZ8y1RIJh3Rewrh9XxYobAsVAsdXFnY9yuUh
5LJEIls0hSJODNAyhBDXfKrw461ev97uMfnnI8JxCll3Vng/x4SQbqV6fEatsWIHCi50CexkOdaK
hjKihY6c2iOG9/uoJsrDrgUwgF/Kq3r6pJl3EpRURXR3nxWKMeGmWKWbxe9NL9wfgypusoKjuvbx
PiVnnELy5DXQqqRgUFm8IlqlvKyr3jx8fXpztYhERhDXGiqIVVpdeYZ94AF/xnblqrG2SUNNF9Xg
xaYbXJ5WiyEbMNS1zT88/hoSd9CORgRlHXe1bQgs55AXdE/YJL7qrGDI8/ihyw6kyfzgW7w6eFjM
64GTl0IGzMNGhNvzwZxbsZf4TXPhllAfsypum3kDTME5dd1ybxEPQ3sWDRzwHkaNRy48xdFN3Ocr
sSckAoybyFoRGjElc0+Jr6Y4qpuosbsP57ufKfmeRY+7u8ppECQu0E7zQk7LliDtph10BisiBtuQ
RIHp3jEhyTpZPWUiUvNCLnouaOUITVg+cynQ8QvFg/AHgizswnN1Ll5z92y+bY5rfA2IQMQ86lTJ
cWKouPP03d3vd1RGDxjslz2PmByvjewRs/3vI1uXUkK7gLH6IPGptv3g84S05aWGJNPb7lvxMZm3
b9GCoWXBsOE2VX7J+L5jiXOq+irZI3SPTF8APF5RMJyR58P1g/MZQqRiMFlFnN4NBaXNWoDO8G98
pYEpRlCIup5PC9Rw4ghPyQ2gLV1TXSEWH0nx17lYcSkbQyiIHoG5W1vEniOi1nPdM/O1gvsFsb7X
j9/hUx0m1zjvOdbmuI7dKRMEXoBk5tvsq3xSopL6Kv91haqISqMnHWSsUh6nBL8H1dJNioySmJG4
NNZAAM0eh9OE70smHekKtYr8WfLr0S6OpGQLnbzsLtGP95fqb/WeI5dnbQzcW0QK41BxbEWijr1g
9dQ1ESPtgE+dpgTMAjMql1/B7cffquzhq1MzR7w+FTmqvA7XR+6mTHJIfUS5y3mya9XVJhxKzWGV
ens6jiCfciipI2zSBemHV0W8iWitHI4CwV3OQFzbzPMssi40p+7xffYAeQIz1mLe9OjPjkn4Qh84
FnYTc3iP3BTmjpBFu0utpypN6snd1FwoMoCkVtCxTfPU0afcq30yiEVDchm93IG221hXm9s1JFcW
4tOMO7Jlf2qtzXq5SX0k4HuJS3I+SyuT8bVekHiWE2jtTv3tso7t+Zu2MBsnKkf8baeyN2Hstj/w
8VxbctCj6yTnYRfoOO6Sf7Hat1H1cyoT2RG2AZpamLsykTdHFDDHHgCFGi7dLD+oib9jHX8C/u+R
2EJHAY1zrjx+bvHvSdByAAB5iZS9oyoTCmNbX/SjX4TmgOeVvB8/XnAk7xcsag+F+99uje61g/vx
dxEzEYQQkHH1Z8oedKySHUju9H0IM9MusiFyUtN+yF0OADrJ9cBrzDTzu7Ug7wnU2y5+rJI8kCXh
beOz3TntCpPdQZDlsGj+dO8s0mFPQG6VXbd2cHCS9nH2wdZgXAzC6mUuQOiUTw6YxAehNjSc54Mb
CB7RJq48BqKCT3nizZKtW6NdoSU0C6jqcD2yWIPWRVBvoiMc41VuhqsdBx5wV2KI8nVPqXOJ5J9L
ejyS0JyuKiULQhxTay0eyiMylKqXY9huRTgU4BUy7AigXPj2VvlVAljhHaA1s2VJJfELUA7CtT/n
3KJ230SajP+m3OG8WHhj2vOJDpUeRUYZ0eelKQLrTuyLN3RGx7G+gqh/NsEdENXZpbzMRioKiGcU
5pXmQ6OygIXvgFb/vDZfw/ZI0ab6SFnLwMHKtJ1fSwg7CqTajqdKfRgPiak73yQ7MHKTJvDhYojZ
5FjZdMsAgI7hnTxoDBzmZA9/5Z9mKcZRKQ6/RYlViKfMSfJ6jL1u3XGqzUcuoL4ZkqiMm1g6TtMy
iDPxzB2CSOAGQgFr2hX8dDGp+4pg2ZAlSD3b7mGUFMDbIYrxwnoTTyYbuQh3p3wE4Fsx/ZENxiZY
CyuppFJfQ1rcFV8Zg4E/BFgsGbGhfxSzHYlQEhgHBngB7UOwCKqvfgBFSUKe9b2TE6I1xvptw3lA
cAYwD4JFPbyxIWLMkwiyeaKBXhkUsDKiM7f7qNzL00dtOj3IJ10BjbIMWKjNDgao8eo5lFO0X8HT
++RCAyGdu40wGHmKtTcgPi3gw2LzO0VDMU0AefSe9A6WeTc07zlZcGi0EQMpGr5LseH/tT0utY0M
Y07pfkV5G+c+ylnr2uBJQgqzgwcc2+o6h1GFHalRF993UsdZ3yFpHuyqeeBx8QTNTlk4QaUqbQAK
3FNRwebtli78YffVKzhcUXb+5te4UUuCO1WKs2QHJUFeoz+nEWT1z8pHc7zhM7GWF5i4C36zIkT/
8ZdVKdyKqpHNIW/RwhTKbj0Dr8OGz/5czdnkTSkW0sDh93Cd4V8ccKOVV5eLH0C8fanXraAa5502
xj9P7n6zO1x4hXt07F9EwM30JOSHlfFbwdYX37iUYoUBHIfR+pSdRF2eKgRVkPoGTDvjZ2DgeBzL
N8zaE+i65seE1A3qzuwz588A/MzXhQOEv3wdoILvQHnvzOanphyqiC6JGzKmP2b0grdCF+1chjIV
DPSSUoslVG2L9XB/idvfNevBaqkRu9Rfoe/RsLXiu8reKCCnX4iZxBh+mHgV6bOIpbwCccZJbG+j
4DgtPxYX3QjP1IZ3/eHov4TPbGSFI5SvLhq2ok0sZG/ZZqa2Bogacewanvesv+CyJno2bsx9eolO
FOYiceqTA4WRUGBbr5HdhK5cY6889QYQWR7RZtfWf+w5tTz4FiWd40XQM1TbRIu3+TIkRP3BH4xW
HBzh5v4nV/9MmYdTrm29AoymseTYEbhvZbfoyyjkPpWZbiAnaGJz9r6BJh3Ecc+5AOXNpJbQul7C
SIfRD2mEbdHX0rfq2onrlWZImHHwkbGwQGXxlKy6IEAC4hSpT8kkzn/YitaURJ7rp+J0QowWyFSD
0rwP0d95PgyHS9oSL9M5HfLiQ9wL+Ihj/88rXazwKF+HpgwGZsMSfHRDKg/zubd4b6Ye9+SCDaPG
Bu350znwP6wzpTpQrOv0CI8shWXpxYOOzBpV9WPOeZGILwKf7REJhm1W0QeUFm9pu2PI86CVkior
Oi3agdhrRHXkWlcn5mhF5cClUfqjmPjeCUJ5PIHetsjKI8FTJik7SpEAU/xRPJxK1LPCrfxof8Vt
YevBbfYv07cbJsOWp9I9ZC/w3IuBaHYzUI3a4pGnvZAylmMkNzweZKYA6eIa3l3IBSBJa8/bsLLM
RAfX4e/5sSCrTqcsT1IK6xzDfrLytpp+eSmd8uzOJ7aQmfFnMtNt5TUFTLx8dZ6BlBe7fMPo4wVx
uxJssY5p7GqHwwM1zFxsj/alj8570jid9lOXaVO9owb/WUcOXqrWOMD2mAo/VNX7oP/ykxmmF+qC
ielvtiSLHktIQnxmbLOBq64a6A4n1qiNyh986dX2p2ltaWPtqdj5vwLxN4oqmvgjYPnPyEJYXnlD
J95n+LgY4QP0pPgWZ/NC655MyjH19o4COf2YdYdWzdpAivlOlxqAQWHabypWMsd7g+dbbzFFE8iv
pAaF91odHDao/s7xBI4ao2m6Nv5u6v9XO2uit0Wo7xsPH08EpOyuS8AhT1L/bHquIpIdWE5fjOMO
T4WjI3S09NLIokzvPq1dwjiPyV0JYHvHh9Yc/L5tO8huQK/xetGe4gQeIfxn/AbyLAgass6i1QE0
Q2oYcdAAAwrsc7RMy8daEkR4rCfBh1hH1f1dDWvKIwygOZCJxFymzXRYB6sVBLaK833Sy9gjHXB4
nBNGA9N/B5UUnhcQIGBCQe1K9oEMgfBBg4FBxBlcnWJl9CE8gwflsOqWGWlB5bFjiukhRBT0iM7y
MhTl9Ju+cV0fVjwQw/W2qVDquzpgrbW08A/oRQ6kw6WUAeqNM29CXF77GN8v7BCfW/me/ZoP9M59
OBA79+oMvdV8kjJtDp6GKR2MqQkzSBHXngEHo9sgp3M+Ci5yZI3QZAQBvdJe3eHqxVkn0t5SjnbN
wzywtYD0aJ1CAb9OABF+aJx20/qMYUkISp3xwYCBtZJpQnuUzguwRtP08hZxpg3Fo6LUJJN+KVsh
dc49Lf9GDJuBEnuHhqIm67eWGCFU507rXeaSgjAiY9+GAcuplJUlimU8WGl73YzBm9DEKay+xlag
qNeKluuy9nFBi7oQb1GnVvMnmRMxhub+Ml7wm2q5lWPCueX7VtZ9MlemfwSKPO4gmz46Rf145N5X
8YfpXEZCpNeMgupLggHO6a8O+1bVzujBRDJ+8PrHL2v//u0WHgXbOEd2wFKxv7BKCJ5t71HEO8NJ
xZp8jWTvadIzJwP//LRbSnihfIJgpE5kK3eqZ4PziTmdpVqbJh0hgXxzru6bgwdsSoWoLRWDjHvC
gXm5MBLKLTlLJ5Jph+xaEr4DHijCIjlo/SW7LPNfz0pLnA33W0UtREFHYxhmPqGeOY4TGxaeOyh2
eLD1mMA+5BgqaWcxWu5adDKhGXfb/9hdtiZdiAUkIH7PFhhaCYDt0j4oKpH10rMxUEi11obtU2C7
T5VZ8AWg3tZ9AUeDz5wx0lkYYISWrym3rwj+b8ED7BIu9gecGnmc4/ULd/Y5xSPB43Uzh/4xsGlS
kt3oKc/Svx6bCS5biOS08/TJ1gdkSbvB6nCDlCGdEmeblfl8emleP8D+4cqhJJH5SXQogXz41sPb
HsljJ7cpgTfOGMo2KhNhX6cQRmoeY1x6iLxnb+PVVkeVS4TSZm5vPysWMRsdK9VyXT+yr1Yk4tlv
YTAHPeDhNV/5C1PG647WJ3fWv4Yef0nN1LfXXDWOTsmbjex07SNpDQOnr73JMb/PX+cFZvJ7No7b
JmEadQwiBmlNUh/viHSIf3Y/Zr8yh/4spVQERbCN0dPZ/BbNvb/z9PIe6f1isa02/pDGXU2aqhot
PTDgQIr6qYe8vgBK2ZI1f9aP3EBNewlWoOH4QuKb8dsicO9wnqvr+fhvvgQAH0PFBrzCutwp929r
DE6r9eJy+3GDnjYgqqF2B3crw8GBV00ue2zpnKwtJhNLWN0xTTysjj8uT3iSVFc4kSj1GqMxBN/t
bLhuZhfZVcWrcbWLPsijUIsL55gOZ9EyIlXtba/i1VM+HqJfqJMIda9E0RhSBueEg4KaLD80Oz40
CsTQZq1GciSnkwlSPgVfc0xmBPFypSjbR/IikqYYpD5YRpnzDNhS34mQJM2QSnRM3oh6s/sAL/lo
ehO0RsfURzLFwtfCFlBAgzC0p0lEhGrc/dNiCKQVw+erttIXLjKMfqg3EpkeMZ6NlgZ26KJ3XmlY
sIK4wkQY3Dx0pBWxnbgN1HkYQ9yOnLGr2lHpP8l3ibWBNPV3wahA5xpI3tkue/v5/dq/0YFlUym4
oZGsMa8gvAWdifLAgs8DlOVoOwkCti0k96fiVLastz0KKkH/Uw1xr+FSnM8RqbEMDy/z065BCcUn
j1VLhawaFIgV4Vy4ovr2wbJdy1omTV6R52n34xuHeuqCo3YNQX41YfrgXK71BxkibipsPPV9PKbH
s9MACi6PKAprI3780MJaJYp7wyJQamVtP+RqaKzyRjINxAx5yi5HCJHBt1KYxUy5vSxIrbWd4vcF
Lqf8/JmMqdnk6t/+VYFqcNfeeql3aktZQSfElm1PRef7sJE3/T9c3fGfUHyxNbAez6qvFSDGISCT
xCbaZcmy4Hnbq6deUHVmD01twnKChU2sYww3R3RsQo82LGiopSfNd/TdqkS0gCiC08NoKKPW9pZl
ODQnl1APr9goI3tlTuWGOA6166birfBIqmAQYeAE8mpg79UxwGKGLs4CzLG6J6l6dF5N13l/MgVl
jyu8+KTCT4IH0DsT87lM8ZQ9kiSTG9WOcjForTNViYg53qWbPcRRMoOvjqasN6iUXietcc+3J9iO
b9+lDGCWeZfuv/KU8dW80kcsKqr8p+kBr3X404vGKHLAYRaXqJ/KZrA7aKnY+zsfy0FmgMBhHj3D
PFsj4qW71O0dTKXRNKOVwsChNWNhxgUOhjrNLKD+POGM825qoIgqcuBoX2wRVm/p/aVJWypPqLLp
ENJN2ntmgkD8pS1jDcQoXJFp6ctlguV4lqZknqSbj3CUMWz/2pRqUxzBvgZayVn8YTCR0JXhkxGN
5t2dGM2+GAYlZrwP3+fqSinjw5wzJNNWwH5w5loIHwY11MMTDLA42JhQf1QdZAzB++k6h11DCO8I
/GtA8BEGjxCAEFzn5ZFa4UBcS3cHIpqzif4k5idq8588gE/I39bcfKGpwhrKuar9Q7/TIR+JjUwX
cEJ9APiMzD4lrk85eDVQG+cU4p6IIztzo/Kr36xcf9tCUSiq6HIdnF41iMioekzSrdQqL5MAICiV
aalvpKBzJrGrRj4qFfViveFN5SgNaCNfyuMhbOoy+3gR+TYgu0T8i2ZjdT57NuuRm0mJ97QDjODv
ZZNKLVjO5koVDpftZUvoGzkzynoTUEimGb8C0jQZ0ay9PWC3qHVS9tvFP0CmEelOigm5wL/1cApz
lDEH/HdJYvzSzdknW+X8JB5nmUQMK1uTgZ1tiORnH5HOEOQIzRFg8L0S3X/vNzjPgsN44F5ZxQ0K
kN2jXytTX3lBKWNuhgbp1Bez1WVEmVMvmFwiEQlrKfkYnJ3OpuGwyuSf27x+WYL8oXMltuI/fIHU
b++tUIrHGZIYnfRK3ctFFsE4+aWi76PjAIMubni8mrrbsb0Xa+RSGqAJyLEAy8wIqwM+x/HQOULw
oQcmFYuVF7QVL6+IEaBO1irLqALIrXLzdfZIA+9hyF0ag55ZXXVHjpowgDpcUm7Q5yJzH6HsbFzD
IefgrMIA3TWcV/YodORe/TZVJ4chCDwsyrszIWimV4435V0eNsS5FsU0SWKLKP3p5eCuI6cne5XC
vbVgRvR5mboK+cgMFerHb6xVboYwh90lNhgYW16/u2hdeb9qfXdMHUGWoE65KrEB1HC6jZk1zf8A
FroxzwO+/DrRT2g7c092fIzUmOR9JSaghPyVJyauzzreFrWIApJpZhbtB2G4BB4/UyekG9cIdVtX
ZlFw/0PeXij0OMQaDmyJktmaworpSIXQUqhi9dvc/kkELezqnUc9XiNkmPtWGndqH224C0jIHqVF
Bo519rVyO5WCy9v42Hc5xCSUl/ovkKV0gsgACp6R2Kcd/4efdw4CxYfDEWYf7FTRlP4iuMcQ3Jke
3SsaDpKSniCaoTnWxD7u63TKxPtipVMTrmHVXAkO8qm8e8URNCBj1ixM+LfEZYcmXZ9isqUwkUok
q5hkg3o1tBCB9WsodyMnTTBd1mQgS2o7VAzrg+jYoeD9eIgRmF54sLcYWlyrZdZ+5KDMe0mIqe90
dJ8C1xb9WpLzHNZhtaVO8k5rGkJll/iTfVhc1aE38SSfYY3GtQlRdXy/IijMSQ+B1SyoojGZMheq
QdkN57HZgtrX3vjaPH8nMbjMHvdTiQDUlrzeXPy/M3BiIzF7VeXX4GtHDy+mnR0yN+f4JyV8xxf3
WNIevmNs8mUgdPfb3IwlnjatiKrTiy7WCfG8OIDPCZEvT+K6hQFmfZHPziGyZgA2Svm9uC/GkqaE
c1oHVu/kckM1KaB4n3ajnsK9M1D2kbfiGGBFGhbvkhQ1sAauMN22Ha75pehUStfPxUbEbwvRVmu4
ZjwW7xHMOAqlADbutI4mOq8DXUrY6ywTpZgps+XIW8hpbzsoqUyDxU7OmZ3MhDQe1eJIl8/ODhrt
gEWFb1fRe+6gR+cvdYHbc3OJ13T7ZsolVicJuxVCXgo9vIPqlSP3QtfkbXvy7qhG+GpSeItywFfG
p/+h++A4E2NdEgJvhFOVkdixRYll3r93XJRW/Z9X+OrFyKUGxnF7qFQMS+8LmfoX05FGOc4lr0VW
tGv+FwI55UZ6/aCVbuyty6Mvlm4Msc8wkGRslqK65YwCdnwRdIdJQD1upB+z4WwFjOYDTmODS45O
2AqxYQtqvjdQ/en6C5d0aEW4ybSgo6JasPOKXcSzR7whM9WetSEBVq4Pmp5G8X8knrTQNvtK9V/n
wJYO0cIVqNMGVRIiKOYe0rpccSNc3XBJmMKOzQpP3ackByqDJkVQ/MaaZSRuq4FNATOKDcFrNPDE
lFODZoRurs4UXnEc65BSqafglCGIhz/1BHzsX+TCODkk2cNkxhjZnTy8wLXOi43TwcOe0qBxX3+Y
PwDw9uQjSKCuTtyYSRafyF91lJiMml2iE/ol/wYcdajCcKLStCdLsF/0lB88whDOoSFhe6ei9idp
REa672Qu8CYC9zXzzo+TS5XJWZiKW6a2ZVpQkf1lzGYnqH06jrDPehXrFfXXRUylcapLM7W8+DiT
VprMnN2oP7cap+Ky1zKKZ3jYpWIG/myAKdlpKkI8oPhUEIWVoanhu1Wgfj78Ueh8dQXZfUjfGos9
Wq9YfuLO5GwCKadNbvi5xDSmBJkqOlmIrcNWobsISzWGJc8tOzzgBpeP18UsKY7thRmUUGF+vuVU
c1sDr/Pm0iReOlT+YEKvHlBFJBq48KJStNUMCVFjMJ6UnYiu/bKtGqDWnEi6UuhAg3pAaejMW6Yb
XstxkD+dJE/XeB4cURB0kc/eTaFD4tMZSKTmZYkAaFHJ+3YDHsKx4XCik13i9LdWz1BNOFqM3noi
2rq1Gm8Sy0OkfEwKwPK145NoaL8YVz/1bueg8+73JfzMUKo/ypn+UqEMuFjxbzeDFcUsdQgDaf6g
ijqeT9W4dNIO4BpXjhI452jAgRe1Nt81pTE7J0i9Z0KvnJ3wAk1vu+5RuX6BAsIlxI7so3+DyjIl
0Y9nZ4Jl50ffJwsp4G7BvtI8WTCMDyUq+9Ok7v7w38X3EuaM6DVPQT2pEqo89vb6DOK+Pl8N9uQ1
/iLM6Zd1Bxrz4Po2WRj0GCL8jYPqIpx30xIQKZZTbZaipWZaDM5GLsfvUUY/IYBi/ST6kq1l9NvK
bdxwVe+NZSmf7VkT92/Y5xmDzxDgvPdcKXljaHeqG5NajmCNcyyKni6apYUiVR/j3W3sWtckzBCP
NtZZ/hbT49IbC+Z496cRJjhnirJ0sGuZ794rxG5+Q3dHPL5jLiV8oWNHDPShByLhJbAR956gEFB3
0qZjOFN+wzy4LeeU9STq/H5tlae6WWigzmxi8uZjrs2SkZhUPKZ6tGRtc4AZ680/7iZeeIO5vTvh
Y2ZUEFnT0RuznkgNYldJoKGdQNRBv/41ZawB88i2nCRn9pLLdqLy7L77vWI+6K8zDt8sNiovm7EO
Y7zlgUk6eJVJW6u1v/ePJewrin9P8RJX99DRABkSBRFTh85cpbZvr42bT1C0AxOUYyGXp5lDNCud
MFjcdmOjnSAOoFTNHC3S/rnBcqki4KVQSnaJAanG5wg46ayalPNYCmPWCW2yFFmZ7vFo0cCzIEp9
PCaB2TMMm39sSxPIG0zqlCVmO9/k760Db6w9dIrd+EVW2/QzrXZ4bjPfh/NpBIZuNZVKUrE9jcI9
+m4Cc19LUEeqXKAAM0QDhFwCvsS0GLwCTH5feH6RKut8mfL7jZopPzIuetAiXb/4xsJa1R+iQOpS
FZuEy0xynoYwLxLB9l/mcaG4+JbiobJNU3sSrbf+9NwwqyPyfZdJOuKLY2+jVpQTEPuUxca03BBl
0vhYsrMVZBYpNYrsRmnrUfZd5hoyugj6H/+hoKO1ogRQbomQmcdHDUbfm//VmS21fvvQog0ak6Rd
qPLex0ZE0SH0d+elLKpOiywbPpcNBwm4+mMbeqE829Nao0MxYnRQ5wm+CxxxgWm50QEzw5956fqx
Vp531AGhVujW+tq/2gmZqIcojyDfEgTFSkBsttZNnVvnnMM8onoav9jcIHUD3rilH8xFcJyu5lax
OEhCDdojxfIrn8u2HWtF3XjSK3w5he54XjSq3/49TK8HDzxWkaqG9XP7/dSWpc6T7cjYUt03bZZX
HA7I62KiqcisY632CZM4mes/MTn+Y/mfaQH3xqsznDL+J03BAPZgZJoJhkKnvdbZOdN8Q15frSf9
nsmgQDs6IEwADu6nKygr2gGPrC7FSRzn6un+VLZoUtmc5/8ITk/rLwNZB3TAXP558JhrRHun1m5D
IDfC64Lt8gh76upX9Rn/pyRwEyZQicsYe1hi5HOTiRT9K/pse8J/Qb/FOsLQyBGd3krJLQbhXd+V
JItSfl2jEZWnCOUHYE/Y9gera04qSdXbpsr0uIP1hLGQVOxkLb6A4GNlUbTCHIgGQQbAygnx3+nY
wNzGAndiJ/9xJIAym+uBcv0VpKKmHYkhYhEvLMaRTlSec1REQerMKoWwCZEFJcJ+PJKexjb+PXna
NtbVUVv6VDSso3bXXlgajCulDPMjW8goNxv1R9NgApjrYZwo3UTO51LkF2b3s7ogz46ZEGzL5tRl
2SwCpmzYwwSytnZdP9Uqqd6B7eyo7REujVf0S7QUs6yXBVbzVEjGkNACyiLIf/YFFcNTyKIVxWMz
cucrSPYpNcUscBMsAvw5d1IiYkbagQNRGSMrsL115owbDz6SAkyXnRDBSJluC1TO7Zy5vJJzGB4I
DiM1kzeK7PX1qhTCfcM2n8vZ+RxIgE4Itz/u3yDPNMuIkHJjaaf1KRi+jjaaO9CSuqWEvRafVK7z
xL6Xpvh1f/JJ/6xDIL0MViwui46ZVXIm4GVyRbawFkuGg1bArJLQIbUPsi7SqLuwCklL1qOpalsb
irbuvaFoGxIzyOAS0DJTutZetYySant8nkFz3ghAXTy65Udqi/2rUP6ayALgByKgbXdYxOL+9BNI
NmCX3YGoyqip4mE5j4c2nrGAd6F0q0vuOBscCgkJPMg7no7SBfnZjlJlAa4zTgUc1M7TmiG1FORN
sDdHIPgcV/WuAdVY7R2MSf2p4gWO3khdl0+vSSb5XcZqLTHKTOrnjZszmukVDLZkS5nQiLhAZjrW
hKUQu8obm5xOQZsWLq3BLov2ZAuskJRTUjgTDb0CetCFRrRJ6kRWlhib6yXfjnGPgHcueyAriN2a
uiHsXXbDSsefUnetN6IUdCb9eYT5myU6Z7fcU+0qOp25EMqajkO0coeROMTShcWIDW/iuwDsTvdg
KsTku9/K92fWDv2ETHFeXveyYuZdwBZiuaEqx9J9biuT1n9lrSNHXWH3GJn3euSad1l26LsmaHlK
Pr2PwR4E90/pV2kYY5Jh2ZM219orzPK3hqwzpRsLQ6rWrtuKZBTb+3Ocnb8CdvjNguAh0OXzDhkn
8ETmTAX3mAmMlfWOBU3+8TvR49JFBJ+GY24c40/tYNuvJTdQHWSwzS+nDRtokdBVB1rqukJMXgUS
YsSqskpg4f84gHPWsrmmED9rmu+dX64OCmlahj5syUkVVkmcLSN9FwlHSujgAHKeA2YwRM0NuCyP
xV+69SlDPEuOD87MrEWiVUdlVWpulzVxXASagZUBxbe7AQ/+gxCcOfF9eAb1l62iBVpbYf90wfw4
2PcKhgEGQQmyh3/McDJWbXcpQRUZ7+Tr2yiE9LurT+4dNiO2yzj8vyjxiwPBBGcSYmS/MD7G4TZ3
svJYeB2HjGoewXo1PHLSly2O4X48fLpE9UvRJCPLwXk+D2nWgqvUbr7yrK3D6Clv/SGXLZ51Grq7
Q1GOZfNTmPWxDEMFYrSDl6lGLPg90ZwiI2Dx1jEmhOm7UjB1bnFxNDTJboEHKSX+zahbHI71Y9Ui
DV38Z/QXVMjiBL9OtzkAt2czr1RDOoMDbJVfLiiW9Jnw/qwrndkkoFQtgS1zbJTCjVbOmJDVbW4K
6AfKW1ssMFMKMjL9afzPL2G0tkpnkCDo7d9cVB9XOGd4a5mhyQW73tViCzSdTiLEl4Lacm6P9/Cg
PjECEIUifSFINLh5L9ejRIRGq8o3QLcEFbqZeYRTlXqcO00LeSdk5Trg+5O3fqwXhIgjo9ggBCdZ
NnmXgq4k6sJPvno8mvpwlhfxA2ge7Ti6tBktYyUqvti/KrlYnolmehacBnJSaq/Lj5NfFp0gpFrQ
9BLQWtsssvIUUcGv5bOvX3wzOWqVD9IiDEj3bRaDmVDviuuwG5XBafBIVwUN1z4sJSSVyVdWZvR6
u46PbFSlBNQsmkdR8knLTX8XFKHaJC45AD9ZUVBRPKkn3i3om44pN1hJQJhei44TICafslRslzX7
qEnmJeV+8/SkYmPiJskNN1H1u6VKVurGyFHsBFCXm87UlMWm3TQYiFJIe9x/OlTgjhW5Sc3AeSZA
PZrNNFi0yJRsgQEUsnY8IeVBJjKowDx/BJvBt/dOjKSzS1v40Dfn+BFoOLHkWM7tmKOtMhfe2Bqa
3WUA+SMEZea5Xr5Y00bq/Wbwvoe6jKYWEYKDp8aVikGos2vcyMWJqnrdqjBIlCfbxwgQfe3Xbu8k
TDogZf3RS/i+Z65ASpl5dgG1O014Ob/hoKgV8XcHgnPJFSsNJIKQfWlCVxrlMiFeHU3WZYTPBm0F
iKnjPZ1hwsE60iP6UeT/QoYJg4RxMBwqWz/x/nGTOqMNYC9LoeV6qlFJTARTAQcBlZWPMm9KmPai
k83jTIHfr2Q/vAV4Ar0SmE1RcInuaN98q/rtn/dXmPnz7GxsP+8OZFdV/Ea71GmeV5DH/OGZrDRb
f3EUElGjA6wzfDPpJ3nhGYp04s1cZcm06g0oC5gYZqQL1VvoIC9z14KiGDJaFhhDrYk9SzQRNjk+
w8Bfx2xM+4VWxa4fDiEKTalP3vj49RF3WZdePEFwf2awp7ds4c1jabKLBpActlFclSriclzjsouv
vJFug6VlHPy+u8rhzBHMVWG/cUuvXTnsj2u431fSbilHtkdtI5tzc/qghLiIg+HKsTGXTRkCLc4Z
y3dsITNygXONN9mD6Z7ArO1MWdtDVo+cAgnKM43LyOyoj0vXGDC2bC2UsRI/W6XCgMk05FZGkMJH
1Wmj2yj+lCwkGZtzPD8W3ISNCo6YAryldkm9qndOn+25ctt1rsvNn5U5ClnBbpVMXnb0oKRdWTSa
osb3jZAgdujM44W+aVb/y/l4EXAa9D0d/gxwz1QjlUda+bydIwZHtSxcP9ZXj51HeFmcVgkg90dH
mK34nWbChzT+ScZhM5jNwSjot5lSJ15i9z1BOH7kl8plmaI/Q2yEC5jkv//kom7Ng80QDeUmzJm+
aRkkwpdYevi0/c43sjJc4pMKeWp6nz6g4mxzneHc52KBZR4HE78xCAU+rZ7NSNQt6CUInNSctKa/
fMrxzZpFB83CPEJpUIOmUD7oEr407Zc782wZ1TKli/MtABV+buXLr5uqFJ2pFYdtgPceIANLPwgq
Bhkwe6E/M1tdS95bURGWnxb0VEmrdughDTBOfSLCjSc7Yr8ecKJJopNN67Y3iyUjI0E7tKA11tpU
su9f0aaUiC7uW6iTJdLotDW/sr6WkwgyrmrKcF9/7O77eYCqY54qHKsQBPYmFNsMZSfvu7aYUcJP
RK6Rn9NTJOmfc+CYwif+nd9xM01fcOk8xoGEfhd2UUohTGt8nkMSYcVoc7qkKjWaBT/zUgxgrE17
JWEI1JOJmTYXgoc6VFeLbAF4t5I3Ps8AAXFdpY0esCGo8DV5ocDkXJPmAXzHPr41WpkrV8+4qPio
wAK+GHUQ9aicvi+AHeSI2qPtRlaq0jvDVrYgJ31dqqiOXxzuT4hTtef1AZQn0lXLSL0el7zhisrK
QHvYURSWnW9mNHR3bcxr9NeBVhHLmIu4cuFYbbSnL276lIBIeStKvNnsVrJOIjdkrUMECRN03Xzv
pBWdaXckweUFH7QsE7W3GpMMQTIryJodbXKYVdyoTL9gCzxiXAJEd3z8slQBdy6Y2POnFJKKJsC1
HL80WJldw8ecNlnWihFj//+m9508RDfnK70kFDTTpfW3ngNAt5rsvjVr+DnX30jOF8IEWjs69ftD
ppRnBg51K6gRcDeUd2xKUa18sqq2gjAatHV6HLKnBUdaMlndKJfz/8Nzgye8fItRLxakGAfFlRWh
CN9s0RWDIYutKWTKJsRMB+BqYfTT2atAjnriAkp04WEZh9JBEbawyJwoZ49WFI8sOZAIRbPyHSyt
JVfpHo+ehqRbKbEsJcg6K3rWvA9LWt+BpVmFClKU0h+hKOfah+aX9DIhqMX8RWmNAOcJpChY88gz
h9Z3+BDw3Jxi8Ci76wU7JH6zcS/fHRNQaFkM2Tmi+rsmNO87C1upu+Ht+SamqmZXkQqZUsN5Z9Lo
yCTyvWHclzS3cI7Wx9ync8Q9/T3jcXReKG7yX5CRuPxWWt7XtRUKiCRGUAYXy4Io2p+YQaZBe5Wz
JVbxMRN1DcfyBz8mwLUyx2kw+X6YH+19/XF6kyvUp3GJdAz8WIpth2xBput9+7jHyP6BM/nMBeCI
PTIsqo2wVgNWk4Iw0pwjbNjgKvc2Xej4Zi0/FM+y0lEdfj+hbwvXDonNcnNYYgitsmq8GnsjJpy3
R4/G+hH/DWhfb1SRP1kDY1RTkBlAYOp7OZjdQcC48nyrckd22BXDUDcW29nelvunt0ozHBPA3AoC
h2DV7Ie0+pyCy073zArkG1wOZJMz3wwlW1Vlb54EmF9XQ4MyhpIpPznCl6RyraGxyTonMADLocZp
lyi78w47PxM3tDXkwT8chSkUYIrNSfGruZrXoPCUujAO7/fXuPZMbHKh+f/DHpy6AGDL6WF7kGrL
XUDj5IjvmWav49rSEM7SnvTqaII0fwxsLPJbrj2M93KrHDVdT1tSv0g0ALKcbmcUFiv1QX93p5eT
pLK7e6MkZ515bWn619dVS6/0XjavLLF+4kG4T4jiBSzo2atx6HXSUW8yHdAlBFFRWLqtVYNL0FWa
iehUJcHVqfcDnH6FKTVVLDDqeAhJMNHjcg3l5v9B+z2IvFBMBMwrNYEPM12BG0wdGd83Ally3vM6
ySfz2j2nt0A4rZW7M7CeH+8mo3gGELjIJT0gUDzWRZL1nMouJNBZTvG2/+slZnFPBiNRmAMQE51u
4mEtdwt5O9gW6lqbqni0rEJjPKEmsnK1vemfdFMxjyGkEhw+5advpFswv9xbqQ1HIB6xA+0MrCde
nbY3+JC2gY0+DQP7lFE8oFbO5ODdYDByiQo68bvVecIdK9qB3PMBD0G+LpvVzYunT/4SIeuDR/wm
H1RnQl+vBmT09oruIOzvr/PzspFOl6nRSFXBmhIidY7d0O3yW/BEFYxoYaetAjHV+AsScAsfFFGd
Z9Wkc205Aj/CvqWHLuk6iimnRhXwH/4OpzWGAo1vDNAwHKL3NOxO7J0oBfjUSgicTEUn57hfEf0P
4NxbHoy5tJqTfWFaS3mXxRLpASRthyCiG4gsEMKOCDtzAjMv9snD1y3gZCHjnOOo11Uh8jmaOEWX
yw962htkPPA8ckIwDRSg1zB9Dp7w/q15DawL521mZWSWjGfQ2xphW4n9/NJ0xvJarzhlsOerNmyG
fttKd6om4jMnWrjCndtrAWRZ/7Sh+8agVsWkTJ+oXoG8EHQi9YaKooOHmbUGsdJp8SrSSvby318Z
5FN73/r9X2xB1z1YPhWBcfmoErKjVqbX13o+Dc8Xy2OfyzUCwqUNWDDhkAPmYKfGU3JLbxyZuA/+
9/bWW2nH9ALlDMKym7DCKPM9YX7hNpKXCRnHt9KQ+KGE/AcL0W+RABDTrVwSmV0VlvgziffpU3Md
oTA5WbpzxfR4/BHThIaGdfm3v3lXTqxqD3bYEb/un47dWNep0QTkq15ik6T4+9nIot9zDLe/8seP
RGewge0zjrQIAUT1ZWyuWHlgDgKsSDpTphuwtI6CT0bUWf1x6Jc7A54xnjLJSVKlAJVJqRzNtHjW
sjz8wwyvqRy3uPdRUT6Umr/VvR4mjpZlv3SWtdhzdFoZwe7bzrxVqmUB/DCzx42hJCCfr3p3XGz6
CfybCczOw5OQNiNiMLRuNJEQIwtxxukSWLRYi8AwE6rcp9Eh7M/uRDZ/9BUtJILd0BasC65hhR6x
it6UokAuKsFI5UFcpdveVnKNkInDOFobT3gYhtVekndhoonSk9j5AodFiPZHhefIaxCFRVt69I0x
mEB+q45ChuOKG21E4FVeTcMDjbdNCiC5DKJGaM5SNNitTkajhrEiSfaBOivbik6+FrVfmNyheHqh
mCrrMKy0iSOh+BLOBuZZ34cGExbHxiup5XWPIP8GLqELdUho2+5JyXLPFZKe9iLFX/J64b0WxqXT
GVebodow96HVko9+eGgCOYGI2RiynF1WtQZmDJxdF6GjoMPTziP2K8Z+K2yOx4f1L/jtbbleQAJa
Kjr2TvaZVnqu8p6S+AOMvAVCIVAdFoHkLp8Mx221tf54+Y5EdgwqNvMNOeDEz4tT+qIfXjNAwACq
TEcVLp5xiDqBLUM9ODZlZ8Rns7ruqwQ2pqJvcK/FgYdaMOSwBMImntsPQmnlHIItflsqTFldhiYl
CgDjUwpJzMFDSFIUMGHVM7Kw0wesVM2OW8Y6g3mPWUX4l/sxMLsAghOxerOt7Di5SToQ92OHoaJg
2nNtU58KIe/hhbmEGNtiNLs6jj7WdudH+N6GB2pvfppmoX0hp1lRtD7WoNuAucwlpT/r2QNAikLm
OGquAHrC8/2526EtYUJJ0JNs8EZFy6eSdj9DA/qENG9b/22x+t5MqN1JTrMyp9MAWRtR+8rZN26e
V8vffc/UWqoOK5isjcW8W/QLhjIHLVtDNKKnbIqgHSbNplYirKBOwRQCqe1N7nohpANGG8lzQfGR
6i+bOXCm5ZBe6BT6KAJwi9OsCyxDOnqYh4xPWXsvha8UuZOIaQcdYXzRQw/WqQgq8mv2RanMBIMa
z6bGnAxqXiJReGQKZNNH3LavzK0kNJ8dJD++nzggOBwWEd/QJ2yCVROtbkLcAP+1SozUWLT7BcX8
vCMTHXCl1tAU8JMGIMJ7bBs5o965tXIZ4/Rt428JIZJCdyDkjJOnS2ympR/5To7mprJsmqUohLAh
bVkDzeyArUs9DScBj7Y1agcXtIL7lmDsfjsa/mvNCmD23aeEsM/TR85PCBemI64LwlZed7dHJXl7
1kVIRlzcWlpTtl+mB+yc272gJLd+z8/OdC4qiZ0QdoytfiB39sGkR62M0H+yMR4bQrwyY4kLmIGb
2c0fIXXJxLEjWwVkLZHNIIsmoSjQlN+hFt3wJ3YuLtZePoz/0OSFnYyfvLEelIRW7mfcLIRPvTWf
yTXf9vya+11BG2780eHnA/3bw7eLMHQ3qaNDNSB5RgAeiAi83fQJ9yyr8N6GOnf3tfT//9P41oHK
Y25aQM5tAO58l51TB40680b5t54Faj61I1u2xJsNYlhZjNKTz3DX7yf9cu81G4FsYp4c9psaXJtJ
FUQIQCxt/6G0qLJIv12rnTRvgjg94dheEkiheKHAQGJFmmb/AYs8ntUpUPdMOcUZkaVA1zhJl730
Od73GBn16gh7hJ+q6SMMhGHZVO4l7GyPUvyaw6Ja6duMOyVR1vNhI4EDC19k6kP3GoJJW1ksrCHG
vF8FcOhtZ0jMtWawQnPkPiJBhbDYB4Xi5dCxRIAD8r9J3ZOqipxS8hCCOMz6qrUnJYnpyhPC+CkC
tjVs8Lw2aMNCUwj9E/gLvz1rQIjglKpbi01aCt2gA1g/zHGIyRWePYjjGlJiqbmyBBDW5Jse5yVo
nOV1TED5iTbtkkvbzndsz/54impuLLVY2/2VVPoyfC/YH0gpMViq5ryCCZvT5EEdZOCMA907aFTt
d+UvRhgQzb/g7BdcLg+w2A0gdD2LbRPIYtTH5hmIUAY46BsAOM2WkUnGN7/EzHON18HQAVGThwl2
Wgi31pexjYCgpls2Cg95q7uLhL9UdoocixnNircLPSxLAnnNh05j4gH5ileih1ZfNKgvBd/StJfk
q4+hvybFcJ6lhGUBNZ1D/oZ1XWE5opK6Qy1uwmpoQG54B3ESGJ6GpGgWI3hacH3U9olqb3fRpROM
Rf5q08y6+d4J5bgniYssXoqE2WAUK2re8GTiMfIK4qV1wnKqEsauI//FdjzRqcQE0PR858KFUsbD
xY2bHlY+HPw3PZIxljgQ0X2Q/qS3/T5omWoMB/vmk3tDDwMzXHq7xlPCgIywc5/aUIqzbvT0omK6
ZZUMqPamKrp1UsOrxXlP+zr0Omf/z7d/xSV9o6LSf5uxhRORiQU2Yc8L6acKbdqxHLMkRskTK0o/
CavF4Dcbf4yy4wAwtZTOomIkW7mB3WZ2RNo6y4jCMu98OHlBl5kIUv/hXHPf6xkI/ov7rqhCqA+h
KPjFQu/bnHW1VA6M+mEjrK1pNZ5XsvGYDLtjOH8b6xJwQP56Jnd2oUGeIXvNPiFiRHjJG4g2bQCb
CE0XONGpMTeFy/YadTz6f140khbflgIu0VYqcQyRwj8Qby/CqrrQFEvGNLFN23z+x9RHO+Lo5Hkf
6AMODbkkMGdGPd3t58CfMpXdSNFsBr7QU2cqdFCuVfAvfjwJtuVqm3/rXgqkxqVItkpBigF5k/uM
O26q43BkKQ7IawhPqkrNFGIrVpLNMNL1sF4rgbZgOebyvmPSEjOn2EjHIeatVuoKJf0//HSMyW8o
t/It2zRQ2vio3L2EeSARVbpgnXqnE6JHPMmXAkNv9f/vDufHIoNrSG9ajsmr+8GM6coqsgGHPjb1
9Elqiw4Xef0sRz0V/ELuUw9ZgqEGqDbPUvF3XoXOi3GKwTzTSluplndi2Sa585X0D9QEgdgD2Rum
WokfPZlnkUoAV6hcAQSzL/eiwMK61Xl94KLnrcIkjC0zTTm1Zkhtu1LSGx5KMi8k6dOcKLgXOWzi
UbHMLbek7+fmT326wJzVlqOjDt0ROmCwwGuXp8kynqNyjdBCnJNIo0UpBOQEReo5ygye2Nm7w001
pFpoqgcXxqVxiVApNiX54yERDJkMuigja5V7/ztBWXgsAxaXdYUMLOSfJbjJFXuvTtZOS0DDRLSV
cEM8Wi7t2mpkpU+/d5s4Z37ru11OsSJdDfP1FyVrTp63MrFLnDvgVPXAtn4TJdpAUrYr4V/ZauLD
ql814nBmUa4Kr8f9KyU9Du6nOh2DKl9En8t91hFvWfZmjAyjWlnlorJU4UwH8vfawrFmA1EGjQNe
CsxGzPHnvMXQPvRxGMkqRjRIABAF/PIeUz/geL+b8kCjnIM+aidUZipgR9PNyYSCqWVx2Ue1rmy1
FsiVtUb7TT54HwrZ6V5Q6qC3VybgUbGBqJSxTyN3o1yO1d8hbb2rf+mHIXnu1BrpQaAVNDc+6S2V
It/+W/zrVXxautRtpuBLFWhQnQf+h3T93r+v0pw/zJAKpe7WDI/e+4elZaFLC65NrXraq9cxuwqi
3l/ow5FngT+pgoMH2yrZMWSEiNvy7wrvkscfPsUvHllWXvd8A6ZDexhILi2gNvXsnBrxTH39TC5s
0S3a63rHe5HauF52IqoMcv0m3QlbfgAruGn2dqvlHsUlcyuGpvmLyqAmJYP6Dychk1PEFAIh+7sI
JUphy3bN+0GHTwhhd7cj817jWo+FEkfVBgQ4worhC/ct1RPGFG3Eg5aVUYjmtZWU32o71f6QxZWV
ksYLrD3lEK1jzuua0tOnlE1bcCcb71bzMzJhj1ixrrq0sTO7JrECmIoKo4o3JabADGPyzoS5PdCH
0vqOF7N0p3+c2ekPx3c9lBDYehz20fVT3zQu7tmosW7Jp6SiKueajIAAv4UoCFkI44jl7RzYD/rW
vNFdkz1OWaxUw1/jHRVWxhNlXhYh573j9JLQLkSX+OUb+6SfuaPGGdkQDmq4Wmvz2YfZiN22FQW9
fOu/yKj00X0bTVUphnQRrCI6U5wyf89lFEUvIlghA1ryZOv8c2BQyJzqNZ11p2PM5EaK4QooBeJd
cSf0/4jjzemtSFUwNA5f3bfTlbuZH6WJTn39ctgLulFEtiS3DfgbdA6rTKVlmQrqxFopFZiJrMWd
Crkq9XXseVJwdigQRwC3IuLC0IY9QErz0XczssDRvDXRtkLT7z01gYVscAY+DwTIFhWLbIae417E
YrUKUK+Wd4Dwb8Cmq9jP7knrWGZZsdP2dlcBaVZK0ceYUjEnCnF0aj/5Pme7Ks3g+w9sWVonps7b
/EO5So8XlM8d4T17550T3WvDelB0DxbCUQjyDA93s+0QvbAcgsN8bFCpvqt/QkAKHCCMvQqRbtG1
C7oSikQBFqmfuGdVaLW7kMACN4jovwAF0eBPAQr9IgYyAr3ro5Vx2M8XnHac2izn6EEIkAIUATFf
DnyYM7PdjydYgbEccqENwyFhfQT7a+oW27JniClxxjZJIcT4i5l+WbTUM6oGLmdmw6/853imkxLO
dVANbLy5y+vMrPxr1MCgmKWtraqWjWtmCAaILeiAUhzcnzQM569TvjRVxIjkqirW5Mo2GhhSExh9
Aqy8cwVJepsSa+8B1hjVSOSAGZiTRjHxJ2K616zlzzIf/0TGTOBLmOxZeUKOnpy5VJbxM1ynrFzC
vnUOoB7oaSf34N2LD9UXA7nsIzFuEhkue1+o9Md1KXwaTWcSzQDaA4mDuxDpYhAnUGWM9gWk/884
kWOh3TwkVcomaRGHVIwPLifmv5bmz5bNIWUPMP9ck9a6f2AwKhrvmzIjoi1Dhj6w7BLTtM+S2z3/
aV906QTq5XDBWQ13U4ugHGVhvvwmXSDFFpJ+d9rO0Tx13n93pAIHOi89WchgQfHK5g6F+C+/t6m1
SqlI/6+beJ3p2g2YTQ4+xVxatcLTMwoLLeJsF880qEaF32e1gemNVk6/TzqtvH8zwqcDQWyDgA+2
SNtZRwakSLofO6443Fsua5NyGxXZMflxjp/+stuloXKVfRugpVxtmC+MZEqRmU1wgObPbOcBKmsu
WZao7h5/Twf9S4HziGrG5vdfikiDo1GCMnA37pG87jHaV5m+ddHzhxwzKU2wYmGY158XznztL5De
BVPBfktN6nt1O4T4OOKrqJGSnbp2ZLRial6epaMzIVbPfjvqxylu1FLwyzPf/+SM5vufwx7K6fvu
1KZhqYRrTh4F+b1souSVTDveaO+sox7xpU9FoyHJ+GGwxnva93yEf6+2+i2rb3pRek2ngfKq3dVM
g+h7Pfiw7bp8mw3p7GiGyZaE6sqbpkgu23t2doly1BPnsOeeof4yRsKS/6EOFykpTfuCCeX2AfxA
dIiRXimkkK7uJQoHqDd1jo2gpga6m7gyZCdUt+RGNoQj/pRsj5mAiRvceLt81FO0QnR95mKpAljf
N+u2s9nZHHADwLxsLLke+6jqON6y/IsW0b+9DCy0mq52SSH0Afr+V4JNLBuaMfd9JUu1QxTaXq3Q
jTtl8MJfBfObuSuHgXWKxINt1ZtCe088w9MAQRiyUCmVG2yVL8+EaZyOdpilBiNpKuTiZY7yr3Kb
Bdl6xOvlxWB7kbNs5eAHzG4Uq28PR/B4HtLM40+W/KxyaLHvNXxmlIqym4O0ixMO5v686AtZvqiA
/I+yn77XYrkttvw8UOME1WQpDxFDROCjfi3lOcRYCacUWWp+AdHu7JBVMILCjI95nTPVvW/Lebks
n2ed2/xOWjaREGbPiGTnTZvOqJwGBeMjqd4UGfprEQ2+b90iRRFVc9+QDNNKRzN6/MFyB58P03Zn
eaTE2rPhMS7q79JlJLeye96814eRsNhSFEZwD5RTDtHz1wYhBJ/Z1Kp+3W595hjzHsw6M/XuOkhi
4PV4uhublCa+wSU4DJLYPzyMYEOFCWvmpHiZEb3Jx2qCVLUbhDj54Vtg+Ti47N6F3/UW2WY53Yft
DEYMACoQe05lwUaxaeK/s2aYrHgEjTqjo1Q6961+lW9r+PZvA3PUYYvG21j4nOfsd9Ac3Jza+pim
eiO7AE56WRIt/HUJnMOGRN3qgFvsjt82lUtB4AMXNanyOp936lGm4R9Sk5QTwhYb/m8/cDWF93nQ
b6aEU0QNt/+VVp/CRhmrgjmD672Pdtv7/h0H22Apn8Uj/QW6u+1N02KhVIjwjJ0224mPSzTDs6MP
MCOfO/DWkLlkLegfND5h3ZiWppilWY95VbJtv/RinteaV2NdPKUzKzYhU0PdwKaT/IRkeE2Z7usL
AIIzT5Wn8hBd/Mx/ekUg24fCw5AyQV5nlyzk8hBW4Hh+DZ9a8XcrPtHn3rQE9EEmpg3wZK2Dm1VZ
6ip2SeIySWXbwbtxPyxj7VeRrGYpIAplnoa8CCp25wxfQUw1pqdmGqpcVlJj5gRGqmnEfeIhIMNA
DrCqShDp4p658iBi6D0/Ce3g638Q5YfZuBHNVHanwBGeqtR2sYnNiQc7A5q30AFFqSeQkm+oXJf5
kFNinjhI+fH0LW4tN7vluQxXT9zKV1BLxZnNNNltA3dkY2QbgcYdfhM0tOf3q82nY2G8558y3QyJ
kfIY1++EE4g3ZJQIr4C4vclO3Bl06l8wsyT2MGmq3kT6NG0iwiNpRw9OuXWzMN6PtMJyficJtJ9j
w4adLj6Y70t3PLOeTj4jH74LeVLjSsU+EvsQ3+r27rAZyj5066qCn10Vm/U/iUg7v8R/3cYHGMNi
3ERZkILMZUDZTnCtVmHkmDCF+U58GBwQeUkbs5tHQkm5HBJZeLV54+BGi7MjhxH+/GvbrVBAmxJC
cnMQc3+aOd1zAyU3DzZLiKom96HKDh5G6FjYR8w9iK9Dk3UDaBJXigFTz9lu7L1inaD6JIBHFngH
B27EGX+JTIKJMc6OXr/I92Zn5YHFp1ftrijTRFocOXdIXP47It3JjgRIcWSmivSuk/hGtFlNwq47
R79RzMkOF8XYKQiV51SbUQqYpyUTIUGVuCiL5F4Vmp0rM3RO+9CbuTDpw7/M7jQI1zeNUyYpPLwe
IF8CnJM9J9HvIvDFr6ICFcA/gDyDYQtAqBb6KPWmS6p3dnHpGx/htwwyfDvZr7LxyQaf5zjJ2PDN
ohYWo6ttKX3ZVB9Ufy3wMTLhkk752qWaNpByfX7sVbkjz8fszvnNlALyTPQ01wajs2O4qGq0xLZF
IfZ9/HGi19G3izePCoU5KBW0PdCLBusjV5OsRu8ZTaPH/IZ4ruMqomM+qPADnoCd478FryBLy5e7
9KXApXbW/aJbNSaDs0y1rPq4nXLMrjt63yC1zf56wpBquXdLNLonuCGTQQA09B/qYNixl9gEOfIP
nUTIipuWjG6avKhJT35tqoOLiglbBDq7QJj/B65pGrxZETQg+7TCUODghS3jWjmDdeIOmHJ0QArd
G04tZCd1leg8prWvJgv2+HqeLZCh+bRIIusQ1IS+1uYx5sJw7yPaUASBkkld+ZSXR5DaU3LxdjsL
Mgvjfc8zGO0RkLjdrGvH9DQPzVBR1JDaX1nxzlj5Hk3Wgu73ejpOcf5f9Hw9beY9oddYO7QnWrqv
cpZ5pmhHipdvyO2j8amjMFE2XwPYCaWCAAZRz6Cdz8VpCKQ2eQ1VlzXKKSKQbGnMo1IDFSkotOYA
40eBmteCSk9JvVhQWuuBEpowFJgCormWc8gGMnkErNWxpA177bs52m17j3eKxh9toD4JbGsdvPUh
k7ccm3ezF4NUGMXrrFDlNtTTXBtrVxdfBnBr8cCkJY2d3D8pKpIIzOhkpH0/i+dDW42tecZ1x0WD
dtWjx2YwWSfNjp3Ri9yuIcQhtYo/PuTHNVFlP4hBJXnJzpY3ksBbOPr+MAqf4oiY6jn5Kf/+i8+1
swaL8MP2QEO977E9Q5+8yhr46sVPm+ISJJ02JGbtlwGhLvICQfj7iTZ5L6qKJ5fiIESUe6Rag7Nl
T6LKu35HK8TbK4S0JIlgRVJ04CDbAQUmFpYOKyFSgPznXtNnxiq0+znt7hsd+bLylewnCavbUt7G
X7wjSrVC5ASWPNG1c5dsAL1O+ibE/Pghqx3LWk1AEDkFsH+A4FzfDR49Z3se5hoFXq/DCDHV0NTe
SjLu+xtdbSN2+l17EdCXmxOyzhDj34ZvDbrOaf81bm+rarqSKfgDYTYCgC/O5wM/dZbXVz5R8DiK
lw7kve6HbusTnqc5LatfdjzIyUGTZtSS1kcQriZ+O+Y40MsFjakpE7/Al8I5fRIlgTQ37ZfDfD3F
ExgJ6RWNzx2zyHGvfBTrJ4tzFqpf9st/FfMu8xPNGw1abiKhmwZ81WzG4Yf7rGSLCpPgyuSuBOm7
tovef6tx8Hw+x+Ugb6UniW7xwhviD3FBgWokYN3B0ibt8xFH9VJokR7I4G7GW0+0g/gUA2mAg4V4
q/CI7MjiY9iMLrFMZF1MvJrTDfBaD4yZcX4c+0vBiLHLF5Y8OY/zyuh0TecQ9rkcWFtnvCrkX7yf
+Er6oZGGneP+P7iT2TB+AlhRVXZl417e6Li1XIMvPBFgjotHUvW1G2b1ezXk/Rdczfkjerzf9Huy
2XIV+zrWsy7KWrDaP3/+AXhvbo77CrLSgUbaOk9MYCMiM6DYzaBRco+1C3S5p8nxBspLoQ0yEqEG
sUiJOjH0UlgSIsYx0vCRIIDYmjiwyHUVMbq1BoPggH2to4OumZFFBEtAFh1NptsuK1AqIq7mAK5m
R4N0ecsakumg6GefPatLcgi0H9GOS+18dAuBJXihKEmCwhyfUgQjUcYTLIc6gerc0eVNgkkK5SXn
S0cyIdT/DdVhxHEo1UnrFrAdo2npzVbU79YGjlpYovlEfeHw8OcVm5v0pHYoFM21ipLHM+L4KH86
bzQY4U5E6BXyM8akhe2MTZ4EzytXD03i8xW0yNddKf4Ub5QZmrbWdmKKj+PWgHs7vQCRAa/BHdsp
F5OxK4iAfWJvm9j5jXQ7Hamv7wDPlOlloVeGeIBf+EqjpM2McJKkdCRQA67mCVvWbUU+Q2Uj4pIZ
JVZflwT2boEgBN5m1fygFt8kcQl1z/4P4c8S1bLOWWjYJ5PYgJL2+Fulg4ltJ1cq59fA+DPyFzw1
gypq+InzrWlgnAHlk3HdEPDJF7vXngoTpIvtro4UJyZgH9nLnSVETrJRaBhQKcba152k3KVHQsVy
MadpJVjIsGRh0tFIMiJmcc0KpN5fOjSbD80wyIBTZgi+zeoYUsqxIYkSuGlwX1ZeK8ZieRvUOdM2
lPpTtU7u9VJ/tPsPNOXCZxRUc/vRhrkLxA7ZKdTL5OcpoABAuk3lIAfWe//6AbQG+HIUamp/pY5T
zwln3hgAw7buCG8FSmsB6o0H4fdp7tlRHZ+fe5rW3XjHtdzJuc1mZ/LQP224MHycuAjy4h9285O1
hG+n49TabxdNjwkFtoqySQH8XpKdv+Clm9VaVqb8LxdWEzRsCQEjREYkiwHGMNJgdOBwFH7exhFv
Jx3D0eTVOS0UOIO4R4rdVy0abl2ymsSnSvDwJcbnnA4UpqpvoxiTc/CJNpZBUmG7y7xpTaJ0BQ4R
ejmM5zGbRd5mRIxUpS2TNXkXm1MaJVSyWEZM1ZJRxYGsJcU+hWNr47TiALw3bnt+u+T0HgZUuNf4
5VSq4MVy0wcA5CHqz+H4MGs2D5NMSUUhKraXXpUERWL0paXdKgPQEVqGm7FjO9x2b3O5y+P/Lipl
eBAZwY7zaiw4inXg7Lxvw/4PfyWXWS1iBNCkSmnxF0VDkuKWXSAJt2Ja1VGEqqBqgLDMx5QzPOx3
ezmN8lSl/0zWjC9wzF5rbMAddJFuvuNI+qxQ+aoE2z10c4ZCdapwCuvKdOr9BqB8F1w/vhDOetXY
YzZschWIeNxn7UPv4rQXPXj1bv33ln9Z0hg29vMpHkiV7aYd+KfU39liSf/aW+eAXiyy8+9hy+dp
Bm3xIXHSpLF/HRPuh7f74o6+tty59TozyaUZ4u1Nh5pJIOfgnfNZtw2qvYwCvYQy1BMBa1FX+1cq
DTJ0XzOXHWDMGfT/zp1Al60lX7QI9fQm1AfOTHZ4BEoRR1RB8YnjDj+iG4lak1quUz2+tZSQR7l6
jQdaPZtX2BZ/KcJifjTEcpTz15ub5+2qBGhsPBPIDShCbjPsJcjR6V2zX5SFICTRFwg7jH4aOW+Q
/mveKETzs6jcP96pGSxQrfadrFcb5mQ4LpifZ4zrW6DLqNbWl55ypC5+eWqD0W+BpGgn96MUyMct
BFqSrKVq8Z1QOsXhh+ZtH1wIuvjlsjUPhU4WLNPRYQN5EzbqFRJ2b5JTnTyaCmI0lXUASp9SMbXD
1mBrL6XhuWgrEHHdqu/p2TeCY1kQzflu6rmKn3S0goffCXyREotrcRs/53GYPggHCZKof0Lf5H8/
BHENkpVdRNAp3EiMDiHOcQMaeNB2WeuhLdcKmmW4mqFbC3ZDAFInqJgHta4SNrvrqaztpt1/1so2
cA1S3NgheHZozq3PuWDx0ubAtAZzg7mS+VQQB7SNh/N4Dct029hNH+hZD0tIxl4a7OsjbILLpIUR
4pr2osPk8b0dkyPUSVTa5Az5JO96Qj20lFWupgQlxxZkzcknnJrZM7NLzENkM4VV8aumBwivw7Ef
MdRoUwXqJbAcx0GROSbS5KOCSekADOE68ZnBMY6h2qZA4lWTtveOb35B+YE/9WHR2skVn/hhrbfJ
5WdRUriUWExiUhfcWisZA3R6S7HUy5Q+Rz0njYBVweMRnGj8cMoVddq2hZpcY11XwI+A7p5B+WL4
ARURI92W1hMC1PJ+yWZIzD4LyEQJM40qP8h+jYqf8BmaWxxQKtSBCMW4RfaoFQPtotWl1qAGL6nA
B26BihYMMn13lNlEpO7Ba4nwoRqVlUixzPY/e4BF+knaKpbda6F5HYIVFc2ltjOH6FeSWe5jBqG8
g9nBpRZ1wPFbFbur04AtGNTqNqwWHLG6Z7IPFHTdrmrDvbGC8XMS7ogqboyQXALPn6KRdnrRnnF/
57dqVMqRbivphiSKlU2ScfwMsyO9FSrvk4z/ZK2pj4pC9fF9lGyoasHmGIJ1D5Y140vOiJQNmKNv
3oDstceQJE3g2ejdiY2iblbrkas/4vANLx6hlayzBJaXg22RcTS8yeW6esxr87bAQjl8yvN+a3Se
+J5o1ttHEBaTPJ17cyQGdefJAepWJs7JQqNIhvCuGb/Vv4XM19W5HYLSZWK3TeJasGjXAnY6t5/8
vcptynqs4F3b617e852rPOa3qPeHehkE1BwCy620CKJvrfv33gW6S5GsSLXL6yLAtw9+Oa+dh1l3
t4yLPFtz29NZfZfFK8jO3Hfd7Yjzebr39cUKh/GUHuLP9rke42XIR1rJiaSzpE4cebu8NPKxXYx3
rUz3mAxCEgFJEao7xNWeqUvsULkpv99jNjnDFOqZOBaMF8SQvnWYbtXP6n65bd3BpkwTWA1Q3XKu
NKuBGnI/TLuDWUkTOVP21fJngIAPhp6gLd1nzZLrQ07JjTJV4uPKPRsy9V044owVVUh6I7dRDOZL
DKaYDHDaptD0XlF6Q0giWcO5+lZ97nvBV39Gpfy/vxq+3SRijavfPXkkK5LOCFKMM0PE9DIb+I0g
eDDg8gn/VqP5z0bZdmbbTeqyHTX8Zb3OHyThA9z6OlXS1Cym20timwAetFQdfTq0Cvs5tnYtjddb
rXuKvwU4ONFbvFIYCF9ETaWDG4WjBnFtCwbcei8SdjBKTVh/F82j2vmzbUIuex9DT1PlgY66YoiC
49FIVdIZKDIGR61s7notq7IVfachq9ezU4jr8/Abjdte50Ez6antIDSD/gKAlpCrKJ+Wos4joYsv
uegxUj0+eGpDVFF1hy6rBDmG/XaulkTgs8/g66hcgDJkLsqn/hOpJat9H8JOIdvPoA3ttEAzBud6
DZiMPILJQWOqgnI6Q8xHitH3TRViALYmMCL3NzNX68uLH1a0tiB2LE/7YsDzrPOgPHN/vv4QwvV+
QiS7IygCExeJek4AZzw1OvJ7NYiwbE6LlMf8FXvcViJGPYnQe9sp9Hba0VG28NZRSu6B1dmZm2Bc
Ek5+Md/tnG34JBNlKeyAyOJoCewuIN9b+XrnqVgVKMyzCVE2iPFJLgKtC0SJFjVO06ISr4yAtmdm
VHzZHlamKpZD5azdkHEKaqlM7/kWLGl+blG8uwFeinhZhVdu9GeYVfGHWTvbIzppIFB0nA9z9Ovo
Yi7csSeI6OnlP25m+rL0+tCy0NY3sXkGglUukIo9fU1wRnbf8YABZO4ZKL1onJvhghhVb54RCVhF
6umZxxT8bL1UinV0KpyZKQLZNlAVyH+pLiWC+dzpC23fTHNTLNZMdcFfdWka/6P0fHrAnzzlWbZ8
nQcjWrcYhSzw1SSdmzHYMkSpe1XWEYYEANbQAd/L+H/KqFt8ogIWZdhjFsKSnusF52Cs9RO/5WY4
1u2qlmtuY/ZtdAJfyMOIEGbGzzNMV6TKSDD3Ad59PU/VG1jhM4mRz+WB76/RRuCMkxZ6ssH1F9EY
kbnXKjkBul0KQT0oOMxIotV4fSLozUpTqxSIeue0cFoYlW3ZTFvhDwjN8cE/4NRakS11+y2VfNcy
/rTAQp626rXFCAmYXZEXH3pQTJthhWGQKGH3ie5ui5vdSDlo9m1M5PF+wtJ5bi1VRxDVmyd/2tp6
b8NvDfK0tQc7XaKd9MRnaLXsK81Thd4j0KswpBQ5CrPQX7iQ55INwqq4wAvrymbILmgB6XANhTga
rfpGGacZSy4Umkj04B8c42oPH15FNaSiJA/SEKl/GKRoxC8C57GFssuYgC+sQC4imj69xNSMAYbx
8P524lPlSo4+XW6cuqlaZEcfy8HwXd/DC9dbV/JjcOQcMlOCT0UAsGdUk1JlJgkl0lsKqKdx31YM
UXIkdC+TsHKkzFjCaR9ij9Xq4Kg5XETlr1RIRI5jSs17H0mqcEKf2KMrWhE2bkwQCnQqKqz+kKlf
8gKiz9TX6SlhLy7+qmCEh4Py9I9rrpxH6fZWdyuoz5Qz3cbPOihlJjEa5XcIjM0+QgT07yzxG3Ny
8s6NLTdQ+nTX2vUFRhVejj6psX2ah8CRyfq0PQFrCd4KsWuwXOVlItnhy/CPlkjS+hMesmlRYpNY
naKeTJfog78Dy/CuUGHTDeDbaEQzNybUptp2+bWuB+Lf9aDHuuluaOUuR4beEKVCpmdpXpKJcsDG
iFDAQkDgVevy0xdabye+0lfkG7FhQ8ikhqysjn4qXrByWMt4eazIftiWnrs/4YUgTCO3D15oj56H
5xWvy1uSnb0D1/o+V1bma4Nz7JQkNFfrl9qwvCHcohjAEj6tbTUoJws+SmBEM9iADn6SjLBeR7+Y
VGyM2FtKUpHFDZaGwAL8Djr6ctOqYf0bRBeirgf5bgJpb1rvznJJEy2wfzsHym8w6NxfZmZ7rhA/
to2ZOAwKjtmPc6/EiQ4YpbytHkrh4LOdhqDkp0nl7i9/VlakHsFKZnVBFobsnsj1QJl3QtQEd9ym
F/Ll8CRJ4fhTUJk6gUpYqIbzt9GUq2YPZh6K80DwpvRqJDclWnDakr2sX4pBxiicAwhRRY22lL/K
Mbp9bHkJ83D0iHx3KutQ1imWH9jkIXqs3F+v2LPEajzwrbEEvITAK3BZxtlbe6lxqzYf9jV0OfPp
EG1k5reuoyzWyiv0zNSG8amuEbGM+h5S8nErt5hDGG9qJeDF6bg2ESTk9/92oPewYWhvl+21aCSx
O+0cpCV/Qu6xSEKr68LG0btQWbiYTEFghMGHh9JkvaCmSHfxuXM+KYdmEiBFQndO8NrVe+X+C9YQ
yoGwmvG27KanwgewuzKhLtviGro79HL+KDGDLy6pmdsTzG7tES8Zi5+luklzx2CCAsPE+Q09IE8A
MprQKx47jsnG9U8CWQjz3CLT9QflQX6wqvXpNwOCeyf6wExYxMlF614oyl6Jm8mdQdRSmKfgrfJ4
9WGC9kabkmCn672dSp3Ef0rH9UJqfu4YfS/lOLFqnRZohhHIRej7UTxFiuk7z8OPBcBvzVEBclD3
mzb9ghnOIGsemcdsrVhSg7yRWBl9PD6+I8jbMB+Lmi5K/vsu5CDrbLurBFngkZjpDzNwtmFzu49Q
1QA15FWsxjSBKGhFwMzbH/930oSIwaR6KX9busZuZYCie/yfnTILVHrdRKDSq9HqKjKS13bjjSLt
1DTXy2iVizknc27ZdvVDU3KvZhrlGC4lyAillz1Z8NA3SLkn6UDiJbwjwcrSkqIVw1h4RPBcpiSd
oOiG2BIShfs/hhg2DW43/k6lgoMa1r0QleyqzptBW5wQHDUMg1kX4MRgPa+S16m28QXwOY8bdhdX
UFKVQ4L4J+tg0qsu9ZRkzb2ecrCv0QBt+5K5SkJk6EUTEqCyIu/vmBl/pZ1RSexCYMuVRx3beSIl
x1G2HqLZ0uh3ot073vw77NEpmpfbfUyWDmj3YfVnDk8UNlfASIfJPjTgXqBrb1F/OP3VPhDvSL9c
UarfOpnJEnNUVPvdlVwPj3BS4+JSeiPrhpAVGFh99WNvuhW/BHHUFbP1iGfuZe42NVfY/kBMbMUf
KDSO5I8g4C8khw1xwCXorkIVR2A+PqwoaBeIoC2M35a5UcVAlN3lpfwo73ecYXgoBVuKZ7OZbLz9
1yV/cXCArc2hn/0GIGeFXFm1/1Z/Yv4lSXhpAh3muTJ0EDr16LwJstOmY6IVoSPc2FW/f1vWIUZa
2zhO31KsmP7GZLEMrl9jJ0eefqfjvaWvLSQYP0ZUYEptoXOoEtN6eYSZge0DBFfXabtOViDAXb4v
GT5bDSXf+SBTnIkiXJb5VH+2SLyoe1dTceqAJ1S+nISRGd4ysKG7myPzcE0XMckjtjNh8lW5pbfO
fqHbIUWZu07wgUZg1epKJtMTOnqk/ekdPeo5aZKo+MvnHqGAgWFdCYRVi0EjrbUJJqg/AeKu3iNB
MKDFc88h4OQidWWQwM0iMdZ7EPbq1B+HD4DDruIZQZM0BCbpMJAcU98PyjgLLxGvQyCPoh+CKpf6
GFMAyFD4HcuBZ6Dhga4ClBeyNcoH0mDchwbMROsI7nsLd09pkXY7ir2fGR61xWcb221ePwuSeGqE
ujc85rb1Sbh0Pd7GtsmwxgxL+SZBtQToixt3yQ2i/0r/hJECkp/ak4CJZ2LyCq8sKEGIUFVn7YUx
GlZbmQk+NLUbiXZndC5jR+OA41rirzOsxJdOIRpQw6BnZN+4LsM16Hu45t8QW+PcINXH80dVYaun
ufBDT8e6P2QMhSi08XqiH2FVVCyGJSoON3DKq8DptNaakFotBhtLXk4skprA/eSLJA1ua+bxkWnD
JwqLdYJLjbA2+LcBBt7kWK8Z3w799O/QmcaSZUYzHn4tZ4U8vJ+elBljR2RhNcl9THD8gN1pjMJW
3PMaYJ4I6g7v3QheWCADHJ3+P5CHIWmX1n2Jf/9yIZaY/Ur8fibvDJm9hDMENiuiKDgF2CJjBWZJ
0jxLRmdV7zIcirDM/+Du6e+J+cZZ6qJsS0zu+TeY+jR4lgs0t/KP+7eL3Jw1VNY/qZkH4YYfm01d
71LpRiL1672MhIsgKw9vImtEhpb7LqqmV3zvwvljW/cL2Gd+4ZqPCfJIDX94vTR0JtzjIIFny1il
3ws5kOR4K2AjjoHnxYUeDPFLe1FlZ776I7CvhV6Rl06Wandw6keZoJC8z69h1FFo5a4+CTw2Ajk/
gNUQNsisUMQsKYw1xHZu6jrk2V4VXpWwPdpW/67P4gIBVcH8cOuJl5nlebzyi2vQ4z2HfopbOOVK
7Srs3hS5MozY9dtfrBBQIQ2Ab85Ow+C6h6/SRTdYj3fnkKMWarUo3e3utDnn+3ZFkMfoQLEOw01m
2ogO++gp3R6LIUOAxNC/8V9nt5lmqcQQT4kXVW8DuMJiDDfa+L6t28rqbEnWKn0f9B7JWiFMMSGT
cVXZljWJyNKzFzrvwX3plTWPN+igK+7vKoPaCjPY3LJixG8Xs8D8jl5hE1slcJ0KXFKgFtr5Y/4J
FWtM/iOEygx6QMRosfQPN/tpWpdzQ+c3sTGMeJ7o/sAk2uLHaLHM5ljEJYHsLPUhPIGRar+nBbKC
D/wwqdiL3Iub9wKFrEyScAKI/zCVVObnh5NsVliuLiPXsWKYQUUTV5o+KFQC69hZ8J8wqZHWdZPk
hMxRG06MKUpuIRCsbR9xwZ0CfJUGzI66Zpj9udG7Op1yqYMDfBm3m+uYT3B6u/hAlcydPsGXO2kM
rpSW6wqVNBwaKM/w1peLYg0Lkp6+t+ZypgValLJIbuHeiI310crI8tPPYVsX7PNGyVXiAz0v628x
qnYWca0vX5YSAWTV7NbpjbHBSvtRdEV3/2ZMFFOtz+RwcsOLAFEV0kiTPoGpEWZWBjZSavwVOTsC
LAciKt6zuPA5R5iyZdxE/c1TCxABdVHQFt2xcOPnIzGUJgIUW5J4XvVZLlzB6tLCIYYTkbtAj/Zo
D2i77gP+DZyDZQVAwoSjPnezKYEzrpXN177msw2JiBSsVrELNXGGTcC51B4r7OftO/xfdYBV9CWD
Y2LBar/ExLonD44qHN+K5tMjCLYftqbQBdg3z+VB1SIGa5609mLXJC/KfP3UQakkTfXKSxgTWS/r
O0/riRGSrgZLUx54rhKz1RXawBGYgnatD5f90VRQKN0xUbk59N73bkdEMK8qZn3Po6Dm+VMF0yaV
aStAcc+gn0fuC+ranGq5dVzTGwcRG+TFEEuDHwUhR+xRRpoe1F1KnGNtCZ9aCkybc/nQdNLHUU8f
k4Bx00n0d9u6Dtd1IOGVPJbBaPwt01KiWXWb8rjRO9eFyMiypMu8DpytgT9+mi+9C84CbaAeV3ZU
laHGJ5XVswBhT94GWzHs/QBwgVFCybHt8Ej25pHhIfX4/GeG/dK5EVuKCHTmYX13Mto/gHEVC45i
uItwSAToneMkpih7U7NgkisS5eobd724IFFjcEOoUIJ6yymvGOiF5rUDcR4T2ZfS3DwSUrWUc1iq
ZcbfeZcx9kyDbjmc2/6ufFj5gSfzVuILq0oF9oVKldfmyd4ke/u4xFSkXX5kTeyqdappJNR318mU
aKywjUx3uqnRdPpaBqPU4/zsIu/4Cr0Z5xX34prbj8jywZir2RB56CJWaqCVFkXwEHKkcFzpKVY5
tzeqP020DnZUfzxisY/QnF99PXHFYl8mbJiKB7Nbdh6M4OFA2HuYYqNlPXB8e7nu+zZI4Loitph+
QQpkUR8YIh9bSwimCM7peH86cUL5rnVfoQqbbSQnkZb/DgOVyQ3stRP7OrofqSU2/dPH8H/s+hCH
g9DTPXQ1w1QJ2UsuTf0UvNDo42BxM23yfbCOrIAy6fboNhtWr3BtE+i5X9Qb7VPrrS8BqakCxvzD
VY/TCG5SubQ8dJAHfBowb099/vZvOUk+GCjmDG3o9yvkNTJovpfw8vxzc+qpDWTNRONWPVvTNHi3
Yx0Q8olE7cqU4xa5TJxJIyEB2bEyV4obIIUCZp1WJb+hcNeiAxczX2oHqmx62vd4Y8NQsiHaATbF
PtFW5dBYJwTXUogWiMPSwIHUZA7ve3T5QXSTea2qst2sX0l1gisKgzRHMC4bwJhvXsgfTZ1EfAi1
i0HUUbPIdyBkdjv9NJXgti9XE3N6tIfObmkl2upwk0JcjX/wPdGBAiAYid4Aub5hxtoOsylNXMek
OG0aOE815Oukmbc7y2lIe+Mea2GZaXc7wk9fU6ZKZjRee6G7A7BBn4ldntD03gp1JNuVTZgKi5nL
9o0pdbwYCpnREpUVhzxxcdsdMu9+703uD1mWTns6Gb1G4yf8ypdrhj5ARS4z9XDr6+Yx++HUzLD/
qT6Wr35WwlDjqg2NdC4HTqPDbVxLrx9W7pkKaUJyClhd2+qTHyzw9KkFtDZSesy7X2nkzQLVSeTj
oVY/lxeLpYEYB7tMQNdiRKvKrIdqgLzMp1OpYvceLzeEdHspKrP07NDm1Kzcap4Zk6vKPF96LwKg
diMZB4zJRLF43tm0KQ+2/CuuOdMj768Rkzb4KntuF8UD1H/PY9JgzzpGKByIvY3gESCxsIk366Mx
TAAd2enbLQCH0vix7yPWRXbphwBkhhCMv2apK/uA9nagparTpna44QzbWJEvCAnd00WJ6kNNJDya
U3w2SuV8Og2Ot1LDnw1w+Je4L7Us7WDVKHUHcbBVYSsmqikMHBbP6+4HXiyggjarVXABxApKmYol
KyWf7YMGdGsDUKrUkT2pQxBqdXvhMEZ3rE3ATh4oThszmlDislYHrzPEDLnIndfnWi1ipqPUeh7Z
qOLov8IXDRF/T6FUa0X0ulWx7dHh9WLN8FPeIv8okOZRovkzClKYINzf7naTPakCYHiuRfxI7+O3
/6EaIkqD9muTSknl6mB4DzCBRLQDR56aaSVm6XzNa3aTHh4TCBCDm7/xOj/96Egf1De1hygzu5r/
v/6agVvDFOO6eZhVK0LPI2Z3CPe5rBTMOJNiWl3qeGVJhU/OK6JYk9MBLE5c+qoCzVLlNH8A+Xs+
sljP9+MX6R7iRr6LFLRYS2v/eIuiSrQTSNRzRlI8lBBpYCLxehkI/Q760UBg/kUfqh0z3Vw3Ixbn
tBgJjJMZJvA7mfZyzNfcSGu7JYlnfSLoZw+L0iGgUGLXILPE0CHn1X7kn7P+Onc7RdG6NFhuCUmm
f9SzdTSp3fhsbeMXaJXhqC/Pjmo8yHToEKJUo+eJpwdN3w0+LmHChDtoF/NEBMv/ehTZhiQ2AfPX
pkSgN//z1tydKuaJou6eBbaFDjq+rdMswbGxiTXh+fQwc8nKFSXAFRduMWnBS2lgQVefm71T9Rr5
3d7W+JVsGGBEzpRiufTJEPydS7V7KKwtZCNILWepRW9+gOZXaiR0mOVx7U4dT+7BQc9OZqYIWMwj
qW9ylp+Kg80ND0Dkb5OqUUYkKkuAjgxIaYv/OI4RAk0UDDW/vthBTi7reirtsbCbjQjZZ0qUiWSF
yVgo2ibfNSAtW1Pmy15ED9cpRd0UAaC3YJHCU7irZeR1tOlqsNrNCUb0o7MTMqKEjJLhwSldgxJ1
yiuBvACVIj8ZScHqvLotfNwGXGGDyeWP3TgMeIgtyElanQCkbUWqN/Gdfy+KZKSkM2MdtY+Mp259
uFTRmJZai/lNzjfkvajF5KGc8W4pTB1zdpqMUWhmJd8xX26nPOk2lo68bQ8a2XT4KL7v7gCZknV4
x6jrR1ZjULM+AMQmmmre6EEpjyc5mnU8Rc1QSSlSvI52CGa4Co7KHCxAGEl1DM1SCOdb5/2F7RwH
hXMn4praQCkF8OyQxUw/++9R7UyERx009Vg2OBCk7ONe/BDEgyhqAfn7aSNYSGCOFaD/RYkrJywN
O7NwTPENmGorRBLAy5U5KIlWRtKpdU+PB2BW6sii+27kiOtbtFObcsID6L4btE7I/Ckl2+xrjb/j
CHtsKp04xF39fmAi2Hd82RAcqVgb4FlKt5ubvopXRZ1r9TZKDbm03P7UBsRgmGAVyxpX+xLnXClI
0Y1z1coMAcFlb8pj/G+q2MzqYCnUKHWam05RbnpTWdEx/1B6OCxjRXGni24v7bvgLjM0Floci355
qxVMdAUuBhfGqGzl/Sz/H+zauWGCVQqTDuk3nYoZlNxZnB6mZ3TweSvXbR94MNRjVzDhZ0OMbirQ
VZjz/GfpgSDoKfH8opQ7cjEvUIhjDW3YxSgYvYxiK2r8gt6kgGuWJf8yRgXYdDh8BhQqu1fIa8ZV
fD3i+uPWIP1miV3kRqTXy/6BOAU8zEZnIHfp3XVR96EQy9aLzQikKGTrR8wbSdKvGok2HRcray4K
F+NGSkFRX4rMDQOphTvQvIv2hoMVpIYhIgfPAzBbTghxwLzuQ+DeYk8APxxXMwLg9VJw/iTufhQx
cyAEqtodHwnpv8OxcuaxdIZ41HZtCTHkMvMyRJDyYoG36HdXXBuCxjPmzxLJAwkymx6L4HR0kY7O
ETvhrOzIrX8fiUEI/TS20Z6wXdMl14j/ZePbuIg8uz4fIfhEeI+oHqMRW5HXLHHE0gXjUhlwSW3K
hum5WLjcc4/ut1Poup5aYXfLEIvcrjHZOukA4UAu2ysodnaOb4+VA5aenR+qZoe4RaYc1M6r7K4g
d58oJEG6/lDp62sMm1rYQLO99Eb8yLIkuvViY/uCJImwof3mqegEEhN0Wtaqys1zvwpRg1oouZQC
aS923QpkEUO7O4rC8xWGDEsQGtCN+7iDbVHlnorEW+6uxYUTVXpgafnbDiZ0fsKvNurQYhRqLqgR
in8CdqBdQGsBQk9QKbP55Bvx3TyHgDsxzkMk83VCbPO0BkjHuAW1hGDT1/tv//fN510M8frFnF2i
EYNavKdDkDUOArTBXF6lStDOUiUbKwLJzNRebBulvSjb42TUo94Zf51P1fs+cCslJFcL/5bIQNsK
HOYmRuYjDqAKxsrzhgTVSYXZ1TejDaMgm18Fne6AZo3b+LRaqbPJtCuv0QQw18sMaqPiptDP9zOp
LI7nLRy3j4BJZmHko1dJN7eFggkST0r30z4K2Zv/zcxHMivWonsPCntvFid490Q/D30NS+cMk25S
O0VTy2OswEOLro6kFChLjwTIrGPh8nDs99zQfrZs62ia10QJxH0vagpRT1tQgy6Rdcmc9TyixeED
Aqa1vja72TG+TtwGqbJfRfw1ka3w8F6tI5VyhreM9Fe6JdapjqYYUoVfAbzcBn9uBWQFNnm0vAIN
tqgE3hdNT05OqL/B0nrWZt0ZTpKfSPJN3LTSzJs9o0jAx/ef3vgTAuWiU8lv1S/UUNq0xVtf7WFO
37XAaUV6hBtqVp8NjF2dQ8ZAOPvPGDoMK7Fy1tbmafNZT25Z7WmCQLJssWcfSTo8sAs0qp3zcWkh
jG3HLDYQBEo/mUPBbr26wMLaFeCmO5EkKK6hY5VlcIvQTEP2Ll53+PSJxwy0YxxPZzciPkZzMtBQ
psEL+05bUccB4omxqXS10+MpA9o9DvxZcKN8XPItHLwbZyzDDR4u0wg3m5MWS9gbAkeoGx4ZXG68
hR+s0Ptz51KYS4AUv45kD/hkoKKW7ZXtVbF00NFzuU7NyV5uFgP/jsp/FoGxj7wiza7nfS5xjvsX
S8WOj99+sGOdq6p7l/k9UjwxUh8VtC1fApdJhtj/MxqgdHSYGMsnNQtJY1W5VFVpROjjJbEICtdY
V6tS1miHtIhyJ4KqEXOkjHlwDfgq5PcVMhXU4Dft3LGyeuANOtvfOlYXVJ8YW3mIcvE9CmKAd5pe
Z319sFFXrNvF50GmHb/DzP0TRIFHUWLbG8lTZSVrEQigAItnVGQulvNuIu1BXVG2f8xyHfi5pktg
6CdvWlOzIpHtgPEKT/WAnFpahJyeY9NUdQPPdm8YRSWWbi7qQmVBzIk0YoMobfYSAfmCl7so89SR
IruxUt0JwmqmJc5Po0Tqt3MovCoi/83b3x7BaTNNb0XcGpmdcj8Qq18UsBgQvP2AAVejYgKVMqOP
j6o6QlssEYfs4howC7MuryyEdZWpcHDx4pI5AumgD7AEufIC+GVM/qKKeR63ZI+q7urGi4v0CQb7
ifJLhRTSeCGk2wGxV/n2vmkDVfYNnMe6fxgISMkaLAUo64v9LDywfKRFCCoDjn2EYPW49wB4Re9p
W9AAOlqJ+LckHXyHULpxRLvNklwLd1GmTWIjZEjMOmMneIVJGI6pgeb02iGby6Uxa7j/dk1+BRg2
/WbqUPHzVw09YDNugsgKYzvMW/hDSFVSH6GaqjdZ127lD0JShyYUrNJW4B08u9r24gbzNiyk7qYJ
9agOEXE74mtvyHqwsikbWV39UF80pHaVKTQF4aesVdUsUQIkm2wzWFC45FoVfr2cp9uX/IBvEQa2
Daq5k3qcN3mhUTGrto6BoRgk5PsHgTjwATrnqUdjiOedW81JvzplBwEiqpD/fCC4gfqML9/JO6k5
P+/2vq2wd0dLzSietxqOtiLmO0WP7u8BSW35RbX1dIzc6hsVlTOyTvATNx2E3B5s+b/P/zPgy6Gd
OPJhB+AGOim07bg1MM7CJHP6qnlAjhmMTn9WYfVtOsQ2UPnT1W9T6OI7E0MgIyNbV+nzpbXLXTti
op4TlVf90ZoZySxNnCOV8y3exWzo+HlxQ1M6p92JCYYquCHj89LTqyyH+VvgpadKd/XxMgu7gNue
FyDOe//zbJ3gaSi+gDPfah9kKSxjb32xWpXoB1ZaUf/JDPbv4u8Acw4ZAHXygjggTup6qLGPSrsE
F7v55s1oDQ5xyVFWUb73+xS62BKzAE8v0gcFvNFVq1lSrjPdrZNxRnbOExbcidMTZHaF89NXvsry
6OtEBD5zqTSdrWvBjICyFY5kzq5Cv9yYwZm06J+BQtccAChtSwQgTBhNIZzvT/3rwk+CXEThsfDs
A7FZfxZrDNPcie3qv88mE4hOI0yxG9suxfc+BZ4x4Mb8y/07fZvAgaRkIymyCa9xu90MRZfxaW+r
G+tcGwXrH1dJSOhj1H16M8T/OUo4x+FiwrLp/6Xs19Af1ElWu190Sm5OS+9NHtsaIengsaiR50NX
ZH5tCWrNkxSVI6gkNsvctMrvsr9LOAcy/UjRleMSpSPeSHYPv8lIzMv5ytWO3pSss6MeTOlZiLk9
8cjytQoqRRzZapeeIAEMhlpPZKjE3ZPJn1Js9zp7adRqhtHBjLd0UJ2PontTG4qXQBj7sLDlZH5j
zcVJCx/F28t9SBLt4VBvVwtlRdVVOL2673R6eO6HEVvIvRoaGZ9ANCCXWI12N1A+/UDIAqakg6BW
Y/I98ImNmp+3tNSyoMI917b7XUXawJZS6bwM8+CjNO+aHwhmZ7FoW5M16iBxxnoZ7rogcFyPqk7v
LaSSSz6nr4bIbt1SK9VSllPwXzS3BhGOusR1XkWQg+hCvts0whzp3eekWbLUxxsNeRKCjguwJnZc
NgNYXpgzwc1rn7GaKiZq2d9mSFvdqOSrhelXC1psEg8DB6pxzR1mWx8yE+yGOdO8IOaDf0SC0IKF
RlVdglnTa6JA7hkSLeNX6xusSIlFotf03sDp2HKOuUS1Xw4/EJ/X5/1BqXDUWfFEVHHWx95PX1Y4
D88LInqo9rDLGfsjae4QPNpo43siAOigLl/X0ZIl6C9hKuUJoVxpf8aTap6UMZQQgJnyri73ojGc
F7ynkka5jL8alq2vvCe45q+9wR50ywXEfuKnjOTA/DnPsNv4AFa+rK7u2q+y7/QW7zZcm840eWTO
2vGIEQe2VX+2YaMCkceDSXeu0am0KNISrZ1q6cSxVTaCmaj8WDgRFzv1h9Nnnaj9FXIoe4HjoGkG
tVifSeUtkYwViM2pJVZWXajnXaoNwO6WfebbHdydxhAZy/HUfeFRrAx6Qhys+/z27oB+X0NA26Kh
bWxtY2T9eD70A5uvJ7ke7EVd9VtoPIfAOcnkOGkiDf/USWAdc+qv/x2szLX/l8FsTrvIkD4DVq3l
/1TmK6A4sdV8XGxyWiUiOXwmphjKQdKCqqrfB+0omRt4wWF/EE3+Zh7+Y6GSEIvggwe4hS8mflzv
jChfSnLaUzUDQYQkIqkoWdXN9W9xABeaYcZ2gSPFYg8kbB7YHuXpB5FCKYgnN1sNd8qw2tOFb1AK
Verb0Gb0gb6+jXt2Wj7b4xiumtrdfWA+qIZ5gOZDbnaVjm+FwTzM4VxK6sInx0zP7wbtal+28X51
+lrkU9MBIekUbHdP4StwPyn9DHBzEM9FrQPnDlz5Ruj1feGn5OWYNeirCf8aSIzJbyoMpGqsvVhM
Ilo5QtM5kcYcItEMbEGMO4U3hI52Aqxw791ajFIlhV6DH2eJ8IxMMVqoJhSX23BIGBQbKwtouKDi
0qP6oPOoZurmg3JP+fr96vdWA2uXDM2k24We70xkvDicCMUwE1k3ad689WkuC13SQiIhym0pYWJw
+hRBd+Be4jpVXFD66A9gjHwPNxOb2uXWmpxembhhZEhFUCm7fpsIgdjS6igzk/C0j6XzBn180lIh
oazRtaLMe4aO0nB+CPEXLmAA9uth1C7r0neGK0Ra6JYAr1JLtWomiprp4QMg3+YSFWe9apnhmxYG
dLRqXHmLdDh6ZGCaIIxu0vJO7X2SFcfMxUdZBXnWDRT/b+NylUC0Qu/VdMzSZOHxmDPSix3/ERFW
r0NL0Ja1aO16J+RhgKZ49VC2LWid6a7ROX2XURDhk8ovIP4rOry0Fz6WOoRt1CEBbtleA3OVBc6/
Ye0eU/3kB9KSr9DrJ51nxXsLTSIYYq03c8cR7/MWjC8heXoGye1zOiqT0NpUjyetxNb9CeSIPOtq
x6Q5Y4NfC/9M/YeYbIJB6fa2F3dmOxZkgrsl83iZSBTkT/Ab7wi5ttIV/knJ497qN4wVUttwGBti
a3ZOh99zPulD4Qv0C+91VWunosdghYsH4jbcgeQvC1hCdL+SH3BmwfexHxA0B/IohBSvViDeBvFG
ygYRvY8FLBptI1F/GefOBDJRSPQQWHckh6f5tzHPZhe/WM4HT26gq8w9FD03BFIBuHQSVAvUccOf
dreOA0UY3YtfxQ9+zvzNESpQOJUIuk0WgRSmsgpcv1Ft+uyzkDRWXSrLVPd2rbL0/EiJSWGfqcOb
78uwoW4B8SfjOWT4pP1UrJVjZHXfM+l/pEPro78xMvCi5P7LpZuik3VVlI5uom/agTqWFgkvoFRA
nQw59LMbrEHPJkt2h0Xcnu+fNfhcUWZylF5EJJutmtJlD/ucYPWg8lXJl42o1eebwkypmjroVwPM
HBGActerFe9j8H0Wo5wOv5Eza/TGYJNUJBi8ZrKfVumo5Yj13rko+SDqimrhM2uoCHNPEoHwyJvI
ftHG2BhRGTo3hQCE+94E3k9Ifiq5CVA3xiUTcPV3O/d7j2tYK7Kez4ZdoTTpxBeDwODXA/7tygY8
H6fKvN/WefhH6I2dTffznVJ8CUpNWiihwTkCvXcIseit3FLYXx35m+unFFydaWf2y5WIKkb5x2Pf
ErgBloke2BcOuMSFxhrffb6ZFr6uWLOko8u9gWRFETJA7Yg2Ml5cpzSGmm+AW5HUVDeRRc9AU6mS
KEgRHLNDKSp3K2xRolH8L9JsqcPm5gH07jRInpSau4gmPBdZpS+HZc0fVM0LIgBOOIutfkd88zCt
Eg1F1/ZgDm8SuWtJiRJcBaMpz/M2V6e5WrlqTinEoqsFcafjH6h6Kyi+eecnSH4U2M+pCde1OuXy
FEl4RYMRfci2RwFnJ/YPmhAEh9YnGgNS/9weBJBZQljLMm0J4LiNSlzXW/yXP1uEuZdHkaK/c0bf
/ygAM3WuBQT1KzsOKrzlTCzNVKMavRPK9NsckM5zMS07DdEfOe1iRgaPWl+RqSP0zsX+srRKvpFn
v7WNrK6+Z6chx28qaxWZvaC08mAYfGjB6/h5/aYOjkOhe3LdomD5R7AOb69WsNyqf0peMEJKHKZv
at+URi/d1r8X3SFtQpcMTJ2pXsENB/hGsaBUqIMF4LpIgGXdoEybfwB+HvWHyZ3zef5/6CCN792k
YWiGaOrDqWoa0FzBs9N4RqILXXzrYs1P+QAeuR+ysaTTplYdffAULPUJuvjsHQ/LE513t4v55x9w
uiv7WNB3fyU4+RTNs/Hh705/18NYtZOFqQl2BnGBbv6oj2mZ5S/RLeFUkVAPmw+jfhrgY8Ukn2C3
IOJO6ljiQeg8e45SvYfSIurfBDJtLKvd0uknn36prHcK9PUSo8fXWqlzNyNp5ACG3qidiyFTTP3d
XEpKYlxuIFoXe8uRSb+lKS7uuyM63uS1PxXkzGHd9f+zIxcSFglm94Qkvj+5NYUQrtRlEdWbGWwP
x5mVlRbQOOp+Bi44Qi4FdKrm1YogLvcWg0MqwMDIRYnvoukOX9mMFKoDTsb1MVkVhFoq4E03ZyMc
Q/Mhs/xk+ktBpytoEMZ8R8kMEqarS44/Y+TW9vPjSPseE1Y+5XtWKydUrQ1NbgMxNXBHEk7p+aoG
G3vlRAlr5OyXxcUda1ny0THNSkKWOdqJOL30A61GsHfQ8Z6BSI/4zYVoqzfJJTVJMV0hN9dHlWYl
dEVyJOMNBnUldoCHQZSqKHEgjGmi05TfBUFbiXs2hU4oDyHKkOePfXWWg69igS67OWHzJAiLy4X9
Bz8j+sBLoqFXKa84FudFptdlB1WRHY3rbHy5FuFUUd1zAL2hwy0LAHwhCRFaZ3Pn5Z4+dsk56NxY
dAR+gb7+viphh7Stdz/39MECVKDNu4Wi6ni3TlQnDuUVeQGAEtU1Tt9NElgI7zTU8X75DBJLF8KB
ocx5/MidIGyrzrZLMFBovqRIxMajc0zxXTeJfMs1SFgaqzg9R/LOvr1wF6qMaN7W96rq38yBBG/u
CzWTAgOhcbNHBvvNvVinhJrJtWeMbAwx3RMlV3ZpMZwPR/DeTcONpoONciKS7jshzMHFQLZQp4Ev
SAxZzrDmDjlnUxuqLYRlS+g1RdEP8X65sbYqaeKGiTie9nhzFoFHuWR8seL8MxCyWCY/byqBsgvH
acN7FD/NpDipC6CRkVv7m9Tuo6RBrQ1wM5eBEzQFtU0x8say22+RizVnNd+GkNnjvIIA//vlU5kq
l6hmlqDiXEZNVNfcE8cztwcpoeVSCljvA5zgdLz4q/oEIa8kTh0MbTFWeBvZ78ZHIzvtA1BXyi0X
BZRdKK9mKuUb8ubgCZ/8bLLslRSuDNW8jwyywq7CYGzRCKY+Sir+0LfMvkME40anEQ+UoA2fTEkE
OjKZBGUPZep0Jax/K7gAtLOtqh7CjeRt13x77sjYg+06latlMkF1Y6/kHnqlNufRmyWuVZMzP0iH
Bi9CVfZoJE50/F+BAPI8ng2SL0tGKbqV9W1AYaUOVStIBiMOxa4ZlVikkdRI+ipIusq27TKv2/zy
TkUEgUen2Q9mLuf1z7ev1rXrziAdwucIMsp+yLpnKCtu1mI+EqmhNw139ixuXrvs7uCn6ITU9nPA
3//K+In8fR8gdBuQdwGJ9fCD2+FqqJeugObY5oKuCoTA/dBv1toQf0Uq7eNOLfJ2AiwiP7PL1yBY
jHmZ66AMri8moiheGJRFVQ/CtcO64Ety+d4VCJVHDnykmunI7zi61dR9d3Iytwl1WQlk1lVwa0ug
LX7G85Xaji8P+CMAvwa/XqicUAb4MCOlyBIIwkZld58YqeYyFDTFlg+Hjl3CNfN4bRUhEf+LuYvg
zR2daJ2JzlO+OCJQi8jgEofH4necbxEwRynE5NPBuNs1IWvAwFCrmoblS24jsur3pLVTV6AuTiOr
ahpYGQIkVlZfsKs/X07h5NHz567x5KMMd3UcX5k7Oms+SpjSD82NvmshNgqzrwLlrsCyB5Hx6ic+
JyO647B6jo+VIX+kEw4YDO1CMj+54C3t1eOVadW+B4CRJlxWZBZ2WmW56qnmCk34KiPkBG4Ku209
W2xt250erM4EWI4Ps2vz5FI2/lb+lywKnUh8FTpANLeRwecjSILmK5wsusCA+94mjetMtXjCOJSB
EskGYsWDQ4/RqZspkvHPSRkVG0Eu8LWl1tMWCSQETQnbhk58+UgLEqjglYaQVze44sfPb1mXhT4w
d9UQqj8ZXmnTwPdvQlLa/oENyVhXy97/VwZgtywW5d2wrV5gacTNJX6gccCr7wgxJ8zsaAVuRgcz
4BB1QA2KHPDO/T2nByhbq+YLVAvnnsRkTyZIdbXTzzuX6yd1acwIDYQbTGwcS3kxDkw0yyzJQclr
ZrvIgdxmy6SkxgEoWtR4BZE7jvPRUsoNvyxBBtFjM9hMHvFsPlgxQ6udPoZ4fSrrNxe5wPRiggiP
WOj51Evz6dLt9IFWM8mzCB7XVp3qGexykQDWNn6l8qzHkjvunwOvcUYU/cKMkFbqlf/D706CdMG+
kOPbU0bDp8VrmYL/9gzrFeM4TwrV4QV0jwQlFbAdUa881dLRgW05gRFqEyRg7Wmu4nobfN/dU84N
/RjH2NImF/mUkox3RolU+HbS9UY5ZlOKJCyE4/4/9+0AbTsHRZrQMSBKFobt6YvNSukuIDqTLWPc
uY0dZP+X+grXZjHxGHilcOwtgIbMuzkRL5aVuLOw7pCDHOLLnzaxVmxMpXIZRPY8wVeeoSZ8IoVp
yLdUXJzZhRSArERHhl9pR0j5ZicSBw/I62iQeofWhy2ty1hyNlE4aTB/DKW9Y4zlFTc+kp8x+X3q
CE6oKsHTX6aAWUE68iu0/kYXlKdx/4hrqPngC0L2qfhSWZiaOPu0HoUJ98F/VZnWDgVWzHwHz0v3
ZT3kRFlB03V4lRmmB7i6/EIxuUYSnmbmUjDpRiXCZ3v8EuHpegPJCxNVtwN14n7OrQVC9bH6hzy2
9EUI3sXUl02IiKcnmh18ZBsWaD3CJP4fmm3yz9Y4zTNjsfpQJ3nXSQ/9ZLPirs+Oz+BY/EJGFX0Q
ErSsGMYjiRI6ex6kHG5fIpjvo4RYv+MKpe1QefGlAgze4PkGq6VjQMxwc8tXRwOyjAxTRKVfF1oD
X55U+WGhXhZicncp+Nw/SJJpPF9SakEiKZV+JkVN/3hFdP03i+lyjwYh46RfAFw6jz32YlqjjI8g
k87uzMNEgyNgLHq8fJ2a5efUnwdnK1gAg4pVAncmtA+yPHZ5d9EFL3yQnhI5rNei1sA4LOPiHUYh
r+o3fEgS+MXHJTwNIRbfj34llpOoCeKyTGyDOcSacV4OfHB5mk2MDtG8akIVYno8LX9M883HrGbq
TmP6Phz0vCbJ2wf2HlBkFXh4Y6w3i1/UmrJhVDoEIxbYuB61choQwlzzm6Uh1ozR0mZagtSmocvh
9zD4IVuXMXE+vhmdYa2MuZbgglrVlMVHeQ1rkLfGi+2iq+GsMfbC4llhGMuqR8m/G5vZUX2iVjFR
q1H6u1xsxIziSQM1YJm9SmlfpugF9EV1gdge00c0WsAVJVUOJE63yx5w+mzuP/BIPyIobJdsV7he
wEXnqMCo5P/c4cfjNfRfv6uNKjvWJkvAciqowxpe3BJFJKKZI2rsQig9E71jWBXqb7pNtWF7jYJh
SdfWBBVjgtlam9evS++NGR0hi9pkmpdT4yxuuodN62uUduJG/mTPAGr0W1zBE/UHHBIA/c5tT6Nh
ABT/EqLd7oosBC4aCeENB4sbEL73EPNAG9g6wqK/+rhZfkthZpRjX7M6AoyBQ/iNkB/VrRXdKV/x
GQwefChP6jttR+9lZO+dfZoC7WaqlQ+q0F1mcSSV44HHXe18PR8YFAx0efCAXRs6JhTOX+bQdV+s
xRicpSPNGOCndZeojuKiL2BTGJD/JBeDnA3VDwmjFI2Nc6KBK3JNuBXW6Xlotpf7Wxhl+QNX0Rxe
FiojcxsBOWuIFZ4XD12oPP8HLE6wiWGY4iOllUaze4aw7CyTOEIHKZ3iE7ERXssz8WTZARv6s2di
p9Gkl1Ibj/+v59rrIKDtxLKq4fCKbteCR9ZWuhEcBAq6SNBsRlIzX95yhv9YThHY+4/jEregwxiS
idME7UahCzilZk7y3XQwys8x+ajc5+GIjYyVkShgdOG23yQwgkpOqrSt7p6arwIq9itIS8HcdTm7
XrfyImuk3zRPJUJIOm69sMO0dCXREyeXtR1YgdpektGAIodWfL3/eeqBRYoOzgw2JQr+LTUcqijY
2t1WDwP6vDmvKwcaB3DuLRCVuUwUKmcKSUci42TWj+ObcvgwYuvF6BYk9M+7HVpC0ZpL25q6C4jr
/E8WrnUhduYEb7/ilgmp33lMaDA5KqPadFOtR4UK7QA+7BhwZ+vK9XgBKs+7JMMR9UIux+7IjW5D
R9TazaYeiny+3nti3yrfMiG8aJoixJY76GGfq6cxH8q8riCJSofqreYwdCwfR7QN/OsFcI67d1aZ
aJmmxsqAT+hNjLGE00D0wTldn/G+dd42X9W9OScg7Phw4/Z7voRlcFy2sv1YRbOVMgE54njc6Lqw
mxGuHatwrIDr8hpBkasoZZ5VQf6MLVABVi/QIIGGc8Tf3ZTtXle8mdYiCruZnYEy+Ku5XN+BvfU+
Nj5NHXm+jLiDDk+WkjoEXH1CAPtxn8IModOzyoaXrm2dIH1wPZkS/iC4qCOp299P2uPp8yIHWjii
vVkjUTdjz1l9D8h6h5K/oNYH5wGM8AOMrO1LsmRr83t536RRfApvgsaAuJ84zE8S2ghH+nm4OAy6
J5Bh7JL2vsO0k50yUkLQv4A6Q8UooT+/dxuPKiUEUZAEIrdOj5wscEGIF9QBLW5CzxyK3sf9aLKK
Pz4HcZFXJcp7nbn/uQmYBhg4jXS4nVh5jp5HshcNtFjGA0HRrC0pvZDaWh/AVOeQOm5pmQGHr0Uc
sWZok1ny2VoDsM4QOMfBDJ44PbBZli+3t3eFj38Hoi1VGvoix605E6e7SyB9eLy8yizlzguXvM3f
IaUsJxXcC5q8Abd28HlcemQd1AFFQifkBJVUf9QUFd3djiFOPD7LR/yn04XE/lKhMy3qD/gWlzI7
8M+mqf8wGtphowzTpDJw2ItHFMEQyeoXMurlBTpU31iqM959EkF5Pq5TQaX6Dsp03JKslJnDNwTx
C04wIr8d3e5Q10cjSRzhr0U9jh39YVuni1sDYKe6vhpLqjZIb3OWU7CNchh+7z9vZeYxz2NdQale
fcpE2JpYeuNzyDdD/6Ua2MS7z4Ja+ziCYGBom1lzYhmpTJsWuAfXQD9xXhdqJuPD/2eNjlE0waCs
7rSHL2DWHLaKbq4zXJGsriDhRt7C/SDGwfNMp1rVUDxh/rDSceUBc+WpMK3U0H/+6ibZBs0ZNFKF
BufkIijs2YBH9UjCnpMrMKzrx4G86KoXT7Qr5Lh+cPYRwGt/lV83aTIvJft/zCaayaATjwLNpYDe
g4lQcjns0y7y4LxrIJz23vQiIdMeoGfB6qEWJn5U/GlUIJvMbZXqiWeyJT+UVV/NLRzVX4pnUMdr
3L3+8QUGF1CqiM9q9FSKSwXjc47ocSMXn6oRA6lPl3vKBDH3sjZagWJRMlcS+Wh9xq1lbRQAIrwX
49uNiaFbUA3FWwvs4QegHb1YaS5SPbXKXFRg1L4EvAEUf21ZbGqqvifN49yt+2m96HQuHBlUDzUe
WimUobeK0CqI9qL05ZimhfcLJBjOYpL3rRzda0bMjsU4tsYTWuILPIurIsbSoiSarNrE44kINwk2
6ZUH0jGxsgLETMaozx3eEjlwa6ntKPCEeEnMnebsBKE7Mc4GPAIfG8v1wGGoFt9VMsxVIS+jpOaB
ieNLNnIhKCbCwlTdfgTzFrRb3U2kpFo2IjcrxbvU9q1EqFkNjeelYV2XzNUR2bVOwSnDydBliSal
IJVyTrzsqW2N+oBlZX+eqgXJWqa3+aRCwkzzDv5tOTm/zgqO9nkKRvoUfS1nzSCwll1D3IqYX7pn
FzCOnPGmu1bLfKvE4FIh/Z9KBfU9U2+OK1/5WYkp0mDH7Gab2CTlOqVLMZZFQVEzrKxcBu9oB2G1
6hCErkMzpwFlu8xGaNGRrDUCEp+OdFKyHdCtiJLI+FFtmE5yLUEnLh0k03PBfww0hUG+scpg2jOK
oHfq8CJCZlb1WbHVRy989o+nPyt9AgtMucB2qaHh7cVeEkvuklAZ8kSbVaHq0/uocpTWiVKCATJn
IiP5v3jtYWLTRbUfXKqNuqzSJZiGs7v/aZZ5LBGEexq1xjxmQM2+5PVOwNCEuH1yeMCN8kQyNQnU
ushNUlsfzP+yrHMhkMg1KYpRQLSZdojLckAV44fFBBmLcyslKynUq8uO0kIjYdsMMBEtXlqXA+3S
wi8oZkESlQPS2gdRHoLSdiPbx3XxhwmYTHD/4xz/D/YuxX3TSP/OoHgKMdZVcgYeM/NP8iVkRVj7
G1AQysb9YJDq28oNQ82YEpVW2ZWNl4/y999x4gqU2qQXDHzKryK8ry8XA5v7KA67S0MiutlK555J
/XH0BhvLtjCBFk/IpDxBi6KXJAfyyBneUcK1RLKhBspQeBGW+UmfvssX0V43tl3PRtvCabk/LfJf
ou7ny5c1JwAS97GjECDADMjVvk7AadYzkEFYkwiLJ5qc4rwMv2yewc7e1LmVj4wxI/RknuFj7Rp6
5EqVFuka5TKhSDNnmDjJ4PZktebLaP+qlEerqELVhNzOhF6+w3pSkZeoCUWmYjSzO+J61EUSUpbv
v1cgIffKnF2ty0B1yVPOfFWjc5DOVzNucrkgSdVFY13cO7Z7yTICai2lqW+sfjyE4drubuhHlCfa
MFrbbV9U9NovpLvwYuNX2hE/NnhHbB4ikfpIAhaIJTXwM11xgxpq/Jb76bSViapEB0s4512ieF5b
5q/w7pGNKNYi3YQCSaIlGJIp+lMWfQjPXOaW/Foz2vtQI2aAVtuii5AqF9iMjHK59s18zBlGh8CW
X/tTyjbEeSQCvttCzAbpgrfnUcmw46Tl2VwV0dK4jFy/usIhhtaSj0vXdOii6zAjNPTOaYO4ExmC
TB/JYjsomM05UKAeO9JCEZ8+nCQQd0G7Ip5gQ96ssTvEmm+A73OAN66bL2EOZrhLVWDMLREUwSdA
mwAJ1dWIqzGeEa70FUIyb52eVdehi6vFZpqKpCSE6h3TkeY1TejkULfUhp0dxrl7HzopF85qx970
1aTu5knR5lE3M9c+jVNwZuGUJQaIpII7gpNPRetJ/Exv6nMEmGsoYoM49xu62BLgNgQxUsHBtgJE
qX6VQKln+Eb1g+6rpmDi5hxcum1cIUMepTduFkUDMXw0YIiFU90oRrLWgn9rN6LLfOBsFB6c/T7Z
Ienny/GLhZsPp8x2Xo3srkHBwjeBWKLgbOE66s2At7epCrngUfmYlPKsaQfsSjaqa2CployQOaVN
AVJQi4GoLT40ztkCGux0xNn0BTT3YDiXKtRqhkBeChe+ZR3feTh+vuvU/EBIXIX05bijXyGZw3A+
zgEYO9TfIrpNlruPbJsJF0wschJZajQasRWTy8s8CdsTSzCqZ+9JJgtYvixQd3DtKIYljSM+SM7u
FC4PlgOvhxeaxLMXu3pTfZDB+9lZfbDOhpSaBEy4q8LGOoA5RzMl3FqLXRZ6jllvdu+jTdPXDaov
PvFe6RqLkphU4U1kj2sAvOjLOgKGTI6VxeFZghWa2q3pa7DPeAT5c541t7dn7HVhHlPzzdzZPt1K
aDrE5VNkXQbWCIUW8gMJJMyEGpt0I6zLDxLAjH5DrvECdubE3XO/t+cG4m6Ixnkk+YUXx53A9/E8
jgc624W+zNJHmmMlPNdN7+alvZathjpfXop1+hyrtCOUYEm3BoYNb2GJ1dWZtzw9tJnx8iyc7XnQ
G4PuCorXcrGxJHUB4FGhbkjoxMHsQsk9JbhtNM+LGBbuL/yRXe7Xa1/Dj2V4fQm3XqrZ57EhYy/q
UuEGcHXsRGViFRvaWD3MIDf0l0uHJP/5s3oLFzqihCsIg/Yri5yplN2hNFdA2lAGIP5x7cB/IDkN
K/PyFtMnVAH5JCxHAvQLnNCpR4qaV1c/EOu07SPyF8VSXqxIOiatbmFPFXbsQ6YQz59REWMaRhjm
3Z/XTG4nPDRKRtPNkUd40Ih1y4xvOX41mV2PruTxlD9TLHfXyT1X12qCn5Vv2YXX6TvlXyMzlmnp
mYfDzhfFC+aCps4eNx2+y6MCrxYJObfzShTEdDarWoarOosf/689Srt9P2X0PmmODXf9nuOLpVYq
LK/B0FuY9fi+ynoUx92mFJvOtZDvIqU01Mqm9RRsg8Pj4i76Hlq06hAFxOYxJJeiOVz/DLKp4Ugn
Tdb9RaAhZxtWwGYjI2lxJGL5YngLbeCwDCopOCuPknhaRwpv5YmmtfTPTIBeZqPsSArRcpWsNIXt
7SD9YvAezOc/fV8/mmlA6PGQ8yMtBuh3iXKca4E+yPpb5/5vXwLTJDRohAT4SuuHLVwN30+Xb0Dt
gvTdInN55Ks4TnIjv2F5iND6clmXRrZiB67va2wEW+2Z3bRADaW00xgGCSrZxqvzdKM2jrtqCvK/
Xw0rBsy2BbV8fmhT/wGCTk0JZne4+LDICgMMmGagNrSUKsuqWanEOSdowciuHNR3EqvMZgCLr7Rd
7p0DRfkqxntr5hj2nI5k5XF88xrEea8R0GJ+xtPbsxQktDI3XsB8Wpxe5qvoMEBROeJhPOLNBUi/
0HvpyFW1V4Yg0Xv5tvnQhf9FNeG/8l6N+Ozd8iMU1DdByAFGjZwueRbhZSWs38IZVyt8z7fnjvuq
PKhlRdh2BnJk9hxQN6ISqQgyh9tfp3CKdPTxlifot/4bYRYsK1xr60o211Z/8UjHAIHhGpxN5w/a
1tPUiL4OhOP49h9y0mIEbuaqQP/6Pe+LcreCJdRwBeFzIWPFsR+9GKD/jAaKJCDodZLPQwerTR7c
JP8P17FFS9jQvTgRxGQ4+9dJIhMbiRco6v1LfIpcDTgfRO2notK4lzUcOEgehbabeqhnHzvAFKJZ
2dMBFJww08AnO6rEzRgwI79nl8unLKuyYfKpkMry1pw+sHcsfG4pnIIy6UyKL3QcnxxgyOWElXBo
Xppcfjc+AOg6heOLO0aqf4dSNQB9S55yot9GB7HtqbuTdenZF6QP3O+TxGUN4YoP084E+/7SRbMC
WfRTpFBqtdxOi8xZREHAwkaXOtaGwv7rsNF1ci0Kv8xY+uBQeqckX44F4aNmLutv1zlswAf/f6da
rGLZenit0sinQbPucltInvD89gDz0hqM6TqS7nmmDPbrAueC5MGT4oUrIRlziYj0lD5i9I6XQ3h7
r4ric1XhUc5If6mmoaqQ/NeQo7R1FV4/oInfKdV9KYblznCP3dUSEc2GNf/URrOi1lYHKEKYVAsP
HFoS7YQ1n7ZcbhzQLQYZgyEQDUTUOHIeEX80YqeSMz2wqWJNwAGCqmZo8Q/2yQZ2Q+fqCy3bP6wX
aeD23KYNAahSWM8Au8Q2a1o33YuJi31aUWhAR0XI6jZcYt2CG3O+e7gqae7Tmmsvpyo6mj8KFc8K
olT7uPvOxi/wNPk4XaRbDMM7ZzaSXU+tH/THV9hhJnEKu18DtLzoJ/62Fg9kMZzqvqeSLBUw+twR
3857lWB8nCshP7y9QTaxXid2t4ypXRYnTueJzmncUg2QbOLsC0prNvTPKTZZjgQgAo2HjP23+s0n
viN/vQgw+LHPKB6fw2riHEyO4R19/dakOI1yjzofIj1cTsZ/DGm/jUAhu6e5BsZyz9icG7jVTYtI
KSBq0qrvE0F/7LXPatPLhstlbOm3+ICR62L8Uf8lOK7KHDxy5ndakvKw1a5EI7YueEDv6FP1IUN4
yIg13ADZ+e3JltmCtVRiTi4jR6rc1FGHGWL0mdvf/mWu/FqRomv8wGtLm1iWfdYNnUv/yRtNxrn3
USAGIFNEPuPHQSa1CPJCT3cNYfqYlewGXaPgqGoiJuU4pK7t4WYWOGMIqfRtSaJQPkhi+nf8oZwY
6wNFXPNW2zG9CDD2nqBNuY16EbsMmdnQEmn28eCFR4yM8Qq/LwhLXY4ncBmClZLN8NFwnUKMxgK9
Pa+Gj/dLQjT0t4plSXwrGmrD0zK1/9SDMY3DGS9x5hc0lpInDv9EYRVpdU2hXET4sE3yWb4BoTJT
7gRvd/QH8hX8ujUFt8IZfdbLwB2m9SAkju3mzgJl7ju5DLs8dCWi/PkAUezckKK8yQsNtvUh+Fzj
VxpDtiqhlIshApyOU8/sBIbi1KtEjne332uXtvOBV/2vuYRFRrI0tj13zqretQhUc1ahiIJB8TSz
My2wLRcmvTYHDC3GkWPAfwuvayxru2F9UAzZ5b9iTwDEg5saVSEQQqJpFcxSEzgosP5XsJHGRDpe
keJvS5Xxl3xFwis/IaIA30KaqQIN4xwSU1MCWS7ChcgBu6ZwdNaQbqQpPH/98OoU0ktHuPOIUJHP
eS1BqqBjtWHnqJwqQC5S7pHBnY84udquWg+WT2R3vQSQXFd9IwJL9kDcDU78k2M6NB5CIesHAW5e
GNHnntZiqFk6+eqlhzfUuT9r/nnSW6m0SACCKt/moxF7npRgittRaNNrkCO1MYYWun7zRbwL0ZSr
dM1rtHi6vd9h9CqthAj6eTPDlIPss7fUSN+nsmNXBnNzkthMbL5/iGuqFpC6peGvbUUpbdsyMFfi
rHnhxfdDQjC8v4zC/1iPIBWMH6oL8aBBxj76MdJ/6nZ66JAjb8ZOAljH9k34HQk3OoZFhnBNh9g4
xdiFT4Ss4dezFxzJDqY6MzTv1Bk+HTFJVVRk8j+W7RpAh2Vo3zso7eRgq5HrxIBf68Z9PIS7TlVj
hzglnF/Kop/0Ha7dFc9vuDsSb3q0Z96BETmngYKbWv2HlQUqv32wFL9+Y0QfeVoBRLRf1HfY/2QO
LgmLxyVYjPzPkS97x8kVYIVdMXZ8WvWRcNOGkNwXmYDf8ExJZZSnxynvfeTPeu+hjA9LXmB1dM93
8SRwOeZqTMoU2NEEwJcHerR0bYKP8KEoqwbG6EVU+jEBp3+nfFqjzXUIx1MUqIKlIkdezPK1qyHh
FFMBBW6ErnWgS4+P1A7bXebL0ZY/MyR+y6gD4qfI28o1EseAnbhCFb7oqWFaad3uvdEVjUaXayEy
Bh4IXV2ZJf/ZrovDn5ptk/dxe5Ng99dDRfOpAw7Jcj/i7W2dz2dMA3hX5TY2Vdpo7CxlTpfLHMht
aeUb8mooKicuh1/v1cSQh/aRk+8Vk8JWoCBqfIumR4YRX033ytKw5uHm4L8l3oOWZFMvdQ0b4GXz
nJMdcnqeQtdQSBlkWxk8Dz7s67To1p+7F1tqkZku5GQPL1Sb9/ihMzOHMfDAuGd9t0e/WAMNKO9f
N/blDPMQ3WNyxvhiWg3YSWC/ZAzxWfcHnnTJ3yksp2G3Eflk3/puGVMP4Ipp85b7FRHDtLXQQVr/
XgQjv715YLVA0cHDCJ+bbHQDhM6ZwsT5/GDhVz3Xae1OMUYglgMn6RXShtdKvcla2GFLx8XWjS/V
/YAFaKB2egduMNRl5rLnFDt8tScP0VFJmDyL4Bez5E2/oTFrXclx/LvZJBzd/9h/yM57darEbB1I
J6VyiyJ2sewucHmJ3cd9Ttav0Q8iZEQLdjOH3iqOS+88/bWH9Kcqg+UDXaTHeV8uE1bvHDGfpz9s
gWu1rGtDoSgoHe+E88Fduk/G7Qt1hchC0MEdbVGHPm/qGDpdptpgtqNY3Z//sEeBj05nEFd2eAAE
EItina1gFLiuGK4mmTVMNb/mQcvrkTbli4rOnCfmXJ3DfkDjn/v7rFhVLfU5wt4KrW5mwG/et16U
HLVc40fmNg60xLVLNEn2SJMWSzsD7DmkSRW2ixXYCYqGwmoB8q5Oy+Q/U0a8gZA5x72xBsfrwdv2
HouZ4gx8eAXpigGVTW8HlD3vV6QRxhr8W00Qd84K238z5/z/UplVhILFXsNVXETtdeMHUyuFEjoB
mZ7KsA7mHUqXCCeBBvLY5dr591Ay/QuSHmH0DAEtTIYyrNxmgPzdtTRqrtts0J5hAOeZRVbljqOS
eBMPn3R24gkN+JGSe868Pg/7FiYn4td92DTjaSF6suEeV377drrvHWL91mpDoP4zWJbMvLhLhyk6
H2OG4a159G0O/7sJlV/+x+Ia8nW9MOl6Ma8LwQSH6peeXpscYCHKz/R1AtWAkOnblK61OQl39bsU
mMTSueXVZRdGLqoLh313fWbkAd8PKVvfHnX9wo5ByT65fEt4fD1lgNpgiHesQaQskYmYh0rc9nuw
pzPgew3XB/jZGX0OIGBhSWqWQYnvjorcFM60SruGwHNvfTPbzUvW07Ko5Yvjh5qWGYYf/H3SkJ6x
zHLqYcyScRfhtqmKrOmCfGe0EMXMvIA4D0gETPlOnYyqE+K9OH0JUMkKOjTjr3GMr+Ed+ytfz9Bg
apxkWAX+bzKyTqtA/jBFMR2DNPeswn8GVEJFqXFOU7Pp8CjCsbwJGfBr8JKsRscvB0Cm/dT4WTof
mzaNb74u/8Tba2jT86a4AfC3q0azxoKBzJso6qMGSCpaWTF947rtNNraq2zNayGFBDO+xx3XCy6P
avII+AVdSldZcHltmutT5ee6dEsk+fTwtR3gVsnn/RM8uDAtMDO3w+A3xVp3mdNA/Za7RukDRdIa
+vdf3Ezx1hMxKH+l3iUir/1YeCjLWHo/6BIb/l4khUQtE/hOS83Va1F+DYktm7x3E0JQE3g4jqSv
wzhtNhoy0NnER1ieh7BEQi5saESAolK4OgbKofHH3eXOADP5eI0OH5FCwW6c5CP8t9eU4AzKsW0o
tudjqYxJ/kLLnbAAbGftSuZDJyxyJ7CHICgS9Fp85+BAQBEku7R/OVLRmv1nbBQ8OS1L4V6vcNv6
/8q/CLFkntsE0yqNnUSstsSzLNyK50DeTyAhg4ehQGSx0EUVwTe50sUu0D4mgSHlrTp44p0xVEw2
9O7oEm8QPcP9MXJGfNbmugL8GpI+gjns5f1WGvyvWK+uGasS+EmzWQ21p15nm897344lO23zi6a4
kWa9U1BrNhCZfhGxwtTQnZ2Zck89C5WU3TK/L6i5ukyFtGk55yAM05E/In8VvURng270jIxi/1jN
JBRH5SZfOhssBCSkUjM8Yil7bZmRoxh7g4l5ytm/DAoMt/XoqdfKBEJNH48mujWZ7da5eAnrrqg3
KquOlvvneZERrpf2/EdSJJ7iLULaHUvTnBg8ZyuMammFmeGVsYOvtgr2YyAbUUe4xzwCHs3vQ/Tw
bCrj/mzdrtCGAYUcb8hon2Rt6kj9Ar0hEdWvtzaVaSCmzeKcXTfUNX4+uf8/CTFgPbcF1cHjG4G1
LegltKQCu6dNsY/3iBFQbhxnL6rccbWVQAh5x+LHG09orp1JousyIAujLX95GQrjglk8j3qO5zUu
iAM7wAnWCiyrv8Gkg4UE1/E5bVbg/3Mrbndl5ILs7FcrrZtvQDcEMMQpX+n/GrVfJqwN2rt+GiwU
Bq/zQJDLWC5d9aV4a1z8bVYoqTm+BkvJjNfSB6sTSdS5IS25m51YXfFcfKBD5sQ1hwcoDO1zMn6v
VVi9Rf6IWZ3hjejzSSiOx7ZRTkuKtpgu8GvEGRAhtJqfM82qRpwJtqXmTCyqpuQj53+e9+AVv4c1
Qvl1CLKYQxtiDMrMT7Dlpp4Vb3imNA5VQ18nu7YmzemznDcg11ALfyvcqEgnhtcpqtxTfPLz9iPf
mHTEigWuNAq/0m9vJwheAJDTXUdrzeQbkgLWuhowDZ03xyUfvXqCKlcFjehA3OOiJp1wHpqD4OHn
pqw0vq0yJ4hnOSYh7UZbpXHpl0Nr55KFStZ7MIDzIhORrhbBed22LIBtxBdOWTR2FZSg7eHVElAk
IMhPOcfVEbHR7/JhhH58Ll+Mfx9bMXTAZaNTWYZ/xWzCpZeK7x8Qwp8BKBFpa3i2qdGdg6ceY4uv
9+ETHKL4dm/cLUqJWKAbbRYS3E6H/vV92hER3i4KtM4y/CpjBcbUBMGAVydBQh7GCt44JOv6ZQO4
Edri+GW32Pw4Gv8o3CK/TL22rVH8x+dxR0g72kuVe9o6Oo5u5BnIJa64DA6NkfOCWLID5gYEvNsX
cMyzGhsnzW0fXaxi/xABOZIpVvttU0wPDbCexDNsvcTG921hj8cu9teYvxwT6CDsahCW6jt1G/L4
h5oolsqq7Vyk6wMmcK6QuXn5ABrgM/MfRUQWs9F7crnm/NkXyZw/i0o8IZx39c8eLNA5Vh+sJPmL
K4oVO1Bhj2sa+K3EiqWjyJ74544uy20LvL31VfTrZtU/U0I2scGQpDhzeoWfr+sqKBmG/Id9cYiX
DkxvtAynHf85mExT+7d0rugsXv7ElOSGrD9d2fPBzM5bxFAF3NYkyqaD7BOYQDX0HjnERXq5Mq5P
AvRQCO3S7hzR1hJtWiLWoDYYksDqpSS3KBk/yJeTyRReFbCrAXR/MEpxtFvO8S2ylnfqMX/J/U73
DSChg2xVFydMkvlKWyMNBqC6ZD9UWFSBeKxNTaaSMBCGRgsgWEFCMBGAI6qpZOaequ+02YhTViuW
TSNrSoqCBI52h9XusZWPdqE4aCQ+piGF7ldCP8d3M2k7LBkfDo7Xr3JDxjZsDRc/j67Hii5gvCHp
oH4YP1vIZKWpQ/sas1sKboWISzQF6+cpAeB/UyImcObbPDVVbntJdCRTLCQb7VnflQrrCgb44g68
DFDlGn83YZZGsoy9cLsTG86qrV5eK6bHD/F1X8CADd/ttdjt3doqcMjeNPDYDTczgjp9OYIYoSaY
YdgxvuKenpS1/hkQuA5jMwyuimJddnWgHIC2T2dMdtU=
`protect end_protected

