

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qyGsKXGf8tZLZ8MO/6NvK8t4R2uGW1SzmyF5tsX5CkXu0PSTBR9S/8/YKPbPyrujE/YTTc88Jf+O
eCpAsF0s0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SRiT9yJC5Uqpf7Myl6ffuoicyiy9OzLI7R2FKBd99DYnc/Ou/e6lORSzOmY3C18qI4YziTtHq0mG
9/kIiomSQZ3NJakbc4u/KKTf4sdd6wdIZ/mvgBltW+Q8Ap0+qgKaXNTzfHyJ2n7Ooz/Tn18T9nO5
QHjNL4UKVvlJ7EstP8k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0eEt2iDjsC9yJcLMh6QKornt3Qp9ep1c6xk+HK6mgFR5fi2UuV3P98/17Y8KyM03HpNkVLTMYss2
6Z1aPy67AzTy6N45W245PgeUG7yY+SedSieqIS0fIFxpZHOlQKRcnMJOLb1yLAb9v+eDvlWE0Bqt
DC6o+3ydVuNn1j9muuqkFFLx2pd7RIg2vU0FWhnTxY52dz4f6uUU2BhdZBrGtu+Cau9ea4vNs1fy
I/3T7fa71g9NdE+G2SXKnMppSb5dRZUuux8lx1aIs0mR64PH9XFHoeK1TPXj3zaE/Opgcz+NH9Sh
oyzibQaDQnD+c++ig6aTpqrU7EjJGQp/bZ1sqQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tf5mZezeOm+OIDtFXnbJOyEHGJlj2ZccsmnwTXc9Lf5eECAxNh05jBGLjHm14homsVnylEfeIkd0
FTR/x2Fa7arDaFRVeIpD76PsHPM4sIgsLzVKZSuDFI9mLQoEjwJzufLxVI1VLrwnnCVNXdnORJhm
IWzM4TmfF+Hx5JOlhkp6LgPD2qnWcpe7woFrqWuJiGRQIuUo4INaMhrQXXkoU+AIRMn8SYGlfbfM
BW1POo7+U3nnN5rZBheCXwp4IIczrHnxpJVCU4U/PKMVsPZpyo6Amt4Ih+tk7bJg6dcOiu0v5cfP
eNQSvIUysD3zNnoO2TasUMvjH92vgoaXcHg4cA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nQvzAt+9jXefqG/QM1RphU5FHai7OeU5Tn31wlHRRHVBwRxy/exmgCmhhWzEGkB9JfWIqx51ettM
u2pDBwcHTrlkKwA+W789dt4WREytRjmkJuAuOhovLRUn9KqFAPPWF61S+HHYBWBeHlxc665U/wg3
55wlrISl8SXBhOUGPVc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bZv/b3M4JYVaBF8S7ZBwGpYrwTNKc6COV6GslrDxCwO4aA1yELtJPTtkKILCmy8IFZM9BtktepAB
8Y/GfP5Zvkffm9OycUg9b444iEC1aylWo854JBsY7OuaJQ9c/C2cMgxojltmNWdx+t9dGUw0q/fP
QSMgjOp16ynE/6iche9QP3Rx9L1p06lw0r6noJ+cQYrK4L2b71emYTnIbR6Zrz4VmUphEvyZRVjj
yRTrT24i7xB/piWEVsAw9DXYWW9C+SgXnrMYe/yevzsro+mKydXQfmW2Dbmt3sY09vHSOMFXZaUe
TugvD5D6QFYttU0YQgutlIEfR7RhTMq7uSAZTg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CSOMXEp+WOvW5Htg+t0c+90atBozEim5hIf3+CSoYdTFFf+wWorqu4mRjDKnMNPuW0VRunrFbBdG
UpMF4K6THmtyXXwIrfVgO9FOmsaKczar1QzWtKCY0pX4UVdiewHwECMjPOr5jwWiqh9q99zvfSCz
XCkYrYqwNKAKI4PXNiBkS0EHsYL0dBSHV48coWMcPXBLrnB9FjLezyXelOQF8LUsbaCJru94RizS
mWbmsFngIlU3c8V5h4cSM51fiLwNFh+r/2AFm1N4ePzurikPGzsWqwEtvd1qTZn7jqg9BI0myU1Y
FxH2Krw+g37LCvEwNT03+jBCw/fNncwPmzHGww==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T9AUf0pY9IuRfLFQ5oO3C+Ff+7HAzyLO5g8IXVyHXsNpsYTaz+tuv31mc7s0mP+bJx4hMUQDQb8C
AEyc6KxMGDKG+0DBKifbVWvlgVuneVHYBy5vDyo2O6fVFQFig8abo7a81VIEFbTDgb4TKRy8/LZY
vdapPIZ1PO1kaTTU6Nku5fWv7YdlK9LCfVEP4uVZPpfNn79aZJmirhcE6rShAYJzcHp2d4fNp1US
X80+dNn6y4NmWWdCX+qRwvbW8B4S7N1i2JlW8ieISjF8kxvZVmEA72fJpAhF1R5m429tDLfth9hQ
lV79mE5RDnoga3gsIjQeqZWK9G2wADk0pQLm0Q==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
blWUaL3aLnYr92n7sNl022vF6ZGJmI4QFMppXGoWIdsoMky/XBFpyK7m3+RodQRO/HelByiysPp7
zQOkPXLiaVvUofzo9m2HyPWPVyJnz5TJZMHXT58n66T9/2AgTLGZGVXJ1SJh0gGqlkzYlYDNApIN
It5vEpLzMakHV9olDytQH2H/2bDfJapFSG5EG4BBJhFKPYPLz9axTzKH+NwCp34SetJ9IEwlcpkf
I4s6/jjLbiZtdgzqVcxuCm4r5rAxcNhqCWQyAbh0QF18n9oVY/iMOKVyOwGU8Bukrgm1EOqKJ5JQ
yaYm79jd9vAhZExjpacnSigTsiauARM2YOZ2Mw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74064)
`protect data_block
5Csz+xdE8S8OQBjRw0uTJta43x0jU6G4sBjNlXsNXyXzJehmN1BkYAWKxS0ppiaeGJ+e2hcssbxj
0lVHIZxQTbKqJkj9kYBSwqd/MR54kEbgyuWkUIY7j2dpwiDTGTmyx55xpym4rPNYe7uKvOzwlSt7
TEdNTmhxwDH7KUT/G1u/3s0tHTRyHcJKlIIHkhc+oUxui3V7xyXE//JlFscde+hU/EsaCEy10L+E
K+aoU+p17p3daBESS8x3EWQWlA1NhndjjJLfommOPyeI4hJjZF+2/8gGZ/8r/rzDwjlbvwMiYa+b
q7G41NQHC8QkVfCO6/cf3Jj1iY/mlAalDnnUl6zOUQQw0QJS4uqYtSzkvCOKM5YtooHYGka7J2xe
FGpU0xcqkwxT6EGP7EzSwBCBF/NgrtivVm2hnwjTRIpc2zAAF01gQdcnV09tVOmhaQKpo00c+i5i
Zi++XSQeNUZxUSUNLhzw26HbWC8ADtJCqC3Rc4unNZXCfzAxYnnvCy16n2My7l37TREzATM/3ZqH
mY8BnqyjHVyGHHONTFTIibH/d19F8NEk9MI8TqP+lB5CfukzNTHmN4+/5c069+QfVEEMDaLstDu5
np1aBraeRhFuZv6a+P3BdaKB3Wbf9m/9Z0pBWvPNBbXP1RM5bD1++gML5jAztJuUd4dWEfwzQf5D
SOTKRvOC2p6oDERG0dciN0w8X3Vp96dDlV1zpipGSX2hS5y3b3ul8NR46fqT49Trh4No4fvy30vC
RwZf+/euEBz5tzf0ZGgUvMnZPyM8oY8phofeoyXlu7Y2J9LfFvqOgk1eeHggcyMUaWBQQ371yN/y
VZB/NvEX1WtuRHwci8sywytcbNzlNukdHbxNQvPYcv59iFYqt/ch9jf7K5P68xR/79lCJ5gT+T5c
5Zygb4rC2LpTqnwRPn6Vd++ww8Ylwc6PT0VNI9MHADmRoOzZV6vIZJrHVrql7UJ6h4sACRqc9m6a
su3xjHKlGzywCF7mWy5k6gjMcIfHTFzzIIaItC3ZEyIJrywxmqorzn7FUeZjWIqNVqZXeRM5jNab
wyk5diIJYv9lYB2z2Aq0rMSDjGkuCE/bYmwgnXw4bgH5l7IUxJWc9tC8klN/nEdCPD4QyWfLy50r
/u2hN9nKKoOvwBwIZ7vILBOYcSf2vASJ3OMNC4L/eKlJ5HxmDEzBt03++oJYE9b/d4OUx6TVCss2
hmLwc3M5YxxSKaastbG3iuf90lR3CQwDMcuh+NNbNuXKea2ui6s13e9mHFQfQsz5x7N7jasyYwbw
TEg/2AXdnrWAVglGKPKjQ1iuuaXKJ9yyPwKBg8boRzkxZZVPBuwjK6qMvWQN1etNDvXF8oWAdHVZ
4ha/r9MkwrGrU3f4IRKw/dp7gyl9PJD22CnfBwhjOjEZZT3dRrpZqk6WiKYXB6BHf9MxOz62G0WM
bQ7RzdrNpD1JA2b1i1ycCCpAQFFigaX20n33alzI5v6FFEV/65b3uv4yit9bngxyJmtVzyg/w2pl
aon6xgaY0UYbXT94YPL4j4Lmp3mHfp4HPEWyyrIP9a0auEww3x5ElSLRHS7SdX/uq14EoUcJzoLv
p3uZGwmvKMDiQ8eTD2xC8T57rE/Z9WwwNTvHEXqjJdNYGd1j2xa3xmJxn2huEDhMLmZwBnqAbTEp
9vxVqjzqk8NDucatKePE94RHsUee8W18RniZOTMn1Gk7YvTYztTYy21+QaaEDThp74Ssv1eWxKyF
C/pdFnACRNmG0kbFrXwdJ9aAg6uysDFSn6C2wCH3gA6BSrZwfjXkl2Jksok5mpZDdk/G+2tbHBCR
e77x9D0C+WwsgYlmWYbiv79jn8CeGTPxGBFTXxIZRvy0ZaTWxbV57iCfxeDrin2gWh37BxuZVSPV
U9EPYWyIkCHuq+iU9G70kckx+pmGPIGFV5SB0Qj166ROu0qXc7EUOWMV7Kh2jEln2WzVAI+Zo7RV
wkfiZky6Is+VEr8ChqJSw+n1dBymVLx3pFVCV23crb3XKF6RJOV3w/wKCUCDWXRPymhgSflSHjom
O1iGdRZ8ZLCPhw7/ZxqNfYkMt8mUe/lE4JWY81308CL3Rms+/qIKbQo/TNQObslO9KSkDyu4Scuw
H7YwcX1QeK/fZm2Vs/t2iZhPOsk7jMNCDpeble4k/O/v7eSEkDhgixaY9gyJG8ELHwSl3adXqVgr
COgdQyC8ckEdevu8ij9JDrXZrV7lUccERGX7OBGWzQuPnsNajRX8i7zGsN+pYIUyujrE6woBguFc
t/TWQpRPbLdSr5HATpTUO0FFLB/1bRyJk8JfvUxlT4bZIJWappib1OKVYo8Bti1pdeQliyXuGEad
h/uzg3nlaKLD7Mi734SMlq/5aQ1MAAbzka1FQsr9yTUfEg0PxHnLfa8hTNSxBS39oZ8WFhxD8yQx
Gw2vTrYPW3SKMl8sitIlOtxQGyLZz5awv2+yAUe8PkC5PoVSHPd8yhbMcDJCY4uiDKF3Rx+1q5nK
JN5z4LKqHzq8dscE2L03wRVYbOXAGEqxBaP01G5JAjnNwlDwGFb6v+Ww7RO1agnxgBoTzstoScV6
DcXQVAzmd8p/zF55BkavBaDxoCSkgjLpCTUjoYHyJwE6HeCV7D19YSm66cpbBb9G4HSpTQpOWjya
SLRVelVupZRVePJahNW1XqpyeWslInehlfxBUO4Q2ETPeAI9lzLX7OtrH6b6o1eGf+dx+2zPoFsH
VTzUe/Bsbl6A583EqmDtu+98TfGb27c4frtMpEBYxzwuA4hFLX9pnpCbz2mfGTBH46tsYdQ51r7o
JJHDPGDYHmMrUMhiJM6MAqJIZVFdLs/WBVMWXXTYKUh9hheAQlaPlEX8HcBbgQhf6aDXoxJzaQUD
aSvUKL+A3LxAM2pW/F/fzj8fyHGulfVRsDnpBmhdEduGY5X4y4XtcP1Qfh7Zanat6ykGW3cZz7GN
yDnUkMi9MrH2wm1ipuj7T6hOC0mThGFIqspPT2BJhYLhKGOoyk3PDuLdWqAYJ+yPVglvLxzvtgZ6
XTFY4Y6ZO/8wD95QFdIPZiAkvQW1KRipnVcMmyogqRhNnZZ95Q7d1tcL6Ts8Eevz6UkSz1XgNRN5
Lvpp5gHPtmwLbZlsQYuIn51tmwlxloznMqExB69sftUnqHzZRSMaLHoxfgxINUoewhODpWW9RVkL
LPLpp2t+3M0w5QifF5gsxhoqKiYfVtQsjAsTySfzozbi+Q2KbwplBpinas5PoRz03jO7ssjM6RiQ
eyFrSPagPvMoHp10MESmw0G6v+z+U7qpL4e7JTiw/eERiMP1/Hl4EPfCftUX3mxjQKLgizOAblgs
pBf+3ZgafPljt9Af2Is/NcbF7uNmWzeBSRmSw3hRoqys6uU3umrN8eYmpRbYHPS655cEunawT6te
UfafI4ahTImYpaZpNdWhLjEkR4KCioTW+i4+2QLKhDzrciTJb3xZWsbn92NSEMuE9XiTmL6Y1yyF
qEo4vfs9iDISqskDatBGxvk2qR1TWCrR4piRasPd5GXClfpzKXPTVp9jqtl3ZNscboG1iv1LM6RO
gryah5/6wCoUECi7opGiUCXD03gLKzIqmimMAkxQyRITZwZKdjysdKVlWmRU7a8GXwCaYdOfJTNJ
J1HlHc8itKTAeDYqTfE448Xw7zg6RSiqT8AAjnRz8RLa4c8KRBcfdLhXu1nDZ8VttT8dkRzHN1RS
SJ6HPSNPmf0v13DDs0KBj3w0egFQqqOANTnm+foqqyLSw1bR0cXKUdASOGpNnBIOI2ESeozPOcEW
wpILM3XEslpuKImjbJo0s+LbKHM3AWjTuuqndhmqD/J05cwVxOF6jOwZsXkGExS1M3XGoPFTtXm6
b0g4i+NTbYbc1LXx37Eg8a9Q31gLWfLmrBZuLt3zZc0xCnlKLoZ8zwEha+9u/M/lQkRQ9Iv52WFQ
BQrYzm4bGlAGaFumvYEwscaAu3rrbBpZHrif7axCDgCPlTvWFx+XhQNwfBonnqbf49PeQfbDZ5us
tVi0FtJFXBnqH+6mQ0Vkb/c7hzL8xoNLV2KdxmkYNxw3OkFFODLKGXeaPIb1wvNS5Vp+gyzUIhcW
6AYvDJrlMUxlzi/YPWuf7w4BgSJbMC9DTh8ojDuXhYnwj3OrMZ5a4XT5NLwLJeO2Qhhv8L4uK64l
Q/6tE1FWuxG5wZb0vL9epa/fNvvTI56dYsYRE0QIvxi6Iw5gVZXSWtqlNU+QY4Jtf5rTjKRO3hyY
l+rakgtCVgyHkoa3WaJ2fMYL1hwdyseh8THOdmNfgRjJKO660U5xymneYMUCwb8YNtFV3qMl6+vv
UsywhVh8/HNvf/ZCf0dJvbSZ+ZSBQ2x5UXZ5xKpkHAHpohHP6GQYgJpJ80TNdleTybV9PpcwFsa0
8py1s0UIwfnh8Xy/i2tSSY73AG97iKfLf0d+6iVlrjTF5ytSVkOStA5gX5fUJnx/0TYJYAWDR66n
O6ZqnmOvUGxub6RjTZlWIyHiFpkrz9IIx9T5J/R+GO+9Pe+G9sfMaUTiNNB2eeLKOvXz2VOyO18j
7SCBA+wvd7gyb5OYzekKaXTgmk8tlqQIB+C9JI4X9vbJi83GaJzJOJQ/IBbVUO2bvNldvjMjCzZn
o1XueCfJ7okzvGAyt+zyBz5TeVg5v64QrvZ1XrPdvTNs0XIgZxK/hRQrnlXAbMLV8bWJ4IUvRG1f
RFZBfjAYEP907jDvtzjd0YKftNC1vFjzniZ8HYs9/CRQB9tmfKGyFYe5cwxzjCrqxSIHGtQtQCbL
Z4AD0GimQWum5CyqYVrYBt6VBEc1iUzUe1SLaIbvqvc9qv5jmx5LTNQ5qSAlJBP5wWUX6SqDNI99
nQmFufokOmhhlta1+TycB99ObUZhzXa0KPc2j6ndmj497n8ugHSq0S4BSb0WYnKuJbjSNdNvuarl
Oaqd2ojBFXgherOQdl+Vd2aYy3AfKBuikIUHKdapNuwtO6DWEl3xVL+BVDLdXM1BC5W3z6UKKZt+
H/adHOR3p2mIqfZsh4/uXy2h6EnHfwJPav9v1bp3+TMpg7RWFQM9QTNeRFlma+fZtbodiE4Sdrm8
KDSBC+IAKbxI/YucI2gAJuheg0QxeclqBSDfE0N/Hgz/sr6x/CSAC1Oho3vmdqUG/Rw7y7jMTUfm
pCDRSLI9k+/+yZubK3svADsw+4MI6j3yzqZyc7rHyUUPj+HjqbNUq5jISyeoe14XLzmqhjBw3vta
e9XbIHeDOnJiOOkomb3zz9UlDxZut1+TncsBwt/Nvy/6o67nbd5IQ3C7g8BLc+79xHPjAQHmQ/C3
JZBGQFtWrDpgDgqsBT8ZregFBZlafbelg81nym8iSrrTmxj2cGpo+kbTdEjuZzdLgYRyCtZhpbBF
vpWaIP9VHTko3OtBmdMkjCrkl2Bh9soSLDhO6E1MQPt2aM5ji0b7hepH55KWtnGln+Qhe2vA8Leb
UfU6tEiZxBUpQsCf/i+ca+WEm+CoeBjlwQetNnga8O8CeOgP77v1lyJY7398nVy9V+fExf/e0Uu7
9BaIIpEjgz4DRwCzcnEIVJGBts/lKXbFdXHCLvBvEeR6wcZ7D/O5sAJSUUT4YA0UnKBvQM6Y/uuk
VDnr7PCK4V3mY6dEGvGRyfO/ejG6oOliGYj5pDl8eu+BtQV7noz08taeyLHcLqqs/mUWvHtiXUWy
9XRtItsj8NFCwQCjKKLGZav+L71DVPkpNU5xFO6ZqV/W+K/7g8SboOIkPonJJSuCDOwcC09o54c0
x99RFJIj2zaywzcE8bqSgH2bYh6IQMcTmjkNQ1F5twniCuLXJ/3BiPKcCq+QDdajPOlF0RLXDnDC
WjnrMXkSu1b7ertB4A9XoalVX9txM3DuzsK/DpGmqq0K5oEu5oETt+CawronYPi/+QzJNgo0Cai7
OlvZQml+HWJl4JyDKMbsIQIcU3uYxX+ny30xgwleEMpInEezGZCh3BumyWqinIuL9fNgtvtK2smr
FqoYhobueMBC6yGKVQvurvQzNmLx6vW70FCKBA9tPDUlthY4JPLPvVuIW6Y+HOtft4unmjMj9THv
r86YsVijoKIun7gyTCxjqdMsMyeZazn9SONOsfkU4JMwZvGMsYxy+bVKNyBcDUtqOnV3c1sTCh+V
kF/GhDG8FXJK8w42ID4mX3eLSOIOY8jlIs/GWkhJ5/PWZVPF7mRmwucMFxNSNHZi91xHwvvgRvwO
FwBkALkbO8C/Sw1DTfh5YOMa85T92lqK5hXpgDRVCu9twxCqJ+la8LlbOwZ2HBtiZSxzo07i09pt
mcatAYMSfagLn/RtKU+RTDZqBpfQlkwtikkvknMVVHGOVnxSzRugNyTPvL9/oOqU6XunU61u+mVX
Dquk+jlA884D+9htkjVrxOcNmhhonumuq/QohfgBwdfpa2TMhTvtL9fmbI3UB0SvXY/tAQOQzSQk
wCWRfbd7X4D7+g+PsvCVQQea2L9HbIWUGuP/bWd/AH4T3mP7jhbQLEFxHgjqP0MYh1st2o11aCJV
p4mWqI1cX1X/ebejugTtQMgtaUAxzHtLV85ygxAsGcDeLys6RCd31k/gktt11wEUz8Uo3HHitjf1
SUuzDJxG6tMBkXpJTL8o3zerEubmNF3ENQfvtVtB/ZDBfD+l+H033yWhFWrs3+mSO4fpzLVQTTTJ
GtpqrDzFf2nO3uEJBHz73Vm3tunO2lK0K1CLa25r/wg/bdA18Ke1p81/RznvjkC4H18DIjxTl5wk
dU84T/1HwfR+3MzqqtsJyh0bwPWTm2gAWnamtRHW0+qIMqmjh0TTpKA797rvWfRblomusX7VPLh8
30GDkhNBWopphS6G9XSIs46ZJtWBRcLYDt4MYBUh5jyiVn2ITB1LoFfQ/T76Dw6cUqcoHvX/h8cE
bcwBP3JBkE9LThsiUQgoXQr72wGxY8h3Pv7BzVyQnO8vwtQ86e90qIUtF61sl3gg8Rv7Y3FkhDUi
eCrEmHh0hGMVGCRarE2tAQ6sD/kQi4rM8JZ0PfDI433KxUcb3POC3YRK3VXuE6CfA1bdqHPeClJU
buVLSO1NtlrRhvuNw10cPnd4nZzQnFDgK1KKZuFVuUik8BUUQmN9QdZparUFKjdIk6O855dyRain
NsiYM1G3WCyIcs5fR0uLj/Ptkz/HepQmMg4YbWaRT74a6wxXMUttVkOw4apJgNWOv4fgGni+2xmf
eQI6JxM5x6vxpsqupZOEnev+58IxNZJIhAdSSu8RHATFRb/OUd8V1GCJLceA3Myrg0FEgX27YHhM
C12/0IH4gqbQrkb3P1kadqvgg4szKysjqQswAeqfWwSjNvBRvyIU7rCQkriFHV5JN8/jVHcUSu2h
nGOthUuivLcnaSrfht7ycDe55Tta9CGlHhbQ0blevWaJpci/6YpA+jrDsaOo2Lap69ezKut4DDtC
YG9QYbXxSz2fpsBTfuQpk1DIsV4CXOpE0CrcvSH0M99kvTBrLLZpJNdLwzTj6iOhK5xci0oBUoP5
uZSsmNTtXiYjyNqFMrWMKApsGgFjHPeYmS0c1RVihTNieAXKy4phtX+Fre0JzATc4X7nwpfKoeGT
qiHArjjUFuReymSeERK3UL3mabXHjc75GowpA3CogkyaLP3si8SDp4LMQcdBt1LttlF8GdQBoZbP
Yk68aNN1kN2GLLcc/zNQbvKWM6DwiT4sK9CZ8SlxyI6nFbc86ZKIKa7KBuSZYEM4Is6FiA7YbqXW
DVo02w50ItwJAzqWuHeKJYXd49QOlli/MNcCXJHR6eGXOxcErauBrBAA3ZTEmBlGKMAIziD2L82Y
KUPn7++wyYJYHTBBbmeiTYVhURPB6qeCQloPZJPOcZVHDIIR9KeLYvuvu+i2BDuG5ra0PQBW9PCt
MvPKqRJyMxJc3HmeJYIGX97kInU/Dyj3IOpO9YUCMlV3w/6rVHecnSvj3AXe8/iP7lSvCDKuWVwu
4lbdiDP29eu21RwewiLcpGmnR63SLPsx0yY3MXxFRd14LjhgtnpFcfUMi98J+qLr+jzd88f8jxk4
ST9F/kCQd+CTWyea500sKyROVbmmVnNXT0wm88AwG4M2vVb28yzoxMlYR7ldpy9Qpd4CPkC8FUIj
hvGoEov4cbYx4M22pVKjvLoW9PobT2+RbtzDOBrCFKr3YVBj2VoiaK5urEvDpGuPg8cqQYAbs1m+
GSP3JOeVDSWbAuq1/tGNtDfa+hTGft3ANbevqFp8vvIRE1J+wwlaNZ0CMBuOUG3UEr6SrVNwblgu
Ck/Jof29N0KwV5GGfjkiGbiUEKfzSkt4RAGUTAYQrjlDCC0pkKUZBYpXseFNaLlEOKazgHyBzY7d
rI3H/vehh2LA6zNYLe9UBSdXV+m7Le7Jt/61Tpu9u0RcbGChmw60GPHisd7yAldl5sd2Kj/KWgeZ
vkWS0fN7fc9E1tG3KGoatX66d5ezVD0u985tF2OpxzqjGgjfDm/Dkl5G5ZCuQG+ej5unwta+4VG+
2+rPRQtJbZAuigObUpeav7lqBFl8POD78FXAA7Y6uhGFKCfN6qXpmD35blQOpuUR0ksx3mitOrJo
KfCjGcGKFuFWVrobwcZm8w7MANdKtiQ4KQXImeVSv6UEF8GTjoV1WLqkcdZh5aiRcc689R+7OijQ
bmKmzMK4nBbRxCYw5sai0i0OMG64lQiRPxC5nyv8SA7V2vlTmhm+mSC880SScpPL7NEzri7P/FpV
7dAqlAdP+M1Q7vIsk6an1Jhl1Bunu2jHRUo48XHSh3zKLP9vs/C0bBNtF0CuLahrGiXdBhXUt/iO
ypTm1EsvV9VfZGxh/JZOBfy5rp3R1Pc60ReoAjtMrxE8yIbkyNstu8Jrds+eP6OMInza4j56RXLf
lhB/r1w/9VRCexzH2tLgmzqhsIjykEu2ehZvURLns+OibxJA+p25GfW47VSRRm8UtqjlrLs2pD+s
DTYizrKUPOQ1KNpWjwFijGRSam0nKIaUSzajv8BV3p+uAFqBNvX1frk7plHs6ppaemZwLMFdEIF5
DSH21HqnRrsX8a2iL5n0j+/dnrj/KTAIpZSyqc0TSq30HeodHBaZdTh9AnN08W22kW+FMMnw6jr1
2X5owiQ6imUTAUBBeAH1o/98CuK5BmC7xMkix24OUi9HzbRtGrLo/9C23rjbT1fJSMotxOFsjuhl
jRQPfV/L2Zzs2akTYppOCxvhN3A1RNZktyaILbbOW5a9MqWoBXmmN3Ynec3Sl3O/9wye+X7A5JfD
2Mzot8xIDVVxHJmZ758sRlgm6xwybtHbNLU6ToUWzPpzxFQAVHS7VGSS4jigXsT35+hMOwxLHZXW
oY0GzP/Fjij13apEmdsCXGuOvtfitn7+8+ydIMYmGDnFQVq7JFZuvSSb/OYEOzBpU3MWB31+BDuV
lS6m9qv3XcIuolGg9xaE3vkO4PKIi7yz/ndUejaQEe0xBclZKvGaSVFouIH0Oq60pW3Cs4eYaUFQ
UbUf6QIRpZQ5ycIl5fuEp+aoJMANE8XnfsPmZ/PRrv0XwHQ3CAc9v4yck7wNSvWKDQcV1f8jQJua
Zk52ra/dmeiL6uKrklazGT3kJCQPURWMcpBN9pH/GTM1z2SbmyNgMaFtwBZxJj63nG0xcuciBajM
Qw7WHp8aKjZ/MTaKFP0UI2FwKaWpQoA5cRWPV9p1feYmhlhPP88ELbKpiHV3o7QdPTLiUhOysp1i
8Hp3A/KQYfknWkESYQf/LddhIJKGQsK2x1FnsgZlO/RAsQDcQCdtWlyq0W9QFS2GPPw6iPizxB2D
s3a8oIBvkJYxPuI5gXYKw99qMzjZ6aMlW5atiZjh7YwVmAArsizpAUlh4OFoUcaP4431rK9QR3uV
2RjcJDL0pDF8H/Ld9m6FrA+ErzC9SwZpuMrX/aMSB2gWGq7ZNUkpooHbxKEQOk7N2qfnALZAEOys
RU9kiwPO4+fZlW6489kdbfgqYcXtPk/jPrPBp4r6c9IWaS+uV/4KhFWyXZeWwiekW1LJtlfIu0AC
knsdSWuenbrMLT8DCw1UvR9SFZ/y1yrM1yZF6an23CwRj52oMstEXvfVel+zwbEgwV0vYWxjDoL1
VjXkRWlWqUq+kSBVXz4WuWqnf8pCLKmQ+Brw4tDrxrFYVkBJSUSae1+keP8ogQpfk8Tfm/PHYJx/
g+ZTGJpvKBU8D0Mld+AeiM6lkqB6Kvk1gh+smTMK4OWLGa4Yu4njLCdDnW+ZnoirMsoSQ5nrLIKH
w8/So21yIopmE1a9a1VbqqDlWbVrm8hAN1jWQXFdG1Pk96Qj7HskedTvkrZQ3yifKUn7vytAicuH
FYadRLm+RtikQbZSViWbzwmmrssQCkrYMxiBBvP1TZw3Z3b71EVFQrWStMCr4m4b06nTgbaCD2z8
QOjpkGZva1LUj5s89HCar7tYVSBiqSMzZTI5FtCwDcgBDBfJ8yGOV2zz9J+2ENRhTJ/9fQq9bomD
PmNgdFTBL0zSKXf92LqhJkaKPI80LhFj7qtRKQj55T5uCu9R2j6PcCqNhs8bcpKaoL3gJhAI8uq/
qqSkkTpubHlaSQBhyAfgXEuKU8TGs2kE7JYi48o/wLzeYIoUvwz5Swprgjp1wJqNHqKRDKmJibEV
zOK+4b31Syq3XLJjPN+TiNzm4hE1c1BqkYaz0V9UGa3tqn5fzrP8JrLtdaOsmvg65uZxTHbVBmJz
E7FKMPgnxV742VpUKr0VgJjOPltd96F1JZpFWVxUG2IprgdQmdQyZy4CENfVB+FfboRm7L7MmcQ9
iR7SVqp+1I3qxsR9kN9A/1A9TiBx6SklWu+oeOy0ScvhMhXeavjUC7a+XU6medecAl8ehvOVJDot
55Yd9sUtCsg2QrF16weXY7No5xUkOG/slb7rb4T5I/6MOkPvJUT3OP2vpjl40IdWr9CzqR7bnbrN
8IticNqlTxHFhsibLpetkrmVtX29Xk40BpZJU3G0QUcqoK27nHKdGujAnoKvRE/4lAgpXVbtgiSL
iDtzAJzoyJMxO8gFM2G+URULMVZ+tgmtCTNeJOFTQbqPz9UXTLzHYiGz7f6TosCycHhfWkPbOwCv
io3rtd2/HxD9VbyosIERBW9eScjPZ5x2APgwTXQ4LaP/Uquv0A/lyrC9L9ETPCfcwhm6tnS4BwEK
f+eq/DB7k2JLVpUXaNkms9i+Jm0i4cp+mJ+xY6ztTTVpIc6LMpJhCkkahFZ9v2mMkhankJfYT4jL
ITDNz/kcFnwapVg6JkeF9v+cFvIaFIwFPOGPjVxVSUAmntKrMpRTpDoMnfgOLWhvYJZcjQF/5M70
ct7+LAiJ6Vxy4Q4GPQaENs4YIo8SSHIDnQjPzj6QZ84Us8MTd/WcThQsacgEWg91nr0ABOxvUPeO
7vdNhB9Ftvqld/xF50X61HmNOohNGg0VzzoT3yqSNZkiU1BJkGhSMXcGgWQuE8gT4OjDIDatqVff
RUDdEJP0NgvvfyXT6NRBsriJ5Od5DOPWwmTqYNRFPTbo28BJFXBifpVj7stBF1CTfKu2/by+iFQJ
lXCqZcFPFzRVkITZX1A3FvDw1m0Lt/QVeH3g2nknbVNxgaO5sHMWtzAXcRPgiyjaeIMOwbgrFjV0
YwnJNSVoLmhI1ZPzr4WHSq4uFXprN+nwr+1jarGaReB4ZuiwQp+aU0dvQFgv5k/3oLQHDw/2GhKO
/rEv4dQC18eCMtVuEDBcmTVipNnn1spKvbHTot05g7sieht3cmyO8ubhN3c2hafCgnmPtbfzD01o
89HKTpeAuo4+p7wyesXwaTQ2LjiqhrYxbDRNJJS6zTYNCDDwbYiJoAccxAkSGieVZbOkeiBPou5C
NcCQD1fQuyLRs8GkfW4Ky+2O9CuCteB1jDii6BJuLQZWiGT20LaGTHMoIszKgczDFBOfFY8TJaKt
DI4RjBepf8cTiLLx7vyW/BwjUBoNWPF/pFdjXLG+q8TCVCUMKNkyFIkJKNpdF6l2METyaPHofYGx
qwVrm45MI/R4KtldQ1TF/aQWXhRg51uFfdWCZdpU2lCjdAOQRDQNzEmdeDm8oVDDsq27KpA6VpPg
XBPbbeRdF05kzUcV5b7syCfI0bsws3Eqba32qas2Dy1Zjrt/SQ+GazUhQG+Xnv7N/SvoWt5R2YJX
JYgIOdh8GZPJ1XF7iUoW4PReaCZbjZhuTEqw2xJBsXT1YaDFLHprKFabDf6gPo8qyb2REGeOa7o+
oYnW7FAzwjsMQlWDB5LZ5//aAKirYfgEJjheUQV5N7tUSEGG+LDT0hIZhbU6vsKfk5MZ2VgA691h
QO/Hw5+AirQfC4Xb5jUgcYCBWxmj3BJ7XP4Wu+4B/fIC2COmxAD82Ct6n71DWeN9JxVhG4Q/FZ5x
pMe6xsEC3ImO9MIjKbKtP9hRroIG9U/DlmELWNdz6L5W3+ipr4P7/hLNpItbrnFQfbpcY9a2LpIE
zHNjyt4V2jbqNm6pzwkBhkitSJ2/FXdzJqNr/8PwctdJQieRrSr8AFEaau8cPRsH7fFA5qG3OcJy
XiPhhxdB92Ql5zLmuHrgPwFxaCqFRPyM/0Pk+s9/W+qAgUIPdYgrwS0D4ThMC009/bKdB7cgeC5C
1KpvDZtOh+gCjE7gCS1tGYG5/la+nNTV1qCwY8LOmUyrJlCzKLHly4JrzhkGijCEm4jJyLDX2i7E
/dm1NpAX9rPsjw5v0s4+JXNsghizdcTY46ziqX0hJxLoe68Wepinu9BE6RxcYzKuBJZmxM7s3QBd
K7TiNTL3NA6W8zhEuIAAG72uTe0cSlwErTbqcPjd9ZLLd+AB7O0k6JV0wiGhEv7HlwvrryhAUYTR
f0b+vRn7J1NZvF6EMmHbI6VfOl/iQSddLeCopEkwmx/HQqNrMjtk1d58UDvbAU19Sm5rmuo1x8F2
QeNXDdABwyGBd4/7w+PeY9qg5jOVN1mOYGJerO8jpPOIvv7kAuj4wBXp6wxLKYv7kDEY79lAU6oM
WGb0biM220NdPOGd4pkjQXlTp89A38BBIpfb8f+x4T7KP5yENSpz4tIgwVNWdvpJkJeqG+elvzy1
ZEUdmeIjf9meoT7d+0Hsp0Nk3LbtjHxiAS70yXAYJM34opS71GuecFHdlmIp2Ob4WToDvYWfZ7CV
ALlKWljaRb3/wEhVnyUQ8rNN/h63+4JYJjM8Gj2+2gdMnfBlBw95FfFhncPUEn0Td+PFqbQ3BMeM
jbyvR1YBJbDjq6FHmM+o8xNJZ+qnTpVhId4FPbltywECen1mQKokv0QgdI113sm19HdyLSRumDWB
VqTYCd4ez1y6/KbV84QRhqtneb4kRxDfAJUUbxhuVhOmbCKHGJexcpDDhhHYUeOYROtqQSBKivpK
zUa0NKMZYxJCyBeZ/6HHCoa4nS9cMelf3Llf6rDPisFqJ03c6n7T2zGXdvK0X+ZbyFSRR/SyJzXf
IVGoqXIfP1FUJnEeJbRiw8bRitOR/E3FoWoWlYhZRB39mrLtdw44s1ZgmrJvatwR5Uf77zN3zjey
gDHhBL7/R0dY1IPsqwV4PSOhto1rmIxlwL9h28mmxtDBAKHyo+jvhxpRpuqQ7HxwVw39ht3hhuhO
8pcxeVxBW9AhKIhh93/cU0PUPh3pDHUcmBgK7M+yl0V0JgduDsD6hpeWfxU8SaBxRNkLPl6tXiB1
WIWVMYX7lg5PyKy0TIJ+ft9RceJkdPK5cQcIKvp0fDEnh/rnBsSSqYJsJV2K/UCY0hqTp2Eoj583
6DLaH11K0Zx680aeZrzKSEBFBZtvkQ0WY/t/ifZcdQw9P3OoHiCOO/hF7RC4HklTMhdDBDfge0Td
QOLL4Bnsj0xxCTLHpOUqGFJeAycBqoRC0xeCO1nUJH7+Es7nig7WxuImm5kS3RRPPuRDI/+TblUz
JucNwQu63nkVWRP5SCtZxD5iFE6rqd1TMnAtNeg5p/DCZJBnslmAvVdJiO1bHSqzPlICJzJkytd5
t5fqP6BQ+lYtGmIjn8riFV5/YEsrLwgglnT6yWyOcQ6AeTXperAyqpSmVdy3b+e2SGQTSPWyJmOD
clyp5g2zhkJ/hb4fYX95Gp8L5yVa0OZLvhghB83vith56PbNEcSR8LbLg5oDhq7DnMe7qL/ZVuX0
+igTosiRp/ulanJwKtcsl8ucXslaQnNbl2XHWTRB0Ag5dl1AHaQHFax8O04jkIZh1+72pG8H7mxK
mI+RIWNjyG/Fs7bYOWe2YftJq270dZq/9TBO4kdcRRPGH5PSe5jdgpMNC4u5aJ+MsA5/NTEHNiVU
qp8ChWT3fEYmyKxGjDzaadOBEAEgZdOAzed1A384KgkRbmFWhjRVQEsfXPiSmBswh0xZ8lOKCpNg
/Vq21la7ERvmfhpcbdzwewtTgNnnMjoO5UJvLy67vp8euM0CeMXplXdAE3rpGP9kc+EIVUYoFRV5
i8kIRz2hnkUjZK7WX8V06XEaNmFh/GDKROY8V3pFarRjOW8SL1ob8MrT6nElaPUEITeA0Cp5XYBM
Ju3HtnU92BKlZK5Dynsyl1ugr9vK6op2kMeM5kP9zS6GpjNhmNoQO8KRjyhxkGaIyFaplban2g92
KeTotNQGVX1GED0iYJXlwq+H77oX1JjPseT8JsVajFoldhkyoMoMNkRI9451VIs/SiKq7F6gjhcA
lFxla3oMkwQ3tgxqn/WKWmJmdOekXHh+KWrff28+UIWKbDJu+LEY8sNihBCENOjpwCvxFzR0Of5n
c/X0OvNpMYUSXfblrVUHCMcvl0R3GL1TDbDmlbBskOebXfLKdBkVZH2DzYhqb6ivBGoKLRy/vz7u
YremcgZ1g7e5YcJj1CkpQlYldRs3oWblJuHHMXw4kGE2T0n47k1Rq//JgPB1xGnE2Kwe5zkNg+8M
bE0+ikv9wVfimjOW/Eb5GyoX+DTxFMVTHWKV0sC2btsb8HojO3H2edx+BtiEHUzVHgPDQo4OP5bY
MaYQlGE8q2N8v/VI8jzpzHlvKkWxpYK5VS0VwoLuyKYjZCcWS7AkEzZqebL7h/ddbf8CyOQC/e3o
NBP+zukdPy1eAlVHTexHkql9bEIehsnsH2dQN3gCwlAMQ0Z/E2oHS8Fm4hbYivUMZ3e/m5wIY3bH
VWnPiZhR8slkD4BO6IhSbKtQm+pwLXEAJtfpFXNQx1o4tuSHQrIGr6zcZcuEK5Np2+Tkq7xT/n7u
EI6XEa6rG57cQ32aOUCiBNx2HFUE1GNaundmubwbzjvWxZuiLULf4EiTWKJSfQU5GKH2i81vSfde
NZInJk0GWgghGTlZY8ibEdnMhh1Qh8CfkyP7cwRWGhqgNIAlnzdbU+V8WRriUuAxX7tszPjn6fNE
poSejQ2e2TlGY1Ke4A5chYVZiFPpo3yoCWSWbjbwfqGInQOKT2yzkiCSXsimCRNpF3yTSD6tw1lM
/yTSdlg/tBShlgOxomWYjL0ZEwsKry6IYGXcZNslGLHvy4GEFsrR5V255EcxjoVILUF89oDCmR8a
9aNHqcDV6h/jKA0Xo0ucH9P4sVg6lBR7LrZAvgkEvF3NmeLDjHY4bml7J6s7ykkBYFJ0D86nLGFy
QhaXtMOMu+KWuLaAiT9we2WOgzzsqqNoJuJf2Y0jzblXZSGOcaV2exonYZS52zCgCRpzI9g5QwGE
Mt2zwmhFcSBCuEPMZ0GnmvrtABpzCMmrTzv3Eq6ucJx63Im6K+BleB5KbULaomqnr1VJEsVbgvbQ
475GZvtNPNhTJ0WXogQkd0HOyPesYi5WWX2vkeqooJOyGrsPG8/kJrLHvZPZiGxMfhmofClXuhhG
bf5CboZu3tN14tYMlakFoeDgBkNJ6MSVctrGpy7+P8n8SfuQfRKPmBzPqqGFGcFnF/bS9jkipiuA
x/q4bf11B1EHX12VP5xO4pCjbD7ftVD5qBOu/6CGlfqRfk/jh7a6IRluLAf2iDH12xT1yT7pcSQH
Bu6c+ued51KRHcjoFRqEAqMKn4g6JYD3sr3os2U7T+vln9qYnrSIVgMO8aGoWAOHimmrBg+GbCeR
O2Y/ZIeOuVVpe7efSP9AMG7LKEieFnFP8poyQ6WwWSahtPYinb2BS9z7gdeOmjsxzBINKVtuwbr3
Q1KeMO+72nUv0Fffy8+posTY1L/ykxtV1qxmKKSwnMRKgP/x2if9d0HPRIu8r6U6Jh/ovlA+wyc4
LaSrlBoW9SsUO8RJEBHPP6jKxyqm6n5xqfdoUDv8Qi3hS9zVTvyFHQATKoERpTbxf4k1renICz0Z
Dn1obwbS89m09CNG/cymnO8QOq4ZufBYU+1NI7aPU3JOeUM5qQRCYdP8F+xeeCZkxbDCYHTFz4cd
jGZeY+wUBU2IDKAAuza9XoLSQps3MOLU8ChPofi19A4Kz1q2D1CwsKurEw8TJGFrrodNRxqXZYXf
s1rbZDLxIqWzjDW890BB3sJYF3sK+6K/FEtYbQnukODMNHaGDRk7kSnf0QIypNUshvY7Nc5Ww7fA
RokU6GWHOwsDYdcDqLb10OkZeWNvHGps93Z2SIrW+AW7gTcA5h5yLcIWF84N6vw0yWQWYsfcYlrZ
yA8MZluZYa+Et7CC8X+Rmr6ghSrtj4bCTc14ktBZw9mQBuyc6u2Cs/TEynxaPyOZ5c5kAZst5ih/
sKEXnA+cFWBfFdPADontVGXeYJjBm1N8slcekVOQuV+MiNSAOvnOnhdI2c+q/RtpCxfBmoQZmhs/
0/RKhcZu6I432GHg+WJYTMVeRqFVjc9YwKDhHwDtDnoiEeb9+tBXdGoQD9d6Cw0JJ/S4QhiC7KL0
zykc4QOPEs2iCWQmw6BlWe+kRROOlq5qNzquI7romtgm8577yYP6OU8sWXKBVpPzCLq8WLELL+1v
La8Bna3GBVFy3hrI7eNkwbZ1+kM4R9lYap/jWsq/fzQCPEqBMX6tVCO7Gxy0joK4O7jASZ9gFFj7
7huLLbYgxdmvpxoqLFQJBRWMROy9MQN2/nYuPeGCfNHEVVEZUTYsvg/4eTehIw5Hb5poSOs3SuML
bwpxhcvDBlgMRwL90M4dx8k6Db3bL6xOD9TvZopHbG/7JBWDSyRv164hnLFpUxrQBarKX/XrqKiZ
1q5tcbN0I+Y512Fckn6nwMNGk0uzpKcznMKJoubSKESDfbo4Ug9ZSag9D3txP8LDk1C+1Oi45AN1
6uyEjoJVrZtP8Sxebict/nxD27ysrYEdk7BX8hwckpT/sXslVT0BK7+63dfwtEtk9phHgDPR+odg
ZOqX/hVddrCvyrRJ5nVLCM3Pot3MXEHXJVujVlES6zBNv8CJc+KpoaOR9FwKawmdk36/mFBOBkfe
jdkpSI8OS7j0TLzVvICYn8EQX87dH6cIaOywFx1oRSpGgNPs0InJl/IrBLWOMsRa0FOO3qWCT0Bu
V9vhbv+V1RECouJR2LITSMpX0egqkkyTSTO7YOUjs4PxuDmj8nNdY7QOZszf+AzYn2oPkX2LXnjF
woTPCajTiYv9itAn4zvO06gM+3ZrLVvenU31g3x5DqEmaMPvlU+18FxF+x37A1oEGJAgONJK0IDt
/u52RoDAdKEikffyY2317jWM/l/YhtDh8mj5wV1BW8rpldi+c3fhK/jlE0abGWw5u/29mKCrvqsT
Quvwc0txsE5mHEZFQskZn/C3QGNDoLeqld6QHBHjp8ns0YBgw4xBoMmPRUMFzVxH+gNZrTONSCYB
jZW00JSlV6QIMNdNp3hwtaR1cw8fGWQoVxXlLiH2diDDI/Tg+qGE2arPt/PAugau9GUtc7ReGeS2
DrwK/leANe6M3czMP/6deZ14XoxxZEX6orsHvLi+ZS/5pcXgtMw/gqBDd4ROWBHBq3skltAZYIHG
54H5qZ8v6X50f0Nt1o7TqVnmhIQ71WFD/gzuwiKKIGfRBAhk8DZ6cBN4LRbh5nLql/fYlVfHdx13
KnqnpZykeRy0uRph6seFbxmtF0sBAQY+S3FqVbZpRYFJ5dt2DStTiYzBqiEWeBSxRsvwOqAasa8a
SNOGlqyN9qntu91GveH08CKNT3I1ObAch63sGHlE8QqECne9rHqDi2ccJamHmdkEKfxfdY9cEEn9
fHk3gZzxHehIMUIUdcwsN5SCtQeys5BlMeIIBEPLfiRH3YMcs+nBDk0TW9PYKKzz3Na5Xw4CfT3u
8GcYvMI0HmxDZy9G4R2YVMn+L9C3meMNnRSAhxcDOJjdIi62mFw+dhFfOP2zS+ZohLS/dnL75Fgy
L60G30FWjW5wJqpe2lCXBUMu28/UzCGSfUTetC16tToT/dAlzDbbfU2Ux818clSlk8Rx1w6GtHvI
k1XTiltbBE7l5FwgJ6rh3k2KxTzkveuSIM9uT7PunMs/lwvGmaK9v89JcJ0NVyqDkIriYpfHi4xI
ookM/ObKK9xWC3dQ5pyrFJBtyM6ov/+CfDaiJXehYKO4FN9tcWosnIt5b8OtZxQq4bn6dJSVehfk
rbymZA6BKTA8iliQ/yzoTNZrJTkxoOx22LPOK6etedSUIIkdoIa7QVDBtKddLLZFATmRa9sHEz1h
RnBexWZtGE2wOY3on8HT9GsZET9XSFa1NISmRSqNmvs3GBv6LQ5ofHk/IHxf0WMexfm45yle6MJr
gwsheCSmhbZiPlgu0Mr0i9TOl7GlYlgGga2jiz9WCJS2C/anP6Rlbh4NgjBgak0jMBoNQ8rIdavY
ebOCzcDTZTiOMEDLrDEKFdQSNyZb3icjS5U+BtiuWtM0y3dDb3OqoW+Ao+Rux3In0PHgExABilNc
EqtzdntBcV9CGj1Yhhre0knNSuvia+dz0ZRHpcSzLPaGf2+9MRKvUcTj6Xs9tjtlAUMSJ70kIQtt
0rOoYbatZADLheICtaWJJ8DUvId8aUI1GMIMhZw8IqOnsY0cPzTpJH8uz58vHa4MEjjF+VdRB5As
Xf0NQuAF8IhOafI9RHNFncPvtcZyHXK+0REXxafz6gg2iDj0DwU4juTTgpjo4op2DzzOxBmVbiVW
s0MwRtgk0wVzlleFC0mk7PMSNlzqcxub0nqrkAw1mwwPmTLeiJbDf3lMbGXPEXIs2XdcTe5KbEtS
DOIaxuIoK3bNbu/yFD3jMV6/BJsZx3FzCQpkmt0GPM64HTyK2NMtWCASRcYs+obyaseTcujfCIuB
dRNOEosbu7GnRLEZ+qiMEJPPoBeA2XMVmNPPP5JMuxRM9uszkQoCJMiyG00gOUAPfupHuR+aCPFa
Bi9aBwXi1ARZSbG2K6jDFs31hUS1SeNB5U+cgn7+VdPe2rYo8yEjsaBP7LWcOE4ts6WZa38ioNBv
LzNa5CO4x222yQ2dmzccZX6A5t61Y87n5WS6AXzzsvckLSjUdTqqrCez4v/GlBhNXPTPLvHjnfE2
Fx3cl0NwrKhJM3tVnKhtVomqkmfkOpEjS5SCHIHcyKRn1JL07Ln03GGCyqyx1PErdfBHpAeRng2D
kzuWUTvYZ5AEo1BkoWGr3fc5q4XP7HWc64NKLWy1iiHg/bTJ0JzzT4rH3sC/Xf2YcBC2z6UhMlKf
DCDITu/0ebMJmBbM9d7yY7v2viX37/hbJb/BFIG+ckrEFKFMElL03kK4qLNq1SLjq4ZF3B8l/jMB
fvCFzmGHdS9uL5cQDvhaugznR5XZndsSQDIOwF3Khxqm1KGG0mBWkfdxSrqxd+IsDcYVYoNePBEI
+oQ7uCHLa94z8uvF7GjcT1rq5ZlflB2quhNrnvQuapnkbxuHqD4cz0a3u7YBwiUjwCqDQUboaeSY
s9CEPkolLqLlgpR7u2hm3liHKOXhdYb8OQMSupodQiIBufFGoQEX9ze212D2txDgpQ1+D2cRpguc
wg0Vn3PtKP7iup8dkDqbYDbrrD+Fx8v9ZY/mARl1AdnseSOqGv6DjkHYMyjNiiY3xRUq/Sg8TpJz
S24+WJz1wqqxAQaI7bzs88rjCJl+aAdbHbTSbL8mnc7OsUr4d+WMcaol2jEG5gAM3s7xyIG44Agu
zHvx5OXsGLmog8XDrhI+0soYM+09ZK29DuBOsulLsUGS0LaeReoIh7U78Uro8xCFOR4s0ybXn9ZI
huGoDUYKCB0xoJJegWow0tPS1yMeMFvZclYS9bz4LvqybU210LDQPaSf6X5nNjCRjmIJFk+cF6cg
xSClfchi517REf+ny0eq4zFhYYqRukl/RQmozGhOJxO0TpPf8H4C4K7QrpmiDeJmCdrPU6iDSHGP
khFURdmLcQwn9zEpXUnxKWf5YQzlw8IE7CxnPIlLr9OgxBwYzEqdu4w2gOwdEVHdqlyAGoILwHcA
0rtW48a4qkqq5iJRCw+2pF/XY+LnHNwdGVwZzuX7lxp8/hh1+XfGpat+9XOuSFUYFcA97SLtufeR
Vw8OOxbINzDKkvmQ44saej+s7MICzatVspSsvNtawJKjYY1bEa3HDNrZ1yqJc7mJ3dBN3xJTfKC4
DN2XByY7IUyYD+Oyilug0lxlVo4fRdkNPVXMJwofQsWAza3rOkb3wCUDJ/CsK1emwZ9SGR/DKQas
pQI0MaCEWeakSYP+Q5PcIyTIVFVNIFrL9lNxp9AVTMAk/9dbFsrvKM1hPwFOCuEKENOSjNfHGDLv
w4JURmK1l3x7tzXt3yNUojOirnMIf9EWJAlGwegqPLkE2zPiZdohen7ZMTlW7FZQkoCuRZiH6IG5
ImeUcLo8NKdPxel8sEMW7+zue99Tyga7DRKtroAjtvSaDZ0aUcExi2fsCpzFL4leUQVF1m60KSv2
ZM+yzhRzK4K229JHgA+iJHy4b5i4yHlX2aJ9elCUIfpGXj3he9+VfU6iXq387bd95C8ZdPVuFpVV
ysXie1ZFLG1K4EZNFAo4R1ht5cPFYqyMZ7yJR4cXk7aBjGJVcb6ImyIn1d4dSnRaQavaScEDozp7
1WpqTT12u2vbiHfQWDdnmtw3Q2KzwRRtFi3xaOdZutxMq0sX5cKmR7K/imsSslt0B5me+G2KnSdT
I6BJxiZFmagDn8B+A5WvCd7WpgP6lXoMypXNmnekiNDxDtVc+apWd4fhzsQrgVnj5pCLSy1X0i1e
jaEAMDleJaAn1oKmCLqQezx8thFmtz28P1OrhPzv4QOrGQMy+AUgwdTXN6nWuccCYg4SZc0YsZZy
dhoWGJ5fMURV4f/bueYP4S11xsHikafOvKeqFQMsjnj5q1pRck+AjjzgucttMe2lfcPsccfSOOFI
ReLI7imGz/jzlqDXceOp9G6zbtODAsuwaShWOQmIpRY3mVtqv7kn7HUD7BfDp3ASdPch/M1/BdQF
fR3OzDEyxifKL/efM1iZLOxek8d4L3JvbBDdZBcyPV6N+AQLJHb6+OtsC+PIxIEpfCm4rmD83AQK
iegKXB5CcelZTiq+AuVSVmXcr2om0aJ6y4x7I9gEtbpbwKjb6i20h5tP+R8pp5V1h7nNrZ9ui2d/
GxO1dwDk3/tdZAEp/+wUW8+xY4+vM0MR1WJK8rnR3Pzs3xTlEkKhl3iUlCeHnyrSE7qh8FMXAnXP
MGxx2BQTe9tCnjJhaOV0fN9mU9pT8K2n31A/5QocQxnJ7QcFT0brtvHKukfUvwUEkYzMbDuCBF34
I/4VluPVqCF2HlV0PzqysT8DGCrK868NuVDQ5qDYqDjw5XSN0JziD8sqImkpPAOsIMB1evcR0tKM
KgNxiP1JFJ72NIz2PbcND0/ADZd0gVeWOY1SQbg5Jog47TaPKMRf8cMXfRXAts9reQY9Q6AyATRR
OXPmhpCya9iaCsGBAPV4HY1Y+AxGBoCFE/O/o0pOlp+WPeC7KtU3Pf1Ql2+ac7+56lbWxfWo/CDb
sOlpR5pRhFmxteYfyjPfd/XJcqrS36tiOF2qU3RpZV5iurS3+HxXC59578/OQCFKQ6sn2PnOc9Iy
+/R3cr+qyvRICYMLQwLDbnVBFDMIsYPd5FtjMv5a9Zl1HiECfxiZNcRCmAYAE4Ukz704qZk/4ehI
VFgLcjz5OULzbqZFngZKFHxpa8oU4INtWVcJ1BWvX9MJgiS2zgvryYdD4LtP9smDB1/XbX9k9Zmf
NEpXCbbyPBwFmMYVKBh+hcWrQdxAthSvI7SkyFWVoRxQoCyOTy4YMUmpFJAJaNxu3DKCQDknlVg5
nwgX6yG1F9LwxXx4/0RiS1qtl0upMeElSELwcS7s/XXMNuMyadGQZp/MeMy29BnN/O/A5utprDLk
QOHY/umQl2surAR8BW+Yhb4Xt+FzUw4ZSSY+dV7vY/q8G0Dzozb7FOI+ttD0lOdiXUZEoZThMn3t
j1+uvLuZ7Z9wdaSWXXTr7NEEbV/7dJI3nybZryIPPu6yZYdVluIxasEOXfqZGqnpksgsfNA1y2FC
nYKxdy4sdcZpvBbFep4Qy/o3sJorejeeyqg4MljQgAruL0AwzAC8MIQ7NzWltdhPRupBhg8iN8Wa
nbFv8pqaMXhuXbu2nlU/0D9wXZcoIHjmdOfqyXX+Omk++XyPfqV81us752rcn+oT8mHxj48kCWjO
Vx5363hOEjhQXdcQlsrXXO6EhXaj56oX2jYOne0IfFPewEYAA02ljt/Pe1u6RVmBycIoWMt9NVI0
SkA14VQJoHSK5gfvG+9FrTlSNbaEqhrNByUKcQqf9X2rvruaI4nE03EzWwRABnOt/kcjVImX3pcW
UAFfGDO2SySvQzIOt/o5Ys15v4azaM6pEkbl2TLBsIcZ+S+A6ANEz5LBXFpPy45vs9p+h7q6PB4Z
wTTg9mTjMc8k++y1CApL+jj/h4DA63ZE5Zt6FcK8gSJfBCrAf0oNHao2VgR0PEuzTK2yzxBAQGfv
zNUwab+TRHqLf4VgPReu7K4VLUw3ZvIS/Ei0Y5sRK0STYV0w9snLLjeUL9JwN082VKNWh5jqT/Mk
KZzJEmXZF9/THuFHQqemyhyX2XdKbjezIZFSPkuhh3QrGpIBQ3vdMUI3ZCatxET8MPoSOkuLyfSD
PBnAKtCGuIUTgrbYsy2SmErdLznMC1ndQGFl+PQbSUV8YSp1yD5kK5uDIe12A411XnERqTMoN0Ro
7T8EBBiDUEumdnvf3ue3We/LwBQgxu2MMGx3OvWwRX0qIjgATC2vLW5aERaJkagGk6bQ6wnN9ANe
eRZvWenYrVacskRyFIxr7VJZeszSGUAFWsBH9ikPqYq/vM2jDaAfPtCBGQK564MGAJFq+D6C0Grp
VS0qH7ulf3TJdTh8k6ETurr4g+PsvmyjxvORIWdJGhNsTWi5J6nAWxWY0tP60y07uLi3rt+eNiU2
zvfOMPo80df2CCDI2Knldib0XFXiE+ToWIyhGQF8myTYZ+yni5C9gt5/XtDY12rtE4y/KCHU5ESp
Vfcvet6E5OJ6GITyNDpzq0Mgf17z1+zVbOSr3g4opJJI26OHEd88WmRuZX4nuKa5EScHbOJAn0Y5
OMghB90PYAlX4iF1Z1MAkAwZncd+db45ANnjFjvfo/QVfLSoPxiQp2Kf0G0QHtvuiddjBzAuTRhJ
kbAVi42VGN0tS4eaXZiVZWvoAgTgEs+fHVlOIzOc6WUz6+lwHMdclaC1k6h96uar+EFepNi3wP/Q
uTlk3uObo07jqO8GISLblP4GbAKlaOpu1H072gcsqknxXJZphOAvs7XHd4JhXqK9QjewqC7QfAfn
gWY6a6NqkZUTaSjQ7f5viGHyACIwxyzBE0/UM/aBdrbaiAtL5sxUjLz9ieSS6ql2rcUP80QPkls1
FCiluO2bUj+wDs1wdTXzqRJv/PCfaUIR5cBWT0HbNptPE1NFbEHozLkhZk41tEHPHQ+kAm50Y8iw
xu8QxS5W5xm0G7MHmg0A6NUdk9J3uSefzP9qZ34vegkmS2V2K3MisZpgvQ+mz/85Dyg/bXNNE7hZ
BfZn78lTd6wwXXUbTxmprIXERdE5e8m/uLhkF8fH5nYkYLfKBN1KzvO6dzOufm413KY+GewEqCTq
WhhRcV303VVTIrrVZ6k3gJNpIyIBjumfk6TGoC99R0bNVUzwfLcfBlfEOD4BY4a/pMl7Ik3y5zbO
c1HMgVHIMTlUkWosn1ll8nLTEkMF9donwfJ4zkRUqp31/etDUcL3PVhtwOnKgatARuVvDtSbfLz0
H3nssggeWTCD0dvm6V9TTePsaTpRxfWObH5wotF/tLHZrDCvVFiV7PACi2HO1z7yA6LftyvY2yMV
IJVgUX/AbzxgaooDTjuQ0Lo2DKFBSDcSviDnJyFnVPGwG3hZqV2UEU0/BCTInbdT41FKDMurjBYK
AZyo0bpvWjauP+af0MXmG3fXMgxUgbnTZnPhrlMRH86RSz8ySKEpFQgsCjhD9kp3egW1q3wsH8vD
AlZZJTuV/RhMeIqL2F3WyKdQcCTIyfJ13hUArJyqNfX8t5IwT7yFcQRldNateM90WuBcudfzWrUm
5luE6vYGx7e/7iPZUKjwJo7Zas593f8WBQvSnoXwqhGIEVL0LAAMkom/7defOaz3CoNoT6C7EzH0
HCI0IpJFzFBfsbvRaU8OfTsXhgTAzC9kqFA7+nBBA6VcjxlaF4E4XRJ81YflfAcwA7PqVn4HQKEa
y+H4E1YjQV+GqBAWD//uGNusOs+49Sz3wDNoYYsDt3AfFiYWR/XXcu/3lcY3DrD8HRWFmvxzq17F
mcEK1CKFL+0t3WeRCnyYjE3rnKtNYINhlUndV4/jT0QH00PsG2WeAxzUm3smgmY0yIclSch6n+kd
SvI2Be0bD6OJZrlAgr4UQWqmMjsWJ0BvXUhLvYunRj7unvV0IzesYddz41ZIxCSWcANUYJm9zrPi
on4XXO7c9vsU/+53t+VwaBYthQ0Tv7Km/rBxRMeOs/9P6Hc25DWzMVuQgIPziRf6gKdzn2+Jbr7U
8y7Clr/Juy3TNZ9adW/4KPzhbKZQxW3AEfEK9yU7VYz1VV3Hvlx2pF7jpZ9NilFnxf96zVTP6eqh
FM4IzKndm0XKqNUBfT+YK46Cf2sFtazxV3PGAHs+d5EM8BX9KxhYfkUlUo2IKqLFhoPTdjkUsVMf
Q6Mm7tqOcsW80bJmaKIPVu23B2LI6s4T6Lp2W7rlFwkK4Z7StfmbFel5czTMSAeAkBOyr8jNjtUK
mFVvBdBQ8uEZpD3QyQ267sY37G4RD8wEWn3f/lhlLE7ukO57HuF7iwooNyCD/ZZ2sfOwRwL30YIl
eusRjNpf3gLhEbySGFZw1KOcerMs5ZNIF4VO7ozrqCnxY+zxqizjuupow2ZfZgDqmPhYWRiT3oJL
xAmABTmgpPU0W83j7lu+X4uSYz/2cf4oWSYEVIEz5ydSQkLnQJ1wnELCVakW7UVFlpOkhVNkU+ES
/vX7GaztO1yGGCVVA4eZ4lnLUbwWHjavoAHWPrIdPTyjbcHJYv81HlyHbjeQb+42dIf3t+uKttA7
yU2UmXfbk2G5yvYV68DqAJVk6hkd2A9VINdszzguC9OSTLc7ejJzZtMJ/CRNr8BQ2WajSoCugrOq
KWab1mqmflMiD37eRX4GclvqGhI8XO5LnegTEMVdDQH/JXZHI6LFmSE0pVmM7M3ysY29KJ9x8vhH
sVoIQj93smK1AQPIIRBOyfYRhjO4uH9ZwWXsz2ZQv5X69zjjPRsYfmAb6JVmK/k3vEXIla469mhd
6GnXDEryg324TFOL34JbNb29pvU+sAl03GfG/B0qUNRNet2RN2UrqwBbYfmE85/Ab6hjH3xJpjDN
RSFOlTHTJRjTwz4W5wcMetOlSWuYZxukYFNfonz8Tv+jJnxqIyGQ/QFrLc0gFIoaqs6zVnfgEtAS
mi/jllSZ2gwgupDzpB4Fs77RPU1J9TGE7BOM8I6yr92IUd2JF1rZd9whr56WWrtbc6iQZprOxfXx
QW0ceuahjnBrLoTxUgVeljxzit3Ta7tndZ5pzvaNM6QoPK6zasOQ4z/FDV2vtaZSXKwG3rJpXQpC
02rXB4ZtKiHwX0SMj6xYpYkqCKksi62PB8o1ntndqpGagqKB01zGkha5HpHH+RW7mFMzmVnDEwVj
nHvRvbvG2p7aHRsKvhPS3Tn7Im8ewEOrZPd1kHUr5Sux9nV3xXnJ5+Yk5tFGDWSF6RsNGs3fF/Ad
Fe3+y3UW9GstlKyoJhWc/Tbj7J13/48mWACf+kjOH2UzhaG/rOh3WtbnZOzlY1DxPCLMexc3ZCnw
fGMThICR/8/zInRBEKYKAE1N+UEoH2AdmE09kaDTSBojyb76VebGYLBYbjGz9ZWftuD9EgL+wpor
+FeB+h9xhWwGEZoCyKGcACRNxDZ+g9JHeU6SWATma3GoS4jfOoxR4BzRe8wrIJ2jg5YNzTWeTh2/
gs6vSw3OM1z9jvB/+RE0sSk6Vqfllu4Gk8iLWQ0/dcgqtLwe0fmEVd0UIIJ0syJ1TeGFJuYr0Lyz
SQAlJRje2qRLM0mck6CaNkeueFZ4t7nwwa0nzZHl9FcBXWlxaNRQMICoYs3GluGoHjWauuwvJwSy
UQ5CrEOMBH4CbRM1kjlk8DHfNuliNAjL5JTRNP6I2VYHNMpWLGolyMA+3QrJJS9W4t5LqpNAS3zR
JIl2VeV6S48dItsiNHWCBE1pIJXyO0r6vbxSBuXAp99KN1zmq6l2z1QghhqP52UIrhvyajkfk0xf
nJUWIFa0xr68SCR2hXQOCrA0HhtqV9IsPeibSe3GC5BiVJnPAuKqWgcxAPxlFc4F2bjasNF4OzYU
dndXF5cu88C8hL/VS3z7ib+7Z1NUG4CCy8NETYIvQ5I/LHz/aMD+bb174RHPxUOTu1VBCLdd9slF
NcZ27+qWKCSh+SiZpV1a1/BGheWaR3vdCKF9+ORBOw/1YkMtqC3h+yT7vNHUXCP9O3UNv7FSBNHZ
rTiT3qbXlinnmFD8j3CJVqD6Y5108+JciEr7Do6uggJx+jyBXw3HL2q3ZIeTaVYiy+22NpNYUGa6
NUtm6xgfxdbZSDxvWGgzVMQg/hSBYbBqi4LtCdcyzGqDRAdYEhKWH0fha0qRKeaT5XrbVvHyLSy6
p87qdESxdRwDzplMjqY9RFXdaxNqqD9kiNL/xxPCpmbhshsdC2AVd2v944cALdlWNga0eMvnhJcu
+Uz7SShEl/Sgz9SppTnpwxyh1lwX8llzocqfqYoxkc2K4w5GN7HZjgVeDRde5JyoTPVH6ISWDbaE
zu3STiYBgpuALVr0dh/zv/ohF4mY9PdMMhlOVNunhpqoP0jMleXJ3dl0kkA9GrlEoN68QKFX6CpE
Cl/pQ8h6B3diT04T07NXP4EQoqPbG3qxlMGN9mvYd9eNV9UuPXR3eb72lucZy1aOx3mWy6R1NNk/
q4SHG4+7tUb1BFHLx14XmniDzcXCHCDv/hjHIjbaWv3Rxuf9lyHrKhUwyrLs+Oz0/Scab/3fMpvh
9Pa7DzE0laNYQbOZR4acNgaSLWMaTk7Eznni/dJSPRrNngpkH9BzW1rg7ciHzjXUleS/lCyzFRcJ
gayoKmu4ayUUR/ENfcE0lALWTqRXH7f8suqs72FcGI8tTNbQgC3WdvJtbW37yYaicM+TZKGLCrBQ
vsz3pT9BuUOq+tjx5i1TlCR3BmgB7uHaD6QYg1xqjSpR2EBk1dtq5H8aYnrDuNTcIsNCp2DEFcun
Dk4jEUZIgkNWYmboTIDoyIto+J2V2+9hifxkFy63fC+DKMQ8WQXJfYBwPkxspnaZjtjfrDFmP5R1
DIpC++rCN4MAdm8MAKdsO47AhZBjby7yxJXM4qorubRq2PsY8Uy8DKUxBUwRoRtK+9zeb7PQgmKE
o+BKS6lUxW/PWjGQ/SoXwe1ZZ7Ix3J91UmRTn9DGdDYcIkbOuYMMOqKxTSsDXb+ZOJ7+fUqwnN2/
Ub3uADs4G1lOvwFNVQwGie9/sARzO+AOwwjE0ZjjLq2GHFGbTIAd3Ah80HwKA+lgr/1b5jCywNQZ
pdKd04scM+ptfd/GFjdpxC/gc4JXRDw8UWTQAvraNjVjMtQZJ/u7xf2sQZGtaeR6SBs/ukC25Z4Y
lqAFSSY0HoOfNrhZQmus3es4G7HhpuEig9RT7KVPaPrZP3i+BNI0xPo15EjS6DlGi/OY2k8vtGsl
khAUD4dTO6S03oP4Y9iWMWR0xs+lJ1/Zs52+QI3bHZugPWHL50rnt3cq0E7t8U6fIml6EsGhj4aq
umaK08Odpic9iADA4L3sZibHt1ysgSCArQV59QElLoDYnI/aoY7EZZn1Y0ICSOkrERhYpOaHkmvc
0Yhk7c41UrP2Jxhwzlf0heKMgRdvYbVQBxlxcCiZKgb52TQaT2QLY9eWOMZ7m3TrJES+A8/Po+SO
TUbpIRVR/QL6/CnzT5yot08+cDTe7Dw+QuWTx+eraoqsrVxL8aURWpEzRkro3UDQOp5bYeTyHrxJ
DHOeNKBw6dUWXO2dN88+3CN39c3/tgXMjdqaKzI3EsjMapUTG2i+RDyW30LdDzuAuoAyej09k2oR
DgYkZse1a5Kjc7xVPTrMkO0JGIHCH8GWi+guKi1v0zGzxIDsGm0T+RG1c0sh33Ah++299QX/E1md
HRhbqbAQeUBnFTYxLkMDj8qB1NCbIloqI74XMLfzy4mJZQFjhqP/gX0Rn+b7YvRcApcJ2347oi9V
MYiA2k/uzTNwI7SwN1KdbG9ULe7Yt/GEyU6gnIkvReVds08xZyGCaNFphLa7pyZtKYu2mvgfZ8T9
R3GIyZDIA3H9MkNJrw+RvDQBk8oA6zezJSL0alBmRfWwFK2iX04OC3mFcxOmQom6iCqRRtiBZZPL
2cP+FNzDZSCF22DPDPwKNuZ6Dj0WAZQGoOGq3VXqQOU2V2eevULZFNPTmT19L0/WbsQgqhjOd1c/
eeAjqGPUneoWPTiJVObhaFaQEXskdDtnVA3os3WeQWacQEx3WwCXzJ5hBLC69nBiJG7aHh3ocLVW
B9f0rUOF+f38FfT+HfUtSbIPgjmeoKXL/Eza/z/CBTzuwTUNYycp1dliLnMyzCX+W9/lZjiUS+M2
ngCV5i2vWKXz4qQuj9/v+10Rq5tioc9xE+eNzfMGWDtgjfnZTsh5d5RPet+6wCyiRUEMmjebUTS2
ebhkUmD5gLKBAXiLQcfjwRWjf4r/iwMIiSkTHh4JlaJPZT2Nreq69Jkl717wnOkmYLnFoOb3Zulm
HQUrqDPMKpXjgqneU9QTSMzgpOCX+nGeGEQN6SuJBm3BklcQYya53bgtkwpzZRb3GSe9rt4M0ka+
xOTs7SE1kLzO2O383yJ5y0J8QcvP+OyhgJvpiSVLcB4bSxv/JatCNi8Y1fvq9aZknXsAeeucandx
O/G+iodUoFYOfb0fjZB0c0NDzSp6Wkdj79JAQmvNLlQomhAJ42ykQZA7q2oo6M/FVHV17fFo8oTo
o+B5qZyV00Et/HErCD60ngHe82y3kbdJrkI78kPaiqhUUUeAEe0Z7xNYSzfIxLFhnQ+71EMzSikb
Z5uOlhOdiaHHGY/vO3YNNxNHToDdcibqyCMaD1BNWRPW5PAdADTKpzLl/ReXEQC7U+QNmWZ27Ytn
4IiGP/zZ2ozp7dVevdTWz8LTE+NiGK/GPlaSbX12JNHATApnLVOIGL87IBs7exKPxYMGnGZIviFg
5wtiF8hZY4/ssJzrTdB9IrcXagjCSv+mSIM2M/DzFEuBNEAxQncy0XL2hn3vgtgi8DFqrRw6zA/0
lxGmT7G26/mgfIlaib1Ej6bFCNWNAek8cJ4e1Gkos1vn+mTfl8vMVyagwBr17d7D8GM2cUKwlBIK
j7uOpcQfR9lioW4Git9lxgsr8KrU6MQ9llmmod+s2dTHB7EaYxLX4GOklLc4EhgTU/jefwKUQrEt
M7+RpxxXIaktOEDc+Ac7iSUdSZdW9NQt8dT8kMfI+lbYN2kv+XsfDO/hLosxhr2j/2URcWpWGUge
sdLn8SsOWqeuzm6gjI9aXcyCSga9/w0TrFE3fqarKZnMyT/pzwc3Fx4L6OOZeq+6mlJkb994ROE9
qiBWn/mXTo0TyNz5uwniAZ0Trw15ylETSrg0lx16MPDG4R6eO+Nyp3bNlFmgVA5znYXGUceJ6ZdV
zJ95e7UfLg3CsFCfoVZzeuEIZft1ExI4RJQR4yXUWwTMpEEUsfzi+vFSvKww3fS3BANnIkPlwcNF
GQ79JWlGUKfyJorEW9o11OWlYNjrKKvWex1r1BzE6Ba8X11Qe712GckJvr2rapn0wkPjKymc8kPw
1yiBMnsMIMi8GPlyqTFssbAMYnjp01BnHOfR6Tj3ygW5/w+603+l/ojRRgM6g7sAM4vELZHfGKWS
M82qAMf/o3MF+/AgytVnMv9TQcY/DJUsuvY+kLFgbJzgGP2ScWBMgKeyzo56reRt7+1MgKGsNArH
SxbZJZ3HOOrfYFct1GF7p+uIcPQkFtNTLn1REKqkZOfFv8xtWsTduUpxwE1b4iPpGx1XrrnJwLj3
1r1JnQHjJygtq5QZ3PQwmLaqoaz7UwGlrHbU8gHqAGMwZgYRf9JxEsxezll5XqKVttjDCTiyAOta
z22nlJyCQY6jJamRlt1P8ZafVbS8UPF0dHkZXF8/jAc9Hg9qBIe6Mt+XCx5754GJIJbthV+j/25G
qQhCGQZ4FeAzecwd/TJ9opMbynmCAd9Y9ORsode94WoiLJ+EcBaueYr59ZygW7GsblFSUAW8t8L6
fpsOl9wsChziEsk5AYij2HGiQNmnDXHEsQSRHc5IowSDCQ3bxjd2g4NTx7vvyH+AwaI3JmwuOs61
srB9CsyGNqnldy4beTAgkMNE3T621dfghsedwdR29hH6MNcXoTmNYVXpWh/GfhzUw9gAGFhpLrFS
GfignvJJdrcC/1keBm97+V0O9An4wzP1xOF7J/YidgzPxtQ8Fx3oO6UaXKfzZsgP12jIhJIA+h2h
QtnAEcVcsNvIwGSjtqrOStXgrIVCEFGh4aPFu1Lhgqz4LW2yDLScQQ3xk3xBJ0GOnFSV2q1fFnWD
2A4+zWNYCnQdn3JWwB0tIpsqPQLj+0mR+2Vvc5zBilO4kxaUOxSIi9PfiqDf0ib2LsEsdYT+rSF5
qGpRAPgJthyYicCf6z7tK1+8aeR0EPfu0dDIDX1eeiS+LIasuLsS4n85J16vxsxR18tShKD3JUPy
XVcIYYUyykbRUczDvzH5/LKqfLEKMXCOnDd+GOURWR8xNPY7QiTWFxIzHFZvfyEI8Gt9w37SCpg8
EoZr5bcbwqO9HESfBSkyfiinQWBXGSa7WbOzVC4a/tonnezmci3qW4Iotru448Rz7SJ6s/3D5sW5
LM5B1SXVPBlMcoMRWXaLvtrob2JPQR887JQgT1OqptuCJS1YUSGzNnPACzaapDs8g2zt2jq9ZvbD
JYnn+YRFv/7tDrShj/SIM7EOe6M7sOtR4cumGYpPhF2hfVkCCV2a9cajk0AgVndbVBTYlkOI4fOJ
nYn+Dc6ysDo9QUFqucMr2Iy7Qpm4L4ksFo5p7RnQWhESPrmqUxPIrlIfPPRwGf2l3y+gsInsGpBR
ahkGzn/He/zcsODc/1d1WCGvcm1HiiCT7oaqo6v2LPNXPJW8GWa0kKsAlajQ4iZ12sR7NPK9nWdY
wKHcJoFtfq1pn3JWhJv8tiX9EQn6a9VnS6OS1SFZyf4EJ4lvway/9Qv/qxwKo0IVcWGONJ4XwZ0W
0oMhcTz1xpNsmCi66fBtiDLx2skC6zw4dk8deuRE0AroHfvl+k1DbX6qi70htl2kAsZer+pS8lGW
krnYk4IQy7Tbe/mKVWCti8S91xgd60uqNgug+nYOimWWgaS1rAnWIn5DlA66KpnPBGAH2psbHfz+
qBQ2SKA4b67SHMAj4MMdSupWYqqluTQyJsPVtDSQa9eVZf+YvMolFMm5u2Nw09R988igSZRPR8DO
ChjrFKLy5dvtyzmwYKqoqsotc48KldBg6AOHcjnbaMrDnbReNp6yapcrQ/pVUKVLzZsv8Sr/v3G4
kFtywCouP2dw1kL1tZTw3vxpGrPh6YeJaIfdxyuOU3hTljTqFoBi419PVFLYdoUNnc/BC30z9TcL
/pZfcxcIKr1QD4Wou27XshyP8G1QlK5HBuRJO7VV/gYcLFzAmrCRj+tjewSxa2gK2eXGxiNkIcSx
zHDYy/5nVOTHU8xG6o7QOGGUwWe9KCNnXTfiQPsmXqDEL9xXnm0cCmMXuMEGLCVkiXv/BXFx/+ur
8H67FcyLADcy+3qOmSIOzx5JMiEsGiORQd8L9lW7fMYbPO9zfqT9CdnaHhLaFJ+q21Gk2vmmiv2n
5lfv3ddwKq10YMkPDq2LrZ0FSACQOz3OAkvt2KnzdX6d9TpI6eELnL0YkURaWLYEAAUogohl7bWr
0jh4jz731VbxavjhuuO+VXczRG7KchVcRsDiy8RQieR6TKI4h5QNftsNbeirTLFjQXHaakSL+IB/
zvHcut4aVC9hI07efMtFG00NhjHS75oa6unvdeUG6E2rTrRFDoF7Qx77lDb84kb3muXAFM5iMmsK
CNpkoRq8fvmRP7O8HpUV7kfkLEk+ws4jMhGiIPeZRbpCmMIxFy/P9oxZsBFjkD1fUhw+p2q6neLJ
nGU7A4lfD/cIaYjoyxsCIUqFmOF96xqrBlr9mgOB1iS3k+6ZtlZjYbHcEWZtT2tGYUNr+vZNocAz
ryoO3ldSQzF+KC2U+poerAzl8kM0eM/+O84R+O/FrUpqk7rmQzpUvEFggWdWIR2D+9N4VcWHG7z0
fAFRse4EW5UbJgHxc9LtLVYTLZViXusYmVarrJkJKBj8uV62iAXhn+MypPedauUi5ogmhZ4cDlrO
lBOU907O1hbI4saRp/dAN9TNxPVrz+NobSEMeg+GuLWrOxnuvSqsDzZNmUkSJBiYo04cpvRGrfX2
zFE+EZ4xXtgFXf27LS2Fny0IXPyZ2KI3fUvlbmVdE+Yz3/8+S2cuAXfNarrb58TrcZ1UmDJ+E38S
20FWofvoxV/6ETV/3TnTyJ47wHfG6meZarrRPsf1rLrFalts2eQrP+ObrvWoycqSdqOSiis0Q7BI
997NgIDqV0FAC420RTCdZim8GZgk0efL8CCDD8qsr0PtcgJOJdM81eEUHgjq/Sn7UGP0AuqpH5/J
qlvZADd51VjoHSHrDgovaAl007Xyis5ciUcal1dYWV3NPmn4metC7YEYzWMnJ1emu/v0rOpmb/3y
IGxX4z54V6lR0ZzVhu4gds7Fp5pdPRK+g6TwkYS0yaN3t+bFqjmFvakYjJfAO+yB7MEWJr55eOR3
5XYa4jXIAUqML4CuINqqVLurowsTiQ6l40ZCDBf5zP/G6fR732AzFR6A2CJ1hREh58ibvaxxDWDY
dz5aVr1V2wQPR1tKTTE8nErQyvuH8u6HCl2LBcxiz6lYeN9L3uMLO33s27/DB6Z3TpnTKcKXa7T4
L2TN5T69dhLvLv2bHqNSQruDGK0PGaOmRD9gFSEsXf0M47cBZ3rZy1TwT6bZeVB69n4nRMwVAKb2
Wq3euDSzJk5RxhNj473i0hKdG8T/bhIrVDDz5fcXsv/SvPxAzv2dxv8T5g0qeblfal9rIx7HvMrL
oxA7VsSDPFZp1G9gyzwb1BIn26XQKbots1BzGcuBQO6J1i22Y86HQh7H+qv7w7J3p3a7fuM+xp3U
yNSDywPOUEdPopEEE0aEX8uo+3KeugP37ekgXMHSJAosQC0eiO4v9kWv4ceUXkJGIorNhcwVzFDH
lbgrB6y7/L3zko7pZuKg/FzLMC8yAlQq77KOZilKPFsolY4YHOVgB5SEytmIcz9LN764qIzaVH9L
4X6S2+/4vVTTn9wHZ9ceHmroAfXMyX8IBO3Ju/JEdrD+a5mupDytgpw6iM3r9uVNhxTMIkyMjsi5
tmyihVDus5+VdWW32Yj1UdROeRoewxnz7EhwAlBpiD8zpVC4Jigcz1oNnv4MjIgbPAizACqTUXo9
LpGfjed8kNkMunn3wUqmwUmII/f0lECJPpByzTCLtdIhTn19/UB7oGSKygSBsD51tYadpeh/yE0T
LqjEg3pq3kX8exoIqmZztfivrpmjAkM2BuY9J7kG5wzV8PesOwxucGKn+oPOyra3YQQ8IN1zE70j
Y/pAX9tSkt8gcdegSWvM4S1PiQYJIELJOpTi6IY20d9U9y967cMfSpy/wQGiPbZS3zSczfhK3scw
gXMzb/SZaZrz/P7bvOmmog89l8abmc4f3LQSHPWwLeTQ2cGt0iXHrT6YnCmF6zdJpdJjDwJKO5xb
d2891M7TWxZtAo3Nxh3IMjmPl5yBwYQRgP1zJVu60fCOtG/9Cq1jddc8fH/oMFzRFk/U99bWrlC6
S9G+hW6f7wVCUFNlkkvamWUmWp9dcUs1JLufGxKPDbf6PrP3/BVehdLE+96VoiYlnSxorDeTHOSl
X3xXMykMJSAzbKm5QJHviHtAdTT1eTbxFNJmPUFaBKUB9TufcCo8jyyDdVIqKi1MsIZfChCcki0x
+eQB78gQHgr+8KIhQNABUmL+RSwqvJIB/Ov6m2zr0To2DivAtj1tPL6mjhXnkj4xZVstcOjqLBHT
yoozBYyv3cSzrHwkzIBM6HX25R5pZP7i5HsfkEoenUjJRmiiUylGxBHSlD2wretKt+tPmImohCud
Y/CZ0utOlJESs0rQ2exthKk0LfoDTHQ19L318HC8acJ27Ts6pTf4SoFNIKWlEicrVtmku0QuK+gt
TdETiz6EfEB2cv7g5yoLjoQsq3C9Bnsm9AluYaJnATkpz5jxvhtYsjup22OedSvl5JR+zzMQNT8g
XzEUOQ1OJ/l5XWiwoNIGnPgdmq2VWNdl6aaalJIrS+IFBCHhxzhE8wvT4HDVyMOqGjUgnYKixgs7
tx7UVZWo3EenA6HTtpez4bV+vYsAuYX26GrIr29AywlYu3PelMUO+lilBsaRqaksQ6AQXtDia1WG
v6NHGW+stMhcVuDWZ6g9VktbguGatwqwBHDVnmIJ1OeZYOvFxkZT//7qbFpfcxDO3UlZrFYQ25z1
I3MbCMG+ohmyjqrdg3qSQnyY95FslOt5RsJsrnz/hOFekc/wVdE6ABTwq57cm6Kk/mX4tlPKdUJI
IyYio2zcsLjnk6v2g74eoo4QAZjBAN+R970LD9iWz0vPKRbCbfqqJ9ljF89mZgZ5Ea84i2s+fLlS
Bl01j8VoTFaAX0ggQDDtNSFPI+0H+iURGDdohqZoox9Wj+4SDcL+WsWVpknC3BbSji8LhrdscpN/
2QEGgJj/j5RYH0o5cgf7uK37DkPS6F/VcvEGC1UwJBO85PBvoPW4miX1hfKEuq2dm0ZuTcsrlTWc
FtWmzPWTy/caBCPmihh0J2nN0LA8d2z/wzPZXoFhHKRIKKrUUkxjHGsx5o4SB90zQ8sP1/j7zF6L
tpZOl3nI2OsTRe5Wxy5lwzAoEjwXVmAUTfQB0lUvmQc0YK0rC4qSIQacANv8BYO/CUV5FiTS/Rt8
2cSAGNBSGzlVXPeAP63mZpRdJkr8sCEJtuo7F+NM3puvVO0W2c/x8pHBbpjtHppPZLq3QPUZy6+7
ELbk37tO+iiNU2ChF4BuXugOUIiM/tOFUAKNcnmHIfiWq+9Jt2knJe43+mAOPahy6e9G7wzD146j
4NyQe7mMVudblyK7+LuCTWcAtvuHQS/xdmpwK9y4asFOFR66hJDMpLGcIdIOkrPDwgMsW+NhhQvb
1Ar6kbkxJLIixUuz5eq/df9EvyGBpPWJ4QsU41hAEJqUK0HkBM3AoCzyGoqy+AIJFbx/KR349YLi
JXaDkhlik+4nuavCnG2DyBCflvai+AhKCONVysi06bRcGGg+MkO++cm4nZ09AoQD52JUnLAxao9R
6Srn+btfXLkt/JnjQlf2FzJ0rcQyvdf+IN7j26Foc8VLCmBr7q7eRcMUzLqHT3QKifIKumSRTGzE
txJCWZ7F94NBum0Sn/TJmH24pwDxEcc7K2/CaxL4rSAEmz/MhF90eFXQ2KlCZAejtg9BOzG6Ia3f
N/V8bHGguhwPYMibuRMAeosWdpIdnWJoIGsqzJnDdQvLecwPjWaTr8XLZZSBJ+GUE9PIoLK0wN+2
JTutRrqDYAQ5difHBpt/JizMRUqeY5zwAgDuY7qpeaQAB6Nymvs0iieMiHoEF/WnSpt3kmjuSsax
VofuWEG6vuewxQFCKWitjisvsOOjATEwXkTG0H2xZyHr4MrGQzQGb8Kl2Vz2oCQRWjjmeGfesNeH
JGXNSyviVFKoehoQa1egKxCggJ4cTqGKC9gnnkYYHtOVk4QvmmRUQRA51K6fFfmO9OYEZ0KDp1Vq
23N9OAMLIDqMB5IDxuDzl57fH9hY/LN11OaObhRCEsRQQiRbD7OduTaTiI4BJtFbRW8ZGmTl2NyN
O8AsDG56TJynPltN/s24sVjk1W+bHyi3ajvo61c8NpmDJsiUKJHWFOfapLCF+nnQdMt40u17uuT3
+DAM33r4Yfp1O7xhjtePSc/0UqPnoKiiemRiBZ0gVhd3QQQbd28adccMmvXvlSF4m2oJuwqveMlD
lP0tvOUKnwcyHIDp8+MVrWx5IlZaKSTb642vcQMrgosn1po2lrE6JvVWGTSLMs0b+wd7vvynr9mC
3YXJpr39JRtPulZx7F5MJgOEttqgDBWWRP3QYwUwfScT+Bl4H6gJZpoy269rMt1eusXz9tJUNS6M
PiIbgzkyCZFJmp3cw0Uk4lppZXNszzmF6gkwfYv9DckTxxQuOM9M+6/RNYuxHpSYBTGUi/cIy65n
mQ83kh7WlKfRzjxsSsu52xCi9zicqYUTglP4+1D8yJFp2S1dRJwdfjz00C429B7ULcw9+1+WTrMx
Z8rZ/e4K7j9hdc0KVEAPa23eGKMWyBODSTxgV2Nbyr0xgCkEfVzd+oXqgyOGHX24MqNd4bbtR9LL
XFjLL+Jo/CgcquluCM8f2AMMkFr/exEWUm/Z3io7W/wf/vMDavzHYyiKt2Sk25sPlDeE4lVZ42Jc
jEgGMaOop6EEibzpfvWPifxfmmXaMyBqYrld9fCmv/AT9wsGb0KSx0FCd0JQ3TuTQyoz2doId5R7
gtLHJvHXDGZKMdfal4SW1AyuwJAhiKDENdPgz5JQTcY5WDbjGOEKNFG/rKgW5PXgDyRCEpNpnEAk
wPqgXvIlRjFTrtLN6nfx9S8ZpANb5QgNZmNVXuVW5cY3ulf78SYSduy+bO0bjTH3uV3Q6YuGRAvO
eHq4y6xFVaApQMbKQlmkJ7pQKNvIYkJbZTgUaSwv4cV6JmDD8TpRVUJ4LuNEaF+9WgQDeAuSsjZv
TDAu9L2LUkZij9Lda+OBucFyG9ualdEwCqShERzxUN/XXBBTmezrcgZrtd4w5BntQNB1ETfYowe4
3OHB7Aiss8HGrkXMvLtU+OTQh0gJIZ4Xkrtwif2L8c09rh1+6uZkf1qH3PaUT2YOxYvOBoH+Wtvg
Q8qA1gnJzBodx01vVUzjrG2gPtfC8ZpiBXveHxaCpahK926vPgY/CWRKH5B2wQi+3Bu/k0rqTlZ1
NLfwgj7IQ4YMYKuIZ4X6GQjwru2IBdmkuZccAIP4kZqSkcoCFxLZCEXfe/BlwKCh/TD2TB57ZcjE
tPCozApiMEZ6lq8ysHBsmtMNvJaR9hI9I/9DUmyzyiDXJzv+TRSoud9a/w/Srctl0RVwxkNHiwWv
n55ZTWOGrEa55NInauP7Lx3LOjVnqUoeJLtTniHz0RE98EWiTpH6e11EIqyfP3SMvEIXDue7vABT
4O33vS2wvG5Fc4DP0wvkZDR+ZcLYW8Tyv39JAI3Xbkmy3bdUAZNBXSqQGIp2NousWFm55zO97sTR
U4/pv70VRpCsJYqoVZHF209YD31yjjudkmLPhQn66gRzhREnTWlxL3B1SGmixIKPQ2he1wBUI+tR
CbtxoNnM1Pxr81xxJ+Iu+IcRd7ZPyTxH64/Ac9kxoOaorKX9PKcEgEKseCHTGIe1+O9OMmkRdQw1
lSvZE1kw5TOCimtd1v060MiEfcYsxdbqFjJDQCDKXGIALVZ0/RqHu2lsAGq0OV7qa0UrqtQGB7Xe
Zama6LpJHadrDblde4Lyfn878b2VQIBcnDEsmf7yJZz/P6FacVhTSmihB6ujPhvjjFMGOGglUIU9
WKExZg9Hq3j2TueuudJ/4Dt8GhcSRbJNmOYbOp5j6KSR91Y/bZJKDDiKWnS8W3/UMi1MxGbQKMo3
dVlbiHW3zd2DVQMCitk0vINuoiVfXuD2BCR6Y+Fe13DXIePHh8dg8bDgEJHu287odZkUjNJ9f9Uh
TZca0b7DW9EFZcDON+lPi1YWBK997Aag95+kX/Y7x5xeCWrYpY7zEw5FTD8WypnNhqBTn72bshQn
gu5jvTSeHmy7zCMfIIIwXpcsnbzzsVjhi4bH+LqvrX/4r/NkUa4Oi1XQh7HHmS8M0JQfUjLvpvh9
tgziMj93nGFAm1FsCuCb2Kky3rCb7sg5F2tqC3F1liZp4KgBIRRx4PW+1Q11rGbAEppEJt/w8JXS
Wx1z04L8k2wmGR1LvunfyyZrIGyQPJQAxRjFK/J83aXSvYd75No/YKAGBvFgMVCegEDB1eY0o3X9
sanPkEa1ov4xPeX+hlqS2sJqPAgPxQgErYZk5Z8MkHKJAqpaO0s6ZhvtH9HSANBJgiVSPGBh9wug
kXoh46WmkF5SaQK1C/ij0SkAgJ2CujtxVGN/Du9D4PlpYCIVPjtxK376NX6Vjh7LV1T6EmXRCw2i
MlUNkH/rH8RmkCbyzttwu3bzZFQx3ki6PQp6UEUy7g2xazpu0S+Y4mK0zgCZpI6uF/HBqHXHV9Eo
anQkiuXMZfa0cVZ0+w+nH7QYWPkoq+Kh0jB/awT9tpaaK5SjVuv2793UFhGL7YPKQsaX9monU0ao
fxofcnFbyPYlCABr2h5loqXVHqw+8v+ZUamNFJbeCsMIdfJyIgY3NYpkM7AmWlzfI3ApvJu36T2S
n9xcAjqr9uJw5gz9uF7oihoImZalkxiqwSrz4WKSFSxdQ3AhUldcqWGfby6ov/4Frep67XYrvCXi
qghNo8OoAO/X9lQfMZFITvMKxgOcMDYzhRGxWyZM4uT479/u64kXctFhx92hpz0WPGFKV8quYdla
3Iv7rWWb5BIqSrtiSmNXsqyNhw7Xbc+bh8Jn08kEb7PYpQuo2tr575EpNv1s9j9+xM+7J7d9mi5w
CUY12iDjyn66zZmrSL+BdIVOsilp94pc6QEUwCWKxp1Lv2RMfvwHI0rgE9tNvvU/4BqrkohmuFEe
zZ5gZkA0HWy8aa2mLWF6guBeVY+EUvHu6lHJryzaXWYEJ8SXKFwE2sMvATxWNKTTqzEG4qobCq4n
dPKivicRhsCPp4rioIzx5jP6Qo3AedPIw9aEGgeTUsZ8SsLu8kYH0u0EGDoMBfBIzzKgy2YCj4eE
UfNJlN8JBHWdbzER6BChtab50ImEZuSzwD/GWSJxxv1y3zlW0qEBlm0KmmI4wtUL+7lInAHk63Oq
Bitj1gFqyxv6i9CdWJVNo2u1/B9f9GIQom6BCdjveXyY1OcYTxqyaQjnzBxhHrBhYjAhligkYGXn
I9N8x02WmHMJ18b8dJsgn0bu7Sd1XpSAanlzAQZ11/eyx9NNlhvL9KePnRTFP62Ii7TKHVB9ryqi
fHCWiYOe0L+wKgHvHSxUCsk+SQspZvTZxpuvWezLAAWUTnyWiGKx57uOAmabRqpG3IFqQNx0Wscy
8Vg4NhO8aLEQZdMlQmSfE379/vvhVNXS5fv6MSEm6OCTSrtfgAEYu/9NpcX5D1Zkt6syOOtaDqB+
Eb4H/2TbihDIcouIbNBw6iNFl7XG260FYl0o6CgYGgvDGHxfuZBTkultGipVaaR/ATY+oYnWynzF
GA8Rfij/ajTRBwaxFb8TCYuh3+9KB1QyiO25p9mJ6KQghAG0ZTJYzADd2O9m17OtNr71eqPhU/Qd
Stp+8D1zEeWCS5yWDvk3HgPEwvVgUTteXU4yOoSm3gWZtrLEkqI1QLi/3H7FiLtL1PdMV1WrA1tp
6IkLpTBUgqCFsUXXSPr/CPlhJIdsxCX3K4zdMqx3D5cnBwzzszgu1sRagvPou3pGikg+GahSXbET
uz4ZUEE4T20uJndY/gfgVaqgO5e179Ugl5XldKLDCyxG4KLt6b3LrNRrKmw6aRAbhXVqy3NvTlX/
tc7Bvb2d7NLQcK8Es3BzpfSP2aVu97O7tR3sI3IW3+N5LkANMMZB7Lm5DdV8+dGeyXxvT1pMLhlc
4kpTUn558qRVnUlSxmKMqiCKAIzYAs24EG2jAqpaAuFc4ULXGePU5jSajJnS/eaarMoNAb2lddoV
OQKPAR/CuLnnlPx6iTddVIgvIxwg1wWy5eGzx0jnpsKuuUI7tZkzZFdcMLpfA2+w9SM+3L4q7XQW
x+wlnaUTUPKC0t3XwbMnE9D1E8tLphmqMuy7D1hzxgUvls1T8T4eCT/ZSPPPmNLvXUHEFWbhgt7C
BJnxjvLjSRMdGgBpDCnNlEZE0r08WqJPEmRzfiNQBRUmHNo8Wwz0TJK0ihjWHt8OJsK0DR0YTMHf
b2okJ1Mn9dVd/CZPe0RtFA//0BXvLVtKiTiNwiWJAR9skkq7UEq4G9IaovGAVZVMkgrXab41KqUJ
wSGuN4NKKNrZaSTeWBYeV2RUEZRmNn4ZxwMYluT+eJWcnglsfJw6tkjzqh0B+53v53tEPVi45a4X
aR3dUKwv84GT3CEZJqUGWrWUFbDEqVxIxCZT3B7ka990bk6dYDdXaWHMueXUS0z7vRHSA1U5WkTw
a1hLtrVQFuyjFoPM8EioRgNSxd1xIIuMoq9pE6kVgvmcUP/KRCkwAQRvcMHErATNGjik6MtrAejO
vRKd6JlHnqQS+UPB28Jx3GjTVIF4VUI7xhj7E2UmXIEzIKdKEvrPI8vaypiN1tEgW7PRkptP1u+L
+BcMNySe84P9I/RBHPzU8kIEfT8+IrUaUoPyvBG6hkhqSh7eqcheQEKqRWqcH4F7zi1fK90jzhH9
PcQSZxkd4AIgw7L7vqQfug6RbMZ2/G4GwmXetrK8C9WkrgUdQ98yu5R+te/P49PPVzi/OkmyQfC6
M3yIgxYoejnuIZT4yd/5A0a9PtLnyozgldzmcvS1wXpz177r2fnaFl+KGRrRHsGjFM/t68ULh8tH
TFEKa0L+wcTK7TD2WdH8MxYeyye0mJc6Lq75ZcVoHacO9R97xWcS72oup0NNIX87Cg+Yzd8l7cr9
Akn4DqcUaPV21mr5brB1NmOz5253i/4KeVkZX2Bq+5KJ1pcM91aGdKJWiGZ/gLebiCjcq7FfuYnd
/G2wb1cSLRAtIrHiheMexGN5/7ssPRquK7aFU0oQcrv/DmTM0kqAE6YGG0wtzCZxsPpaB5qMU2UE
kpomStB9p+y9cr4uC4QvO+BWDDtXqFHr9RHKvPLZObYNQxZWwuoveXWd4cUQ38WrTQsU9Bnkv0jb
Txm/T+nv+xgBDGmlCHu6tvk9xka9cezCb34ATUBROQXbLTeoSocDhDIn4A73TwxjDBOCQ0yDRtax
hOmB6Cs/PD2DrXkQZRKHrZRANPTnolj+PtDPF58sFYiLVHQSUbZgSf1+wnrqIQgFslj9tddPGuSt
ovmWx67LzMvNZehuX64qUKzejkO58l8zldLYZ6yF1V7F7mMi94JjVgqNpvLVHvImvp/EU0Sgmxm3
dX5qYiL6L79zNm9lYMBoynH7BMazVIvZCGG8bv6Z6j6ovLBsUx+Ipj+UIlNKyAxQDWXmG8595Qpd
QLJZw2KkMrj1bAHTDQlNts3BrS/bwudG+aBSSMxhlRmpe3x4bFy9+mxLLjw7ypGkiwobWpOlIrmA
fcqwDcj9JXc3Aql524nvoYu5+FHGUnZDpmWeNodAiznwQL/C1Rh2obqPPZ/rG1JmAfHMz11UlCvM
IuN4QuHc7pt8qGvrl+Mfl8kkFbbxb8tmUNA3D3n6mFDoo8mzunVDotV9FfzH1WDO7ZrMXehvtFnf
LQWVC2epenZqSIAK9TPMaiKPf89cxxId4cQD2Pk8TBR/KdyLidSQKTQ2lBl0+zZgj/fFploewXqH
xQeZRU5IbqsZBwmNTGLV5SlJyk7pCz135aoC+yiIo8Z1LSNAKyRnYQ+Y1qvl5dlFjE2G2yMa+HLP
POK0IHbSiiCSTDo901E0gtlTqhWYXuHqBpOiPrIVTzWd6YD817zASvNFgq4mu2Y0KPaKrvAEeNF6
gqR1Jum+E4V7hLNE5ow2CXvey5NCRlwH1h6Cm15XqCUTxJT3saMedINw4fe/TrnJA90o7L9DgDc6
YQJcuyQm2cQDkzvO2d9H+UmD1WqiKM7w2nxvY2Rt05S/Ud0yLXVAy4eQazg6Zcjo6ARGuQLFQIdd
Pswdjw43Jik9aGuEhJuPtq9eh+Lde06eVW4fv5Bj5ZQ1L8aI6Z/78wP4QT7stfNJIkjf//nxXNjF
xCN7UCqBhHCWOor9+lXUE5NFqnuWAG9luf0RoBaJGSBjG6BNs0XHf40EmuYnYMUlWBvTe0qtSvDs
I+CV2RANPevOZ0mdYE9ReaFg8IAONC2vKik3eJDUt/+N+9qeZU+K9uw7DxB4VnCC/QexztvDYhI4
5tBL6wWpjM09dD9ZqpAd+iJacPgp1+Ihyk3r0sxxWeQR0+zpgTjZxLxBny+x6ipbJLrM2H/hnlpi
r8WYj8KD3uEkUuqBfCqQ+3SB3SrZS1hFyB7nHaIsuEOjvAZbMdsLGLB/Z56soocFVMWrGaTs7RSI
tcBN0SQupmQiWZK4hHvD++hGXE2EPYXXhD2p8TCmlyK3QMM5ooDWM2I/WCbQY9M3I7zBdLme6LAq
sgB+pKskrVzhFtp3xppeJvQwpwgXN5cWnchnXhjrfv4S9pruvIHAUv2rrie1fRUfMEjxLwHoOqEz
62NncUZP5B2PQBasFWZnLMz7g16EhTJDBc5c1SNcxZSKIIfCrB7YpjOUkzWWJkGI2RIa5TL8RsOz
vp4GMMXqUlFj+yCq3pQgrKLrCDj4UB6ytRlbMIRXrAteoWO+JquQPF+Gmd0GnQ33KCkSporhiTnN
d64G+Qwq50nYrdM9nrR3+LYiZ+brcQ8w+r7dFK9qYeH9ddtWSzl/EokI5FcCbraKctwxVcrsUyfb
vGsaMsVOgCb0seFAwcwl8VGYncyr+N5nKJ3kJobD0YCa56soXopXCiWHIwzpttHg02rZ1qjI7O+q
ZNrd7DJci+JiHZyH9nFGDCiLq7iAiMYlmunq27gdKqlM2plJMInd88hJ7UyXXK1rrF80Ip3Z6ysL
M8Jey8HMjV1zOUTelT2cNLbZU8OBtB7BAoyWSTOvh4wDiTAr5j984XFgC/mIWvxB31bJg0vbpFYT
5MTybHc/lWCW/I4peFcu5Cpg67EFLGgxC0FbbtcXd7HWgJWhFV2DnkopRoxis6z9HPlkQI2oPKBM
qQyyRekti7COCRnDyQT42h+rZ1fUi9mx10cWPrYctBuh4h8+AzIud/oIJmHYBA+VI085MXlqGHhX
1GVCoh4jwpt0x1n7nWenTLQ2+wH2FkVqhga2HmzQZWvI7lCJsI8clRvY84gFXgO8bhOdOpR0D79U
8lmIcKciEfQBTE3DW9/HirvGhes67/KlJK8cwq8WtrZLZ4BkBvZ5/Ws8iAO5fXMWlQU4P5rK3WTW
Ndqegntx6oKEJ2zYMn/U5taCnUjuIEmAm0/UzrgqP2E1+eFSW1XAtJQSBLFfmbTGhr7bkEEN3SK3
QOWzr7Ra/R7qt87PSM6fDdMFnJetHPkf60O3H70KfXgtPTAawm2fgLM+aP9nIvBLsSIkZEHpeMTo
ai0QVoItU5lcvJjUzxQSHxLSiLPb415xPTM3B7ltylrK8L8DCHM0peN9+eSl9NRcboeehP4j4fNy
5f3/TDCUyx6m3zzgYclwGc1tSErI+j0nlEWQv72GcJnhPDx+tOv/ifwp+5/ChJbiieZXtugMwZ3t
/TGQLg8I/NY39FannlfTrN068QsSDRpK1ohOBuijS5mQrN+VX+Oc6qA14m6OoQlSCowvOtj5pcJK
pRISpLlgLGXlpGEUeJTKcCfcCvWLlsLWC2f6N7fn46fK2TXB6l72AUwyF1F2XHrNgksSak/Uv/aI
WS2nKjhHtTwDWyt7ZuBw+qL/Agt4s//haPZxMuiGpvhob0TjStfIaZN/8nLVQYZ0FRdxhbP5Ti8o
4b+3tlugdsAIzdiWonxsMCZndEE3j0NTTh83W90tht44/z1iH1+6a2+e5tTSUaBs6ICnxvkfhbKa
PjlVkHet1pyCZRZ6ZR8WyDZUeF1YGPaFkMuYRatGb/nbyvr7/3I4sJMpHuHvOpxnYH/r+s5cinIC
bFQ+f+BcqYXkb71LraDmdW9MVHiIKz3WOQSRERtVvM0O7Tk1UUEN1M7PYCSTGhjI57y532e/3DAV
/LcBMn+s92CWhJRdaVFMjfvXefCTWMffyURQgqh5d+GwHULyyhzo/SW3jxvVND4rMKajuwz6mm48
OeJnqnV04OINba2uBDxF2V9uIhhXDe3qhxtGfpr5uA3UU/EpqLUa8NAi0q9g8QyypEzTmTOuiC3z
73manc7po9cJ2PfDJyAvLr1/bVlgVt6HWTxSYJ/0oixwTUzSTmZU5TvQvzsO4w/e9t9vDv2Y1kEI
kCJHONC62u5zabxI1ea/iJgvQ6umakKNPLofhm3sOVcf4RTfQ4f17EoS6YghavzFqtXXpRfv1pDf
viypsAojM5xKjcCB5rXjCKyGMkHHUB+unVNYxmkgo86/6qk8TpzC4Gq3Q6v4fD+LijBmDm4f10AH
X/kbfP6wexZBtxo1DqMwBMHXlzA5QNSm1ibC8lkoYKoaO9W4T9MDjZzckepq1HbxCKCHMonHUYMt
hVrMx4gOHkD8QuVvum0UWmmK3a91jEv9bC7eGpRQ3MybCUI9mNHF0mAyKf+4wmOUjhgWcbyxMiEJ
R6ny1pbtWwPY6lfE/P3qgOZ3Xrdv5wy4t2UaXYDth3ogLSb4gwUsykfXFIqL2gLnyN3PylNlfHKk
ZUgv661zYpU2tNxZkLzNhsi+9u1aq8hyHZ4rFyfsHWzUxURWVQ7ob9dDZxAgVyy1aIMTacrndk28
bAtS1ilIKGHmY5echGRQ0p+ZAryVOEb32kusmkqyAcFKPjMeZXZtllF9dyGKSDvV63VzyVBFjK/J
48KfyDVWwJ171LyGpkqEfxG+zNADo9xMtpj2GMcNTjrit7Sky4UUUNkpqcmytpAG35moECUXcTdw
sVuO8izXxL+xtaNI2OGueyCfzuQXH08ALisT6k7GfAu7kL5L2q/aoVqLsFjWEWhr1n+krwsnLZId
cXrlzHb74SO5cFU5TWCSc8ylCqtWiDqussf6KIHJO5SpMg0+G3SeClLTbWxMm+EhX9WKshRoXgVc
jQ/wCm0T1IgcoT1RcT+CeEdCGTuzDTt2Xzkm4HLSaEkvZ3jZnY2t8XzIEuTobtL+ZHIDUkW31hmn
krE/yTnryGEpvxFsUp5eG0ib43NdXbGf0rvC0rzXGsy5ODF5jFynR22EsxyKjwJjwCbFZa0Gfrov
bG+JMM9GdF5i+mNgz4XDr4OzXWZS2hxXfLgJjO3aSw6/f7TAxF8TfvcUweTCG7Uisely7gE2egWo
o1arzsLxwIeCtwukmMVeeFANZ+bEotYxzXzTZ345ufInwYcscKegwkjR71ctmDO1fsnrExUeoWxb
BqYKxS8cEoTFZUS5R1zeFRm6TIOuU9dfeDxuTcZy3YTXZDYn2CvSVbnUzqcIP9gSvf/Vo23JLyHk
x0l6vye94ng1m5OkL1yrLUPFs6g7ZMw8hCsDHXqe/mvKtNAsiYqxvGwHQEcSaB79oMglsoE3Xj9V
qEe/QtV8fnweGoNdenPxsk7RdgqCCQn7Z5H7bxPmI5wbr436ADEykmPuoejqHtkgjvWn/7RsksMi
CSyXNNdLK7ivaCcoEfJZbK4uXyoNcIZ9uTlJjy/4wjPq9awcOtgbxdyd2W0WDI4B4tzwIIa3Gse3
8G1xtGCgKdHoayQrVXZUyBtbJq79DPp8n5ivqWX8sg3f82hTI6HO5BNha6gmm170TUBJwSDNJC/x
qRGm7XV3gJOu8Ka5C8NOclKNEp6hdcGc+hSy5OXmG8ukJpHxL9dy0QV2knZxoCz3XAIa5k4/XaoK
tEYgvsKMYbjS6zABsB1O21xW2Ry1egf3tfTfLqRc/Dj41tiLlul/bWzj1DnJC2GZOOI42A8vhXwe
rhef6NLBp74gzBbSEX/S1OxzcFSF1Vlb0GFI2fNJNn/G6cEWE7OyJP6wfYaxXB65esLqKeKOtAoH
5pXZ1ckdu5lou/hDti45YjGQE/WhIDfr3hInj23gewDFeQfRC8jptwilyRbZYULoUbxRkU2jRsn8
ERKnkTsBMOJkBttzoxCzLXLWEwn3iyt7ZKAsEEQ9dP/iABteAqCxwAV1pHOz2AOp0LIz/c49T1iU
/bbk3QEYmugwDOjKlwSbT6zKHDKCmJsENaKot4m8+u7sES63uYMHzxtKfb9XQ8YVkqq+xp1NNtbZ
SdHgipHnGC9xED4pvfFf50czFuuONE1IBiT/odHoTQaWnEbNJpKy1lcODiIzWwFgBvv+mYu3NgAf
wCA30PqNfYfX8+5NBAIQen4nH7ZNfWdWUln1REc+UvsvokbwFcMkGFbGM0o7CARzxq5Yw8vx2MTq
kyUUfGUXjHBKcDIjIGmaUvmtn1wDXJh0HTB6769NSHIecNrEWNLHp5IDaqpHcqL8MOqaN16F9jr6
LJvrVrS5Pzhu+Oq5ZDAwplwg9cEcOHQRAb//mTqstJdZG+FDaGz/11XtITr0a6EA8xUOEe1iIyMw
PqbMQSUeBUZCKFpU/dhmtavGBxCEP6KMBgsjs2Bjou+GV2XpEb7JkE9533JhClkIcmzE6VOb5Bip
+EEUt6pE6+tQQHmAU0aNpmXnYV4Z5cwtsoVnNV4YN/vXbxSO0mxqm/UpJ+5NqvyqpG0E6KsBSyzN
HDgYn1pX7OtFOa1YxyTFDmNhnXY0ZB6Gg3iKxETgNssfv+09pq0FFAZ+vq2dDPg6+pdDTJm6D3W3
DlId9ZzTBFQGgzdPVLhAsQvb9uWSq2h15Xpa+9sZzcz5wOoxIVWPo3ECkzNYXgRa54tNMVODlgxn
Ya5V4elvDEQUv8XpqsYzoqL+VlCXCWRZ2IAowZ5Hg+GiyaW4ItmqBn/PHqsXb41i68afRn34Z3Fs
Yd6YHL1otLPDznMjhJ5NY//thu07mi0BbvMU6fqcnGJQoCZlcsMmyorPvW3iztXVqBbVds1Y+gcd
nbagM5nswbSiz3pbUr5bTJCub3U4CIYU0LEtciFhNHrm2dYKaZvHhe58Lz+7VHJHIyoJmXzmCp5X
FlL3CUOZhVJFiKmRKFyfsmq2U93Efazc2yJf/3jd/57Jzb1Aov5EkyIlm/h2mdSr9CF2VShQgmKA
DIXGhmb7gaPxMWyiB6kTZhcQF9Uc6ts/6HgIQwHTCG5ij9vc4mrxqE4uKx4SfhO87ASGAD6s193p
7GsFeOwPak43f6Hey5dg5Au0WZ2eWJiu2CPtWPcgpiM32+t2CpbF/3EL3SkWkvsI6kwOYuBsOsLJ
HKDt+XosUkdYoIqkLYGTYvmFuHZiIKFkTmYJuZNSfy+8TZkA/lNEYRgHClcBF6MlJtggz2A3J8SP
HU4JayzLCxaTBRP3qFepG3Oo5xp0RGLYsr9/xKrH6jjBILTI9EB6cLpsf4GYReowfTmBXnj738/z
MnMdWSZIetcXb2y85d86zNcr2aB5OXGcJmYXHDv7c7ffwmapuP3Gdc6dXU8X5Jc1Sw8ljaA4tur6
1xL3aMx2QV2zfLyCVMnJTyycNk8Dl9eovOqhkH69MVMwAzUXygudBsclYKO51Gym+LVHGku8Pven
OSJsscBj4oS06JlcqZmoDexWCbK5OkcNJMa6V4YgSLGnztpeByJBK+W5cy0YmDqoYurUmxorrvTr
FmbsOPQvn0LrgWjVhiAOZ4Ncv4KZaMvh47EMJyLPX5ZAl/VKesfY/ZQiJzBQzkZMvzTl+dAxHfdu
+1htUKb0HWTpClgsA7sxwFjUSuYS/cMG15iwUYLLd+5EcVKkph3F4gC8m+hD4m5b/PljdPXMm+yi
svI5IEYqKvGOHi/geIKuZHxydRsGtDEJjZr8H1hLtdOewaH2WeToEJhubFptoo2R6+4+Hf3XvuTe
5FkmycTj3BzzSug5za/MM+WizvdxQs8i/5n5CjxviGDp9hD+YCUTeUOqGJ2aFRKugUSbAaurvsQc
Z0gF3WPS2gE5oqclqPI0s85xGkCLPCkbwWnrW3DCW7qzlXoMZNafb+zOFRKC+nE3tlfUv7V6aS/d
1R8M/HpprGfoMRqo7HzNoJ+Wjm2C6ekmgw41Az+MFXOkI4aLf2T7vX1e2paqMdGFocQFUjJePRBz
xrgcfvWWnLLvVQ7gcAo5zNUVJeuf35zmFgB9L5eo2ogqrsx3rpEmtiphHrEOwwGirrbjMb9ctRFy
YX0Zdth3E2GSYFhXB7WsVVXFKge8OTduuuGdknHaF+M2ym1t9Le9zocnSxv3Yd+uFbofNhdNW3ID
Zx6ceBh9cixDh+Qd8HpQDYHsDGXcsaegiuWwpAHjXVYubWv23ivaUP+TRiSXXDTzMP1if8K/RqpL
MCrfGHbRVHH/c4tg1//6w7g2jEGmH/0Vg8twGEIq6jkV23oktUmR5i3pU8RlUPfaQBpHrL9XwMs/
fXnkTekA5XzW92uokn1XihkYx+XKhbMhTzA+/kS+5pKliI8pouJMBd4M/4Ffdf1jSThaIk97K8C4
Dnbvq0yG7N22otVznnR4TYlAgzpLqhzXoShb9iyWfEQyrjBhp7k+tiA/QrZJRGAfSHWT3XmtymUW
4+1vsE0nQ7hBS5lM0FHAt/nemmB5gAawhCMhJwKb4dnR85vQj6uiNtbp7IgTbp2Z8tA0RHA0HIxi
wUR2f/jx7CudIsw6hlfLSJMO0Q1JqsCfN0K/XV5P4edEy0Jhu9rNQDUcmCrXd5E4WRqaP0LEHLGU
h6QEwu8R7yCTLEhasi1ciIng7QCxGvjzIb/KE9MNi28aXJJn7m79eL0n8semW6MQ/B/2CvaQHlVy
CpjpDmQTNAz7kbT/quqaoE4OnAMlWBCHkOzFSnTBLUlk/6o8OkgnTZ617oUnY/InPpJoYvTKwHBw
mDHuZ0yEJyJrellNSYAiVZhAlFWxsB0gFakYMUOLNJvC2k78kcvFg1gQG/76We62l56d/V3UN7og
RKmAEAJhDrVSgUHCxpqd5CbZTJ07bOaDwY/1wvr4Qun1veMJ8hsYrzvxuF+XhSWpYBCPmTVr54zg
E4k831pMplPZMPiMyLZENaKJYWMwPJ41e/50E6RYCoz3rDm6RwgbWDO4TpkCCA1rZdmOtp0NxhhE
touAWLPW1i8ode3BzV566o9LOl8dmi5m8Q93JaG0ccMFmq/vESfs8W849D+Nip4C+CMYc8V0t13E
Sc3b6wB2BLOM2lTQMQ9k0+1cj3l9jbokJr12URzpKUauCGkYeS7jN8UX/BHHW+Nm9W3/ZiEWgQ5w
rtb46Dh7kde+CnZQWln78ZCIdli2Q9F2ZosUSwkPTLNTYe/w57sQtk2LkJp86XlNt4NTzAlNGyiO
cEXs8wa7yAYcpbSbNC90NT9bRh/5oeOk9aB+chZijB90Y4zksAPpAqbznFEex0/qJkpVnuwsxjLl
9rD5rOXpGBMrKaTNPDQK87MducVJtqAA6BlKiBD8bY60R2i4Uvt44AwhPYfj3Ac1HIWauSJYEJDQ
GvSmoKA6f6x886nCjQobERyrjtnbceCqRxZc5CaO7s7igU7K6AHopGMCZHdhjH/IEAx3FavIYXdq
SxCCLINugVnab0fgQ0NHdZvUU8aQFuCCYL1UfhlgdpPbTg4n3hah5Xa3qO2pWratlHuLp4xDG+RP
XHEI1KigCDZsDsmwSIYDujTgXK83A4Sqxvl7B67/466fGu3vFRbYBWs7bsd1HcqL9oJP/DutW74D
W9+n/Q4J9SiCpXlknlndHU9AlcKXOdM0eoAFSKg4An+evgOf+M822dX7LNcVqje6+KCxGYYHSV8B
6bh74veitY5FctL1cWqC4dGpLUUGWo3/WaoKbV++cANJGe04BcdKRURussmPLeB3KbTiGbP0LWqJ
FBmMau8ifjQqiFWLZAVszaRY5I8zKi6uTB2t8c7rPHJ0LzqmrCF4kOTUTPJtYUofxVHeOhH9BCb1
UEwVvn7Gyfudc9opaHjbEtqY5+6y3gv1XcEgR6PEwX3BphkzeTjHwNsgmpR2taWp4zgttghg7DfI
Ohk7OyUfZUCoYb24+epjJw1plITNO8czGCyIG54B3K/OKiCwSOBNLMERM69pnSHVv9hJ8YMbVwGj
7gFeOmlI0yofv0PZlM/7SfYJP4cF9POL0jQSAS9RhvGMkZkfRl+IwvxcWW3sGuBDVulznYbEFUMl
gO361XYL0Sy7qv/oPqdoe8j54KhLNpQYvbz58aNz4yJaRA2lOUJtgjmMk/1NglyIvX2U4tiLaynr
zTC0OfAuLeBKe7Z7Cw0JcW1pldYVYPH3NygpbWzMv3RQp4qVNNyRIdCgOkEQN4froYVzWDFDbRAQ
Dxtey5iGZNelD2fKd5Fld6APjB8rPezc8scBEaIKxE1stfrqAdAgLXsbBL+d1DM2mNbO5JezcyJv
euC948y5mLZbwj+L4swZqrR4y/mVjxoEYsBQZT4DYbNH5expf3Rcb0EdlJypX5HFM3tF8AU6kNSj
kR4coOLI5bt+5sjpjoeRQkRZfdyX4rlZhZqhcenRXgSGB/hKSODw2UD3qJ7aZokaJifhRkLu7gW/
wdEOL7NyE/f4Fhp3ht4BKd1+HWI4GKRr1hOCQFa4rcRhQVqW8X2m/MY9yHidWU6E0Ey4wj3ngqqT
eoUDBUPsmOWIqRQeqT4xud/rlsoxwluqU4d4vsZgUk/XQidOaATcrjLvOUKwDdOPdih6WLp9N5NQ
s0TAq/y4d6bGUq6mh4FvnXKqghg+mGKOZ5VDMcBdj0LSkfufzGby+2t4tnSZ7QmK/k4hBI70ydL0
Uu+QN4LAa8H769aatfQitmjaFf596wO+AqydWf8OS9rbZ6eTP4cphrhjejxNrWjGrJsvihWChulh
EDxREmeTLC5chXWQUeURxxzYa71E1Qi/4cvJveXCIjAZJIzQ0tChy9ngjYbF9a3CW25hyuJw9gDb
T0BDiRyBx5xaPoM2UiFQ3o7b5xAFu9Ibevhy962tBYBoYFopdg3TbP141AIsNenDcmPdn47P38jW
oFRXzXRj8sfIj46CAdL6t2AetPSMokXa3a/r0ceoZ6xPk2wPGcoPkXAlxEq2DQYE5lc19JVE8QcR
Eh3UTMf20jaimkcKHmoivp+2cqL60+Ra4V8ABMy7f+0OsCt5tHgO+Y3lrBgjk5tFg5lqTGeU29vV
C8QyqcrFkgdXzaBUEpNmAnotfwCA2QiykL3M6GxDQK+GCl7T3cekMD1hJGHlCi++ZnXxoAyF1FOK
X/c0Wje/9k6Yk5Wit45Ef0DUjKCgrhkxRfAHJar/OlUAPwKt/Y7QjgYFEskJ6skL6TgGWPRzjSpG
v7B70oZmDgpmFIOIPxhLnF2D2IoNUuGCQG4oy26yGqW8GueVm/wF2c/gBFvV1fSoG+EVOrI94q2E
uNUreMAEpaorpQQT0xI5ILxN1vrar8g/y9jBkBU5JMRmrGfoFdO54WLvXi2LCZkX0jpe9Rx2SHXN
mFOfdLnEey6ZP+9LhKYI7JR+hAOd7hHRLQFfs8Wan1p5c9UJx+H0B7AP5f+UckOlgknc0B7/mk8H
OypgUGYaXM1EKUtLU9g6F1Aybv0YUzLzXoeypVsWeTB78IfR3pU+ZOgLBQEf5Jmen+lvZDu1fwQd
qS29F5sWhhGU237J+y1OB4rABHC0IoHLw2PnmcIBTsfWJDaAFnyHYNErZTyPj8+317OsKNE2xdVb
PtHbRyZPjky3i+tn9uKe/qJ+8tABetGmFqTSxxELqiVg1dDs7hfkeR2qxKv78Sfnb2U72z25k/DC
yn/Y980ucDctftQzIM1plzgCCo/7FxoL3glgGtiuCAm9lQ8DlZvEqpbvBbeCoRwB0FmihIVN8L+O
pFmSpFseko070uG1/5rs5hLShVwWVJtfAqqi6+TNec+XDKAOP4lzzKzDNfxzCe8eiVaKGn2ew5o2
VysxuzvV7b5Yn8xdUC6Q7J+JweZFpfOdsF544VEsrQ/8+m+FEU3ut+eX6oPvYa0AuqUh9DWdRJbL
WvlSOOjHNxp5F65Hs8EiDGp6Cp2i5VjeeYKhoUtpo9J7W8i6JNG1ptGpm7LbMIfvJiBqtZLj+wAY
mES1wRuXe9cSdI5fhT/TRt95UCmxgTc7kToPrNjmmVFLD/ReRRPV8CF1fWMMbPX/N34tclykDdmJ
InMb+e36Dv8VWwsDQeUUV8nEhjH6626iyXIuV6goNW+vPx6CJfJPfO2UasoBsPJvCwtmO6BK/gf1
QIaINlBfMWQARxuDdrz/n6Ie5Im4ulkOg/ts4b46+Vq9xuGDGuwdK8fn/lVLfzvdACEz8z1uZ+ga
KHYTbIA8WK60KACsWNtTnw8E2gyvYxzqxFZp8/aiDfuOzfmjxjCXN52TZhUM0lVsv7QUegR+gzqx
ZNt5DsfPPNa7/2HnhdNy2s6rmzgwcqYQTs+3VvCScaxNFn01D1hfqrqUUjUMhnSIr9VAfEfY5hiS
s66D1Yrwqu1lhRJW4nTmUrYpfzxqro/hbAPyN6k0w3mmO6ERGRXFearPt3lqQdO8ZyhqbuBVhJQu
+GS65wo5+4QlinLu1ZQJrLguNjQxts419CoNQN+AcpK6BX2lKgFZlOnbtai4B3wOGqkncdi/sDeZ
yNNMeeHIZno9z83CBesfKEbIkmtRvP1L+b9pWANtdnTKII1Bf9R5neEA6TSixbM7BqdARiBuxT2G
E9y4t4bHmZn7ZsL2MqgCD7QTYwl02Dq2FBIRNMZH5Ah4t17q/W2x9qS9wyUmY/cqGQRbHBXdA0E2
eDqi5VSQ1KNwYSm6HWRMtqVJ9Xvb0WpzsKrZsIgfUtk4JTjAmImm1jUW4DzhgLE8YnpUgPnrxftW
JYYEJpkryCEnPZyBiotQaw8YZguo2ytdVuERTNeAa6tpFloF9XVhgOKl4z5qkoCt7WRysfZK3o95
5fuL5DTmkZtQxePU3R5RUWD+XBKDBsWx14gY8sCcSGH0vcbRzjF2WM78jok/p/UJtySZkM8Hs5y0
QEXMvXRrCUD9tphgtU2OG+glYtnKR8JxKBYNiKdazL3K+/qsZEipqUfyLPOiqN3mOVqOLDVfEizp
Ow+l6P9EPErNu3t/ISU/T/G0PaXMZz6ZwT9vWFsReth4LzWkoCw7jR7RL559leEnpgXMZ0ajQ4Ib
+qdCLu3wC4QPJ6AXGT5tHnuGYEvWQj2rljOu3yE+7KAwMt/r54jQuIy4yQYewO80CFQaYiTtu72t
I+EE7TtK8P0r4jTETsLO80WSPMeImOm7Uaxfq6VnLsIbQaq6lmn4XTFKZTWW+x30luZOC3b3KTwO
GamtImTjiDhqQO1K66T6O5x1vJLSJzBUwHGqHnn6x3aoZYetyG2QzuXXW/gfQmGEf2hL8jNnOAIZ
i/bwx0trsmwl987zu7LudmRpW43R+gmc4WdyOePtIxFudz1MORQsJT3SFJoacToq8K1+jsZ1tezV
9FlIPf8jArf8+cPWqtU11Ajd8UupbpqTDuXMzuBBAvHdHvWBco9TERVjesgb20CjW8QmQa03Suor
4N4G7X/ag8YoSI02OHuvli0pBkQ395lwF4Se4eBDeS3SBOMJDmunjIeQ6tnUR41NqAwO+OwD56dW
YBZXnFIE8d3rSgoMbN1evBqAVeIzHGdlaxcrNuExfy2P7B2wSbqM1UUPLeKe091foKGf95e/fitF
yDfAnESIJlOpNCTElZDnl9rukR+C+48u7n5Xk5D0FCse0TPNpqQlJEf13FB0ZgLOXIrcFFohi8t9
CdhHn5jkbdt1AvzrI0AvOczQvErDAYCHtDLWQ6OgKazOUW+e0Wrk2xjr2jX6w6xqneLEbGEWWusC
i5Y0V1Eqs/p0Yi2Mma+aiS28H/90x2ho6r0zcZPLnm0PgB4atFdrrdm0Gz/0xsauJn2QEcbdCWCY
IF6jMmpbp4r65Wg3oYVx3jGDXSnud8Zwd5XGaSR03NhUTVc9/8RpTgI9eJHOhQrRssbV0XADhMRe
nnzBEyhCKLgEjgsdyD9tilsq7n8vUeq6EUpTFm3sxeb4N+/8xJ4dPLA2K2L6+5WRYzm2T3GcV8m0
h9PMTunHX5iEADzPXeAmTmWMJept7ZYeQtswIhE2mOMmx5KdId05xU7BKrOcUtJPZjOvr6a0/9nm
VNr99j7wzAkDLa6f/GUG1TMjX4jMeZsYVrWUs1H4KuvG7DPmC+6iuxnROzLxlkDl8TT2dm10h1MW
i85TLuby9AKEj5gsYx6Tvd3rvRYlobaVg1IAgmSBzdv7sE6/SnuKPh1h66v46UcEZH5oLR+Grmot
R/eMqZxKHH1Rol/jWBlW5i32GVe0VwT+xe4rKvxjJDH81IWc327b8sX5a4oqSixrKZE+BWIikiII
nYRWXIj7cB6M1zTTTk1Y0Qj+8seVJU5bKnIFJdW9YIfKewOXSkv7SZKPHgaEI2x6QeiRAHPnxHAQ
K9AI67cn6zDPkUebhj2bsIEClJl+hz4uffQAfvDF1O15YWpAgG8Ix3lT8M6zI1IhIlQO1jtM7AOK
WEm90he3NGgtbu1PxtJf/uKjajdKe2WOu6N2JWlJyGkmCNH3xFT9Bwki8Dvqn3mqjrnKQuhZ6Q5o
IjZdLd0PRXwBFKqMt9Ij5RYpaPick0cCJS4tEfi7sJCyebcJq7Y4usDMmPs8NkVrXMpW/caNl+jo
Xg38hYlewthxsHwi/lV3MvlHgSKEZ1l+mwOZtW2T23Agz1q1ZpwqfCoGpZVvjThyCTjAlnbwmAiH
sIDPGvi4nqAgcn6Tn4B6ARcTPUn1JDNvTE7eAt69ElZeV2xx7O18FUlnc+2inwOeirf6dYRwM8j4
JnmhtuXGsw6Jxqhh8r0acGTwUvFn5hHeap6O7x8dTUN6/8imDXA+aTuO/R25oa/tS5/gN+/fUIIJ
Zvx+pmYz03AdGHQPtrGFXktr3HIHjdXv3dwO/BUFTpRPxfxqX7betwDAUFzf446eXFq9U/ZfySCx
T3kh0Qv6gjXp5ucgLXrUWLbhFD71a8RlNJZ1YO8dHmlA/Wggd51h25O74WIcgcFXpRzblBTb7JxB
1aivD81SqVANqjhMM5vvJhbk6KCS2CNV99ct7iRtZPsXb9DIU5AVuT39ci1sMxLDVA57zB7CRllf
e99/NMwpOhclCIBLU9pKNiJRPSoiKQg1CkSbcdac4gtVAdjWviEDUDYza/SXOrha3yb2Y2ffCMKt
tOrQYY23pJgI5vkpN5jVShLji6TASozlm6UO+hGs3gJacoU0m+cS+IQnfR5Gy56dmCgMhqSOrEeS
uIF1Iu9+3+D9AP8bb+tlfOBXXcL8T3lexssrAjmstkhzO4NmhHbluqv7FumKD/5fNWm9u3Yf1ZkD
7SQoInPjNvWgCiNemUfavTcehILFqUu2W2ehbGs6iDa9OLFXl+kAZ2su6zv1VabZ4A2Qe31YHPzr
O4jyMWFDUtwsjB3rF76vchiC05ExX9DEp4bKVV4zbpHL3nKRsBD88y6fr2F/lURo6OcegM5ezua6
bINyLRTqZzEXzAss27wLZ+w1Erh/QWBLiBqgeeCDLD+Ic7HPJgEYvK8VOxPlV+hht8i54jt4VKNq
+IXYlQzwgnyqzwhoVmvniLpal/tBZ5F6b75X5yVTnZu5rnxsc8jCg3PZi2cbm5j+b3q4LJZtS/wz
kYLbgRCpJN+iNl2yBGivPlw361fv5R4XIQ68CbIbm9fn/6i8hjtNDS9+UCYL2S/3OgxD1C/NnWOY
j++q4BSAcYa59K/w4ZvWS1bj5VqfjlbL9pjJz38LwN78A/PhX66e3dw1asJ0Hr+UOAprB8wliXH0
KVqUK9IrhTm8PbVgvXa2yd5MQMtOa+OWIAciTwlYNMslrBc40zovd18o/Lsbtf+WEv9XqHhpiDmh
Yrl0aYxI5NqzeENXzaLP/j/Kcop3ehrIgg+MHw18+xjFvjX0NjsVKMqdMVfuXV/QC8GJRs/olA6d
e0/dg/huoMKGxeMfX1DV6N1XqgoL6ToDpfnPkC9YWrh+PusJX3Cwka7lXCTP9gxZxETQolD9XNq2
YxbhFORpSoW6q4imvcqrPIPgkqCBdGpHdRdhWa23x6DOz+T47wVZundGQuwQskS2Hw+aaGsiukHi
O+uSWBtU+V9N0+xTm8pg9thf66aIx/nWRC2w6n1zlu+r+sN0N0Tf0JLy7cZj5aFVOD+z7A4xajW1
Bx4QCDRB8WH7utWRZfo1S1CV++OBxkvs9c0MzYZcZ4vHAsRUOESlZgfDOcJY30UjtR5HuSaddg9i
A4ARDE4hkMllptzIPx+vO3pM1A6d+KXHr+fYKdeyufbrfY8mGax2pyGw4fyTWIYSmsTQJwPoyUMi
0OukTkXQVaD4P6CC3bwSkMyj4UaG1KmBbROYGgtRgDb2n1ZSMtAHv+jyEYjjcJsLT1HXGM49Vbbx
Ke4ZDlCbmeOmID5EitjMS+v1Dg0dkBG6Z0EM9c7phIg6d9s3uyJ8P6Zp2GTzlS81Yj7g7vVpkq4j
9lFczYLDTJxhZspSkHrhCxDCeDQ0rTmnr8Az4GTdaKsMW6CEyNceDJjVZjjL4Ec7sccNc52ak5y0
jQW5w6nWBOp8i/ZKgWdyCDdnQqlx6e07Kt4ukj8e3hvR/PqXp6JUwWeq1++EiZA1Z0ikNmIEE0rM
qg/f8p3YrqySYz5etOo+ZlbP77/O7Bzpvn2fDDqYa+ENtqiYN3ZENudTA9poFh52NNYD7S8rySam
IakrXCDlNa4U0jd+O++7C1v2PkfO0dQ2kJlCtJMcM1ULygRo5HpOCBH4feDFCWNFGYEojE6fZKQe
/TzLydGX0NiiDGlHLZi/VuIXLaRrP9/37GDCfn6JqmIDwGOn44QD/akjlI2ob6kKxbt+WjmIfwtR
yBmcUyi4llFN+8imqO3z5si1815TaHjmIRE6S0RnSTJ6bnDCGHzwlU2OdV4VRRmmxoGc1Qgh+4YM
S959ia3cmLJewOyb/uraDBN95z8O3a6XqP5jkreSGxW9kWVBKwul4blTfjxIU0e8OsLR3CTUynZ9
v5bKOGymeiRkBcHSThhKOOKepO7DcTAre9EpNpk2aQHHv12CMLImpxIlmN9wVF2zwuhM3DFnCab2
2DYpQKow0zzjaf13fVij4Q+TrmDv3p+JkUAAkSG92k9VNVGVsGQeXZsI5BVAe7g+yACm/O7IP7Pz
MHEwwWFkEJPvtO+USomfGlYFp5xrbh1bXH/c0jaYNk/+FcSxKzEvkdn+zQKhnqC4TcSn9mfdLqMw
dNkrc0HuGiOcWQokZ8ISwzei/GkLgfFnYD0omqXSs6MxuDZydJPt+4jjBMP3k7oTuET6LMyI516B
sEKlhwgIyyVCxrEX7TyhafUUCvr3HpK6YjM48mnXKNXnHxvVwcvcMWTmZZJ/f5lEKPevmaIRlc0c
ij9AA51ElEYBs4V8ww+f6Du2rHGevYtSaPLRumhEDB3VJBrSbYv9ahsvC+jq1D3zg/KLib+HU9Cb
ePnSEOZkfRYgfK9sScjFzsmV0ueBffZ+GqX/LNKBIqc3P8gCHGZLkY5tzNSdfTFr2e7IYGirPrd2
i776ZzsqU+EIqXDNrZhtR4Yik7YK9sf+Ocfp7UgmCdDhEc08VVAI+dAnZ9vhaXZ4gJV0ZxUijBiR
5WM7isCBVXr+BFyTViwjH9DgntDUNWBIT97u/SyorPY0CYsOBbjQFhLaNqKmahEMVNwRwaM5POAm
y3gjG/YCHsLGOqRwTvkC/yRQijvdOBAmFJz928Z3rBmgHbn9NCdLtpMQGjtRR4BOCcMO17X27XsB
4nFEz23WvMZQeJgKsge1ltgGlFEW+fmH0isSl4PSA+ohz3WeEuvqUU8g5QQgTUcxNkY6DnyT7FOu
B156uhV/umImtLNjcU1eFQ67j2CH/Hb+tsm5vrQymuc99q9+7/OXmGtPkyOIT8OWaRJaxN6TpK5s
xkFDlcWTxorPwFHmc4Zuf5tQcf/CsUyZdQEawNdev/i3e768KNHOz5hKPq9HHjBsHkCwR0xpeVlP
lQGqu17smP8MMnPh7EkuuLkQ9PsEDCnuif9u/Fdsk4Ivw/HAgwHK3TbygA7FBq7Qf92SmU5tGljS
fHhPHWEgxeqGV/Dj4MDuk9gSfj5ycTxzRBybPpwQOPhRk74PeKJh3Xw8zHcBpbvcAriYvgSWL0C4
mYc3oFf80V+tqh/ZxXkbPC6tVbxt6f8uTitB9hnPELQk25//ZAj856VAfLrhIIwJZgJLoC2DHBEZ
qfxhWcEf4HI743Mz3RTMLsyuuHTgzOpDXgaWMk1pYaBTUkCPs0LbkWrNS8Ui8iha05gzxtM2kYwx
z8IY0uw/KT6H8+Io9aI1lXA215XhlBXL4ckCRfhBlTGP3iCki5kXEt6xN6W9/hBCURDRzaEje0co
VmXBxk1up9LtkPrqO4E9Yi56w9Azvzo5+ULvKoGsMVfayWyI92adKJg7Ty4ZuowDUMt3XTGSF2Qs
5wXVypR1y6LNYznqypnYYV2kn90gbb0EOv1xemWS5dRizgKaNZL8C9RqHIuXqHR3WzmEhEq9Y2Fr
lqyxRF8cE6kCGYHV6eHvouxweEtPdO+hBTaPLEHJDfj5rXEgdP3HKDwtFawv/5Ps0LB/5IhEV9JB
31puFmKM9gVK/auFs2PSATfSwdxhDCH6RyeRTCk6IT7hIpaBuIgQSCm+NYIaXrHnEQI2JvdflI/U
hhMMwOr3jmSDmhSgE6mT+00J9w5E+ZdnrljeLdwlsbk0PQOzxU/ETz+iPowD5UbpczKUGEHCfvjI
mmBmVHh6z/uJjO4QP4LMhqiNvC2wUnGzJtaOXRDaDhslvTGBY1JpwzWmBYz4Vlr6Y/A7CHeo/B+F
cxLCPRwFUJ+7bqdPI4ws+14MtbryRr7pXZRRK5H/HsOVmzxbb2m+vjmAbVE4nXmANHTzv//4QbvT
zY9GGo211MBiwtC+mroJaEn7SjQhIRPNG5v8X7AsWi4JWVFIpXFQSIi1YdWBtUF6pJ4XJSgz5GDE
qjssLYkMzV9cLUsVj2EplN1owkmNTMIZo7L6yaywxfUdNldlJmj6S7AMnlrOyy0OH6TgGXTFXTpu
uXUzWftiC6EGHGrKpxPUzxwlNq/e3XER1H2cDhYfEcv4w3Lgb7l+WRuLkjFFuno41OjNg8B2Vty9
em9X4bmZBTpQiWCh56lbz8poTT0rCDHWJ5YskZK/J6WPYrpyYKDDC3g1JtTeavDH/B9Nwf8JYks1
7uN4L/qELFjmMKJoQgTHKqs/cVTSdZnkxv1zaWASDLFvBTsqiKWIQt41888VfNtrhRpKwT1mC5kt
rgB7q9RDPNYE+jMKPR0aoeOiOQQHEGEGLyPvgrvc9qm85XHpKw+QV/54C7LnbGOHJV+j6GXIpwUk
N8gCDwNpEud/l2Hvh+VNwNwm05xqfpvh30R1u0Roh6wzfUVaQFlDFddcJeRp5jKM9UCxJRLwx3fP
wxAImcsqsq0aBiz6i4s5G/599H2+5l2i9M3yO8zsnJ2BLmLUyRBM6JnmtDu5GHec2ltkX583o6xP
nQnqTjxrFI1VUjDGvpmU3xE9QEvJE9U+uo6Rr6hJmD7YxvbFSK9xoXlG6hBTkzSs2R7SdMEFNSWG
Mmsg5pqNS0DbCgP1AvbD49TYkkdYMU3wqy09Cc1dd3eAGlxuq1eFtqQrQ/TS+vWmXBe8HtDrizDR
Yc+2e4zqHOeWMeicHU0UR7KCFbnO/2b5kR+5ct/oNMK0vekPOjUeGuvcPzLwCCiXivcmbuIpSO2D
cOMyU4RMwqKnUsz3Ol/VP/4a7eymeyuWa9JH7VpulKINTtj8wPzEhaUIJfK3vZrKKjXAKu+RlnPJ
eEKe81t7zgFWEPoL1mB4I9CKVu+uPR0lVtcNnVZl96pkiTkrImrbHax/qFzc9UMXma+xAy0el0+c
l5cyf5gVcP5HXhOswPx2pgYGQUO5ka0+iuHorIgyhgDEevcyy6pYuDr2j67u9Ms3CCWZTgy5lvfX
dNHcIRBC9++UNpwiNQpJqFUV6e8TSjPWNTOmQSC3GYdD1SD3RL4/5eGdmHNXfsVb/8jxEXAxDb4Y
Nd/yH3in0VblojD5Eu6MVz0JQdwHwRvC6f2Ipji1aaxa6INqpLE2FDu7FW2DZCvQ2E5hFs7LQDyA
Fm470UnZvBMBxk9zR2nEH7p/cxXD/olVCfIf1qO1mOFy3Nompdqmuk1YPYeZ+Ywy8w0LZK9FTQNQ
boRE0ytvwILIPBAKOGUnPluMJsnraS799Zg3W77VbHfSXSEfDPtOG7vI4S6jx+tAaxzDatSvhr4x
/6FEez8YJAo03p2nAQllKu8Mm6xHd30i1x0OUJ8ZfEmX94wWxeAZSkhdc0lIJObU6jd23y7N8A72
8ab+Ro0LZsTus3Qdca5h71X9tms/WwMSaTawhk06P1Rs4wj5Od7hsSXAFO4mro4U5qK3MrZ5BXRj
F4Z00FnwHvLYXlEeTMbscuBq+n8iTiD/32m56+dUXIljWMOU++bfxrnplJ/GyuhaTk7I7OVxPZ+B
1AW3lM0QldZ+zV/xtp7bGKc2VNhoTJV6W+iY/okcZXjrny4fMbUfjcBhuI/gks3sg2OjnAJO/roG
hqXv3U9YXsCWaLyUG6OXkjQMBO3wXQEINS5x2BKBd38YiJV5dlW7uugqljCRtr9XXNB8pVIMgJkp
jSCfvdR/FM622VkbDeb6pIe+Xfa5q0QFQn8MpCh08G/0Cy2tdxXUReb8i9AY+92zTD/la/srBLw+
HGnADZ44+K9TMwWcJYquhk16GTKgIb0H91pqgja67tEe4DDcCsizxw1CKBgwD2eIOvExF4Ikghmh
Nj8J+8nPgVDnXZP1aWBktXm4Bh2ZkOHr4T9k/fG+uvlup64uJX6PV5BZcQhlwOXdMTRZnLuOdCX2
nV5pSwKS6bF0a+c6O+eTBYbmsW3AkaFSzJdyomD4oNeV+mcSSPGmpjqy/wf1vRV3JrjRhLGDBliC
VEztwsLAV84AP26cHXvdp9qMmM96/MA5vruFAdnDmY06i99n2GKmepTXweDsA4b+8U24WyTnNag8
2fQ3BkJr3pt6DbVY9NLL7N5P5YZrYx9AM6UXQMB6nt4UwE93fKu2UnxFvS1GP9Aa9BlzxrRN7Oay
z5rnCD1YdbY0ZdHD285zG53tC7CJ8rV5WAGqsGgagDxL5dQ9rp5wlkdGj10VWQqJFp0oLrxwDyHj
cxKa1r38sV6pqaw4D2rpY9/Fyf9FUg6HNZLZSMCDURoONh4fhj9xv+XD5jbZSD+yRZykFg0cuYR2
PBVivqpcTu1+YhLLtt3B2HCHPL3bh5R2NdfCp8m6vf2d2mbfg/d1lQ5jnLS0W4QC7wWzKniXKRZp
gJfGF8yjCdNMqN2BVGyr7rw+6kU9V6YR/ag8q2sKqFYmdi+QEIAuDrA+wtOFPLpOWGE/xLEu1GkA
pGvk3aQx/eY9anusxhyPdp5FNTmawkjgx4AW43ZuNZGjvkT+uXVYYrn+XI5QBp4KKkGjnfdeamir
411a4m5c+CGZ+FXtcbUXANqhKh+V8+JEyZqLKDrCtkZFCqD1Tt6N/96KgYFSPiC0RB3GcBW9v1Me
e6yBgGWx8CG8nT+0hcdoVSYAWOZ85OFHBfheupstPLcbrAXYLO9oiQSX0ER55roO46nE6W3i7zly
E7DZsUS+LuQqzHKcU+lpc8qh82k2MvXmY8+4xfjcwmCxUYQpLOmiSpyRYPlkzpHo0MtvPE8LOrNo
8qZDbWiuuCjo0sxZujqhYV8Ysh3dM1ZdXVxq1jXA3XqfqLy2xMqkNU3oY6o6rex2HGjKcFitoM57
+FYiwX+RR0/ZLWQ9BVRr7O8+aUT/fqprFSOGVLDRx17THVD7WtSkUT6F2XhndZfhN2mUTkXuoxFo
q8/XKeRVd7WbD0WjE/ivtaTRM+5t5pJQy5rYwU3vYYBUBln5ykZIjy3cQJ/agUUSTE2yUsqe7088
I06vKEhLe6DvFJGMILGNbMMxhBQ3e3a+fWQvj7i8Ulr63+3P9fTOQB3pEz/fLyTKtvzyriqmFILq
x4NmSN9yJU1/7fHT9fD1v8vyQehzhXxW0r7BsC+peMj5uYscUOv2zz4RPSzoquqiT7X3qHw4oODs
Vy1dAfqFI3jyUK8uF1BES0grh54Q9u2f2w5q/0IPA36I7VI5SVUY0E+vJ6e1+ES4ALg0b1C+ABP8
bBybLgkPreIA2I/dMYrMF11/f+944ZrhF8HnzJfeT+S+dNhAEMUGfI7tbNOJq5FaW+2xj5z1fo1w
SLHSQ6vjoS1jbi3plAulB2PZAWHJZ++Uzo08quf7mPjLZBTxeS86OU5nsqtS6k14DxeVa5VhnQSe
BZIRXoUKi+nk5rYD8ARiw+JydYgNQCC3itnbSrV/cBVyTGQUeqFibJIxIdZE90RT0lisLUaW88I1
ejJKS4o96B4yvHS5ZsXpV2otLb3dt7ZOfTB+UZNTdtbVqx05+3YXMSW1po85WGI1NYtATz4L7nVj
s2QUbKQQjGrUghx9xDvGxBMjIw/YyJVgYrKXxgsp0lKkikbs/HxM3q4Uj7r2a3ASN6q+WErE1JGQ
/mQtbl5FnF5dmzXIkpJKIu5PmnlswC+bk10Ccbl1tangIGTDbKF8fsFr433XoFJJNy/GdCWxPjBY
Lxc+x51loY4T6EIn7lQxTMxWNOgjhaBizbgmhXn9dJJ/sketd7iAT1LHTFvZMHDsiRcWCKnibRvJ
ojGunRmtaASwkgcaGdFnD9r/u4opWbJaVt0XW5c1N+OULeUtR4Cqpj98xzVCxdUcUKJx8qAjiNE3
qFmMelHvMgp77eXs1m0G2pMhZkW1y2pIIHImG1fiiqiowBxANctq9g42S3INjwKlJlEedh5kTffG
P8Qyjrn1Gjx3w9QyFnfVjFexJxBW574F2TBf8fjIW+V8uYYiUe1GWAgS5PNzOPPMI8Q+NKgajulv
Bg9MVahDe1XP17PpYZhjVN41Jkhyz/+S+weoeCZ+ask2N1xRCPm53QFfwqgspn292vYwOz6OdESD
EykM2HOWmfwJMhPFFj948wPGch4Ti7v6TOMjJ+rmz6gd0QVN3LYlQLQCcL2lNfuxbs/SFNIrD3gU
RCCPLn47GJiqmlD/9IMeTG/B37atJVScl18p2OA/r3g4C4PK+oKcjCSuUhAOpLciNMi2Su8dLUwl
v2wNLvB+JZ1lzoHMGEMeRctth3D0ZWrmKvYNRWpcPlK3v/IEGXo7H9elf/UaJoHcJQeTVrgQLH07
58VTFJXDSRUK0C7R4LZPLnAx/HNhyUOtDARRY4l+m2jCoSvu6/waYxUVbxlmSlnOC6KkLxGFbO8G
xm6O9g1jiRvnUOfnN8BfLlyTTL0C6/qkQbyDaumm9vLF3CXANwdFEbuEpVWN/Jzrqrmx4X1jC3Fr
e01Z407NqIrWFrhSNtVHt6QoGP2cGJPqVyhIuTNeK01JW+fh1kNYhoWMwQF934xU3ObBSQKc4Z9T
+qMOuLI4U7g5dkr6Vf4/RTUSANn0B7TNFExisbbxXMIl5SEHdjm+fZ56crPfRCtj7EP0N5+CbbM6
YMeYvgqyw+BOsuiea0ntcdUkf/pCOeGpmfQVzdGvkjUTbFMNuEtc6kt6DEfdyn/l39r0qgrQOlCR
xNAA2ME20yUcW77myWPxh5FlCTs+GgJKCW88YF2437phFywlMzBm9PbWrELTD4ohnqGUlCFdSlBq
AnDr1HvNA4SMsRv8rOwarKoNQMZVFXlaKFdZTTFn2PwlZ2ZemT+vL4ktPHGVE6fqQYu0mrWOKGrw
ftrImJmtrmWghSkGrkkSHIg4V+Y4X74IUixbieT/02fymudWqsP3wiapMgYBui9StgqIOIjP2We0
sI6h0B8PqnBQts8nt0FF+7ehYZbwiXLWjCNKHNapCiyS8usf0GT7jv0jx/KEQbtwu5kaRWJl8IJB
V550KT2KyigIXQ7k8CibZg/o9qYi8BLAF/oZEUbPPGPTsCSJjBrVR0TwnxuMCb0NtMsLaBWoAzeh
o1Bh3gnHPbrIryNHnO5H4lLDR20WFrzNvb2JCvWCWivsHACJD2YJAC7k4ShlZ4ohBfRj0hSxPwiE
8Vn5LAVLB7OimRIZgr0TMXqmpRIHMz0oWvLq+Y5ctv0oLm6XvG/rpXau8x2/qGxxthKBrS9ydWs+
S/92crVvLFcA3AOn457Sc8d08tKtMXboonOkawh01RbMKpZmlWn+4S0TOMe2bb6JUZYp9mAXAOlf
Jr/U+BuESHV+CmC2LTbw4boOWhxQDPYBnfaNEIfzFg7farNnf6VxzisaeoYawJya0tXqrw3uTeNK
6/AOz5EkbA2Mw4xydTLeN5IdDqf6oaWZUXTrIUHN4EGgs+OoOhaW23HEd+UF6cPK4A8UyySXo9LK
/PNyC8phMR8AOJVHBz7LoVDUdLqTH3h7qoSmgLmnunFxy+uuIHomk1AvTQ+ryp7wRtHgwE3qR3/p
/yto2SLQ8Fj5WodL2j7ZyOuf92LK8p3gpRbczCBJtaahY6l/wVc8RSsIGqR1JbKVD1hM6l85a88r
Nzre8vh50oiLM7PuTxNAiVKtAzzgfphP2dmkoiIY3vrJ69RgHmx2r6XmZMkX5uzySdNXx59343FU
Piqtdphhuz9rumCeCuaMPkJxNKkDVmjCI5EnYiHftjx/d5gSx8BdH4T1DTxradY12+JJNP6waR1G
jTeFg/jh+TOsRHmePLzDXg2SUuRD/bFK73pkYPPYLmdvcMCkSIdotTsaYvxtkJCj8wcjfniTsr3I
9hSD31zYK9z0li0w7hHzNK9OKzHnuEi8/P8fAPwP+DqfUMVAKPSd8hQqSI7jHq0c2Pa2WvhTXZjg
GAxckTbvLi3AerBm3QGbDL85m6sGGIiJRXkLyj4u/51quRSAxG0Hd4Zv75jahTtF7yHaIBNVhlKp
fG3FFa48T8hsT2ULSHS7GLAvSmlz15kSwJo+5yq0C+dYkpshoCHUoVTb8YWjXtMRemFr3kUisXPV
WR5NlUmNhJ/b53vRVHog6/iSvzmZTNNmR5ewkqhz5AU2ZfuBT3hLBOTzdBTU6vlQJncYBVUoB4x8
VIdduc+xX7CJ5rto9bbADXQds+hsGfH6d7f5aVIxNb9k7vyBcAdAo9LGxeR36lwS6xJhrv0IU4ho
M2GiwLwVUkByuq+EWX/u1VKyyXx8cWW1CTl/lFSX1VcZvLIBbyZv0e4gTj4N4hbB6ypt8dlaRmbE
La7ivQyypv4kMfC7sPXvoTAXuzjJxX5IdZ1l9XiRqDbONxWQAhiyKlHOweKQkPGFhf2NyDoYuUJB
U938Rh9xdg1Af0OMNSAU6pCX+H5/LXKvLqB/dZoUBQyFNuwlks2RUJnrfpllAK3+h+knQaFO+c8K
q7AZAcboNkeDEpTQf/wenRUZydUueBQp91HJXQXBH2tQxMJfpTDBa+H00MG5zOsX2JRmDtih02Um
IhYHUs6Ra33TCYP8+oE1a/2iJPeeIJRTNRFpk1HPAzw1jpv6ZLpkLf/y5z8GJxJJaeehjG69eZLE
rFMExxBs8JyF1HZj1x0c+2vaifmBjcli96PvXQcd5DUZtvVTgNsKt9lN0gzgsN3TK9c7lBebzRiK
+OnsdgOA4WjVHTxM0H/wk9AkvKXiJpxrBrc3xNsjomUpctcTRIlVJ7hogqNZFTy3Eu7mtrbv0jlD
NpSW7ofT+GiTnXIiXyP6KITYsIUT/fwecYPeASFF4cgvFGVHrL8f/05OZK8wXvPOqt6Cnduc5r0G
0XfqoM1cGyqATNYkH0VumKgpvfW054H+Bc1efqXnMM/c5K6NuLIYNEkVKUeABwh5FV9bznxeRED9
tOpr9cxduIzBbFdMwZUDDCfO+E0Q05A/CnQYTUL5S3NJpOmMBCh3cCFXNgSikfwjV3p4Clnd2IRX
BEOOUoFg6OWy6E0oMJudROnyzzATIgHuWArVpsTVY4eheoJO/tWVW1B+NGSmuXyleBskkat9rbB8
x5lHkO+rTfvnx8PvgCP8fzX2dSMzrGuO1ES01M24yuDu5ekLq45GUVwfHOpw3Rm12t5vgSRxUOpC
0M6c9+PUpGS6v5qkeGZHjaJNzXuzs1ZNntlv1BU5XFRgNTtmoIFAeTLQc4qR+V5D/FhaKOavumeg
OhCEgteA3MRG2Ntl5pHqz1E2bhTboqmy1+ALWNnCKTeNgPbw6oPUv8AO36iY1oR3OsRH9IZ3/WMl
AHrUsEVPhOsfvkUrGKfsoy/28NyOb7dqgIaQrlWnJHVZkiodkUdZt8+M36vwLvOiC6FWsW1H+6Uf
zOb34bPWPvcDL1SQElETsIC7eGtsaz5YqmJM0kEPNP4En6wAPddDxxGVj42jscyt/sxVK2Rs298B
FdYQzxVtPDAkj/rFekwy8q+Ece9W7Aq4CVDre1PiRMjwKZgmYizAntfBaFcwiuWcf6sBHqKE0ToF
MvJZ23jlO+crJ83SxxCYNwbXbH30rvadBHPIufkfnBCn42b2dWo1UDUr/P6tAZ0WUuWA4wW0Yc25
6xderCVfmOVNvfDIdhfw+9U4gSDNEJ97ky3ymHD1e/wb5+vlM2HeUyl9t1AvvMGlgdIZ9qzo2wMJ
m4xJaTbDWT82zTqFDzgnIPHN9tbSSqDhtwchSCU6EovPgqyDzWwqzBIlyzJnmHc6+9SyBl5KHjy8
dEINmgHdmSzuiN4mGknwIg5dzY70Lb84WsCfQQnlG/YaZ+8q2104FWgdWVIrxEJ//jsa5EzmCGWp
ykgfPdPc2Nj7NLPR9nkwN05A3J3PHKK3+DtJtXexrq0UaptJxeSmgaap1588EA0E9geo1M1MyV9g
LK1OX6bzM9Z48oGRqJbJLNhiSZPTA+9WGZnrLPpwChxqmgasDmNfMqryZd+oQNSVY+cIRBV7zWHt
jrMSwU0yVj2ToPyqqsTvctq0yc4qPd4DSzi5ZBi20PQ3vEbYtTqlVSn8iterk9aGEs7ivZIa9+tD
fWvGYCzmF5fMp5DC5GNAyTlgGSQ/8UOS/8gQTpykjfnekGBuRZJJoyh9Dpvu7xspe/VmtxocmV0Q
1onaHnOqSGnuHP+nNTm9g/VmC4XX3L08hZG5fiaHVIkppNdQPZ/g6Jmfh4iiJAUpcaSmrvvsDex5
MeqXcXqWTj5rw1DJzM0pZvxOh/GxwmKQAC2J94pfHNpbI7nAv6wf2+DA0Qzx5MQohQ9VweuevZYp
wb9apzQtZTbAvdQXuT9nWDhea5jsHEUp9nNqxWLQmG5k7tK9UXZmXIGUpP3Nn6HDexghE5cCT9KN
xZfMS3sPLpqc+K4+QrEDYUsng/1ib5C6CNvnjyPlr1nTjcP3N8Ddc8Jd88savrr1YPOC0UhjjqV+
KrONalG4B18KZZJtFgbBch6WUgCGdpVctWLfHATT14fWiLF1VQhBQeHi/veZgOIskiQO8ldAj7a4
/FNju8GK6TFyI2Qel7c/omNFA+cSPcCdyl76u0Xl5843XOLojIwMhrZCpj/Vx68Nq7jsCDyGKSZh
I7sQ4YXdxGYKewpm37WLQML/uTOxlYe1Q8dz4aNO+9VVjetIyKeSbZJAQowivwcIYhy0CJwaeRCk
sb9SiHCJU3YH/2Ac74QvlHJVgiT9zSwmrQVDuuRM8G8wPOOtb39SXbIP+QBx+LUOOl0i4cf+u1Op
hf6EEThuGov56rziOiDnw+YHMv2aEIdEdyBit5BlB+/i6cMHrUkFPKIYdXgpF/1MopFtFgzTCd48
2JR01ctPmprZVh/8/7dSF5Nj83pGTegzuU8iIhdM8pdSZCPRcA28/0P28h2zB2IWbVI1kFSbxTaw
d+0Kz3fFWvR/Edy4J58ehGvNxU9ab3nYFRJLxo32EUDEwoDkDP9fzsbj9ZufdpOljF5lVudHqhaq
2ncQ1kXLtuC+/g80fkm9ejVa0kXjiT8L/J0s9CbprzoasTZd+vuGGqFWnnY1oHlE7EQcAhtSCvsj
r6V5krroeEiSiB8O/gzLdKmEDrCCDO076+Dm76IJerYfqnR4zn58myTOkfgdYWb6YI3zDrpf5J0j
W6MSDK10AG8WYcPPjUp1dQcjka4qkJJPct8iAj4tsWerL2U2cXkN0MCa8iYi6lyBp1dQPnNY6GDw
BtQ1hAvRQsXpBDOqL8s14505MJ4MTWHShrHx9MCouvQpzCICQP9jYm1CqbIPInFN19yb+suN8J73
fLNeaZ7MR2piZ++F/hA+TrMZc528/w4MSSRIHzNaRGdsp/I9J5A/+oMiMaCeL23OTp2P81JSmno1
P9O37oanyqGG+bgZIfmPtetKKkdHXXBMKxpZjDQoeJb9Nauf01fRDKVMjWImwAZTJuu3Qe4ZPR91
TJPRFwkQ1XtUAT2I3Cmgc/P+hWHRYM7PuytMnyfD7JV0n92crIa+zYoa7YPxblC8lgFXXo8U873U
dbOCI2vjHd+4qq7dqMF9/lINz4Dym09d06DKNCHqa40etyyaOSFRcdeVH77jC6hQNQYQqjvzbPGX
bk52cITteV1vOquiFsILxyYMyqEBhKko185S+G8psHnPx5utkd34Zns9Y0QGowfuNlA1Z0ZRUI3F
/1505CDtpny2pDUuHmTcMz0u6ZNk0S/JleWkM2jjrO6S3KaRAIPzNhiCJWOpRkA4BvU5TeJAKUf1
kpOC56l+kO7fL7wz8J4PqdRwIS+90d0FmdYEQAY1++lnqR5u98x3cRJF1tvfTzeNGk1d7JNZB6lR
gQOrMkt9fykWa53dV1S7Q+ox9os83iVR4llMH0INyFKCrE0v8guQ0V6kfNf4cumE191t18VJsRo2
FqE1usqFAkbwPxlpU0jw428gEgRhNWkKf+MNeX142pWX03UI0RbzlLaAlkB6iafgxUueAECMroRJ
1I4Nft6/5Xam3eem844tAxoY8hWl0r3SmPUNJ1XK8dZ+28fnfTBSkOAUixxGX5huaSfWtLAPkDWO
hu5PdSEqju3dXw6lZqe21gPaYrx2ICYZIuL08XNwZxRlptsKhL+0WIWsDhz3Vj1En6fj1TnrkHhT
N0aYfS0OYJ5xJt/DtQROuDecDaGwv0NmwPWn+Y5OLFiAHT95K4ryqJbjN3iXlDhPpgbLU8BBH2XB
xf/j3tyMoe1dfrQZv0NB1nAti5QvdsP3606g6O0xbD8PwU/xY0XbbrC7bDUvY9bvZbER+UoMAZ7H
6K181XyDQwZU/guwxoZV617jDuZPC5cw6a/vgwSwxRSabbvn1dFxGbnm5ckHoR2YjFwLRb9ex8hz
b/2OQbiiI2KteLiGGT7zdSZwu7TLkWnrWQwqWJV9MVdjck79rkEXcHsQfWGD5qI36MT7Zqun/YQv
TivAk3u+ZHXrgDNZDcvlbe5imjAzwivOrUT8qZr/h9mB6eyq8fUkDp/R22Rl0DtVkyzO3r5efSJQ
YdZTJhqCwV0mpqD9TbhsW6ZTGrKcww++jklRbJjXdZf3P3tvjSxIAeDsTsYx9cY8r4TF+HXQKBfj
8qzllvAlUuy+P4awBKuwMAgoApHkYi6ZeAbVFJeOuH2J2Dxe3GiWpkUIfk5FVudsCUXoIfwjd8t/
iS4YoZE3lB/ZZcv+iiWkf4U121ih/7E8XaLX4BPc5Cv3YnJ3p3CueozCMIYpuWAohZx2dCg9F916
NTQrtQzBDZUeKb3BYgw3oCFH2GiAO35Dw62jpafHFLxTHVeyEGvjLYOyEOSGx/kCk+ct0nBB16Z+
aBaNGyXsBhkhXg61pQkD+JKUC+Y5KWnt2Ft5WhUNPGX6GrkMAv+ezcflM8wxy4j21PVqnya07wUp
pWM0IBx9R5ocb+Nsv9KOOOc3wLDpm8gmuf0tP2d6M8A+wXNtscR7+ZBMYFqDQANwUET2ehUt3mGk
i7ZQKAqJihjlK2+4LHuOXfbK4JKIxX6WdRbbFPaaStLRlXnbMbV+oIG9byVRrnghLTJCFJhSksgo
KGIpgAla9zcbL8fnSXYYaLjEIK/vCyP9JHGZUtyXbvIAN0XaXQqV8Jzu5pEwHfOdyazx96p6kIWa
oTig4lHM9XI/I8BDsDPjS0cyoxVkC0ZA7yco8lZL7eEY6xH4ioiq2I6xvmwE3J+F+8MmhOVRwABw
glOUMVkNmTJNr0qUYKaA647xiIp1IFQtYpJaCZQw4o1IE6+pZ715ffgiS1vNr3MdhQR9dQLZD+EE
jNWqT2VIynEbvEV2O2/0sa5luO1Q48mfGmU51bTxF7vrd+IIpOVXYRomoOhQoQsdyTPYHmBWZWx2
2Res1m25KQibSvxLGolVxd3D1DE/0g7cGy3z+2d/hv+1KGPAEYoYlkYkE+b0+FaRtRCoOy/y/jGg
l8Ehc9BoJF8bizKuswZbM3Rhf8RB3jSbMDyPgaWuvDZ77SQ/exvZrUzxuPSZGqbtqvqljOYHN6f1
hvx+sB8ScXvcjk6FLXIhIJ7Tsqs0bUPacVAMaAokvW9gEjZp9Ek6WS0FIlgfzC0UPMKJDDx+0oJW
ubNoC9ZP+62CT5DPIXX1bLfUJTopMS+WNaiKLPJAyoBCa9+cafdsEw/0oo7052IvCqaKuxTAWdRs
9lcOj42YjMJKMER/z8E8lGD2tTdFE7O5xg6DMRUp0OGbTUgz+G4a38YQFsymQISXFZvI+pbeQYCB
ehBomeCLKYikA9zeIslpRs/RflpvzoShij8ogQoyD+eLveikRxuYuuafn2xllMlkyzE2k9j1/auk
CmuncZe1Pu1PoCygXcLZrwms8vPqoT6fFkOALPxLdMWpcB6h5iaQLWBTgrLiS1yZWghHhWTBorG8
WXXC9pPjiek3JCCDND3oCt3o9EVY6Y2G0NhJnf771qPrfeCqMtE1bKpDLddItun5X5peonaV0bMe
Uw35JA4ZLp3xJhAjYkqYZGtdWERxJ5oymZ5xq0PZ26Tmvgfv0v6UA2vmoBYG5fmNB/4E5JXVPCHj
ABYgcJj/ry6JATNnuwfzNxv11eAu1cYlatnQiCfySq/6+F842gGxqt4irQ3D1HPlETinW6GSnkv7
pBp5jFUBL4ydUIDPdKrQyC29MQkjkkQ6go2hPPqaypx1MBEKdKdhNhe75NiSxvcMT6AtoXCsL6GJ
XuXcalCxKgSLnwN6PucMxV+ynow3nsZlKYfvMobIpKx98EDKE40iLyaXxxcTbkG8MY4CNi+T47Ua
5oGSDbr8PjYiCkEl4hGy6WOAT+sz4ESd8AL9sp3eFNAC6IuyqMJTnKj6tAZBmAnWxgQANW+myHUI
bnkgECia1Ohy0U+XoysCh2Md7AP8qioUVI5XL7/uxlei0F0o6UGIHixvEG3LUbnkH+vBwHoxr8o6
qZ1fG9mHFLG9Ipv8oPE07TAIpGgZm2AvGTNb/Vgepe5qQt/it//BcZXSjkGO3x9pYHRPQWu2Wn42
Q9ECwWbMDhvjAZYJd84RY40h03IJ6yWx7fqYFUIosoo7h8rYKPzn/cvImY5WAwdyiSatihnjhuvs
znhU1PMuRKFI6EzcdBqCJxNCu/cDgoVAFW/512jGCCMZhLQp8sFP+xdxC9BcvNVqCyfxmRWsZrXF
XjO9SyrS1Pnnf1SjGUO2IPBHEvZUJ3G9iAwv/nueztUfoFe1C5sgrEZtKs+L2aIhKqsHF2hrgyEC
HrXPiNkj4V+ctshJ7/0jGTv6mztIMU6l4xt4Db2fSpvfBW2EfZtp+ZyhiPXU07dhMqnUA2NGpMT0
T9+EoPQ7sxKkjcS+KDB4ERcfTcSHR8uskXCxaahl75Ox49cWv906sVs7fz/OjMlxN5ohAOkrFAsc
FMgYndmPZFptnik617kS6InrbKEduqQLhic1nUNEGpCKBFDaYUB78w34jXQ3Ue7Z2+r0aAbQr6qZ
OiBLxydtnk4aBNzi1p2gAhJFNwKYz2L4vSGFlpFuUfzlOGAnq/MAPKHc3/1UU+NUh5Z7Je7px/jZ
/aefMC1JyxlubGxiot/yH1T+3BcfFcwNxgHlM5p8qmMKTMe7mmdG9pk7HLv6yY5zrPXSigSJwi88
pw/+ZvsWqA5fAEtIfAwQ3wyRw22bCmxMGGcEKPjpNMpG0P+sX6HYhrohzwPhF1Ol2FKoS9NE6iDs
eBJxWUS0Ay4AAoAGzO/IaIPTKr+9J6bn8XtidhbLxAzet7nsxmAqwkPtTpg61AuFFKPYzhI1+iPN
S3fABFTG4iOmTIReVgNOOuaCCy5eRCpF5uf1u0f7yC47QRhS2p13+ogYklXu7M9ppKuYNMPa4KOE
HhgumBbPSGwHh/PbqHXmPSO6/c0qFQbkKWV6EZx+SvS0nIvlmxiLij8NF2NTOALBT+3lDxVESsYL
Icz2SuwVjT/sMzXXm2He4AGTcg54XykGPaKEBjiDx+J3jo1m6iQ7xhMf3DvRjV52EbPnbGatti9g
qG2UPfQBn+KIn0CkMrZhYTA8xPx3fpK+Bmcm6IO4tHiPWvwL71MErDIEsbClSBToyWKCp9rP3haR
IWS1HWj8IjdTdCbSViFl4+Yn1Ktm4r8THg4ayK+ebcX2NiaUoYHOySUWwDb4IXSLFYbSTfMvk1e1
rm1z1Gc3tNzrRpmwtuCmw6K+l8Kq3uP24HXgjHEURHl3iiELhpgNKpPyRWYGl3Mx1ggoaAcgLaDN
sseRlyhnFVbljhaWXK3FGNVI4F/i1HqadZu4AXYy86PWedqwIPITu+h8aEAAvQcDe00vgrs6L5BM
IxoTqrRwCMkJlLFCbe/U/Y9lFMyOgXyNm3erigV1BQymxE0zxNszwmgs0heNVgQOK5UCl30Z6jxH
7XGJrMtyl2yD2IgEVK2Ja62yk+67J859ruv8RgK3CBjw77cGxdhyqlw+fQQapaL7Abm22lzCCiEn
A1h3CGsg/yHBl/8CPBJp8kOdKgOuM3n0jt0ZWcw5UuRIuObl/3PT/5z72G0mHCbeipqCXAZUdhee
xNdNIgss0XdNdTF5W+1YKtdjaxVnNvGohBboGPyaiwUi3bYM8i9/bs4CtzogeZ8jo91zduLGUocM
nBJ4f/V8hU9eDzCBGjDQaoDXbsai4VVbNDLc4iJ/JSCnyzJK+3r7k5g/P7KPiTyeAFzO7mvBTB9w
Q/ev5S9uUrrRN0LUL3W/Q3YWA+rITa9/Ho0DERtvpOF2IOBjNW4jSa649ChP5C7D12NgkcvQy5x9
FOGF69y6iZcGSV+9F2lixEQW38sVN2lvv2eO4+odWU2GS2fn8BAZ4k0puPEWAp9n7/vyS+qLPqov
V2ZEzsBU4i9kqpdNpNh4PKsdz4qiCLz26ugTv2Drwj94IOWVSW0PmjL/co6YL7iPewYM9rmpthFc
lpBlxDtO3ef0KEBqjvqJm0ZHRCdSwgj8y6jsSgmfYCkOeTYIuO81RQiKPNVd38SX8dOLlnbp7S4N
O+1kxAmllIa+/ru9EqHg3KgPOZemsnlFR1j28mfCDDeP1dTOcdUOhrQHD4EOjZOxnFwyqnO7Wm8u
6YkbyhwQ7+F0r/jo27Bb1gr1fiE9TIMEd5DMrLfKDUETHCHrMe0sjA745H0suztPlRTYNvzqfp+M
rtoz4NDJVtY7rHmyaDNXJBUWmvpecp2rDaKXuN6G05K4lEnaAN/rG6IKNDuoTuUToV/Fn1frXWs9
hXMfU5ZuQf2pc3CxDiJhN3BZq5Kv7ocHrTh7lSQCutZTlVMcejZJTDVPkx7rW/X2xUDEuD5JQwTG
i+eb0kT+H3eCMCspgTitHjW+5GJvG/GCnGb8GPQ5KQOukpI/aDiYj3EjFL21ncRziqWwlYEIfV9t
k7USKzhECdeouZx4LlhOp7BAM9J/k7o3i5DqyB/q7lrubvIRWLFTst3DDzefKS0BGMNMM5mr5kVa
FctZx/K4bfzApTmFsX528Z/x1PKYsXTdeq1JEGZslEcKRzjzqWGnn8HHTZzjxf7/vm9IEuAoHaia
dIxKlaLcjVJrz0X6Vr7o3ViZewxJL4G3lD0vIXaD9SOtEXRiphnnFYrkwFbihdb8wMNL6Ym4heH3
2d2eGTijTAl5V7UEcKHt7t4reFBmklP1FmJ49l0s3Ybrn2BIq/yfFb6dRFv1Yf4yaw3p0pwSZZc6
iwtH+VliVyctVe/9k+pgulrXfjwR/ip74VLV/3tp8T6nhmUKXoYo3fZrYBn84SpUKb9bt8Sr+oBn
SztVtYhbDdy34myp+COwhvvGQLOLy0aziz1KlHMssRMvW8kKxXzdDbLph5VzJgDBa8MOjqaFZgCL
xkp86hiO8q/oTEtYMTj3BFai5/rGnfQoRlgjRyuP1xGqFBGI7UM0lPIT1sEAAbAoX1iWG0yKxAMJ
2BsTEXJ5XCohNr21mbroeAgXl4A44Gm8gRIMcfte3Tl7LycqQkKaYwQO12NV/IK8X+7H2LmEWYyU
yufdTiRiVtIuy04r+5Hk5OGi7ECMi2tKiFBNLP3h2Xk0X5rS9POvhwmZresSZ/Lp8G3oGgSWHoE9
NAbuuJLlqR+HKrJvHtIyRR/suImKEhhCCzj3ss2ULR6i1twOpMGcRIe05gCAHDO9gdt2R+ZvE0/L
onzRBZSTxsxUCshN7if5RJIinospMqg9TkmqaMYfWgBYkk2yPXKpf4NPOYr3tob9MIzAfCpULBh9
Y/IvdiVuHd5MjGW/AYlnPtG9wmPqEn0LV0I353fqU9MTX4uu39kxLuivBJRPGJiDPcOA0/UFzuOz
0cvPrT2BDsN7CBzD5xh8G8dp98UYZX/thLNTUOY4mgWau+0HCxPz78+bgZruyYkPm3duAnw//HzC
L27jDSsg0y9DThEUGT3ZaXT22Ge97FFd26rQsLBufl60YgZbuxYl51rf1lOjc5xmmHMEifGqcfI3
GU99N2dDkPdyTNa81q0cKLzfPr6nzQgRVMU3MLCZO5HmT25ocHaE1BGcZOE+Grn9HaXgkgQ1tq48
2cfAUipMz1Ghjq3/dORNn46q4MJWg+d6BWxcH+NPYmIP+rEVv0ty7443ldIYxnXcdeHsUbmYjeMa
H2WHKCR57rSBuBJk8ikf5VrQ35aZd+jBmmDu1+kOGs0idzdtR16rGyzWcbtJc+OMpw2iwdct6XLi
YzG7wzvjaTMKXcWcSRbvsOCNIIv+PxUJUVfbO9ZfuFiS3zvFeKIiYiMxM6kjBRSqpy77UzsPQwlx
TWdRRTSijLwJinGyk1yC14kHUvASVJGaB61HeXwZtx7MR0pm3Y7CVvVKgqcUqc9xZZSli6HKJDGi
1a0dIdEGF8u2ndG8bOBU7TpmOk42hgMwpfW7ziHxId5LIanOmIaUzopaXVXAIYqNA9+mQqV1hpPk
TrWJssGdrp47SJjzPtUSegyxKhHGg2iI+3CoVWoVcISw4IYXyG0Sw3eUapiMsu7l/aye0LlXshJG
/AVIR08ur7GD14/zX5xgRUzR+8IA5xTRmD9IUB35OW+oy17jQfI0+cDtwCMzoJgabqbAFJxV/QWR
fhJF9KllLrSoPxVuGWj3AYX9pG5l0X6gJ+lnw+qFKWk6cvHhQm20PLIGDrenPjHPXnZBvp0T0YlU
2eNaFxFfXF5pqpM2auFbEGO9QYxZmfiGmn+i61xHD41fiS9dOc2Fx3F0Yy5QT1NJqLoEwj2VlNN5
tWb/uethvrkoeHx0UTuQVjL4r7vJWT2+hJ87+i/emYgE3XIpb25mKysfs0mtNnV1bOLF3tDDEEFP
dn8tmxVFxjZVAQHdUbC/CYwvddbLwHppGAQYjzOpK0W972Kgqe+BH+VT04JrU7pioEDi8TK3HPoi
wiSLK0WcMBBQWocdWHJDTNKCxZ3gIZ/D+zgDkUAHks1poC3rQdIc/oyRWa+RbCiqDk3quk60URgX
TVj18XgiAVq0qnJWnT1zOVPH9CWF8X6Z9LQ5anFyQz93w6Y0zaO1fTjamPwkMhSm83DxQRYeYAv5
JDkJsy4Ig1Ua+bm3MQGROfbrIqgQoe5WLPgM805BpODtjAZqs0qN7GZrSAuayV9ucA/qFfEWeDxH
lTJW2ORpQXdZnTI/76Vhi8KyWa5HWLMMAqHt9OFyOzdc4QoHDDTSJJ4289qkMRirvWg3grISmMnw
cpMWBVbVse5rDN+cm3Z/AELYt8ccz15GP9IgairGAZ2AhB9q6IXTOrQ1iGIcWNOtaZYd0i//pV5D
XxYyANNOBNdS5yYDzQJ3BZkqvrcqhbf0WnKicnNL5TXK9yw5d3jUNPX0pP4d2SdMJCEVSB/B2VY1
Yp/2SSN6PCWtJGoQPIlzxHhqof+i0s0RkZkHc7xp3rUiM+OxJkGjVjKRFpcLlMQJFdbnwZx/X44r
KCC8fVFNnveOSR0JyFLrd7LhK9+lUsTzpd/qdYHgFDPtItETiE4rhxKu8YY52tcvSg6XtTIPiyvV
URJYADgOnDVHGO/OOcK9PwIwvPnw5bYmAVyGzi2hgjmN8gCRKXmC8M7/5gXMS+tvMRRerahHv0zf
+usB1nmXDXn/tKAdLmLAqD+8m5fHXjG5CJ7NP8cghiFS5euwQVowfscQW4RqdX2gzk7xn9HNMhdI
Ll5zwOslo3pdVFWjeCvxJEGmbK6tOoas1FScpyIrRxsr5EbysKymYJa6CL6Lu/BAE6ZQ6WMU0QDz
1Qyc0/XUuP5S7GUtHYZdAlUiJt97XfLB235spB6N8gXnw+7mWCFoakaNb3qSbLNEgPVW+e1Jdynk
FOfUmdoRB4N2HdADdFJrB69zsVXXZTwOkx6THIoX3J3td/nXVkBBIjZct2CaxsytTOYR/nF6zsrr
2YoEr8Dv7TCREvG1Mx5uYCnfa4UZyfq2tUlyvhYT1eg8vvB9wSMkwguyrLrpy/GT8FevI//G4N3m
SWoS4s89THxB2woYDlEbPepjdkT+u1EPyGE1NCnntKb+k59lcmd9JuC9S9IyNqGu6hnvaJJghxys
ozs6tLXPPFvW5SY32GzZhx8Xl6e6JWgfP6/NYZn0Qh5PMtcsdxW3qibMHU5fh8PgRYXnFgDegxxI
pA/5iT6MaXu5Q+R/4ZWuhb8TqZ48aXoBedGeOhEzE/CgGgpTFxZZANpmVTAQQ+LOqd7pyjqhnXCX
g5UIfxvYcY+NQJrfaXRgEq7jMFcQNgQQmBL+Kj13+hlnqWw//MYrilaiI2X2JqIZmThpOH0lYirq
ITWDsOSMUelUT3p8nHyyVq/8lAjC9NJar1jnjF/pWbyIv2nf5gIpxneiMBBS+IJmU6EFxJ+unCK7
NFk8PpjC5h0g5rj9GwhhHGJD7sC7jTbmTA+cZUC9jdU1jIBfuVSzIglLOHgOWMOvXbUJv0oE7A8m
yBCUKFzTq6/Pr+7MM4+/yPH8vvdSayLkBWK3ap3M6RXMyNnYqfyK84atVGvT0bWfqRkwyTIasvqT
7V0aaS4KxqLQtMsRoiSJwpV7PFPtw/BszGv/n9AdL0dhUlr6CDXJj2uAJA0/M1utbrYsrdYwPcsM
n1brDgSAq35KGAETYP0/DAZ+RUXh3zEm8AYDGsdYCnaBq80ejM/ijhkYsEFiHrr5dHw6A2iCh6lN
die7/a1jgptEs8H/dVR14TGHYBzIRJFJykR9j79HiFWp7f2Egg57q+yqvWRsjnfxnmJdWISyqqZV
Koi/AgmidnhzEhkE+EPRh4mJYZSBhT4WDzfxYIroFIxGvWe9/7L3ylaHmQW3IW13pvToyRBI/Z55
Bpjp9cuKnZ2/NEhmaDNUWsjLO9bZ6GbaxyeoZCER8NTiTrSu65USN9prV+3n24VTQyMTSmYknS3k
MaBiZvc+5GiIdhC7tFVGxcqum/yO4EtN5dlfC9XGY3alTOuGwqiAXhP0bJoTW7dvQWKaq1T1n+pJ
juu0glzCUuasMAAPsf3wbior0St9z1D2Sv8VUsDvmwzJ0oMMC/DpN2lRyJy76OaXI+3jCrjNbFjk
4V6Xlh+mdUI25X42U4Cr98xhVxvSMV9VOKhu8Tayy0ps507+HkPMuu4PbE7A1+c/tVPsZUtzIouu
OYohF+lE7S3bGyeS/3IonbXEx+xsbZGohHYd/eyTmzwdVRujx05wy9LAHb2fcfUIhBvkHoD80/dr
+pLYP9T3hqriIrFXBDF9D4IEeCyP7vH6zLToj+H1hUtnuvW4DUJGCC04UFJ2sh5c7WzTAQuyKPY+
Tqon7AsBmjNKij/QHJNtLnYA/4Wsd2kR7HpE7y+TjAkv/P/x+snjZsLhGvpoIXrV4S+iCdfRP8S+
ucCJROQZD512Ogm1aTQ7RJFM4VV0j2ios+nykotItBE/9r+fLHv7z9g0Y6Frke6lR5GLwrWV+ZII
OwMUVBFYuLzJSu8+YE6TBDPI2/d6EAptSKjnSjHco42/Nv+k+0qP7bXm90hUdiasChyWFEVKuEHr
KyuujQ8p80Qy6uDuXeMgxgEiwYPAY5QXAnClaM0siUuEaL0Xuj+AFi+7BZCNOPCdEq3elQdLUYgX
tO0YNNyDpcv8obsiLpzuPIluly4PLLj+UIH3+WyuTGzGbrFaLc/b43mCQZX6gDnxWoci+PgvcJB1
/p58YC3ddMhHmZX/OqI0yiDHJtwewo/pEhwOL5MaaLtklRxQb0mshBz+39ePdU4eplX/TEXmtPaI
z/RYxXCbXqsrFRJdAlNkNK7url+ojzHJVdFbHndTyhbhw41UX7cfuWxNsMYZfVvyo8JwrqCoM42k
fR+oZJRrGV/6BJJi/15p34GfQc74G8vazgG8hbuF055iau9hE6JN+BGdBj4JoholVhq/XCESmyaI
w4toiTbY5HQgt12UWDKIVuMzNSqUz3PKwHuI6wbceoWDyIUmqn/B50dSUIlFM/F2djd0LRL1nESu
mhp2SAE01sZqov4CEFu5gvYeuoStlr7TSTpPmSZsUdHRHG8tWGPPQTXMP1A5HnikKBzbtZaUxuV5
6Dhw1ZCoaFCEWFdhvUu7435Mw9K7G69aTsfUBvFrRD8vsX63HFBf+TxWsyfbq8m5tZOpwaZmWk2a
xn2PMEBwkmLS1WBehW5tYgqSpcryKJejhhW1AJJrG2ezsM7lgPLfADWyS5HYUb5WdDjwgeaacFdW
FbVuBX4SWOe7ZkawiGcZl+zqQUwd4I73gb7W3aEeQ9oBMmtH9EaxRm2UbjhH7kgfRUslHU5Q/Cxk
TkjWOzHC6JxncpUSJFzHUk3uhoWWCwnM2qE+6squaiJmRHk3PREt5WL+E/GKG9P3+iUxu5v+lpSR
5EABN8nkDCQC8gQXaNHsq0Cie543jKbQ91U2qNekv7egYQesFYdYi2kPJcLisAiYiDVEKL2rKcz7
7jxIpAixjt2Barr1Wjc66b5hOGSzeMB+NFfl9xPLno0LJE4hFFfKPYgjQyrPPNpBSoL53tcIMdOO
XDz5WVd+MXwAbvhZNkuAL7vnsJ1EUw2JFR4moWD+3rJWOltgQW+NkdbhPpAAFSp2ObdCRoOWu1/D
Jnt1K1B3tYx4qFRpYAq3XKCaG6Hvzb4gnyFLLTPKw8zMf5RROkTYpsCVSgLKTq1JbR1ErRg2noPw
dK7d96z+FkQO5pbaCqgXmyfdHMoz3lAM0hWfNj6+GXYn6NAHxeqr9zTXk8UFWfY16brJo86fEg6y
bRdOiDVL1Sq3Ka11+dBHgoyf1FRUP9LmPevA2Fscnc12PCyfA6K8P1EhGcSudQrXXo54KNeBFboe
9UZZTfqKmOOb5jHEDIy/1t6bR4G9vTwVfs6OrkburznxNZGFKwItt8rw66gYBsYlnRWVjkUAGC36
b9pvNrxDbhqWRplqXrDY7CBlci03DvZj0D87yd4P0yqTSiW9pXZi9v1SMnwSV6NAVAnv+ttUMy2d
zzhAJ2dwg97OQ1hk+Ei/JKIULEsHM9JZzK+OwMPSc8SZqz+rLsETy7ImIKtlJ8odyqSJMbyGQ760
QoUQfO4EL0rZZkpebf7+SfkCP6/3bfsC+q9Y6rytqA8UuWz13rjkW0YMzDphNCAvC7SoMKca4Odr
yEPGMG1xmaSuztH4AuFNvvmaIVEB3DwJJ2OpEiUAL08uwRlx12oqDDhLzkaFaq+aITVjeejFlUH1
FzFxSnVEZVAGdUsunDR+tzpIXwPWHvj0Cw64mFXlco/BSNty61VtqhutEIuRhRJonp+dcg4tVvRk
Rp/f7VUtdP2ROJiR3JcqfM7Wvc79t+uPNAWwpO0dK5sbHkfCfdHE0rM4aP6isHJGTMju4C9S0Trg
IQvxaQOitP91488NnGICh6eLNvlyDho392iCOznvXlJYmBq6HzhlUWfxNUVNApzuADBZ8pRCwEjz
KKFyQTpUxsWgOoc9J+gMy+VMumAR9Dnoq2V06mzPmiwcrqA6cDd/MGLH/FkfJtheqXIK9a6LZUxp
u2zDTdX4+Epi6/Qc+11nR6mgS6CoyfCy1P+x6JDqC5/WibfB5IvWI4Ov9Qg9xhWBLuAsQ/Xte4qw
R1IqlVejXFjRq/zebscnm6I47ec2BaxnQd3Ved0Rj0jZDASEC3g8gzATKNQOWMQVWnh56dDaIzXR
2ebPHnKMY8F7ZwLzmT9I57viauTeE5FNNXJO5yNyDwChd2jtWVbnzUu5YGCx9r1VgDw5hejc+wGv
yeQWs6Wh9TX6UdI/nAPXJj9hdLb8W49LFgWSy4kQaN+/FGzYzm9fqAnydmK7UW4gsBAoFQdNiwvr
nGqTGrIl4LnhadtFxEV1s8S4JmUTy3nIPCKWbuZfSHds1Th2C5XhuGdWvRUpuKVwtT79+njcVeHt
XkHslxJrbTdQ5T/N2eXOTUZVArblSAMH2UOJZ2nXiWRAPrZvcD3ykZw+6VAjOfw2q7FeTMx6Ng4D
ovqltmBnWkoEnBcp1U7Nci9yQ2Aftn7Mdkux2Sf5KxubrumXfK8TLPU42scqn3Zgo+0PRMDft0pf
Vj+FDREoUqsHuLy+Lnm9Mco1Tg1BScWYH7w4pgzwCnev97mfEv2cdAvBfd+rHSFcLqYfR3IM1qjv
LctmeNTVSMddGo5GF/medRHrf/KpVYw0UeBMA4yVvDbv9FSzSaV8ygYxcSjBoStStJWuPn+XbuDE
RitbfHqR8K1ojfMl1AmHP4Xg25FUgKIpIt3pMxfCG9bHm/FCCaS8k13Am23aKk36vNXQ5eBiDcjs
PnrrzexIkUDaJZBaPxynUPitTStqGj6WqbHQwf+xWv1IbKPCnsnvWWe4H+yrtnx7SY4xlVrDVbQk
kth1SGoz/P86eSv1XICuD4XURcVDb7x86rCDNgVDiWKeIczrfHdL4fYjScYrNpY9WTFktfkEQf8/
ndj8UFZ5l0Craj+hpk9hW8dncfV0Ul17hcwbJnyGR6G5bZ13+wekR5e+aMl7btrAkIc2NrdPFRP2
jpCtqHOVKL8rKGzEIMmBCUxcYsU/vHSTYzYG5S17C1FSQ/8SHdZ1920eowZ93XMKeg3NpdOHE8AX
tnXO7hWuCBgJuvASodlmJdBWg7ZCn+h+Hsepe0tmibowj3X/2idar5NxZPLOqRCqLvvVMn4iCI0U
FqGOsiGqQKVu3IF5rhDhhmIqybxUVm9La0nDjdTSTnCWta5RxOVmY6bSILT+FHXTIj+YVnApqe73
zoLo5OiQ60DF1Cw6xZNLBDmZ0AZkh8i2LI3CMc7/C/wNUIQnTrL0j528669rT9kJxaTnZORwexS7
5HQoH6h/ssMxcKqpGmgIumYfDrYSptUpspa+Sfs9m8U0MnRVwTuSm4d2VCite8A0wAT756S11n3a
wqb9UIq67bnFj0XEXqiCHatup04UWnxJ5NYc9epf4rlEB93cjk9GZZXlepMvRvVH3pTbJhAwOItR
Xn/OEPEsHTuT/OZMLZUaTY5tAZxg2NgpyPFFnkC0Z3fCAv4Vml89C27KBCke+Siq1Lw66QbLxA0U
5sG7sQhJSONVOlXWPstc1qq9iZjC3qiTxzBG3603g3BT9QQGeRAvy/9Rp0V7rc7zuy7rXVSWWdFJ
JAaLol/5V5U1tMNPBUVKpiz3LTeCXJme5+yp6rO3V6klJ8EfkkfSmcM/isok8AXXE1rJ3Zwn/rgR
Krwuql4MGJ0FMfMCIRfCCSv7NDtyrQf2ps0qXifa5ddCcORlRtoFC/vVPFu+GvsVOUI4Qge1/DsZ
P0jqxW28arXLE99L+13ryWRRKlSYi4q/RVZGwO6hHsyzk++yRw46SvQHVOybAxdzRm7KDlbqLBpY
UYDnsvE923PbLZRKntU3XdF+ig+pDibLOmCFiUjglcHUncX12+GUXjxcS1/ExDP/LKbUYEsCrTMy
GzO8tFUbEBsr0NQ3S7B2sQgejMDTCFYxGiapDaIgyD0WYln7gx0+CVrSe08f6u7R0+4Nz9J27OeC
rIYvdjZciJYtf2pzU3vuKO+tbDJs/Lk0ypdw7GR3T0l7oreSrunpk51j5tS8v04AlbPAL1VvLI0j
2eoYejH9LjLj9gYDERcJg2yBBlV4u6s93zrs35SmjkdozFr4KcBBNhuE/js2Tjxnpzsppshf3MqF
ptYBzOcKayTsoCyZl2qcP2OHW4IgonYhKuWf5ykxxV0QoNj+fNwyrKGGOSdm1U4zWTtzzXyUmoTL
YGoGHe4NUYGQoGJqqppZkw0WMIBWOqSUV/5Cr7CHQ+zVS18F6fhxopDdAV9t6jQi9iMIL/jpq4ci
1o6V0nuSSmSnqvfKMeO+f8q/voZa4yeZbb+VGQtn9eEAqvtqPOY7xsol5D231pjdzgDdwNvB4P/i
kiKvZpGw6+Z23rsu9OujO2eRNyj9uCaNfBYBXDhbl2WnaK5T4EggeLROT3j2Ytn1gMfciMShizUO
iD55oQHm867qyGfCO/WcZER40qxZG8GFd5bGz18DMfWpTarUv7xUZgKK3toeEv+Yyn+tgSUhS88z
AXU0L32CGJvsayEqrPU/6R+M477zT5MhFKWQ8z0WtjUxqUkvNic1UIwBGOXLE0VZTHKkJGo2AkL1
tMW6HJQJffuy3rTuqrGJiR1MkjMheEE8hIxF76yLma+2egkIeiff091rfkzu+KQOvC9igIiEgk2w
4FsTpcLsSmZF0yP5wkrGhu9QL8GZ2gGUEGwsusqrPzjJvtJx3/B5h79/s2XeiaC2ZkysUmBXNXWH
kzi8Vk5YVNbcHLe8oNeMkwB/x1mFCa+MJuhR6wX+ZC51Utn/UsQIqUpFcV/fOeOX2pwPPlneaRBR
XSQyB4e37wBOZu+zzVtDcvvf0PiD8FTuecO4NaC2n0CYNkmF+SPQ6qxRgHXhgbFiT2zv7QNrY9vs
e13C5E41WeoMLFP7EurVlxrGcdH38OI6ZeomffOUdu5SmLyKRTJUAeR7nq9jl4kAohceZBYPYRg2
TyzjjAJ+poeZZUXBaytSaVt/jrHVkdgrhJdz2KlOA1N85sfZf4l1vKTnr8i24clpPX/HA2PhbeNe
KGtvvZdxiwX+cNyVvXw8xPZ7c/yRwKzitlI/py2q7qg3WUC+EHrACW81tO8uN9G47eJ4zGKgKhyV
o4Uz1BBDQ+1oOiAuXhhzL1ujrVSY5FlA5k0afkvsIETLL+hQ37b4PF0/VT2gkVhX3fSg6v19ht87
Nt72KFGOxkzfZ0j5pg27No+HDJ0dxcOb8/Ocl6lFIh6iHlr+k3iFu0Qtw6dxBTpn/3QegbBc86tQ
Kg5zP1CXQsCxileKgfAbp6hOO3TlwROFPxa/WDTjcEnIukBB16pgKeH7iLfMAD6WEzAZNjkGlpRV
+WMgv84SHE+30NFxHwE1KERZ2vEmSJBY7thdxssGvV505uHQft1HdO0atjktm87AVwR+/OpuUd9k
VUOtd7+Lwp/OknsZhcVMKFcImxy+9egcK8uw7Ye1ZWOeM6iYfTU7GrIJvrRHJHoOkk4fu9RfFllN
2E3daqu5wkoNBq1qdfU6qeCece2/iCDA+4SbL9t5KPOQox8G/o+VldZFK3VxIi1qiy+LC4itW0zZ
q2HvmwRkCTkpMglj1z2QKO9Hss9Vcc0IWW7AOpeniGx1kXiLEq2xqyETouNw6ey88cH0FlHUdt43
TUNMzStnTSBdw9EFdz4gpLrETwRyn0Xu33fWrMUs246h2gV9yCt5UWu0Oidm82f62tigJp5PgQXn
2AsIkWIRi5oYjWyERt/qM4o76LZE0uYkS5ORycHlw0Kn7s8z5CQk9F2xlo3uQB6ret1rMuEOyIwp
6q3ctNK+1Oubq3zRdCBdh0TLtGmXkwUxMVaD12/iabZdNpMt7+yzU6h7bkCgvGyRfHx8lvuwEPEb
vJiclUCrSFqbaetej2lY1Q2wftT85lrwft3kQ0+CL37f0PefQx0Him5QvI1PAewAvnZ7VLEJ+No3
IwYUnuKs1SXIk+/tu5Gy6jOdQS6YHQ3uUKVj1Omk3cmjgWXpFic6OfIvw+UBkj2bITAHOWzRf/Es
D1gYu8sIFNO1zs6obDnj4S0r8RWUCsVOnrwY5w996jkyQyQHK6P9NGCQqm7ZlwYCeOy5wxO3c55h
6FqrM4AWWoJRl002491WDdY8AwxRKZmEht/uVkDSWRt76HKJ5eCakWTFDukgikXbz2u+jWDlE+Yi
PHufUkXfq7hx4yNd4bTdpgwmp0MaXPY5LRIddvFxir7Xfe8WkwDfj5LPIf3HqFKX7M/vLHYe+4qv
3ZHQYGv/eV8gSBw8joqTIg7pCejpgIVWB6l1OqRGn+8Kw8f55bmedXPL7wCUjSkVzE2v6LqhTFq+
OkUeqVx8rKM1Wl2njibnap3/Jc4B0LHV1Be0RoT/LT+JPI4kibCvZQFDsUYXe1QKQFvIjbJFcssu
jV1+OwylJ8qsGkHv6AGRu5aCF9BcCANtsFJPx+wB15If8kB9nH0CDlCvkTvQeZSLJCyl0QbcmHY+
3S9adMYUb1D04BQwaUSPRj80pABm9SA9F/Vwf6+VlPemdX/ZcTsMgpUAuR/EU5Y2zCTe3ftUC62V
c/zmsRHQvnDwwp5jZi2OJwhL6Ij+KgQk3M+XARWCSdEoX6YGCbypEju3e/kne+ekSGuWsiZLZjL7
j7WYpmfdIPnS7jhIs4DRH0GBm4CWGUrZgHyo42Gg3kqAPV6riyZx2z5rIEZxLWRm9iSPyjvd1+1m
oNYhRnAdvE6DueylEhLTfnI5d7I/ofy87q4OURcG18l1VE1xcEv9kVC0SrRgxpLZAD18WiT0tUEU
ZmVgNH1IuevfDzQfCQoDNlyg3MSACNDrdRP0T7cWE+c0pK3jz+YoHYNLqYa5TdmPO7EidAxtivAA
KsD2E9/ov6f2Y5kiUYeCg/KKkojBiS0+1eRKCs9eBcWW+xvcVyg6zZnXGFJPZhLF/aSdQg3Wz/S1
hUluSD8BAhiailspsCm3xaCaDLqhbmotePx/8m6Sp5PDjvLT0BNN/8K2l8Ki0UymweSY/ScoQhdu
4a7sVfkQp9w//n5xfZbR8ls/bPXTert5crZUi6OEDypT8uPw8Pe5ldfchZ3Zp77kYmoyZvXJ9USY
Hdoxd6KqNnWXEQhEqCKp9wY6uzUYgBkpwxLsJD0o3Kd4UB9wxB8wMNg4chNgHYbnqOPkFg5p6UOe
TUGIew69cY9ziaHOg9yIW1RKH60TnT9PrcIC4UBgdynFfPotEDG2MTIG2GKLH93QExv2wsUk6PK+
DfDvp8LNsmlPF/solBb2czn3RbM4H5uAYLO+6jhLGfwMv+8SItD7GSyNo13GpDJXFFF7nH1diF+P
rTt26nS4jhYHHR6+Emad/PUZ/9+Vk36hfaX2hxD027MyYmIxxBzoKAyi9pGJ8hV5v0kN9LszUBdc
3zPSP6qtDdoAmQ/4OvjFta8RAJX0BMtr2gr04bcoQJHbhVJllavrK/RDmYqckQs/J0t1EoIMv0fh
9FtaELZqXrLrriXIzz88LdkQ1Trm65ZT87b2GThwb3v0tgFpRF2yrcFHXQABJswzvvOm5rsIDD8W
yNh1teJgTKYnPpZJO5bhJAloHYoYOaEgxCiWfgDhz9hvQLQX+INt7Zlmld2KmY/BsP8Do/vTyQ0i
FI10ELJWx+tPZCd/sJ0N1M/E9jdSUziP9VtMsXRZP/St3s562pVb+iiSqPFBNXryWq9Deqjwy68X
PMOeUewJt8owzJyrMNJKpuArdEy8F1kIQj16hXgUETr2BGeXNA8/Tqa34PUWZZCN1CxX+ZErIVbX
2a20LJYq2Ma7BXjDMmgxi9bkPxl1nf5xNuDdURNTsBQc3st98/zyHB60D9ZMYO3Hv3YsbqQb6Sd0
Okw9NtapSwYQcMH0OKdBY8xoscovSozymOrow3SKHUydNJJMETrqLlXxqmj1+b0HCBpveHuPCvTy
1t0lO8WQzoUVuZqoLdf6Krkk9EUWHVSsCQlygk0yL2OqTJJ5Ws28gBJ2ON7ajbvprCYGWZg92B1G
c5kiA1+C4L5YbCiYg621XV05rggPqnjZziuBScCAevBg76IZQxzfjed4EnCCRfj8hTRmxNWRLgvx
s1G/IVFyJbxjZLoPuDCVCYAFM5p7tgRbMxXXh97Qu8Y/TnXV1qAnz+i3w10OTPI4f2lv0iCoK17Y
5AMyYPSy8uNzp1AYqnmGvL6n4tzZezLaydiveYoVCoq7EfnXSx45M7XcJ75g61/yxluR79nLn9WQ
OTHMZAdIwz7mAbusiMsGV5vfASVuRrGj9V4mkXr4yPyVxbZvt+kuLepBbchg8CgvLafw4pjrDG/z
L9qOAoBbr90x5ox15oRNlgQSbNIQAOXu4kgr9dKzDSpbZIQ3tm8zW2xpkUDUc+DWD8Xkg7aPq0Lw
dLTHYl6qJHD0jLfa16I2MPfjt5Qyo8rrISEU8x/iKd7ToLxty48qVv6utvnJoW08uz+2L3/V14yG
jsfmUuY5kugrAnBXS9YRs02jEqmZiUATlwz1tBc4nG8UQr0DYS7hVUlkhu540JlH1e65qFs3AezX
zCDlTgBqj2beR31gftOaodiQbjul5Uz5n1l2ee2Q0O3vn3EFe6pTSLhQP/voi7SlZJNnK+M6ioNY
0m+MyEszOBuIKdK86Jl8QR3FeXWzX8st6U6MR0f+yjXMaGNZE/F4Ar9FG4JKKKNPYRqipIsUf2YF
vHUIWdlaLDDdjuqXdevUfH71vrcJQb3enfDLuCtDRtt6P5eoqmEyPkqvCyjJbUt0gw8+b4EO3BBK
j/3ZrM9VKv+z9FZ5Zb7wT+7JeV6ZQafENGpPHduxU6trY6KKk9ATjSKefFxJmkZPw07s/ugdpD9i
rOEWPLRvtzuFdG1DD7fu9+H23lXQkheA8E9EIKZOGV1W/10HPeaUFT4pWkHQZI6KOuz+bMUIhwbT
49FVTmxxvzBjYskNqW2g5AGtuIVULV+KUjLNOQrNKWPgL2L30uB9QVvOsKUaFQh0MOcNfaWuf3NQ
xmVVmRSERkYiNmGisZLy+jsqI5GrjVk3YTiJbcFIQ/KcC8EVn/NUoNGAIHVv71YsB9mEE32SzgJg
j9yQ4CgGeVxzSQ8m3Naj8/HovfaJnKaZ6ktRhp9S4MiTCcgWVB5rea2Fg+iAq1Ze/l8sZin+MYfy
fJTHlGApFVho3SsGwZFA7pGVyapFVTL9/9rgIDptLgmGAgq7oqOJjf2XGH05VdDER9gF1fDYA9zh
KxckK/5bbZ85y+feytKGuoEGd5dF6GfCI/BzgW2+oxjFkd8KdC6CaOWXDviII2ANDn+XTosqtwpw
24hDI9PG2gux4DEdnzl9+2rX8ODc6cznl2jF3OEtT3XkyQoqnBa2/+njcCa+tg14WHEQ61dFT+HT
DfbPBbPA6EU78hfy63YkhSGJa9Ad0ZaMPW2ge8L9VoYVA13CyMpL/iLEkWV/oKHwizIt/yi+q/f1
fzSPvOU/P2TqpcFOGyvwkbng9zfsgn2MeKrwkHLaS4F90ARLAo9hGd9tMtK0HReSPXe9K1qmYmwz
5ZUwxWmj4XP82cTtQ/iSb8g3GWg0J6iDPaE6EgiwXpBybiA/KMAijT+nUa0mOcBY3AYgCJKZlzqr
jSGc89y8jSS66KoVOAJWZmICh8NPZEaIg2gdCY/EzDcKa6FdvbXih5Za5Dk384n/h7bTinDQoDkD
Hec0MLMBigHkjaUDrMZdkiu8IireE3J6L1VrcXC+7fbNjAGWzySPqOSfe5Q0q+hqVsiD4iChY9aA
TshdKNzg6GryMjqlD+6y7fJGvImtemcP6IJtZCO5ZK10tWBB0ee4hTA1XlfOHDEe9fkZPRttDhlw
YmxT6nuZtJdkjkidvPiGE+JdQVRw5JZhLkcQLSWN7Luw1YCotCyNbEdzYpFQR8vgNx3SX6ZYY3JI
UEQ/81IXukW5Qg5gCJITrP/3IMge4rPwJDU9axqjZQmKmrVD2tp8Vbb9HJy6wJXJWjrFHeSFEF52
/mM3HirpBQBzlfe9VTlE6PvioU7pta+WtYWlhe5+BYRGdaoLv1dpOg4DDiLHPFjawqwTcIBtzuom
SvbF9ndBkKj+6El22ztkki/C7cflrvX0qJLBA7UgTPUcGSXL4ep0u/CH/AEUWvyqziqKYmP3rQ2i
j7V9tZZ9FMhFmFZawoNB4e84s38Gfmc943um9YOXrY7aouhhB6DhDLgE6Yr4qUn/1kl83DWP4ZKP
6j+RPQpIQUGBVZBBeWG3R0oYR8m9meV1+LjyCkLirrBuBDmEopduLrhLW+kKWcUvKkquQtE2MDCm
nxbtPY55trGvqJzgOa7ZjTb/TrQIxh1jN245PU6/fM+CEgbOEkt1dFzuBdklYGeUBWfIPStl2Hca
P1Rh+faa2m1gdG4bmjljWNsKi7PwqoXnNf4XwB6lCg4TPtLbPGhO1ZBs8ie6KU1AoP43p+7Pwo5i
2nkpXjf0WkhnVRMRx25k0bq5wkzT7CVFye/Oj3njXdEo260MZGpjBjGcKOpmjnBG24k8t7QGKPwm
vhwVoAHbYzqdYDfxrNNBt1VOj5AJ0imIx5Y+MimXQaEEliTz9O6Vtfem/59LHwFTcuEimapvEXmP
ec70zGK60AU+oWnN1ItS5GbPXGf5jhv9gGxBlY4x4uCVZOChxYwUDa9kh4wCrJJtkFHNZcDwVCd2
j515ShiDb6envr6DUiOV7mqQR3Omdu1W8uromeXk2P7qbwlqFjyXyI6Mqs3WHNXNw2zzkbLUXB8q
7yUYHzZMQKVJY2XxPHmEwlgU5lcNYO1yGjZ5jNu6g9Ew9Xg3ZcUo4pVQa76VS6bt66mBa+OlpuO1
R705rENXQUPDDfVdbU9WZb7tS8utqbJVQEr5eIiS0dxSF0MPYxcTQKO+ull/4X9W4t+YSM9N247Z
BVr9w+R1rtKj8kP1un1omwMVx+O/reti/ezzx+avz3IfjZuPOkfDhBHDAZOaRjyyq3Dwl0A3Thi/
G2bTgjozYBmAijAWD09dQaLT3aAwVG60xB9GkwBCjRQ/7D85yoXMJjV0F0vXUWn25Nh16AzgRZY3
9tb2VZ7cuI9QofEqhqZNxlDfeBkQV9NS9B2qybqg2KCEgHJYm0K69lIGveGy169Q7JT3xUeuYNPX
6ev+pzqKusHqZ7AnCVmkQfbq1U3tA+hlgB4Jp0HBGtPr5m+h7+q+HEckomuARn/F9DU2VFNaF0R4
81o+LdkZhkbFm7kOt8AHm0pfFuhpx8deUPDfwYCbCITs1NmOHLAgGWvYDyyZMG7yDOzVdygVeFQq
GhfIh8u64mljsChwBM9ArGB+ExM/J3aEuourFPnUaS6zhZYKbQBwt67eBOoKimfiDGY/pCkxIPvm
vugEex/w39z7cGtveJBAMN8w7XLzhlo4tygXlJzgrFEFb/LglQwtdTyiADMahMI5v4+yjgPl/yvb
Ni0HwpdPW2RIiTZhpij7iPxvBdM8dRmDIlVDyAFpJYXcP1vP0V756PLodcm8NaqqasiCCOkp2sA6
Qm8PhQN5f98XkblBSN3qJNFkR1xtfyLZJAOdr56x3wX6WmftzGVCFH1gsH7Y3V1XHeT2FRkm5iGn
l7p1NdAy6FqqIZpnpEMWxUl8WYz6txbTNxgXgvJl98sQGKPNikcntUa1ce9rLCS4Pn+NmLJS3AvJ
D2NZ6YiiaWyKoKkpqhO/xYlYJU8+Gykr4P0pRhMPCdH4iju0Ma5jytQxvcIG2e7bhibCr9GS2gXl
63Gttkp840EvSJtvlD6YMsZJqfBWq8o480+oG0da7dWh3h2ILwWHEUBTF2OgGRhnXA/7LeQUHxdA
MiAD7V7xXjj43XYSFr6jLTVVJevHOdv60Re1/EMVZn8aVm7hJB/NasVy3qCWa7JGpU0Idi4+Rlzr
LZfEJLsBt5ZouGm+feS3wtMRg1lhVGljBXVpTM8WpEIRLGS3Wb5FcJun5cwRShdkgJTwVIJT36J0
xXBwx2Qhdy3EjMZHkS+4UYsvcuWtQyP7Qh+7U8mTyUBYSFCPq8VYJH8QWTx2CaubeuLA+oe0BJ0H
YKF81cKQUIBrTNKo5Q9t5xEv8Uxb/el6V2fRqe/HzLld/bcQa9hwmxCpjN3LTjSqvCZFvIY0PDxv
EVLstC7oUwGYeqfKYy3CHDxCz7HcRMPdPPzVE9O3UN77iAdLWQk9GLLMsfj/M0vm8SayIHNesWRA
AlFTJ4mFU42GNjb1dUWqPMuCPWZ+bchQRsWROvZyCb8idDYqLYHbU9Oob43057w38mWWFIOHresK
Wl6gXArP3G3EcUI7vHYI3/OLzRzJgclFLH2m1o7Vo7nCrjQZ8Fe6WPJJZMnhgbTi3NdnJVKFvKHV
AamslUL9konMOxYkdxMbWwxS1qLjXcgZ0ezOHN7Z5ytYV3F2/IEubbhg83UGnlpUNziaKd+LTaKk
jK+X5MQevd8tLl1HAcMcXAp3SiEVFZKRsDKJrEGR9f4Xg/C8whCb8p1OlkJGvCgcoy0yZyvXwjrI
BcRll4jDQNZF0nTxPm5E1k8COy3AQzsTDp2ny7HTuPasqPDBPQ7lGAwR6rJdMEUCK4T7H8zgiA5L
Hr9PpkVDYCDAZ+oP022tCXj3j+yu1SqW3JoM3oGwn9TwhSghBQRGeo/2Co63NuIlprwPidfHZo5X
t7nwCrGX14I509AHdzQS/Y3rRHYayxLr1Xsz5GtUaED21h7NU3b+n5ywiqhYUKBIPt022HEPickH
86JvSa/EmshXJmpydCzrtJZvzNpGtFyoMWOxKwWzi0GU90rCcWUNtPgWblXjtPyPdtD4rXsNlkfN
Cm+7KKbSSz/LdIR9A7B+FFzK3TbwiVnEIZ9QdtWxsKE8mvy3aMRNcTeaqQ8mQK+nguxo0VhIfiRH
ndnhCqyfMmskpcTANGMoLrPGB+eHZYZW8xk28iXFCMz8ivDR/NtDT5U31ToT0zoBlQErmfD7kN/0
b8GUVZcZr575ONmQZHoMvZsqRXjij2+XyFed/KlhLLK/45+1IDWuIajvs1dr8wKsGfajZkJDYsHx
zOGUwMy7Fvf4XVHPtqc1SEsnqX9OYLnbL+ye274UsWMIRIr8r3L1CO295cSj5UHHhx2GvxAZs+9O
2FO8hC+TCPJgJXo34c22PXUTRwzGLg9Doyek92DLMZpuSM64jiXG98VuvjRgCEdd75UoBchWYNXq
wzI9jl10deDLMioHqZrWQsVxf2wMldawxxa9966ShJ/WKS/3AavTJjUUeWjVI+bEafzdtd9dENbt
nLW/Ib5PYUMx27vC+DT0Xx5lS5lJib23BrVhDi5+1lCRN1BKhjosDlIrlJvOE7mngEQJm5Nw84XY
KV43+23kuOk2IJcjSVuOKjzIcKXs+BkdUefAAQ7fubFLHJ1iWQAGXbudYktC+xP1zpKnW8SEn3J5
ScHd8nEf0N3dAHLK5KqIRbSPAVnl8seUlmRPdutTnjSh9ZQ6wRLu9IkcB7tUfgLpX9ySGrr74AQ6
OaK62kaoHcru8IOcU6H4+C1YAdeI45SBVp1gcKF5bSgHyxbVIgY76KGaEOnjNFi+2aHd0C+YQ7Zk
ptmdn58LWrYuGYunDuCNGj4JmN+tbwHeEM9geb8gzDv4KnE02KrxdgmTi2gnAZ2mvDWFpxbrh4x+
HMrMiq+mL3c3iDon8dkEEgSDqRQ0s8xW+Fap3gEr0SroMObjJVZTnUPVDKOowkWHHJ3agRiFsHSP
ugyLbmNlGQ+N5yU+uz0vPDv0FjfZ96DeIJ9KZs8uZI3Gu7B/fmIYw3fAkEuX36oqKcRxFwFOlKZX
0drYBplTg6rgvc1mTqCXtK9HoX2gBFkob3UVESudsolyucIk3iuF0Bo0F+hmkkwRXHHZ8SPapeKP
F9mqVbd+R6I7/ax6GLLcDlmZJTRRaRsEGnjfeuyV/Uc9A2vDjeLBTLEkgsZdIzlm0GpMmEPy8Gni
5SjzaLamV2Fo8jJwwTE2f1EpQN9rv+v8FdOHT3/POZRzdwNNHBZrQCkSqwHFVG5HKJVzbeYZjxYI
gHJVQQDe1h3zA4n0g1+AjQcGAbCnQqEJNhGfDAxavS0Ie5oJsepz27jrS7vSCpMphJ5FwgnsumWU
Xz+tueP3gxXHHCEoZsMzHw9tiotQl4nLW8OWnWQjKav6tlZrEw7QnIf9HpXJMQD4DXtW/yTEMpKD
kMM/cJEQbK9yRfBfY+lmbxnHbnI0truFdkhak69YdGz57Gbkh1NCI8aUCWHJeiAr8nwy2xJ0cb7e
AQ13Sdy0i1q0hdRYfi1JqppZq4xlqOuvKNy0zJC/ctFDp9kKbytT40UmP1PJ1HrhaCoAXaZCEI3d
tKgUXXINmhxFRK+IXLgkfMiSTOewqagt9OnPqeWqrb3N/WTuAhLj/4IgIYn60U35xCXo5g/R7yL+
8WcC4AqfXExTCKxSjm0H/7vF/98A2T70sOsZAnsY1Yk7K/wzpvqqfB2qirVwxdMfmPM4yPS/1mwE
wQvfOM03v8VB7rMCAFWByqJhXfGzAK1N2gV8/GKcoImuWifyxg1BMqqGC3bI/a/DkFnjNRGbjhmV
fQZkM3YxQkFE7ZA9MGA7Y8pjrRapM6UdqbsPz56QWu/SoOx/1qeLFiHilTxoB246QFAmG+AJN/YN
QfQIftVN0v3769sGqAtDYDJdWpjxtmw1w+u1FWo5efQfobHmsVEdvyfEzIzLTCL6TQVkNDcUglXi
3TfWIMer/jQcEFIEQBjGR9ErvDwMU6ErSJJfH1IrOd0t9PUILB19qvKaYuoQUffeHDXCEER+ApjX
zA7Tv1WAN+c9U73C2tUs2jDmFeekZJ3mvSnQkKlv0R0+WaEem5IZ3Ie74laLMjyx9cjqORKmVV70
LevQ3yEn7qA+VU2PD21Mjoept5zQfKXklS2tWPRcRlQPNRo0e4EWnB/RhHuX/LoonD3BzjRIx2dF
kcYBh+5VcGgfq9hgYvaG1uc4/GFw/z8PBI0LtnzPnsfRgxkhd8Sb+TSf8qwQE4zTcpQgLYNYDaH6
PrMkBSiEqGYgpOc8TdBAKRcqIbwr3LHk/VB7NSg7ryC1EK02ACFcYk7vQ0XiC/+nyWvrtAvEvKkh
NtItzzj3QrGPHftja+8/zXuY15rsDqMaBMDTudRFZcARIWllgu8wm5CT6AzIteI7sYIvE1iF9GA6
OCC/cTN0RaqJMPgBP1x0LRXL/G5/ki1pN9yltcxDAeIN6naS6FDdpxjOrfZG6nB65Im0iEdp76xh
1GDdCh53Blf36/kn8iNuYh5Xq9MtQtcUsJXDi3KmmoGiA7mx6G3yi7sv9DDFxBG+Zp6dxtLJz7Fu
oh/9Ou/iK940UHlu34eOzznOKpbcLXJWumNTAkZoijxcuXEQR0ijGOYSxmZGwJYVSBpqa3S4iviw
pFGzajMtvElJGc0O1GItSrsjkuiJ/HAwFQ6Dk6yQHnB1Q13GxLJ2mQu3O3pRM5g098jzUmIyrH6h
Zx+WP+onDWFxyzwb9NVhRfghX69zFWReQpGGL7k2v9MWNT7UWqztHZc0iFNIHifu96ouGfCnmg9z
RZhte2O7PW5hooeXMC5+qRuNz6lgopvZJL5pLO/kwSQ9GS+sjf5izm0iKq46KTVfq6nxueHjW1iz
e9M13jiLna/BgEIRGI6LohptqOCTALfKxh618DGNH/qFXOZGBs8cKc2xUE1ebSAq4A77PYH+2U1r
Dvb7lKrVeZYQuDOmNMUrMUPyefe86Kx7TBqJAsoyPIpJNzcjmIe3TQnYPm9OcAO8bzcu91x8OWJ0
O2XjC43Ew/yis1cgHa0FEWatDOm4NBG1UtbtOqI4hXoe5F+QVNDFQtcXl9kB9WJhxFZtpluCiB8G
ZzTg85gyc2jJ5MtwvbvjaHV0M+VEDInmaaUw7MPFgZ3rA9e0bAgnIh71s8JfzN4QOIq9aXK8B6Mw
jqPpb2QVlGgXZWvxTeuNIuQO8qw6Ic/S1H7fA+vItmBUv/vHyFZYGeZiz4FhheP4HilJvZuPHj9W
Z4IrNDGkaRr9+Ux4282awAiBJWarcf8JDVUYC3kVzG6vHbsRZcFvMiR1WqRv46Gw04eQkW00yHuz
M9qQHeSoLATuaIu1V/bfNf/w4R1u2KWQlgJ6DBU07G1or1a+zIwqNQOxKOjxgKSWp+r04pAUtFDJ
Q/3fRr05/2o5/4FtTIre60KYC5CVSk/JitTXlgjEtb6bP3yW2cyepZnBaz/j5gs49FY9PpdZpiKm
u+CQT2ZP5mKIUZiVZ3KIzchenyBRcd7InvwKM6ENWZy7uGMzu7w16LoTeDhjiEYPVon0ak656qtQ
XA0DjZbA0bL6nTSg6Bcnykd9taoCHlxq79ZXDLdkjbB0Mu4xH0gZAnN12HpZ55gRmp2sIss07YTb
P8YexlvV930hC/+2xTqqiKglI3Bz+N6wBKJJWcWMlxe9ZQbCIXrp0HooDX9UE/lPRcLzT+U7afrw
zFvrTRjT+kQFsAeM4fLtI1SXvu8IySQM75MqIOsS+wQE7pTgMnr/QfdqkSSg5UrTx0aaneoZZdLn
8J8N0kqwzmQ29ndeYITpTRM+zyEJ+5xsv7/4BnlyQIr9LiDYrde8ny9lrE+YH/npQLJ2qCrVdN7R
X2rIkrquN0NWgqQA0ED7uL1/BR/vahvHmTu17jVd9yf43/L3l/zT9k4yFLpCncTq+OgLePR6gC+q
e2Vphi8xIxS/nWt0JRozff2/AMLMio+6mqMWTzoW222fb/MzG2WGDxGPY3EcR1bju8clX9vR++Gt
TYau7iNxijhdhAjM7MgIv7PlgzMbfhxZwhwBskJeMqtNCabqP1L80K9PfpWJWuFlEqe4dm9rfyXB
+ZTfuvaLyvUioeAxGpgMG4Y5Bob743VSLldOpBP2NV0Oa88C3H0DxHMLmyiH/Jazl0fpBM2OFiJw
Z7UX7pKr3W3k67uziA+Hp76LqI42tvsuEMlTo1b6O8IAweymqAl2T8W8eXQVdHgg4sMYakSXc3s1
A0g9oTX4JU1JZr5zJxcom6k993RouSfy05+9MHVec86hfv65yvnfNHSM078vyLejBT+277nhjFgH
KF9U1AD4VaIkYsiyTGfJ59hW0Zme6BIf81QBjY9F4HTyPDVbnWfWiUTu7xwa8k3P/q6Zrlu174NZ
ylZcjE8GsYkhh5hXHEpTthc5WJNQwC4dFRaoG6qi63qLUgFHZqMSd2AllJdgH0eMjsoGspJkAWGt
J/WbSOFQ5XkI+SomPBxF4NuyOvZyWy5S0eMvu7lUHegjVSDkROhB1jTEuM0MIFoulAvdIL183vcO
7Eusq8hywCPAQQQzlVc05Vov3RNOTe4okT9zt9hMRcI3swo6s4YzIN1r7gN59ZJm4U8QQtxQ1rIb
PWhqlt73rr5AX0IlDa2wihGOUbYZ2PMW213trRCtbcOKYmRUpA7hqdLsF/OUz5AChuvGSsUjK4WZ
Qbh08VHTrdEvEbSwm8riUp1O3WozScOMsLGhBmJMGoiMq0OoIczF7TNcBz9SlszoDEvlt5mguJUu
hU9YdVZnZBeS0WrUCkmwyZPojhWGHLhBL9ej99v0oRqwpO150BybfUKrdYO4sxoP6tyES8IKNRJ8
fiUD3w7GJwj71BlwoubJDy01vWJE642IiM5/SOR/WOwy/sdeNRt48YvVlAksRD+3HFr9zf9ZaXRk
7puQ5Ep8ownqGdWkRqnP/3a1Az4H6MNd0W0po+LClU61WZcDpb0oqLWi15l3HOwmASMTnrsCcyoL
Fp91CW5VSsRc6ssw7LFYxkHH73Eibph6ndjAERpCQ3QrKT2AxKpcL+05+mp6zeXbxVpQO4zeqwpf
ouGmP26byAHqXkr5aJZnhHpyei4wvpth1pDSfQX3L53XqCZjpNBjfbK/jgr4c5jvQblDWOzEt+3k
bRoLvCS7obzI/KCW9FqIkpdFVg83/pRFSmGdBKkgqWsROPC1PxMKv3CRHkGDco5pMQ9ioWmeOW/z
bVd84kPoU1ZF4L+rzJXavh72SeEjEMj1CwyEx5BW3Unkna59thgBygMnRUpWK8V0X0FShy8ZiGtB
14ZlndalkrWH2orvu4vSRedf/vACgqyo6Sz5nTpYO1pAbsM35pZQiUTZYzpTdyz2co8LVsAH0EEQ
qRY+CPB+B0iTnsKIGpTORPVccM3mN7qBCMK9kVWhkmresm8ks9BfbFhx5EZ5Vmedb4P3AGr8XO0l
nDn1sCNoeFEFVwilxzTtEg+BqGYSVXqdJ948arogSsCB6goEqAbc467vXvZPZW7DlTW2J52EYYl3
JP3+xczA+TaUeXs/WnHrE6+7BGvM7YlpMB42BBxU3J/LGIteYIvzfdGMC/cfrCfF17UJcyYb8XHS
HQ/bGUPdG9yFzZtkeOKiPw5iw3jzLD1l2RJ0pApuEgCdGxjDK8idIRUsj6lzyTAw+UFmDXG3L2KJ
yvjO0cgHIkhEBYfpOJahSwhp9Um+y6d5PZALf7WJhP641buh0zIYtbJgwK7mR8+3qlJb3DX9hNf9
9N8+/XHy1lFT1bsSmpt9pPSUOCsDo2y3ZLKM1ggVE5E0XBsWO1yKBzLwd2f0vcEdfFrqly1O/Kf3
AcjRa2xB8zStO6V+UooMetxf7BYCO9vq1nlQ3/pmCjKLFpFrFC5vnlxVghTBd3U459LfGpLbJwR1
JArnmTstUmRysCxMi9Mcp+rJ8ii+B9w842XZ5Vdxesfv6DRSNupXKrWiJn66xkYsWbJ1bbG76vwB
QmM8mk9dOfUNBWpDzAeHTIS/KcfSo1OFoX45sRwrSUhqvFoKnIEfFNYOpV4YXodwmjA5U+llps3T
hcaLREf1XX0g5y/hKtBCRluRpHRh082pI1I9E6XYt/MDjeX+9DbtuJ1VM2z2O9kJlQ3o3kkocpL5
zZ08WhSlgOM0Y1Rw1p6EudQFZe/7AFxWeMFXsAOmf1hH7N1bYPhfaC2eRfi9gQBpnLbjTHR8RAAp
I8umESV7DFsfGrI72zWNrLWNRlYrz1C9K4PXhkElaejdeNDeLoEGXZg/MPVbKFOHslTHfv0e7tpt
3i6dayYYzXFKM3L9I8q5ql0D1KWV7O2lb2l6o6Ab0Ds6FWc3PWtXjp0KrBa7oM3wk71uHNhHe1Al
uzvMnV+tatbY8ZR6aJPrleO6l30wRyqA2kBRgAoa8d/qKz7HuZTqvKJsOB5hYk+xMkNK5QsQ8sQ+
VhBFvLDWHucL4RQFD6ZJsmeSwcNxG0vUyQYBGIbBWKW9He19tTBSGtYFpI9fuZ1df4uXP6um7Zpg
9BBb6Q29+1KCQfrNNax5MinYogmGuU2d/vKFr6suJTIBfmQLN6m3eK8GRfUyRl5bOx/orNwD3Oh/
/8wq6PrU4ipeGUoZOemsRm+CItle8MQGIlFRSUBbDigmK5fvAZ6PteWZ/V0WZDkPTKTo3HlH9LX8
lmQv84t+mJmjV5U2m5eeWZhxgHtcx5q8aAnKvsH56p1w6EtS0wgd75e8dsHI2qvT/oHGaycvVMlo
fFCp0jVtZiHJNf0mZ2cZOydRZ4qeLAZ6CO4uGA+e2eHdPJgpLkXYL6dkh2LQ/WQymrVB+K9QpFgb
cgvi6aVU6OG5pPxd31aWhMc7BrIht/42qgTaJNDLPMzTjQA5tBvM7zVKB5z5SFp+j5peRs2YQIe2
zNO4fCRqH9atFFKiGmP99ozW7fyBQzlvmo7Wk9MVx2Tl3y2wlOsFPHEaAikj0QDJAKzgSVvXcgvU
toqx88XWMkXTd7FZh+f7PcB2lWVJINJ13OgFoMtLx7VQKRS1yqY2t1oo+vTfTkfsmPoSChaY26Rq
FrqdaeqHy6Sn0vHfhK+NObZY+8FTf63yYUOnHA7q1+dmNPzSDW6x4mgUxft7WU1ow9RgEWwRJHEN
zLy4nG0UnlLybWD/ZilT8rbTwcuqVSXONdRiaNWAroXRXLUIbZygzSrA/em2mUmsMyMmNoKrDIm+
XJ0x1TZOtnqQEDIC0ixACGpwASD9+fpie9X7ICx8oX0LyamvrlQ0xg/ICA7OtHJxGbdb4v3omPZo
AG+OseoMpe5z9cSj8LzGBL9EtUyHLRlo9QEkr+0uOphQ5fz8Yz5CZWnlVNwNWB5SgWqFVVlhm33f
jLzZQZD1GQRwHaoBqMNqvTSy3TTcW6t3KQE6s3MdyACjrW3n4mGWUuZQ/esRQ0vFvJlcAJXuwznB
K73xTup6WFaxTxWfgW2shD0Q0RRh
`protect end_protected

