

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gBBqHtY3Bunn5h37HpCTrctVa1SkpXy7VKKB+BLoIpekT1JpAEXVRxCRFlXm11bUuVEv/j3pO5ho
t9pTutZSCA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rT5AuEipXCjHo8d7Uq82KPZlLJRMWXHoM2CEgdCzb72AUhqeRT1qBpZCSEtuISLEowB+OqwVoPB3
zybnMbwQb0oxhzcN21zHYr3IRmDn/uWaTM/MMZ/bnwJHAXofyVKi6nJ1ZcQvvuVCoGL8KZKn2sQY
BUZNn2IeXewaklPHIeQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ddHO5ZrB/psVOnMQtFAGp/GctaRakAwKZKpb8fZB+TnHO79YBQYZi/vlr7RpKlgamWNfGsIyviHi
4DIn7nUd5XwZ9QHp06khu4m91TFepB2UCDybY/E+nqujVmmRIT1MbkiDUkGmGhdlaRTui9BlBtE3
0V8M0AdcuyXLUOGcPYN1g/l0n3iEvu3eoNOYYP/kCy9cKfwaeQHNoZehf77AMdR1pfynz4YwSujK
w1CXonssc2+GvTDEUoLQ4/Q8xeAeoZGD3iG6YPZW5ScawzhsAidgis6DgRGKTAhRGMtozCJRfR8G
WFjtcUsenGju3BFqb5waLMbDwCr9/0sFXCYQWQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hcWMtjkawP0pEAeHRPrwjlkoAY/aJ/OE55+xUYc5sOa68hwNrmj1qF2ncvb087ShjKLuEH0jfkUo
QzvhJlOJJxno7QOxZuWkvY91+e5UQOL+2j631nFnpoZE+MloH4Mb5itp/2QKWciAqiwm0+YgSi7a
rgZJsggXf51kL5HqrmJUBWR7819hS9n/qP5XtJ8y7FDBu4ElmV5DY2JVmGTJzFc00gGCP6g5ZCbZ
x2WaYEa9rwkMAMQIYDPF0j3AzZOJf9BZ7TUjt58OKt3LANApygtniZkFFlRSo2PBSQ3No628n+ht
7Do7iCucrGBsrniezp+n7TPQFoCS/PsKj/0Zag==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M9pROQR4pNGukvruDI+JPpAyg6zBwqv+kvFvbZWk7i0NekZFvWp7FY0oY1eWZ+XxMsuNHPA2Plg7
MH+MJl6VkCL/cJ2+knD2NcU1AoFbgFqErwcWRYVepmitEaQCaZwfy82Wax6bBGqHKP4X1cQ96V7q
2rHMe6dFzQ6sbZJDGr0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YmZTg65xAenvz/Kb7OqoEnjCRgOo02BX9BzONEy+LExgkp5FbIUmzte7VnUBMqyOfrjbhR1gwsSC
E7jpY1rpbjcIx+SqgamXNDfuW0JF0+C1zkLYSPYugbcrMUXpChGH7bk6WesFdUAwr/Ktyh+Urq7s
BsO32fxnO0rZxYMJ2voFB2hV9nZov8aL7baRr4ZUYDmQxS/z1gPpjxqoqa1AuT1OEpW954ozW8uP
b9TWRqViZmVvgktghhAp5Woa6dttGplqCv+T/yd6WcKv8U+Pc0RzryU8NUKwL/WxrBgu7Ba2LvO7
g/WeYyKq+hYf3O4ZtyuIDfGHBhcpqCUnRRVPSg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XSieXGZEsQhOJ2iwjK7eXEWDvgXxCQanpoMe8ioBhtE8cJi/QGFtNn5ZnII+9PCK7NrWxywdcuIa
c1zWLFnxppl000eGkfeyNxHN6jZL2+ZFu/PdSDS9iHl/x8HlFh40DjlqTkoxZLUs12OKV6MsJbnz
eVDzsmiGuMCtnR1GD1O/ajyP4J0vmVDwGm5WTY8NXRuJODjlsSgGP9qnxTANsE2CJUW/5VjwahFd
lnQc7QKxVYFfivRIxRpjMPi+njmOySEXEEwVklTwOXobxyeOZ6mOeReGoAhbJivQnsxe34MignfB
cR9hfUmEkcVU0Td9FY8BgXjUjjeywjJrKoW+WA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KmpD3XZFpLe8+sD1iGwEup6bfACKiedaS21mQM1V5CyQMjx/p/K/npJNenB77Gsv031GbqLJWf5V
fbT6GSFj7BtI+Zci6hRlAkvZnNNqCaWgoXdIoDE+CXp0KnBn5CaDdAN7GUQ8EPx3UkZWDjZ95/80
Pd8OG/SZdQpnjtHOs6dZDthcXgcestj5Jl3/O0O4nevBH+OB7KqzA8UymTcf2NHBnCx2s6nfDbW2
C9LgfejwT0EL1/dR0i/f3AwiIwwTCQAXxFiE5IaoctK3kg/KtdmAblRzXI6FOvwjGAZLCzA5JXkw
Nd/EAOBJn0Rk095M3rpMJruHjbzpAn3t/WzMzQ==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
C+FB8r/tMxRA/SU4aH6F/elCSsnz+M7jAys/z8YFGgwvumpGQFigA0D8dS8S5DvMgxfak7tlkOE4
LEte3Em4KJ2VUGOWsRCSJjerMYy7DlhPZEE2q4yhdU7fz4hQsYWnnuuHt+uEzyFMESj5KBVKmURm
a054fsL6z4UkeMEwHG17eluOnEb+vJWan2hnHekSxUgqYY2FX3PUgRSO47TX4qQiQa4pdDxOB9Nb
dtmBxXkxa1ey15e+nNZf7ZKQin3MH0JTFjnbz4n0D/ERFnXqnTG4Z2M6RKyohLnj0TyxBL4Psmgb
cJ53Tx7rODwX3skEPgU3YIBRbnoh03Sc5Fr2cg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
HvV6M0f348fbm+2j7xJUTkyfhlC3Qrk5Ciyyu5KYgPHztYMhoHwe6SFbeN1mUxKewXpp8nFk1tUT
TLIVnOoYO/V8Ex+0QQt3jXbZeUC7jq7qNW8cVIGLhtFbGXr8YILPhHsG44eWLMB8gUmcdWxbHRyn
B8O6abV9svAThlpL34tbuhZ8mchpTXLqTDf8+nrvZsMJTiE1GQQlmtekq6bbt+W5AqoGbuEElHlx
mqdXqt//BHeJjjYA/z11uZapFqeDg4i+rbJgU5KRggRL5SGXXqu4FwlL3gO1o/QwUxiW2DaeWoVP
cihoOSpZOegDJZrtxB3wdMfw48ZJCFFE5w1Y30wDYKRrE9ob56d2KByz9A/I0UtcJDu75teaivYn
0mOVX+D6Ku/XxlRjehpp4X5x+pcyC7voiuDYCxGy58GVfrRziIRIyrCy3dyW6I41ECWaNsNMKWW/
vjtMOx2lYSYrmN3ic8krpNGJc7hQYw29PpvOckq4+09/qcnfsPit+OUGbzkJU47Hy5xo+/lrCovn
aSPw8cfkNWwxw8o86zWxMBlBzBNSPC75PX6QrHO5paCa7Q4HE/tDCB8t3m5oU6585fWxj3i2ZdxT
dVPVJXJVPhoT2J4uHBltcXzi/B4480oAqzfUDXjo9/wTSeW2tyiOFUeBAAW0Rq7qI79k5jKEPgWT
mHuHfeZL32Ka2ZhbdlLsI3lWbsfTgQlN+QJgTjZ4Aohpk5dbUe7yjiQhAcD17jkS4G9R+Mp+Tsm+
nfhOXHwF1k2HiTuU+UUV1QX7PazWo9ZZSiMJVVfvCrZgAmAQExCouIW6U8RdnWLHR5rJKyckvDjE
T7LwrWuRqgyUXT1E5cSP0VOLkapBRBsUWzMr71vElaxtuJp+bhDOWlQbH54C1ZZBExJBR4c25oq/
0KvUyxgaA+BlIa8FdjZh9AWN8pTY7IJ9gMsO33tPnJ2bOxLvSkU8IJ79Y4EJgCE2DB+NzA+9neWP
TexEoxIQ+IGb+k5DccxrBPFH2XNHQDbMAxRuvuH3mLll7mKlsw2eyWr4/K5OMRq62InjTSd1uem3
dfwNrF2NrrkDTjRc8+DL2a96U1dRRxG55nIiTNWF4O/mo+7kht3muGYJ71BZwh5SLWo6D1OY5wF6
q595YKDcg2d6P0IS5ZkPtQMDFquEVcdTr89QjDMdUPQeFFpEXgLyYNZckMMQsRVk7PDQ7KE+oNGV
/Yq9eOdbgw9Vb0aNufRPdEudUry7qrzVl0hAeH5e66cdGo/iohC4M9E3ub/ZzT/ZG8rnfQQ2Xvdc
BoytAlSk9sgzqZ+HW1vuZgfjsgOOIfBncZMY/zUWlxcpuRLSau85/R3XFmn6u8ENdHwCQqvkxCuc
zwc6/gl7O94oa+ax0qgKRjuivkZpG/vhbdXv2QOmXUwUcM4X/lljtEdqdDc16F03Mf6KrSG6qHhk
4/KcC4P5w+mZlx4DZHjtm2W2rWAJJhSt5PO8KlYf7vKKxQrXzhmwPrpZdTTnMSUqhNQbFB3pS68W
kfjvIhKZo8x3nNYcRKSJm1RWUVt4VqAk8/fsjPLH7k1Lu1iiYdhHMSBlv1vRRul3mgWJVxSdO0NW
DruKmEOemWEt9YpohPw1hwkRKDdQq46Hlx99KZTPRxRNxtqb7qdjKuHcuIatBe3ZV9hhEL9ArHD2
+7vmDuVfQWBe8Exnlk+DdYIc9D5WCd2mQl1+ZnF+MOQMHhv+G9u48sC9w4aN7OCW7SD9G4kdnitj
8utbtk9LVimrHWwZrZ9maDWyolw2SQz6h/XYAAj+K2xP+nrO/qwlNTNFUliyeQnyqZBTxcua3kOZ
nRaejFSgHbQkcjcVTkuJm5C8G6+R/lvk6x0tRlLUZyLZS6iDsOaBtL0fOBy0NEmCKTdZMt8BI9SJ
noNoHDaXnQnJ0lUxx/DVqIxwxoD2kL6ahDaKOK2paSX6oYxp22KMeL1KjweqLPC93jh5lmsOzbU7
trkDm6WcBgDQ84NquNPdL1BzmoQ1v8nAx07ywZVTwvUshzmR5i8MZUqjliZSb5lfEsWniudBd+u7
7VPq7AReiBQxdahAMiqfG4lPEBZ0BIh4FAHilrcFNwU7mXbE3z32IisSUh1GEGA70zLv2kAI3+EL
ozUrEXq2XZjM2VVi8/49RtApKFC9+tHmF5/pegx3ifF8/sN8C6UXi5wEq9lhBZT8Dcr1eKY2Ajuj
SlQvVkBVn3Aohw4uJsCxmzBxNdGEW+ZBQ9FpfYmfRy9kWfbbnoNM8EiFIP0IhWeEPPIfsjyLYZxM
2hkcGKj/NMaI5Y9u7kF5wulqqBAo1f1o8lEdtMzj+NiUQ1qq3c2lbwCKmXakw+E9VtKr6ZiW4a4t
mvhI7idx0R52gVo7wfomZdTTF05+V5Hgfj2h8KgvhhB0K+wf8xzv2DQxYqM05c0O1GAIUSWspzAA
/MqDwVaMkjoL+4OqQ3d2i78IZuehz3cqaCIs/jTSm+9uAtR6J9UqwvzWiV5cLojVpQ5TKbjTh1v3
e3U9ViSg53+ZwgQOl0p7CDui0INAl5UXuqF/aWdPWjSk54tmjGMeb2X2eachD/8vdQouso34pgqx
/vm3W4/QyaYU9WJA6A2RtjMgoUrvx6Xx/DtOON2xlAqnvuZeTnh4ndHBylIEecogqe+Tk2Y6mWdV
Ue5dg3LSvIpfXo0UXU703rX688Dyec7ZJ+dy9p1ya0+uV0tx0JuqY9Jt/Q2MAeTsc2y4O4+BGwZd
Kz1+PQslrsPlE/wY7hH4qSTE6dRaKAkGzKYE5IqmzSycMwz8yZ4A4L3whL0QzCxkw/tO4zCLMI5z
DnBBtRJUcEs9O1UMqhvkxFnS49DBoKJu0LpIi9AOX2Gdn73uCJRs5PAZnv5oK48z4oD3E7rEenRx
wllUChuDRBBuS1EBA7ZUk/IwUQxUKEfk17PGo3/qSu+yHHf+KC7s+jH6TSm45N2MOuvSKpdQgstO
Z+hUjO0jIgdlQalDBUcn6q2Y2TkuumLY/OpYAUhUquxB7IG2QJinuLK3GszY1nV63pfWNZee8UEA
doErk1v5YBc8MAz/JVgFrzUXnhiM4lCBpwcdOZBpUVEYJEMQTSVqthcJgBqKeWHpd/BxixTaehXp
T3jht7TyZhuuZEX8okyOPyiRHODeXWFVGXvsCQL2IhJ61IiICC478W8DdTe7fiwbKHQvEdDc0cwS
NBuONQwAoHihkmzorng/3C3Z8JXdkb/8xEVH4mSEYPRCNpjVK5qE4O8M29B64ktb4RyyBvXNqoEp
2/Bbbsa4DuYYfmVs0khWJ+2SaSuojX7F8S3xWfX6j+YGT93eoQZlcaXPXx7NprCZeItzmR9MD9Ba
Ou8TiXPgZHZk1tIRuArxYibY8qhfmdWJU9Xhfw4w5H5nOnhi5Q0yidTafmSIzr4NIsiJBhE4Qh+Z
MHmA+l/fRbJ3GZQdIfUvGGP80FE+mr1QXFjA9cGZruXv0ynEDX5Q8tR8M2otbv2yYZIqTC6SUbgN
JGR36sQpcq+RbrPVDZ1XbodxCZ0TpHsteCjhr/71lCySMQlpqrSqEjMZbJqgKA4bTirsk24ntDzL
8sWmQ5QZx2zV5sFH81Su6FdpUCyNlZKOjKTRVg0+GHZsR+VeFnxnM8rH0dTyzoag7Ii0lNSiEq9V
M6oIQBwmJRqCteoGV1YJoaZ++xFUde6pv2IVX6/pToLV7LVG0CypVsiCaCKToyTFLGOBmKM1E3Xv
t+i6dseOA9snkO/0cF1X8Hb44tjgRd9RD/+5f77zNjK87hwNKVnoXPMTXXihxFnE7SYO7IHlpXfb
PqWoZ7+3Uts5esmXzFl9I4u4h/OT/cR8blgRPz23ecwLp8HQxMQSb7Q0hz44HevNL7q0VRxZ9g5b
7O8T51bNnRUwUpLx10qNTEO9ikzeKmsMbRlYsWXb5jt5+S29NlBrZmnMxKajr8kNpDlAvs7UuXXz
L9qLEBj3D+o75zy530PKe5I12PATozwiiWQJ7zb7qmiUWrfekfCi3Yp7ZJqbsV5yce/CSylG3gc3
+7a/plU0SHCW23QpN9NnE68xl//uxvd3HgiY+75fA8WwDIvD9g9lUSW9Nx2Xa0faUBJ6GCpjOSIa
BTwNItdOBgk4ppMu0Xj9yg+GracIleksnH1+tLvVl97IfSxAX7tPRYLTaTBH/rXbIAJIQoKAJ0QI
h13lrFe1sXc8z0enjlml2yp63eU6YVcA2X2STZgmwzRH2TCP+G+WjnBrPTag8B4lCwih04yce1Xu
VomdmKQ11dUAO5UMQW9FcnfHDHG8iFkUvjw6ghRMsf0mYMpY97YnokkVt1qvOn0aK/xdKc/WZGEm
Y9tMVbKQoOnmgjLrgkXirmcw4O1rL3DTeDQ9QdwTyksVtgivDDs4sPUE3gxMwuoxXSZea27mrghX
At/kWNLt/dKXbryzdvLjT90C0zqv+GiD0bwQy/SAYscKgr9N7RKD8X8Q4jNe+ROEYIRAcAzuLeOh
YemsgfykvN5coDg9I/1Gf8qzpztO5JtWSmbpAWQtw189nkjm/L7s8eixTYyy1iLig+4LTp9960AX
EJleuYli7rBkhKa+vS42YSNPreaUQ8VPDORSX2O1WaAgeIZV5tr4oFGyuqtOf++u4ttT1w6bCIzJ
/MXasK7obeHdcIsYkMA3UAA5A/K5iqRndGe9Wk5V9l92h2mHiHOr9fsED1vEleXKES/yHWdsHX2I
p63YAaUhqYXh5MzmzSzVYbicY76M5K2BtuLdb8/mncKvZ2CgUNBLkWagw26WfGI54qmnUGAjDIkm
09CiCA7Vl/MpReAt6UhwkVd1CV4qr4K8a88Wf8XyP6kKaLYnGfLhXQAk9o7aLBWJJRcSdSZDqYeu
EstLX+FyoB+IrZVdVBAX6rl4OO52pU3qeeKy23Tv7MamKcZrQ4NHUotQa687LXeByfRMbutXj5+Z
kZj3papNmuOL7obW7lbXJRmc4/EMzwL4sxZDI+dn5qAKsS5IDBM7Qo+bp4fFHhpyAn1StOXPzfvE
pUHxBHav3u+1cEXelzi0uF1RtQB41e6m9+lmq0H/Bqk99TuXXzNhKT0lfMS+VSdHURX0KuF85hht
Ky6NZJms6d+jMHuUtoN6CUGM4Ad8ZWjtjKMDzmr0HxmYydRDODOn+xr10zJr7qsOZ2d4u8VhEbnw
jerM6Y0mSU36WNe7pZ5NgspVEyWQchTl3L4w8QD939Ixl4oGRxlneyeu+s96/OT/HolKepWdPwN8
LIUk/OI6HwktoxGTWRJiHBo4PF476wU8L88QDUJ3EDXNkq9dGX/Lh/ydT2R9qZAsqGdJq7ugCNxs
FCq9e8bltMM1x/asx9XvUrHBDyz2g5OhEEvFBtCEtHPiD9pucCpzLGLMX/bG6X2r84Q+8HCVjnK8
oZ+Z7kFIh1WFjrcfc1EOF48VB3naoW6tuT160mnaxKdV+I8hUKmBS4ij1i/Blt57CVzQqshIIhtp
Gy3ZNYYese+CAHTgvlmZbwPXlYyxSoGhLvpwyLb+Plzw0V8fer86kO6pUNjSgc55HbeYXuqM6Uba
b9cwzI+3BJvBGaW9OUrLEsqNocR+hdWxu9PWrL8td83UqwxHDIzy8TFHPfVGwdNeDaSdNzTCWUQT
/jd9Xs+3F7/zbA05DS0yvgvvmsj4ZmXnuYd+FlkM2Jki3OMOmN67m5KybjmlrZpFkCF8SVLYdXsu
mMqLyM6l0J3T49ZpWF9kJisANoEhuLfb3jhBmp8YESEbm40FXs83JZLsL3nRfl0G2oEgSGphJnjM
fY6kxBBjkWBphWcw+16PShfsfZtMRlA+kS7T/q4zXtwcA5b725tC0SF2Psb2U9QlvCyNumW4zeSB
irYNweIIiBBYR8nrCHeF3DoE4ratoB1p/b6NGlT2vcF9qMvyt9GhHE7dkys2dRYThUhqwcjCYoZO
s4ziE3WVZakdBg/bW8cuykWBLuR1b1SBChul8vnJxoebeIvP9nCGJjFJOJjCP3Mip2bAK9sqQwWD
XsRFAo8Mpb2/ntFxFaeldXUBqevlp/P0WK9KPYJKB3wEJl1bDT0suXrU7lP7nrTPMGPQ6elnUDk6
QxBVgK99x1ijM8S0KN4xgAwhjOM0mBW0D3GYYzisWWaNSKZJ2MGvDBYduMypiS1yJY40sttvytzL
ukyYgVkrJMl1M39MdkSG4p+TO0YZHFqfL2AVZaSsWr1UDMz8WxJygLjy25NLppMiCC+aNe67diz8
jX2BTCmC3WXEHn18AYJIomB+7npMFZSSshYaLVawqoAdU59nGrtbkIUOM0UOG52mU/hZ/9zXNvr6
dBdv9PG0GZjLlSlfjL/3VzHiaHIlXFkG46ge/oBvyfVVqDPl9VHxyV0MqQWRgQ9oF+pKDjGFCZ7j
Lf+Rv/DhCsnmBNmLNOCx/907bUkotQ+bnAn9SUea8crKZi9x+lgUo0ZVzfp4j30oBM5OC2KTxHi9
LiS0ImFM1rJlmQg42lh3PhQmvA4azRobGbHw2JpWNi5gJ8QjHD6zlffWBswdI8NHRdDA89Y0jlDg
iprDtZsmT8v3sKKdsqg0H5KP4mq395IMZJZcio//h1w4tZRSTEO49rI5ZQiopXkI9Gs2QCZ/E5AJ
DjnmzAv3DFuM68tNIem5hvQdS9/j6iNfzLEiWQOMaqmh8nFL12NC/vZ+7SHZSAjHKh4v+yTuICos
pMBPtxr0Nmh/uE21y0cGCrSlXlMhcjs0KxLZDWhRbhfifHo7IlpQ7ZcFTPVYVSpJbpp0s0gsdal4
hraf2g250HXwzrVqKOqLKjpthpzSCwcvbP+L93jAoOYbq8tuBZVZD9yKjuUkVsVQoKcTSbPly5tF
4uOhpDHDExzJNpSgF0LgCSO/7AQIDVevjov6JM2Pg1QasaVMIDqtyaHIVowWXne3vE4JTNrOoZHx
qFOw9AAdTjWALR3zwi4RIQCPR3nOg5jkvs9MaYb4Rwp8FdMzq7aytKNELZR1nJxzkRBkBdsKZktu
5mu06V4+nkSxpPxTa7fflLNEzw7dCQ+o0MzhmGX/xFrUlfmgR94NOt8smptHWiYTlt/WnRvwgTIL
oYClyWHDSNb5/UgPAkP/Dg9s9xoQEXSNph6Ks4+ddXNs0Uvq1a3OgpylSfWBIh0OSYbvHKPsob5/
LXQzHHp3KSnx/newQuWHX0d+5Vs/wMyKWdMxUlvDhwgTk8NcFBehH+EDcYCvwE6NNPeXmMvApvem
DCUsbm6reN6CYcTNMy+ZERc4mHAJxK9/OjtARty9dJ3txdbeH30/roasnf1Xv3iQvx0YqFrOYxaa
KLxS4hE6Ug4TTKdgvXcS2POs9eoDZp4le18nsW2LYH0IZcqYOGOFZ3SLsuLdhjJc2R6e2T1CHUoJ
kJ+gvTTRiG1tT9m/FtQcbvEMlO/syP7m5fsyeRhDF84BFWql1VCBS7QlmzlchL2ANAPcYe+nQWhx
wBl1hWS/r5RNYD40Go9ZL7o29IGw0nfD717DmPIlww1iR/BR4OTYax6CWx4zr3+gR/etTJv6Dk09
75KiPUadkbaK8qkpLP7P2B8K408rVzEkJGGHPBcugTJNYCk4wfe8coTZAyDkbg37Ie+++aWlUS/p
gRCtK9v5Jc5GSszy0FgmdJHPIZ/jCRF9gF8lE1IrFV/RjN7/JQrs5HNMTk9rTEs3VfzDXLqyWzGk
uQlq0OhsLq8qqGhS8AAaE9WVg7q0JMijL/QcLHEGVFomX7ARPW+nskmGNIkp/WAoE7uLAOd0sjoM
GcIBb6Iv0gQLtB7cm6F+n1eiOY+a5msp4PLPsG2cJxbmwOThyn9+Vk+nqGZq/EbFe05/EmPIoJDF
IOnmq5XESVkDllXhG3+yYnl0gBVRoItNSGTBm3W0V/Rd4IqAP0n/7DRq7yMnFUdLDHVcx6hFiFpd
4QjAdG2K3vIDX3ESEU4eqLHO4YVIi4TR5tge1s60W36deMfXp2hQGxjG4wKoMWgj5NxGEM2C4HUw
28a7PDwBx625YYgKdNwDLeJIF4r4zFO02rBWn8vIs7TJfv1VvP43KrtVXr6/DfxUbcYKO0APxMhj
q+IUxcPzdm53F1eu0iVswp8MQ7QYVi+Sd6GEut/tVJHEKHBhdwWyCcti4OkLBanwjnYMESJaQbv8
+4/SvsHIJEHEzQIpdpo1zEU1aXJXZPZvoegnS7dYb1nMG/eXwXCz0Arn1aBHLEuj+rzb8OX63MxD
ZI4Hdr5W4xzcPyXvl4bOje+cKx7utDV1dmWMDjDMekih/V8tvt9MI7/gZEmUK5BdodotG9ptupRa
20LHuBBXxLAq8Vhfk5IsgIZDXekZ3hA+sL+Mv3COy2XHExd6LHnN0q2YFZMA/N7Hqy9FvPozAJF5
smqmlnZf+B9m9sxiHKKU8kJHFkXwXEGgrDclHa/tYCjld7LoY44zQMa0vRLMziYFDOLSb1wPDsAi
9xSR/59+JjcVlrNao0UVCSx2ZKaJnc6EK1kRzuDVwZgGV9VOOBDcJq1fGJBSROCXd3BpLYc9XNsH
KIdKY//tJnBjouPKdKFJi0VLEuLu8QWcegpxhjaEJGxkeZ+U9hKOye43KzSzd51tmwv5CRYZLzqd
IBMJGMcchqUHz+kPS9U4f5qt+xuIdab17H/ROykHeWeTiDrWyJM+rvMq652dv7AjbKLhLx9+GqrB
bVlb3p0bkAnOKgTaJ8dOE4wHgSPva/NOycfKYgR0MwUpX943Y5Kg5vwPYzMtGj9UqbALgKfFEPSG
o6tOMRCOp5R49b1ByEfu+CGmtCLlC9sWWDk23lCR3h3b8JomRNHttKAiuTlueCGsVojk0MHJlb5p
HMgByuw4bjAVhbsGQDrLtzxMMeT04opvsZn7a16lVyHEI2KVuTLHFNZGWLUuhheV8QPYXvFDzK9V
uSfN6QY1LosqHcqZoqZIeCD53L62MHyr4pkGsTpcW4Te1VzrWLLaaoKTjj948RW09cyVVjQ1OGTh
61YbbA29N+LqNol/LpByqCy5RHGJ//zAa1Y1ZCEgcVDH82phdlA+3pDbsAFWn7gNP+TKczDcnmqs
EOjujYw3p+sbVyFFFYWLJAGMsvtNlSh8y5MUq8WU4AME/BlKOJv1ew1sPd5iSLoAc7Ubj8sAhk5O
fA821TDUb+Z/GouzPltrtpY8w6SxyYuXk4Lq0JDfBQEx22v1hteIndIYt9y24oRaWr/CFfimOYtA
ivOzWtC0GRz9yApVp6bdaePZ44/uH4PnXM10MSZ4YxjiC72TeBmG3RumHv/jhjjNzunhENVzOb3A
VjXOVVg2kTa4aY/EoWesax9ip7hK8Pn1MDbEkr+huilv/mgRzOpbonLg2FUJg6/I59P/Jqwzx1J0
kj9BnZd1hNag/KRYd5E0V5tEA6yMS0jYh22ifrxn2vfyNxa2eCHGdeEyWWENMhtAOlS7zavf1vVY
2S8AqkiTlZFUZVx+UeX2PRTucAkNa0U+UbJp1Eztc/jVQvarkWwhsODtLYlb3okW4Nq9b80jP8ol
UdlCGqG3pdFLKbj88y2on8OImdPDRjGZMC1SEXDtnruqoTQpUsWBLwfr+H5n/uJG6U2QTEafS6UZ
yh+NSQAxF4wDg8Rb0LjmXE1VcDchQHOqXppoeC/YjpnhpEndROjMvZ47kDkDCwMyh94NajUho3w9
Qt1lF2AXksLNkLns/eV39hEA9tCFZApP8xKX5eSeU4jI7aNkKROgGlEjATxZoOHdB+/uOlgrTe2G
H4SwN4yhGXRGZj+jkZMCPW+HxgudCeKW6fEz8QclN8xJgL939AXzH/u5/YQ05J1s3xjcaKK4m9Nc
lSKNs8WzrtJb050ue4slISkIvPK6aRQ0sgL/yrUhJ2/btNo8K2vyP4GMZfch1CU3G0JzrShTNDnH
NU1epdky6PxtPK/sJtsalqCKp8c0AbSoYv50V1cZ7+V1Yc6WNsyvNE8wQaV73LuGw5UPUnViJ3eq
bWhSOK4IUQk100rLLLzA41Azgnf1D5RNBu0UksHwaaywFI/S+ye/+nf/XUz0YgRYRtmMui5bCkSw
/rWbHq6oIEWgZjXq29rHa+3W0PhGQWmy30AldB+IYEn2tNQsPDSGcOlYAZ9syG1YTqf4ks03pHXK
i/+NhSHUGO4aQOVkFajGyxtnPcEPRpjD9Ox0ALdmtPUBZr41dLzKX92oXDV4HTpI1m1JypLmmEZK
RsLcn/wzy3qLmXaQVkhGDBMR7s2QY5L5XIrJxKSD+hPW9VqD8Ov8zbOlT9Y1qJCzp16vuMETh5zz
t/FxvsfA3lrovEqDd6I/eMraurVhWSX9H0HBRnRaTWU7l1/ojksdGAoutOEC8gNkuaH+Vr5RK973
agZzBh0kwMMvDt+f2NBi65PvLM4qojPPzKpwxwA+7pJpt7MzJJdXCx7zmwiNDS0FyQ/t7UnSPzSh
GnEaJaQhE7mQViAiwZ9dEHuGoWrC7PEX3vzpHTdxaJU/vPLHB3mvmbUSlxWJtq8I1aqUN18IJmSo
xSQMVF+8RCk+62WOY5oZC4hZprx2Tq8YvAO01g3bGITL7DjuvyKe6JxI2OTpWMI5qduMxl1/dod+
WDI0rjOHRZi+lhnR7sVt7I90l7U/5Ga/EWSEUl4yd0UB1t/kXt14IUAjqTwr3LmtUfTTjuUY4CLF
efrWzP8LdZKXE8UWh4ze4Zaxf8kmd47Z9VzU23f8qTXdxwcaAKG+XyI/x0UgOYqIW2OllUr8d2gY
GP7BjWsyFz9rqzMFLRy8lxoUvPUB6EqycDm042gDXFmOUtXtDdnrvZGM0Z8oxQ35qcCuDAyuqdX2
XX2vH8yhNCzkkx4uyUUBeDKpL7GxYiXEtI5FskiB7uePUFVB6gjgeYpZjsd7ZVm59Cr8N9M5KSoK
HuiUxo6qPYYe1acfvNvSGFYPWbFl/2q8tB2YMKTftSZYOd1DksC+LlyboJyrx58vRyFcwGLJm3En
prcJv5XsSuOvPa3i9V5pcEwSGjfWsXnVA4Gd3kNGTc62xtbA0tiYn43LTVlyxksJtIf4LsGrAeUy
14w2KMEFY0Cxul7+f/oMnBvSgLj8U70WyIb7nuq5qfP521eaAZHTJoZLGKR45gGWcHt+zt2706Nj
pxcELu00OVd6huHlhruffxUjqWuANz8Mffkdw8AnOSi35I9RjJ3W1FXdyG2CiEKDfSgpsce2ITix
zgukbyJUrthIcIKeUTHc4eugJ80CjuK77RgxuuR+IZUIBcbPTwhMzD3VQl7V1tX/f3LP+CpbT4yF
2qVVPCyddmptM1T/wlTmzJq9tD/DJaHs+ZJ/vhWkxW5agQMfLtHFpO0JeZtFYkZfdKpmAaFpXzBW
4bz0ZeJNydZ5n6h4OHYylezLHgFHqOU/fUIF2JZNFrf28quHB7I5gYv2ehTcKFUKxGzjetZHj630
9GIYpK5RjDNBeO37k8fwn6O8Y/xp6clHbQ4qIa3TpNBDWRd6Prt2qAucCBCzVjSn6EfztJIL/4b8
dL+WY/plxGGmJtUTgbwGNu9dwrHau/IWnbq+X/V/+eX+sR6urr5uOMiWoITS9iZpCUxgDSSEsUZR
wjjS4CMveLdg7qvzzY1rVA9MNlSg/mrrVIWwYGrsH34M8C65aTYsilvS1KKw7VEr5sO8QCmAknCE
37ucep8gYiyZzwjxEf+fEbANild3+1SgpZExVCSvUsg7MKiK4TVF+xcbTvS5X4I+TP0Sg1xiuBJ/
UWaN9TihJVjpb5J8F9RupszRb25V+T4zJ+cOTvLcols19qR2nzSbLpXGrRWMOfRHlA4hyvRxqT9O
jM5zZK8PRePJFVR+vO6Z+BEomV/5qbRQcBT25fg+RXDo7MLloIspuW0iSUMMSSHYbbbteENO1Ze8
JEM7fif1YHH37uBU5WsXiC7GFVtUhSX1TrH27hWCcHkFaQgUbHWDH4gWMlmxOAeNCYAT+EcN+x6i
VZRqYfYOwDUdOs/Ay/cqWCu+3kBEg4bL7AZaQKBnBJqU9JUdj0riaWdICq5Bokv+g6TNZXBEXMkg
UI8NNrZNvNHPyL/fjVXgfXLirtQ9+ITQxelWU89mV2ri+alL5mKPWTOIpzyhGe2CH4tJfSkARKo0
BUDZKSHoJTgM+F411H5CxQ4m8j/rVgkfvpvb926fo8K+wmqTMKhvzR2n9w4Iw8EscB0bT1GSuUnV
iKPXS4HLMs5Yohjdzc4N8w+d4k8a8c61MMv+dIpQu6M5e5QdqoxlmEg9x0KcPpr+2DkdHaWLS837
eR4mACoAVoolEOkT7Dvheq38uTg7hO6A3IvBSTUmdnUxyoSYeneBjAxAjp39A2lxjnjbIj98EIsy
rEHuoAGuQpcr+4yIT+ytOuOLPVdYDI/m8+E6oj9b9fOjPoDo5oq71ZvGyiSjrywEbiym2KudF20C
/ZzelMpD/N9A6CML1yn8LkgDnYYtGLTTHD1A5U9GNNPlIi1Vt7jdIn5tuh7z1CfMdDw7t6SUnpk8
V9AxtKXiOpQN64Y6HT10GxSrrpZtIcwIh195N2d/aqR88BV/pRAE15oGJILryl0ac/Rw3f70XH0r
ihaTlf8/mijWYEw7z0B/eSBDWRTznRIJMPz8WQQZs7Z+HWBDyV1WjUWb/jFzj/hJeN86m/AqgfLZ
vdU+dvM0M3AdqopYY/W0gtZwhLvRokLeyqhPAdtn//Y7DSkiKRCavILtcAUGa86aMK7y54N68hPu
V/UGXpJIgI0XGwhl+4sgqqGRraexbcBTL905fi/WOr3EcF/eUYPoOiSYljzKeY8tGiwsnsymp6Sp
8lX5Pj0oD44KUkjrrAD3pFalUlfHokbiRunKt7MQP38jnZhP2LictoaKJTTDBfL22wY/kIW+e0JO
N2RhAx5o6esMJxXIXydKvtFk5RMafFmSl9hNqxX4DU3Uw4DmN9bRnweQ1fgVlJ/qs0eAvisTs+AJ
WWDDRL8SmO2ebWNRvYqQnnq7zxzYsPwAQy4ENoCGNDA9lWa6ljhGH0ra4Ef7Zpm8DkGMUk/lv1rc
qvqfYpgAGCm1iaxnp4+TBEnIYvOedGBjMHVlmsRBKadezem+2gMBovi8JoNjZqRrI70F9neEM6zq
PKzHlfLv/ZmbLLgY+NrvH0+IHGC5b2T3FkCm9SJ+Tn0EOQvuWaQ54s5b0PDvb0wzpFqeOfXY6rAB
7XIP2brN/L4W0iq+TXukM6aOh7x66XoPp9wqFY5ehZRfCLDqqIW1Q4knvFdV54/NK2D1AeRLnQyc
UYTCnNYfJR3ugGXT0SXRhDzMzZ2kB1SktGKXq3rE0u9hw18ln4RHFf291TIVA13unKwVEwhJfwO7
/i32cMtvaru0hemYmHSgZyKDnWYcheY2hMBFa6qIJkz4m3zm4gKFXBM0JU00WYTp9AqUG8XijgRt
FiZ1iijpsc7VE8MCT05HKZ9RoU/F5UGQU9uN7Vc/wKuoJdQmKVIkyWh37GtoYh9shc2wAvBTu/mM
ZitGsMdKIcp9UTKyEI/INUPT2XNvpKkW9j38VMzsFzNA7Gg8JEX07gpby3j75w+oMgJSGq+EjgPR
O/WXCF1vpNdzP2Y/KlQyYQtCEiYn00493hS8VX8MFwwIpwsHTn28APNFZEpdAAlL6UvPtHVVIWUV
6VZWDGYE3yu3XUi+BZ9Jwot1I084MO+NhENskAZN+mxCftkrYh4HJyhwzioafuhVe7m0GTZRi3dW
qAeJZHNgme0/aTzQ4VDK3qOycWv3WOH+FsLt7xeT3vUUtkxEBuvcFmQZURcvGxffgiPXfXnPZJif
SbtvOYvoL+32GtWQ4MnyVA1b7PylB6q4PQR3PXhgZDIZGoNXo1JDom9x/f/M2dqzC45+WozWQ63v
QuI1aBUshgQhmSIWjO9VDpkQkr3IhvrZ1FGcF0Aggc93B97r0xsRvOcxRd7KFxQezoYYo0jZA851
CRo9yeTOszvkv8Jr06GXRXUBodzYY8MTgZgxgbq3R1zxMrOCh5yRjBFE5GZ5nxCwI9fW6uiM5e1P
4OFQo7AKfpCC1MQe6lT/rIhVfkKWE+s7IClYAch/+y2AcoZl0762+jxCvkSgjB79djcSD1DaRNzE
4vQijB34H5bBbuUBlhylKrWKYQShKVmMB2xVSKRhhP/YpME9dL6M0lNAlEqLbV5pX+RJxjTisYLP
054Cpek95ZpBuRwfGBVK9ONYhIaWkFNmfGxWREaa3FcXYkRQrxoq+QR2kRivetmQamZlJ4aFxHBF
daTaGHa2Wwat4sfaaeAsAIifJAlB7Czvs2olOJeeYitkkqNdmiLIyqIL+NzfJGFR7045OudWEaIT
yL9DTp92mdiXaIGxSyKS68g3cahSLqrZq9I0mAC5HU81rQcPdk+7GNQ0ceZzDR8g6O3Z+znUC/Nr
+bjrXFK2NZo8mi/bLBFygAnoC1zhUBSn2y6UZK85R0U9sKjWXm1DbujR5IMTIDADPoJkp1lal/AL
9j6whz9whlOPNwTNJOFxf4lf7VN5T1IRqOSRfTvrt3l0TOSpPuwDrgmmFhMDEQHn3LYjTlhsCccX
hVtjAvxkTQrG/LJHRjWEAmQQoUwKrjFRDOhl+udcQ8qd+Hd00DMUWtLyGGpahkPxwePQifG1QAa7
4KBaiDNWWRBFJlBkvPs18gPGN8I3HkJ+NERkWvDwFn5ymBjlycnmlcY2wTkZJ4vmOBtj1hZ7qowT
RrSKtQyKZcIJ/WLUC0uTomyl3o2dozvQDquKEe+uXVtYRM9RKN3Jpse+nCh/VW8GtBFpCt4Zyzyv
UF4WNcF2j61xwZUHeFq8rvnxXJjR3g/5cWQPgCT2z36hTExu3vNekKuIEYG6WpZNx6D0Zt1k5oeN
Mo8CbQ4y0j+65nt7KlYlHVhks4wcOaIAqUV83mvDZZW6Z5+9RGG5zl194thssF5ghUbKC+D9+E4J
vSk6leQCcVrianKgK5o5NFddwDnLkMONYYREa9hW+uAgxSFe0lDKlXaarz68E8kxWrfRPSfYM9Ov
XLbRKVba23MgN1k6Kup1Ver8UrV6DThySLSigmRKZ46FqIui5VjPj1J1r6vhd0j06lgBslUnhpNY
qXf3LRuU0VI/Qx1Hb1x/JvEE+MBwKuEmQdyUsA+1CCRDQRyChwg44zBguqF9vWqo2MdxapijQcLw
tpRwMSzLpSWiHdJf/p8MeWC9CiOVotLcRiaE5TtEzvy5c9jEyWPQyq4KUqTkV0fLAB+3JL4iJsj5
5pOGWpxQqVIw2OXUr7IDdH0Y8x9Ez64d2B2sahY78D773D+WUanV22dlzQW4HU+ClPhzO8LrIstW
QGtx8MIrZnLX6IiRrf4a6DU7tJg78MTmtFrunpe1A2cTFGYbAAiozCgCelNj1TVuWcORL9WlkUBK
oCJfoMBTHdy8cKttkxiAyuGyh5mW3/0vt5MjEhcaQnhkypiTabuy00ly7Hg1HJ+8BDm3AW+lcW7q
DM1EAYgaMtt+6yV7VQLY0L3YykhttCHWBnsgoe3r64J31qCOp/F86WL3Zb3gxtEJDAgfy5EDAaKO
VmXISZko29Hk0H5XG8fttiSR59iEHt+621GcVY4kRWY6rV/q7wNQDZQcKvOMGs5HEpMMRy7nlvKu
1U69AT6MW/DchpbctmCaGuw931j5bP9RIqACwxVmJagSIHddLGuZngrD+v1yO77LCi3ejT8kEc2l
ZYCReGALtylnnHOtAuFtwBdvRytq6BNfQoS0u8QaOoLjITXDY8Yc6SavOMMmf136ickeAA4T3wGN
vK0BYiV9eikV56+Jsu2+wJDvv9/0lSRQ7LSFnMSGOMmnZFhxmoc5jbSfZKuYwGKH8kKfl92s9ZFy
luN7b9kMGp2ZK0gZbjjDAN7c8mwqMVeNy6pKfrboB7V9rXd1nw75zRSSIge3vmNKOv2ZH6aBmY7X
GdBYNTqf/QQbMpxX9Iscj44qtkiG8BZm2BexiXzTrF6KBCaHpsIDRSRp1HxESliJMR0bRdtggf8u
xC6+1ETpzrom5J6u8t1mjRjnNwraU/br7hn92s3qJkL4kGWQ6aydHE3cDVh0uQYjVdzUIgjFFz5W
1cP95PJ8eaCsmGAnKc4MTXSFnnJnlTXHuI0MRtF4MhWlHiWNO7vdt5iTw6oIc429GsFd45e7nAMG
N+aSlDGwXYV/xxQVVd1X3wJpa7Vn9D6T9TdKTfRuPD+MgwpgsZgrKcCBZaEk+idlWVVAmIgTTn8d
nGsX3SYj57YUYTkb4/ufdwsvtz+YV22GXmvWsKX+gwaTYGkPIw0XNDu1D+HcI/KNJ0I7J+9iMQWJ
JvkpObhvHCCE6rGotgIe3A30HDeQOXHdl04KKNzkNy993F2p/zqn4VVgpFAmjYwNar3Gz0cL0QFR
ZHVvxGmUPDjCh1MDc6WhgPSs4mm/TRtApY/Hghvc0TZmEtY1JlOuQ5/l81NeMpyLN3BTdHruxKsE
ev3sL7zwnsYrFGJzCwUNLlboLNh6kQmv+Ex/hAHaXbAatZgNt2Prj+yDMTQU+t5cT+uNk/+J003Z
OdKEd+IHgrLib+O6ZgD1/MUXo1O5icjs4fCurnqJmMOqVqYx3PgSylXne1QyG3XpbH0UEMwpqan+
nZm8IT49Dp6IhmFtZj6mScRYhtU54SRxaLaLs0Fj07lkhqBIAVWN0vD3MbHwZDe3VddgppSC8C6C
8/nlAt5JJ0hLddcrcxO7z7rLVfWgsMQTCtqX/mUgSqJIysQGw+mRnkNDgIb6jy1LQnE0n2Oy2ZvB
YLVGAh7oDHsPGfHTG4ONpKjmZp2orlPEQgtA0tRWpN8FkHa6YETDijL5WeqlmN7ny3DI0nXTM8Ve
/H3Sz253a8uqVhiRy9tNi3MRyqZ37W23Dxed3sM2jiDu5cHBl9KfGAV3YvhlgFZBNAq/ey/qsDVL
xxJLAIc4SDh7i+qd5jtqGeOJT6/aExWfI7Yyb3VKK/4sN31TFxMpqm+cHH+tPlQ1d13uNDH1725q
9BJOt4ufU8wBUHr9fXWgWCEaL7NuxBMcAz714AszXFXPU8RsmYDahHHGJC+BB2gSYrHkqU8XBGbY
o+OwnGkRS5ZIYu3bY2S6W66GvKXPhvsY67OQeP9xrmUt4fHBXa7+86hpPA5vi+4HebePT+7Ai+AB
aPoPcfoDz9DuWGfgJWXKeSjWrPd79mLr32h2AyxqfurqVo3Tt6Ox1hGgfkAmXBdcPKmMYK4cY9/X
Em5LNF+Z06ACNUi6XG7bElxnzwBTOBcyYAE0TA0Ez/XSS+B6wp9GMhwPicWhcOjN16QUhAPkHQ9H
cwQkCmxfWOww8uJlUU7vuIkFvCPHsXxNcvCRIVcsl9e+8lbpBlLzMpN5dhQnCCz3kN6pUvZ8oqxB
PCOLmTQcObHIr1XjWz3Wa5W/XacXqKDlKaRUmwNpERn2DCp272Em4Gu7KmALZo94EwozBMfw0Ilp
cp967u72fbuWzJl/Ztb+gMgISXH3n/XpCiJNV8Q7N64GoFBhv9onJwRkpT970Z0bEgZrfPSuszyU
voFTkUqOhlievxfe7aW+JuOOdBUW1tHCKOjn6bqfQIlFBckPO9AX9jeEZ2GWmLLgTuP8/ZxDzErV
o2klW8+FhukVbfp91b+K90icqmFxCKhBuBT67KstY3yInXf28PfsCTN1kjk/Ph0SdT/EMbt/59PA
xnq1hJf4oVwcw8UutC73K2NCjMtqo0qqxkONgwpL60oxchMrfGmMAp4wUcuYzElen1MpXJuHVC5L
AsKTS6B0z+Ap/1qIRophuzX0kWdYLgbpa4rZtr6g29LzZiXCZkoL0TVODrW6kIe+WyJl2btUQJ5O
xFUydUwMPQSHM5C3FQ2uRmFQJd+aSwK9gPMgrsEMw/jkIKTmHzDqswQQ8vzHZafz+hEyeWMhQJDb
nE6OWCa3zvvdlSIIBWvaFYkMeDMXDDdGDZpqW1lt5oQqL8imqRyseuVE/p+akICdl7eYliKctN+a
aDBNTPRm/7/ISvyvXQGVfkTKT+kQuo2HyCyNppKtEsQsMXedsRxQVTwlEsUfd6ZZa98x7kPg8VOp
lSJ3wSlyl7oe/ADjA/ZQbK9GHhmoYS9Cue/5zXKyBktYL3md4py2a6MzxC2GY/saT+99KOfvK/z/
NpVnQXq+3Hp3fw4dJKSzo9maC9dTXENlwwGbFwNbw5geoStRx1neq9EiDDD0PQv+t44aXrDO3ygS
/ju7wtfnh9IoKZ0JQ0dB/zUpuVbN8BULYBw1GvJUKJuw51OMgUFx1GgYROtDHBt7F6RvOGSBFYET
Sxh372JPf6YCVBMrT2PDgu9R4jZznXRaohuDdX5JKqQMP5bS+bcAL1sLE/3i1deQtgQC7v85bvjW
bElNdboQ6YeJkicxX5JHnsKFMx3e826aoGBqt5+FWghwm/kZgCZMz2cBM1mbTiDQd1LIANO3I5/F
+ZSHkZyXVB9piMk8Gt68zpXOHkAGHSpoQRTriTT2uSkqr/giLrozcZYlOGL+37wyBNpn+U6lbNSR
zkETRX+33pVivZCbu2rzAwLkBsJolpjCz/lmrBXnfruvPop2ovUAYN27j/EYwJGRFzSd9FIR9Uv6
CvR76YJerdvRsmfkqMfRcfS7PgQAL8reIEYQ8zS+V06zeAMvhzXrvArrgiH4CwuVeL3diY4TprBm
0prd4ucvL5mq4CXQUlb1UJn8PJRfYbY6+S8YXbiyGx22ug7kTgh7ALfbqDLmLhZ1NRi46Sx5/1Hy
vLqMrWmPZym29gfr2JvWUaiEV3fvHsD7fdU3qG4wjvR71oc9wdBT11eT70D7NvDpmc5Lv5e7ExA7
O18gLnU6X3FFv6EXFYtl0dIRowW4OG0VT9cyPiyNb6SmVNQZUsWzlSb54dOPPvEyIloIjW6EXtR8
32iz5N8WwhQIQ7zexWim0LnSCd/dCcZPYYxOszNvOpTrtGnQuUddtLog6nblFiki1lWzMQpRDkiv
F0yOHy3l3EjnCkOqL5aQsgc6qzqacFqJ7Mc8t/VsXZmTViUkZWWKwAcwcbOUiDowFKuFuhkO2GvD
Z9PWNJTEZrZq6voTpbts8RxsHEZzjpkc9sRmAtIqSTkE3CEjhczlCcCgXxEl92q8u1kyjft33O5T
9GwNxGoE6x8rOCYyJJDVF1CIBKqMrA6ejruwfrm7nUkUYAWnq3ZDKrOyPN/Trn0yNlXEEQ+1kjRb
zvT/LamJYmX/PqwuFQl7w3iu4OvQSTvB9xvsJVDOSX45Esuv0gdX2I7CjNeErhnFdYiSj1ij4ba9
o/m1Tl1pjhVC1BhfJAVPDy3lQBsxkrpaExR2EPng1RH8dlTCQcseoz5moGfu+U8YtNfpLL1xGiI6
51+uVHU82I0OuvHgCr287c6qEa8SEenxEflYrzCk1B7SFWwfVgtlOnTkB/sdVLYesNTSwDeSsgpX
BQtnFSz0WrGNRkY2XmT7z8qHTN9AxW3Lab8OSkyFKYM8qz7pc1ZufY3t8imoMFI+AeIYvybdrdYP
iOkdBcX7SDAy4ehdhV5qs2vIDe1wCVElrSff48YJG8aKZRy32vEL4yop3nzLDxjaJ63NObQTluU3
pmQX3EJtTsWV0K4SM8lI0cNe221WtClPePXGMu3Syo+zsj8m155ah1NzmtxTBg6i7QD2N/zlfttR
mM9JBNRo5ihzPSn8PKpIb1ZSVWQaRs+uoImcWgJjO6xpP5hMjaB03j9+Yc2xV/tgh6y9Iq9WrCjs
lMzy7kXja4hE6spA9CxbXpckx3i3KFaXpk2n1aEbYHljcUfKupknGdCTT6OLhWTFXEdwcPwXcJ5M
PxYV7pCzPwwBB4MsQ/fuhyIINmlubMqvOFAcXuu4BinAKfFUkGCy9n0EHcn5DGz3A5eRoVL1QxT2
bz7sf6kRsxfeOKUZImT0WCuHwHER85KaW1EQ2N9U7YRnA4OsepVIduO2bheiuXCVUrRIWNdmlNfZ
0eOthmX/eBlNuCv4WqPP8uhZu/2htgV4kYfUPwqrUM9UITHPZvkA6BapM9nxNggTwfXY3A7780tI
otUnAniM3WqSmA8xVSatvMvg/VKX1yvditUrPM1h29SO1f/8J7R7Th59PTodL9buk3XcWyYI5crq
P5maP9lRsQvYmcxGUOMfKHUR9Wr0TyTP55ZpRiZcOHzl/zkv6PneW65zbWWa7sHw+Z2qy+EEtxib
gJshE12s95OJYTuZ2w32UBLyGMq54GboaiOu1m1YMRw1O4BhS+j9yzkJXlDV5o2+CGxwINhyFENl
hL8a63wbtsyPD4H3qygFnQ6sRLtwq9I9UiysWU88f0MFwX9r4DfxYTKtsfeRIuaOH7It0P6c+hcq
8VWhc+l2c4A4yN5RnHk53wUIQ69AuMFqgs2u79ebuQWyR2FwQBbprMof3rBkrVgYQYuB6uxGjGye
zro19jafzN2V73H6L5R0vCrmEk2p3YHJJBLpeApEYFR+gXSfMIHPDH4gfF02uLmzaxu0oOAm1ic2
Pv4hrD4/gM/fTVfE7LmUU2iPz7JDlApzc679Qi6ssK8ENaUW3efXFwrL5W8Qappxtl31e0oad2/T
cU5pan7KTwriTFmrmcN6sKL1awMIeXD21YwnmmsbQEwSEG0dBWZLhBkz+NI0giqPVg9MS+2avRYb
+Gej0EuaD2yFsATvAwCUd2Ps4kR6845cUUeSSNDRsdLgB0h2ir6pSHbopVMgb/3pJHltBUdc88TD
F6AF3zZ6E5ULv3AoZYAAIb8/C8qU0Y5/xVxG6puyJxoSYhVx9Kw2cjt3kMp+/yj1ueQxTSinzkq8
WuvNTCcl/YQFY2Y7GgueL2WKvnHoWHzzmY7ftUfX3chKJd/E+mqr3yhE3YLpsIsHW9cbYRAnUl91
yBhdQZuhVCvEJIjG5m++j4TZcSDIwOTQOt1HxSFoio7alqF715/W8NLFEWl7jrSRL/i+m6mL0zQz
1hhpAhV9gJGjaqM+IGqz+HdEereGhW9ck+/ipd+VscnIy2PD1gGlepIAEk0Bg8GB7JCnRYNuA8gm
sA743YNfdALW5F1m1WBkvTtHAwD1AmdMEAWf+pR+imnF4UuoF2k5sEsjFBX++Mn4tPBS6GCm7X8G
OJL6xVkcVIY89ZTL2Ljbfd7L3LcWevxMK+M5ac9KSR9WTEerLu6lsoJrheR9wpxMR6kqUblkONgN
PRETQQV+OnsSqa6OtvOCN6khiZe070sJI1FgO9M6LuX4qwjuYzSZZy8b1ZUwvPhGbepPkq36KBFh
WyAzUmusOp6ko5DqlfHH94Un8pPqzWG92r3ggTkyLenIK+/o0/yewKUYC/UFkq7ELIsqY4Z8k8LU
msbaVrt2p1kW789pNkPEHfasqcjMVPymM26FHlZsdSJl0k9dsYAzTZLVQiwgknaabA+ccJodq4Dg
Xk17QEbgWKzWmBeIUGKR+jIqKIpU6LVQqv5P5cpDgvHIqv8eUjdm+ndxhYu3MPTXCk3JDhOIyUyE
jy8WAfaXG8z4UJSTd7LQzglwy15M2S/oLH58QbvXT4x+AcH5NSAf5qNrCkqOmw+kYO8DX+6Z7fWP
5tleYy7ir/UHl13BYx2drJvbtcp412CSZiuik/gQhH6RxoZbsBSHloo35LPGLd6nbdhf2J857kMJ
1kBBsV/a/w+q2Ytpa2Z2/8wFzv5nQLF03AsP7gNlciHL3fplThUFn5jdAYq+IQe1o09driGV7KEJ
MDE3WXojuQWb8kLoIYGFO3EhAIlE0QsW+oo0tCemwaGCkr5nXmkMfD9o0Bnx/CtgmITv73LhNpil
fFGPu6iQ74JmCUJaguqWi7iav43XhOqtmxi0d6qDTnLjBAGEV3fc/DiwhZTayCkc62QIqpyP+teO
bos02pYqu8yPKfIAy7rU6nNW94DBYYV7H15uTcRcOuzPfcX3/si+Q2S+p4JINhkNS6Y0C3YS5DHe
VYJUsX42CWTZOsuIRExtBRWtiMC/rh/kqX8VsatTdn+ReOxbgzXUvkQknJIBbgRkD9fA7SbxvXM0
iTGmhRyjjQbV4oVmf5y4szDOcJMABzMcxcTEFan0+MGyxXBhu+aI4IgET/xfSoPB8OYHgvLLIyjF
S54QBYDRMEyQkqBuf8PMAoeRLQOXDsCAmWNVA2xNi1CpgmgeYCLpCLzS49z7seTOGtn1aKj8Jy6v
cHoSboS3UTSQKhBTOuRSSQkI3hC6c/8aMTw9LtNms9AqKePF13QW0B88jUH5U8n9jNHpbxiYWYg2
2bbBZyZZ+TIS757m9/omEk1rC1qXnF0nqZIiCSRGoi2L4MLcaQhN1akp1PzJxWSVd/VIylmBpDPe
fhl9cZ9hFZBUebQMoOGL8RgUm86bViHmGbw4w15BulXQlSbHWs1j/laj0HVYR6xLh6UjfCEnpOS0
3NxyPwj9m61DP9ACkmnoX2Z5Tbbfk9xMXyIpfutjMXl+l3YQvYTL7G/uI71HJktJyI5Qd18glmzN
JkGCYCi5zToOqBGDNZtTA9n8N5qU9xB+kjmLyIGbtKXybG5hjftBUDCiqu24KNDfuxUQUMGMLTSn
4nWKgo5ioD1XfbuSwxrCMMMNUuO/VOKAQ07jW0TfBJjY91wc+FaAu5OnBy2mcSSfA37thgw0lggo
84g6cWKzAMxeJnEE0E9zMaRzVZgT98eWf/Zw/OFJKu1N6s9g7mXoDtHXRMIyS0c07dPJpUZvx9/u
MI55H5sRSCpKMDNrGGkClmLJYugpuHDqFHSOa0/eSkcWuDdbja3FnkiGngKi8kix/pg7ag0R5XTO
yPrh/QXAyIl4neHfLd4BNNsuMZB4tlwCrRzo4d+K4F0H6oPAjvsTHoavmVR0MiGpryKgQqGmtFSp
42d3YP3KqPNEFPu94ED67PLCAhxkdOr3hihgzemWppeRIBRMlnrN4ebzQPyTaS9uHIiSoy5KiVPz
o2OBdJFEuEQtbXyUKsf7yJVc517arqTK8q0C3SXR7A6ZHxiDlw904Q0yXSTBotxoA92pGGyRYetm
vI6EFzapLvvDJfqhjuGNHeVWwWRvo3hME1RVJPx3FfpxCTSO7yeuf+Xv8EMIkcIwOIMkz7zrpwH3
079roeETe6fZcV0TY5T4uIcZaoY1XiTYaNxBOS/v8X+zl0sih35fbICK5gsN+uExz32X7hnvqD2V
fMPinNqqxPebid3f9VF5c0yDrHdabbf9Gsg3wzTHTMsji1GsbV2rXCIy2mV8DlMgsHBCq844ErBn
pXByFCi/3ObMJqJ6sSeuyjGgMo93Ct+Yq2Da2rLLiRAM3UzRP73VtTpWQhH8kHoTvfS7OZij3G2v
QnUrUud8WqYb+RHse7itSieFPylPUuXJQkU+j7tOoD2N6Md3g87MjqtrGzG0mPYyxgzhX4Rk4ZsQ
WPwyPz93tGA6JezWNUZbf5VdYetUYkWxnI20Y6ZdrC9VCN2WO6E9wwdW3lRZFAwm4hv8/W7POFZo
x3jW8hGBTgO/gTYJKlnzX7qB2fvb46eqYh27QE8OQWwDRaNM71SIuzEyVXXsY28X5CKMiJHOHcB5
F22OQuuV96yb6DmPJKGYqJkmZDQRhA245luH5nNCBbmVE3BvmoIEKioUK4oF1+98J4INRNzusHvZ
LD3e5I25Cg6mTzrezZJQnBxivezC0dvmgnEVRafVfLsum0rMEDVft4p/IPiRXa8cTjjfRokOYr0Q
444enbm2EXSuyn60GsjuvfPtj4TZBlC61W/iQObr1fUaoqOaEebpS84Gr/Nj9gQdDnP+6QJkUEyR
O2aMelPwvz2cHp3WHzDOx1yhqj2sEfBaMgTAnIln2a8qnJ4a6RVrwmta0ZOJ9h1ut29p9ztP3Roi
tX8k1Lh7dkWFbpxK/AFM3aHq27n7mwMbKTFiDTaLr8xckkH/xJKVA/Xx1/NDni4aT8ICfQ9s7Y2F
41iFvQWEbwFjCtEyEgo+bphlfWWdkLD2wuPNdm+XVUl/piBfJJtujMJ5WW6GnsOmt4OC3rX35L/D
ctwtCoc2Z2eFXmQkDXk1l4Rz/pWrIn9l+MCl6ejoQR6u/3fj16qKIZlLwhMEacbyKOpOmViQUrsb
OfVGJrYZMtxPg/jlB/SETvisuz7n3UM2nc2dP0RpL5jE4PGMAJdHZl2xi0SC7BExFhgnooYnE+2D
9v5Fhx3mKY2Tyhj+Z+hHiRcBU6hVN7khkjAJVQyie3N/joH0I0pArbz8H3ycrvol5FQ7DVaneFRi
lrI4WHQc2GnuEn7SHBA6spD+4qK1PP9Bxn+YEiO1GlvqFcQ0LKtLwqmJL47svDyoWzr+eZWotaOg
fSSBQklpcsxCBq3R8b2yA4XY7KAxGmi4EWsGYnDxWiQirfZtH5s99yYHYiGxHfqvmECnO+/dIN8H
ELqNdK+eZMrxrvINdRfhSS3Z1RQLxFjQ5ziQjj1nQRaxnSIxo7gXCOHBkp3ahqj66RFwQVG22Prb
SbyYjxZ/S55oa9VCN9azeQ/JlE4rVBjrYFxOzxx/Ko0Q31FkSUXnesQCppTZNu9gX9zJWxM2v1p0
0hj2/4tB1yHHI4/Fsm1Dq5AQ+uINkCc6U6Td8jfhjXauYUGsQweuw95tXM5I60hIRb3QWo7joHNr
uPnazmAVb83MF8YPngk0ZeMtcqt+HKNO3Hyl1dRspJMe76WW4gm3K1Q3wjcBX4V3sm++f+7xQ83I
GtlU3/cXLfEniFD+23+K72EPEgOXY4z08nNcsoQhjrRrVEvOS3tcQ/huQsSFBcnvAAGXmW42Cff9
LLjKE3UXtEu7ry5ShRoDlNt1uoK36hWOWYuFLim220LiEuStd3+9mZ8jAuvimBB0DSGb6oqJ9Ep4
/7KMqV5h+VKqi+JndXAXW08GYghSKwxL7ibiFPQA7kHSpiYesaxaR2Q228RsH8lZvbtSRYywZDw7
h4daFrHzbx5pmI1uA/FS/YZNiYHEZiINPdYAKb8j2Eexb8sySGbGSHz3Cs6binZcnbKiyS5qJZc5
FDpaaOWDf2pBJ32P8MwsGZUhY+v9cDVS3K7j/11q9cZUxP57xjrUKHu5w0ZenmZBLwXIrV3E5wHY
ShmLLCRjaliBQ+H4SiZTMa7YT/QBACzP1V8aL92zI+XsW9865G/16yla9stczQSuXSzNjtRwGxFj
reKsDOxmiPVjoA1CDcfq4gp3gS+CYU+To2TWsTmMCWaAYxLprxrMm8lZICnxMCX28t85Ej5hZLcW
ZED5X09/BfXkGpAMQGqegOgiXZOmuhXgW/HBjDeGD70Bkz18I/5QQuFJj3hzOT6ZJMzu5xzEHENf
QexPcX+lorxqyK2TgfAV+fuNhpeki+uRQGl1jvrR8G5wG2w/3Hqk1c+GQVN3ygXalDPrx0jKfMhZ
MB8/WMkYyCxNlmP5KujIR3GMfk1MnyoTcJez52rh8qo9J8LLY6DovbqudG+wmd/SmB3FLcIF3Yo7
7pEa5YyVimVYBUfwMIsqRgNnyu7IoGx1nOnLet3rGYDZNOapngcbmy3AsVBRdfuBaBPiq17hZIH7
WUYXCh5DEdUIyKxUYioj2XM1FhKYoe2sJutKK9+DRqnykaBoo7dYQeXDhcRno3U9QnpStdGpwahF
T9wJFWzIpQOAEC1vK2sJdVoAHi+zUvtrRMiOw6o584m0vc1V+SeGKQYFCz6pWu/eocDL4pUiZrHl
abStY/DLjR1PF0ur8HUTjR/ZXfp2t0jZWmW298rOmcBLFy3TbpFBAvQjYGp+YSrBy5OQyRLjRpmg
r25bDBq4TbDL9x8xJL/4uOWo4o6kUPVMpkQbPYvCcq4rBz59WIXQ8dlTKKZRBm5Nx7A6SsAT2u1N
2fEW5AtvoYve8lswBDMYobHN/MPSgkAYDMpTKAWXY5T25+Ym4aqnRX8TMzw2jIifqPz6NMUTvxA/
zkyLG2zfR56AUp7KAcbpv/e3atZafC+4E+vMhZwVWgv5YwIQS6Jt1YbUNxoqt6QTszcz5dHKntor
lb2JfU/oNrPDU46bmRqZX4kq4fn22oK1lVI7CTJMQGaQKot47JT/JWKRYdlzu863z1rGEovYhkSs
bSHl7ZxN2SWtW+ntpssEGn3WohTVzpHzFkICiWixmF4hZZzVuSSORy4UtEvOW+EkTTiYiH8OIihW
vK05r1YDnVhvndiEhwr91BbwnFcF/PZB93AYMj4IYv6daTXC8NezqbKN3JC1u6J960q2ElvjVbph
4zrC4DUQAkGLmcQYrerM7trktVzUC57n27X2uW9DDAxCK89gyNKGPhdC7kxNn2Dk1qT0/i5ua0S5
/meh9q0RGqcF47cfPIUULW+FbRfuq+zxknLEOY4kEPRy6zuZFfertKpHrIT5AN0g4Q1cyzybXmkX
WQJQtzj5Qls6qZJw5hNNzkqqsicGUjtiUnA6MSFM9Ik1nRB9yzOrOttNvd+e8cjyt9/OKl7Ja8zz
xWqWtEvhvquQrOtTuyhrr9SOVNJqwNoPdGiyM1kQIk/dGZuU18j3wM2qtoHr9790gLftl6c8ZekO
Y1tAqpzUqsvV51fK6LKBgPzA1hNnDheGOuafieKdvgYdM78PMb5RZjvKY3EMpUE2I48dh9X2b3iC
tytKkOs4bg8h754DuY9YOngVUbBPdd1BMtLTT3qnHG+qUlxc5Eu8UpAIJKFjy9f8yAM+aoj4aCRC
8u/9xjrNsm5idDeCl8Y8IRkuo+CPqeRljA3kM/0adBAes74IS9T2t8cguQjRpKqfbncrfLRJjdD0
I8gu0vi0CKk2S/bpUGtYinB4hUT5Lm86a+u/DI89GFT7OFFYhGD695Rna+vh+NdJmE7A7l+O+WlI
SMD6yPsHADL9d1NTG6E/6kia3y4GeMqEKgLrUB4E2LpEWGJKyTiitL/F3vobbkGn7HpiZKHZYZ4E
W/cf0p9jFA==
`protect end_protected

