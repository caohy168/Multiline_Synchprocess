

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qyGsKXGf8tZLZ8MO/6NvK8t4R2uGW1SzmyF5tsX5CkXu0PSTBR9S/8/YKPbPyrujE/YTTc88Jf+O
eCpAsF0s0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SRiT9yJC5Uqpf7Myl6ffuoicyiy9OzLI7R2FKBd99DYnc/Ou/e6lORSzOmY3C18qI4YziTtHq0mG
9/kIiomSQZ3NJakbc4u/KKTf4sdd6wdIZ/mvgBltW+Q8Ap0+qgKaXNTzfHyJ2n7Ooz/Tn18T9nO5
QHjNL4UKVvlJ7EstP8k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0eEt2iDjsC9yJcLMh6QKornt3Qp9ep1c6xk+HK6mgFR5fi2UuV3P98/17Y8KyM03HpNkVLTMYss2
6Z1aPy67AzTy6N45W245PgeUG7yY+SedSieqIS0fIFxpZHOlQKRcnMJOLb1yLAb9v+eDvlWE0Bqt
DC6o+3ydVuNn1j9muuqkFFLx2pd7RIg2vU0FWhnTxY52dz4f6uUU2BhdZBrGtu+Cau9ea4vNs1fy
I/3T7fa71g9NdE+G2SXKnMppSb5dRZUuux8lx1aIs0mR64PH9XFHoeK1TPXj3zaE/Opgcz+NH9Sh
oyzibQaDQnD+c++ig6aTpqrU7EjJGQp/bZ1sqQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tf5mZezeOm+OIDtFXnbJOyEHGJlj2ZccsmnwTXc9Lf5eECAxNh05jBGLjHm14homsVnylEfeIkd0
FTR/x2Fa7arDaFRVeIpD76PsHPM4sIgsLzVKZSuDFI9mLQoEjwJzufLxVI1VLrwnnCVNXdnORJhm
IWzM4TmfF+Hx5JOlhkp6LgPD2qnWcpe7woFrqWuJiGRQIuUo4INaMhrQXXkoU+AIRMn8SYGlfbfM
BW1POo7+U3nnN5rZBheCXwp4IIczrHnxpJVCU4U/PKMVsPZpyo6Amt4Ih+tk7bJg6dcOiu0v5cfP
eNQSvIUysD3zNnoO2TasUMvjH92vgoaXcHg4cA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nQvzAt+9jXefqG/QM1RphU5FHai7OeU5Tn31wlHRRHVBwRxy/exmgCmhhWzEGkB9JfWIqx51ettM
u2pDBwcHTrlkKwA+W789dt4WREytRjmkJuAuOhovLRUn9KqFAPPWF61S+HHYBWBeHlxc665U/wg3
55wlrISl8SXBhOUGPVc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bZv/b3M4JYVaBF8S7ZBwGpYrwTNKc6COV6GslrDxCwO4aA1yELtJPTtkKILCmy8IFZM9BtktepAB
8Y/GfP5Zvkffm9OycUg9b444iEC1aylWo854JBsY7OuaJQ9c/C2cMgxojltmNWdx+t9dGUw0q/fP
QSMgjOp16ynE/6iche9QP3Rx9L1p06lw0r6noJ+cQYrK4L2b71emYTnIbR6Zrz4VmUphEvyZRVjj
yRTrT24i7xB/piWEVsAw9DXYWW9C+SgXnrMYe/yevzsro+mKydXQfmW2Dbmt3sY09vHSOMFXZaUe
TugvD5D6QFYttU0YQgutlIEfR7RhTMq7uSAZTg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CSOMXEp+WOvW5Htg+t0c+90atBozEim5hIf3+CSoYdTFFf+wWorqu4mRjDKnMNPuW0VRunrFbBdG
UpMF4K6THmtyXXwIrfVgO9FOmsaKczar1QzWtKCY0pX4UVdiewHwECMjPOr5jwWiqh9q99zvfSCz
XCkYrYqwNKAKI4PXNiBkS0EHsYL0dBSHV48coWMcPXBLrnB9FjLezyXelOQF8LUsbaCJru94RizS
mWbmsFngIlU3c8V5h4cSM51fiLwNFh+r/2AFm1N4ePzurikPGzsWqwEtvd1qTZn7jqg9BI0myU1Y
FxH2Krw+g37LCvEwNT03+jBCw/fNncwPmzHGww==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T9AUf0pY9IuRfLFQ5oO3C+Ff+7HAzyLO5g8IXVyHXsNpsYTaz+tuv31mc7s0mP+bJx4hMUQDQb8C
AEyc6KxMGDKG+0DBKifbVWvlgVuneVHYBy5vDyo2O6fVFQFig8abo7a81VIEFbTDgb4TKRy8/LZY
vdapPIZ1PO1kaTTU6Nku5fWv7YdlK9LCfVEP4uVZPpfNn79aZJmirhcE6rShAYJzcHp2d4fNp1US
X80+dNn6y4NmWWdCX+qRwvbW8B4S7N1i2JlW8ieISjF8kxvZVmEA72fJpAhF1R5m429tDLfth9hQ
lV79mE5RDnoga3gsIjQeqZWK9G2wADk0pQLm0Q==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
blWUaL3aLnYr92n7sNl022vF6ZGJmI4QFMppXGoWIdsoMky/XBFpyK7m3+RodQRO/HelByiysPp7
zQOkPXLiaVvUofzo9m2HyPWPVyJnz5TJZMHXT58n66T9/2AgTLGZGVXJ1SJh0gGqlkzYlYDNApIN
It5vEpLzMakHV9olDytQH2H/2bDfJapFSG5EG4BBJhFKPYPLz9axTzKH+NwCp34SetJ9IEwlcpkf
I4s6/jjLbiZtdgzqVcxuCm4r5rAxcNhqCWQyAbh0QF18n9oVY/iMOKVyOwGU8Bukrgm1EOqKJ5JQ
yaYm79jd9vAhZExjpacnSigTsiauARM2YOZ2Mw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74064)
`protect data_block
kVqVGY1xILkXefhtPndekrEaIkgdFCks+t4fw6uazGGfIUEfFILghDEr5sxEHrW0MzZ2FDegJIa1
t/CRkt1r9ct754Q+UKFG/ZSaJpjUDEEQA29zN14RRCT9UraxdwCJLjZAKk0xa1oPCWIcaikAmv1/
tqTHnwIoTzRXCUcZMR0YhGmkCSAUiaGfqc+rGkdOZjdNCWgDU+6h4b/pEVVTLiK8GDcJGpeHq0Fo
7w/uuUEm94ViTLcktERSIadp3Uzr8V/Ob93Q/ZefLhvNwWs6W/IDJfJeHgvIAOludlMfairP1FOI
udVOAcBJez7xFlrG/N5Pl4V0UTXmIA3OWz/Hae3PP8ODAFyUqQvdpaDz/a+kewrH6WGbMukdwBCb
/teowqYjSVNJ95LG/dRHVtDwuEwRefODhUC1oG2mZAt/hoMwMk4vdThFcYuPwWE62aG9HNN3J8vL
tJpyE+CIxh1LV9O+/MNucLn8EI1FVpokHcD2a8DYffEBxk6rL3tFNDkAZO1az0SLTv5m7T6+QoFd
VuHEs/7Tb97eoYTxA4oc/khXneRlUU98ZT3ZSLT/FITy1DeQX87fmnZZPfZFgZFzMURfJkhdDiq/
dW6ZG42vDXt8nlIfggvr9TB2KS7VmCGmzVZJ1ggSWSWdx4b4ox/ip1GDXQIUn47Itt1efv37rZcj
lb+3kTZoEb3lihv+uWSzO4heV5+W+C6O3NlVbIj+K0kksDl4/0jvKm+rNyZWGcoE7shaHuvbsRHZ
MJApT7vzhnSMMgr62kocuupvaGQkO2gCq+Vc9wJcGCmT6HbOk25nDErN/Hi/bSSnWLqYBmZ7PYJo
X/l67A4Rd7nNQ7sxp8PV5GGLIskJfslJAQ0ZKWYa09KzRQfMyMqsyVQfS4ofxS+Gem+jbEXyNAY9
zrCHjNK3wTr0UrPHEv9xfHLe1sBtauszvoPT2G2tbr1Ad93vnPUa0qD8yaRhTyBBGr9ai9VKgCML
WxqJXiyHuR5d1be9NJd2bY+vGCoTmdDQNi0QFRF+7s/PLO3nvNWv0SRlWW6GaLFh9KjBtg72DyVP
hfeVqdJbOlKVdJ6mubAWZx9kkG/O+PiYg2kIZQovHJAHgYtTHDw2ZxLg3nHwKmJKDapf/R/ovyqy
cy2/JXU5M0qy4zB4pBpsKYuNcEAHJxqyKRdjf2C4u16TThB/pc6F74iFx9S2TYO6l1rD2rmGgU5n
E0zMLCgNTyOXt5lJa2uTF5BKByiCKiUshrr4TDXMt0w5opQNkJmdAty7nzqIKmzIXDf5ITH4XIzh
/plgzrjrA2mvJH6Lua8tuhyYXQedkqvwpZoEdDy4UFyntaEVaHHYbcWiOA9y+qLJZf/lY3K8SQ7x
XRSSdrWn5DorAi4Jybhsifb2mlfp/s9oIrhPdcJts7TpfNWZqna00gjMeeIY5599dPqacmBLW2XO
Kgd7PIG/UkEn7vTg3/7lM2e1NDie5HqobjOpf2riFe5/BusRh+5GIc5/MGeZJyYrmtNjdtS9D9un
BVlRrfWGYRe79i1p8RnwvLsUt8w5z6PIGEuCoRaNDPgwAO1S2IzRE9Uk3dQxhfuCw8VsxHHOR2zT
W4JWETB9IUgVmhxN1Q7fT6WutA/Dnl+y4YYasI2sFhKv/k0GB8ObIQcG51Bz/5MxRMHoXJ/pjsMH
shto/N0rzXQIAF/LtykukTKVjiTP/jt7Rc5Q2y/k+faLDhUFT/HI5JA68xK2AZDo50+7JBpKBIBh
lnHg0LaDyl5gBITJGqZ7gpXB8jsQxfGQn/95ypwMJfaVWr9ymW87lpKa+SbptBDIOZkPlsGoErWf
P2fTwz4rItDe8Z4IOUm9cB0Y9AXTaHOnfoUvwr9mZs0s0LpwmICxUlOT/dak1dweWa47rNP1BdtF
KfWosepx17iWsp5LhKN3s4eRDb/V6HxmqbUT+AxyxWHKAxe5W1PkIYON0BsF/GzbP58BS4NHOsgZ
l9XESwivZvhOCWZy22D6braPVooRDclAG/74CwW5R5R0T8B2ZgBfT7saSRT3fwAAcNzJE3cVtSq0
D4HtXRJXn0f987gtlaK4vh6/HUnIV+QARQtE5TIHOu5QIfaA80XeO+bRhUmXppMao9Z7F4YNNV5e
yOl4aPaekB0ngMgI8sDsvhvoy9yEhQ3ciovQbQN2Qx8dSwjQkQJyPRHlrMXKQPtdJPvA0Ix5DelX
4M6qiATcQnIBtLF2i8hFTqLARuQKewqLW/C3KpnGbLfqntN0xxd5+0JVONR1PDLifACSBa9cLmBj
j3sgf4T1qOyjkmdcmKf9TLaufFphh6EviVLHg2iKPqJoDf+6Y8SZ/k2yBp75/P5J6cbK4tmHjiYr
iErHYH+/42fL15lLBTZo/P/2otxQIeWZ/MQusglPUcO+ORzN7ZtPnbRweLioELQJc2wDDHWWQ+Sr
tYhVRiNfvf7qVPy7qZd6WwBcj5gaAFVviIkXD9yy+0p7VaFhWetvdvn0mnWVZL04lvuRpsqlWs3x
/0lm04dEt8XwHNYRix/rT227PbkW0l00J8/MsXwYEKh41JpzliUG83iNgPk6ZWOj6dS0CBK8Tgkp
mBGcJvBOmSPWRAtqHXuNhA6WMi6XqB+Tm9cEgm2m+Dlc+MhUIanYDQ2MbsMAqD1BR78PLP3yPa7F
LbYRkveeu9svQXsvrDOolbnq+02sCIrzXDLKoINwuxqQVDqYdY7D+xrLabzjCg6ZB+yB8wtw6cHX
Y0qasUAFp4a5TtOZh85bqcQ1nCIzvFY/Eeu5M/KWZ0mpT9eJtnzbeOAcGPlJsIGuIQULmBUNisnb
NqJ6KvQ66c4JrAiSa8lk7owI3dXMptMLfaSV7pDNhIOiwY6Ucwz3eFWxlZXkCFCzc9YWMlmS2QuX
yHIDNkgRE3mwb0Q61WclpGQQu4lzMuHeLTlj7QxH10EGY4nej8YKrOJiwfRRoKa9ydJswlfZHZZb
0GClaXwIP8LmqMIlZv1Dpe2j65cT3FDdb795/aCSPHLio8DxEXH+ruuDBTiXU8+ydsEVaOsjgG0s
+5eiTilYnmKDlWRbgpKzA3ughbWGzmS93ImkMUAwAxkPJ44sBDuMQi3rgwqIH2bOoo95WpeNIjk9
0TeaEnNN8mNN4CKQ2Z8jwxQnD9NynJzWQX+A/GKBzT0yT4QBx1Q9aYKW4A7PVicmJ6SUpifwXOWM
q33DC1lJRjRzkM40zQEdymvuTj7UzFDcqdfP8GGos2Bj+SBdJpuRpO8ntlHN3/RS8h8cOJtvMVcT
RRFW6R4ZWUihw7hzTaq/CL57K3m6ofG9AgrUNkbc/6RLtaZxH8baNsLLNi/+phWCUvb/xJ9OLi1m
FGalOjHhrC8bDjw/bExYEICHD8vqV01rOaRvcXKuybIygd/xhsSRExAOyPoelukSmj8MGRMA66AQ
74hWmkjcy2O4UVwBYJ+ZNdE7m6eNfrnvZailhI+rjZM7tQubjBe40nWo7v2DQM/wbxphlDxElgSe
Hac5IMtNoEwHt4DzKnyohQj7gFy8Pf0RFxnmlgnNXk/co8q68JZHgxl7Nal6NJyEr1DB7bLt8YEE
V5ZLooREtNiQ1sI3gzbFs5aIdowrDsedBVSHc6DaUualycrSRfR+cVyuZP3uQzS/i51aHY+CwZw9
vedSMNiKvpybljmFFVxO6szomFawwlrnOSjWF7ZlpuF/7TR6Uw3ZYjW17km9cPutrZp45CMm3dXO
mDi0KjPXWCPWcCazq7t7fO5xBxnXIHP4c4J6IsXk9jXdnW25JTWcGnptQz4z3LkGfWE9DPcZlNDm
6uNNGRprpYeS+i0o6ZcCULMfJIX5EVqu9ROubPXpUKO2PtNzkYGrLH9xHVTz5CM2Nusgh3F60tip
crqJl9g1EGeUsu9rud5RQQJkvLEDIMo3hcL/ierxl0ACev+AXaQiRDPDFCmDu475vg0tDZSyd0GA
Sv/DdV3RBtafSNQmDhd5y6FMN7+vD8qJcwk96G1JEI9LCKzLsdxnrSsoTWtcLugUIMqF+Jpx6ucb
IODUqssVx1BXOQJAzhq7SkbL6UmChey7G27q3X3maSeZL8OSxzGpThegHFraQL5d1Jb9lmvzWvSz
YLm7AumSnSAiiBacHBHxwag3OwOmPUL2pmsVQHH9pPFw+1AzQDQvdCeiVnZW/1yULvWiPTuouxcZ
DO0/nlcBmzO3boBcdkNjzdTFiLxLzVfJLEKQ7VltKwwoQLokvfQ29UvG/4phQqX3D3pijS6rvhux
MiOLeAP5Wh49mIyCj7df98rM+EK/fst/WmE5O4KRjTj8i8bK3/JQmIwe6Eu7syE/xXUZrQAWjqQ2
szgMMYp1JvzSjOhmqFU1l+ZToo+eEJ6KhC3FShIflPIhi1IXpxXU0LZmnb3+U+NDjMNFn/HHmnmx
4y33S+MIDGl6Wc/ZYzWq1V0UhrD6Ti09RcZ0B83IFcergQQWpqlpIr+c6qG9XS58PWMR4OrxD522
zkbVx2iT5PObJHyCHY0mNimc2bijVMm0mna4WGUCa0OiyIU6BIUK3cAcFHwLNcHUTz/LWnMZxsV4
cqbPt8NfZ+2OL4ZDhbB2RpZhxQJ4B4ytg1tn41FbakZz0VCF7UzvPMkFUEyB4leX8Q+ZN3nxyjM6
9Zh8xO6nRRSy3S2m1X5N2bdXY487X41TmUl8icUEmZ1xI8TufC53Rz9QFZyZ5gSFDrU7VCCIE84F
Epg6yIbDMZlUYuVOQwFNHPCyns6rt/Pb6t+EpMo3rMyb3Bqo3QK++iAk4Qrj4QZ7b+wJ8b1lJ1pg
0RiqH5L9BeAb0dEQoyx98U8gAD9NBkotomRDVF/2Lnz9Uzx2Ez8/gM7QXDpOYx1QOEJ5c7bkc+8w
eHol80zn5mq6y3nDRVQ42KfJxG0biAXvhl2Tb+LZnHR0TW71ce657f1G6qcR9m1jf7ps9odBJeDe
A7tBWRPyKp71wXFXkjk7jTweufHAzr2FVfpvEErGTjfM7jJOFQXey7V8K/NiXAFjuqI2HhvK3yQB
+hAbFhGFyeoHH5Jd640UuENy3Ta1ptkTVUa0Dm0uklNUBt5ynS4fq268Ur1xIj9xWm+BfvTXtl7z
n0Cc1sTfpEcsoikI7CB0py0gQgGL7DvY1G4n7VnbGf/nbHcP9jXH7qdQiNADlv+tjDX68byCHP35
5RKknLHCftb3Cz9YSpQ+qF3KLsxKItwN8Yi4GHEDFxSk2KHDOeHqhsPFSq/gceVMyPoK7HacgHmn
px0PXTvONb+1HNi4iS6xfMcR7kCKdISKuZiQguR8fbbO7EXIlL7UZ+27WwaDb7AIfukl7TqoXtS1
PVhh5lQal3KVmZeAbxqkz4F3popsnI26w0tZd4tj+4pOUtQwlHX+HLfnA6ulpK92ZRMboKyeOQnt
dxpJTciRn/B6gDxDEyhUa8VMIb49DBysUPJ28P/N+vQf/h0NWX0nDclotgxPnSLskOToaAyBjqvP
azrv78srmjC/D8+DSVvTGTuI0n4kTTBAaASSx/q/YqS+CcXESVG4s4kPfDUvcnob3458TUi/IYfm
cEYj4hJvp/J+w016V5CisW3Dyg9pkApbdQIqd4zaXpmJZ4S8N2DO+txyQzHIcWSkCVmJ8RweP8GM
nNpPr3MOVgAdKPgtVkw05OOTrlzZtHg6AQi26pSzaEbnQHkSStZ/fNAnNF7KDmj79b8LzCDhJ3a5
cjXZWNGYAt9QcMkjmcACWByB8t5qHs3uV7lnw+fCW6eOzhAhT0duW2cvAxXuBU+Vy2S25D7qmeXA
BbjP/tZxzaaRraN+6dE9SGXM5Fc6q+u1/4z4D4RSVQI2F1NNAxKHfpWzpfWOpMO0D/uERlXCuSok
1s3Dlo4FJcvX1wPopf1XWR86HVFyaKms/cXr3AV6SjTjTlpRCvtH5ObPWu0ewM/xuNVG4sTn4L3V
E9cBOSgIQVd8876mUJ143TMEq+bh9zYajsMibt3eEwoX1uFYLxnY5Myplxo34iLOa3vWlREX1dHR
/hx3uFD4mnGCcBrbxiSmPf0pi1M3mIxuSvg+eijV2B8McpoPByVNfagUefXO0H7g/d1jVdqJBydl
iLcbPJUsI+XEalV3rrwkEdmINPbEdFLV4fnrZwK6V3okTAv7MWIEgPFoEi5XvZPPlKg1tUjQcbAg
gB0cDnPowYY+dCPmAYedpWnU/HOzlAZ6obO1krak8P5b/pJtIC1z5hgksE0frhu6GtktOHWs1/Cv
e577pAb1Zl/L/LfkL8gWzsdnM+/vMWoV95OcR3I69oD18m5IIA/vrjcvCSCHpltzDlBWDIwEqLr2
QwJo8M4WAzrvruuv9g+L7Kwjd3pmwu9HoZlRJD0zBXcKixVXAfseFtoQJoC35fkTf3N9XQw27Crw
ZExALqUFKrRxlN1o6zdHjUA8VIhYbviWC1Rx0j2aTwgks+NhdD7yHvOsaEkZs9iRZmERzt0Kas99
I+/8aAx+Ktjbi8S62YRY7m5ZjqE4LpJfs1wgTYzJAhA/ONaQmZ29IFQhB7zot335M7MKhVlsiVk6
98IHqos8Rwe/857Mou6g6c5WFlX08Q9lxGRmsvCGpclXYET2mwotD9dC3SL2NyTkrN3k7R7B3wmk
ioUq+3P4aJeuqLhq0aTU7IH7sOnkgTELirXi4YmBCHvTA+jyIW7xGI4CKfdU/yoIlWJd3/Y9NXJV
Yn02BnFo3mlXPS61AuQJk9zoBVROJkvg86yN5AVJpbotJlzkj4XgtuBFdA082wgx+/I73dZbHZLM
YMUs9FmZuEjQ916VDg7H0/D+WQUq4oUaFBEbHM9Ju1cll9b7QllKPAWKR7GjNwsS6shbK1o7zeAl
eBYgxiZ2YGFbBVUFuUbxoh5GCj+aRHnIxSwNZs+hOfd2zcJm3dXdetqlGIIDbUUkugkFhH5Z+kGL
J+3AJoQtmS3pSIaYZS6PBKUq3b2ug9jAL+ofbCnAul5p50eDxxPBc6aTExGPNfpRWRAkxg4pEh44
ZpAQgZtm10+eAQtrUmzoEgDwokVBlU/St10Z+/LA3dB+Tc4lOS7F7tGtOFPmwa+qdpbsCp0TRDbD
gyAV46YUdprifwqABZo8gENolG6Pwj5Et8xyZghG2uzi+ewq0KU+2/CKzX4u1za3+xMxZXTS6lV0
Oamq0ZUlyVtr1K/V+rwSU0VsCr4byRZ5dgQsx4BEDfbqdtYlnWceJmDz+IvwMxeYWrxJmp2XykfP
eKE+GPDY01mW7jczONQ4lmOpAW+sm1HsGEb2REZn2TEzrM/WC+K/CaXbIf+iu90bgWw8Z81f52k/
wayS6C4MIrb4ZZ1TXxiVMI7YUKsqJyaMl1y5x2eXQirLzcQ5Rnv4gUXnlAVveZ9IzqXgvponH8qt
CqvvKqi5g//UqAk1PWnjz5jpnpAJ9oqUvhKnm6ZewBZ4VAxe1h00zJ/9vm1QTix6430G0cXJxNz5
Lm1zhqc5xUikDCI9kFk05KVKq2+/vfOFfEvVdHL0JFJ+8xhCkyxNCpqB+XUovzOublaCDY8Q3fO0
gxuNSbD5MNCFelB6YGGPZ1Q+NJnPsm3nUOZS02PqZCR11MzvXf6Yefpsg1DU6C+AgpCw4pCFermr
1poW02PlXPWN7dP9GYgeENdNYFmjnOVGRbBPQrx4cZlAoW4a2qWVcmiuhIi3AI3cElRmho/dupWD
WDdTVgZDrO9KjLRYsizco25N2THieIgOQ/gMEM/jwr0Yb8ou9uwzPI57gtjdpzRR0eD3vu8qjqEI
vtq2cDmf9A0U+acQkHyzN+LJ4KvrGdTNSLvIp1SjQNEIv86NsRv5hzpss1X2XrJJ7QBlwWsVyPI1
JPxNP18X2Q6kB64bMkXK7J41AGMjK/sl1eSeLG1J2HxhBxTMgkl7NB8nAxIB9ODqo2LSrrzXduM9
tzk9y5YloEd+UZtWcDyaZU+lbqqUli1TdMH6bAZKcw43csk8+MvWdQqOVOYsOasxHtBsXPzkNES9
zq+rOOrzrarZnGbVzUI36Illh8kTlm5hck7AoyNd+oIHlzupDKV5Q8QPOnj5KloBr02R/3poXqYo
Jj7q6awGHqwy6oh9NrHfWJ6ejnVlt+Z2LtR7cV49uuSTvIo+awasMNvoXDltnFxKIiGs99ETviS6
Itfm1GFpZzHBzVh4opqNMwOFa/mDKAz3k+uRfXUjzEFE1Ckhg1ccJHc0WuyxZvKKmbq5Qo705a0q
MtzYTH4/tehibeFwb1QGlTm4wJFq5w+jZAGwZAdfDMmm2ef+wq/aGHVwwZ/EG23OPeNQOBb2msKT
GnMJ2TB91NDJ410NMMJQTJRAXOEJyrETqQrPY157FC+KEWGhL3xBcb/52dFaZIxjfgdXS8OnOMAd
E7U5lknj71oYZz5+jrFifdmleSAsJopPSDbqx7+IVXAnuhF2HwmfOAckdhYNTd0+J3iuFUSqSCTP
P5hytxeOKbEVtUhQ38KZJwLSnbHAt8AKVDXtwTX9M2pMwQYrqz/Gvx7FeVS7FwtEPi7V9zlNohUb
Vf9ubZKk3TIYtn3X0gHozm5i9x1Kt97tWI0c5OwGw0LbW7+9ajYUUskbRji5F0A5gAkp35D1u+Zv
rcI9ZRQ9gEoAFMvPIgwhUh65QMvZK37OlkKWhYUlYET3AKdl7TWGgfYvIfdbUFDMS3h8YrsZbIYs
Tfh7S1f/KpUZs5j/3NsmGqpi5KknNmtu51LqmZ++PFpKaqA4dc9GuiWxWnoi4Z70nqCYa4dT4Bzg
R/H1admkD34dUdrAvEvTK75aNcuyWCYuHqhsEbkLBeKt7QfNNUe6z1oz6jEpH28erG6AX0SmBzAz
qQhuXmE5J7uNlTPgoIrxtgb3bZHdIJsZoWKCPX2UHtNbaUMoXgtC5PAwbM0q5RtcHHyLlBrYGWtD
1DH++T7lTDnZ6pTtjvkeHdvdyPV+KhRLVXHKeQ7d4Hds4eqjaSHctXP8Wcx9H6u9i7AHVS0O0jPz
lBizaOaHbRT4J0OQdvSqVJhPuzGC5P7EjIzPDhP6d0pKijgw3kIQhEGfdUFYqq2MNv401MWAndu7
ZbZ7YtNmlO879rV3m6eLGIGYsE+6ElxPvunTuSE44xfxBHT2pp5V5LWp6wXNYQBbzjIjg1Ns8Bgq
oYtfDH/s2IPZ3A/KohwuveI8HcLvbTEhJYLudZOdmLgLNiWA7TlWik+4kBNAvzxajHbZYemlf9DI
Y+nGFpyMAtAnezQVYaGjNn3VMTZLpw2JfgOiE38yDY/KFrZu9MlmXYD3FEYpAFHLJkBVx7ygfYmt
38m64AZj82IAvXoO8GIX4+Zjg7hvbpVpVRYaWrYBkeTscUoKP8Q3z4h36LtCAXK15Mfix0NEDIR3
GvHzOgGfVhKZDEkvOdljwMzckKgHhtWhYc6VHbNvbZO1epquLVVg6SrSAVRK3Qo9ZL1XYyZNRjlc
YFq6z+0d8I0sUCJN5iNVDTV3yc3bzoElsl9kDnsTcY33KUm4F9qH8Qu61Bd2pk+V1bws75hWg/cg
lTLgUHChHM98RL+aNUCdBoCEvFC7G6jE/2N+z3jrQnh6NWzCGurkQ/OsUrwsPbTrCCgR6W7tmKhh
NygtMe6IBIwu1aBy7pt7s9ALrI2cjlyR8waBaaG88VYATRh5NeJ0jfHVA1A/VxA8aaV3YGWhsuWN
F/9Td8g99U/IreVGzH8kdyXkuJ3W/NKcXrxqfWgTbpEfXF5dtecYzbwAIfbEV7vT8E9v2pQKJl89
rybOdOSVdqRCEp9+iPbd8Nhpmlj77rhd9vcFE3eVDTdUs37+iUfar4hSHcuCkq/RwbP7Ax1sgxS5
P8iYoCDlRaT5m6I2pj/9t6He6ZcdLBvg5s4jEpSq+O9Om9LLSEf/AWnJU6mUILXOIiiBkhqjnH9Y
QJxukieRx1cLxXIH/RGUdK1Vw2QTdqUHTgZegiw7Z9IrJ7g4NxVU9Xu01o7o48WYkh54hiBKt5Go
4HZ0BaPJu41LQLGOO17z0id1c9A+ntI9W6on+oQsmqe/zZh0qTKpDpbxE1rUxFLIrK77p53g1hIc
sT6pZLxv6+jdDYRIwKNoH89sSHYSSA4LJLarUTOl6vwgdvXoxhgz573NSP0ghfYFYVDKIlv3qIQc
6GpnCEEplzXdzGojDN8PVpTZFpuHBivoQpq7XMm/JONzl/JKnBd2GMNr4iUHYKkC+SQKhOzx6YI9
Z5Vvyfkq7WmzgSaoB4pG7xvnbBYEVurLHjW7XKX8/JnGwDbnbBpfdIl8B8V/lf4rT62b+NvBmDFj
fAoEQmtEEigekkJkq7SWcBEH89nFTkC9+ThwirTlV8PtEZsX5jM51MfWcBx+rU/w1EZMc0fXeaFw
zVuurZXcCRSsKCPe+0xXKqfzASTxFh/ZKxeoDgP1VNIFbTAD/u29m8Y1WdBWPRY/ZvxQEveoQW0K
zhx2xCslm27fEwEFYTcu4+RmHtkIkNsxQOB6U7M3eQvysB1b4YSRd/nYJy8FKHpE6s9lR9pdQEDL
7RIIDkZVyABgVQvfp5cWwA4S/KfP0BMfEMFpj70UAwBg5WJ9gZH8efUcRUzxpuMhHue5e3H+FwAQ
iYvOIvK7ju8JS7eTC1+tfB7S+14vKVrhkA+lN6ui6ztSE0dR3H5X+LsaqmHouAKq5GvmBrn7s5VK
6xEPW6cB7zQNcQ+CQxp3i/a4+4fbHkhkdTyue29o60CM5oS+GQt4C6MAo3qEu5aA/a9zdCLqgW3b
6s3601aUZ0Z25LUUghRiCiIwpmsuzVz8rKrPWBYpBan5uNNS2md+n7og9b0yjvyHGhwa92wXJ5Y/
JzmRaY6q+MXvWi5IvrN+Uh6Pv0NkLNUbNzKaqo5ajY54r0KeHAS7NrESsVzcE8KHoA8HK5/gaqN5
tTILD/+PC7VnHLHtsB86+JX97llOvnJOv+Kh/675QNB4E5vwy4WjvXr2YX/upZ1aJ8ILj4Rg0WRo
CC940tDKG6M4b1TsCZsf15ZFogRwTxD7pfb7AxkeiPn1pqISy9tigBpr6DBZfXwXhQ6BX80Ck+1U
ejEhUFo6hMO+XNt5SpEVlkmGkvGzWum00W43c/KKHcT3nBkDcBpRLwyppxcy0FPk2Rymji4Eg61o
qJC2bAF1Vaa2y1HqLI5R4CLZ7zjHjHb0DZj82ftCpvgKS9Z+ontJUyFCaOfVYYjvebhzrg0SaxgZ
RZzK/rcYi8gAnX2Eou1bLFl949KpWfwE/mNMhn5gUPcfN4qzg4F90gDBjVWt15mfQ7sTmm4nRgao
khrvivet46222/zWj55xM4i74dyyZzJQdXGMh7nHb+aSVaifqHRqH7i7faqQyqJJ82oGukqX+leL
n6Oj/JtSrryNlwOMSoWFfXYoF/YswlF79UY30znb4Gh/XMbIGG8y7KcxTm/XGb/KESfroG7+qWDG
mb9tsFaGtoL5Rs4u0HR9lnpOFIZ7w0Q90cRqX5ZwmLz4kHd7V3axUXbgNH+RBXdqziUMOG+0JEOF
A+10MyllC9cpUJ1Om4mBOIqTf0wvDeQixFzQBQYiatO7P65NaNTQ2HoTckrRR5GhjAr71lzu876r
nSvGpedk/21N/p+0uZB2SSn+j8dyqUhDqEON8wEFxQm/+fTb6XJCByk/Fyw8fNzHKuXNDah+sA5C
dxPBcCi2g1tcsg6WE3Fkwg7XPZdH6i0JmDVGdlPcasydq+eK7mOqQC7QECBX+INbzFH7634kZcV9
1+u1Z9YgcW7laLaYGSjWW6QV6dPbcVIsV1AzzHHu1EzzFtP/Ip14ybHch0wFl7bkOCQ3kCFHdrBV
8+7m/WhUQDCa1ji9BV79jqo+xznFKWg3yVUruRUv4HfFjdIhtSmv4iQBlC4lxOa7nZ0c4JOFoZpe
CRxspCdQdBPlyQS9s8VUO8wdUwUDY52XDJQjij201RErG06491JIRYqbW/4UqB6bmv29wYvALD/O
FCvrA2EYf0uD6UxlheIfSQGlh5oK5EALlQ5w6ozwHTiHWtpNFLlBmBhdQ7Cjp/8GBo0C8V1rjxML
36GYY4lrrw2/oGmCZax4Nsvl1XlcSP4SuwwYxhpNgKdTW1mBgoF7hoouCWbijgtR1MyHTpJA98EL
du0EhgI7NZQriF82CyiulFPGaUvVLiDfTr24CM0IidfgAgPf/oEzrh0txirJXGvEfq/Lr7aS9RJO
FGanWPQZzm7KGTndRxYLb3Ho0D8dRHFKjjADHDxRMhvVaoXzCMgUTy6/u2+SxzTTD7pWlmwjY7SC
3fgJVYCnezOoPuRXOWyXCUs9jWpk9JrNmpX1xXbEP1rqaM+iwf7Dd3OI3/EvHAO6zjOdgR09RLQv
IUp7ZxqoEURyUobbdujbmI7QqTJ0uyEc8wRLX9ekyoJoOdd+9tpiW8i06zhNvGsYgf0rKi5m79hQ
ZZESOwu8j6jHvTxBpfRUxX4Vs1id5302qY/kqSq0Qc+l0FPe1flFBprDjJUggvQhntpi5rUo1Ima
wjKjMX0uCZdd1joPh8dLtwUZRg3oZBVhFcHjZZ9ookd9R8AZ6oZKLQuYvd8b2XakXy8E9wMjcXGM
5wd48kn/0sqAi5klzACXqm1oCgjg/15o8T7XEiBA44OODLJ8KUlHXnrjwOotfGtZvFgb6suRiTzw
R2zprbCfRZEg5SLZQX8xosGFpjodUOnpnr1n+cimoajtTkqUTpNjgtYOmPUf3MGZDqQPJ+LDX8i5
V/mkYQ87hahqsnARDlw6PI1IDcOqApg3tlSG9TI5s9sDcKN25PcLSjYOzWHVwdCFGMHsvev0clvD
L2nbTGSP1q6auL3J4/KW14Bk0jwJBw5vScZoEXskMYN3EGwcwqJUVepQIvzbcwU+82DPAM13tGzO
aNb/omrpXf5qMoD/X7CNK+p+MONVFXf7igOpP1NjvInOgJXQBtr4zlCqqJgqbAY74aGp1FBnOtrG
sjDVOt/8hsuGcdL98QXXZWYCgRKZZNlT9a2RGTMDBdvT963oBc4YyRKMUQUFBp6zHQzLeydCkZ98
kX+xv8m04il8rOhZcWJdFprMnstR1gPn6vJHrw6jtrvNnQfZdnl1bQZLx5NSIhS1XRK/zXEHdCzf
6cTCjkgmXt1D1zQiN03bT6mYlQSPTGGwM4s+VpuZ1WNCMFtviXZvBU+8KAb8f9L4iU984vZ1wYn6
6XNC9OEe7romeeKheZ2eShjJtGEPedaMYzleJ+LNNxLHX93f8q1z8+nbDNMLq5wVRTorn+4h41OY
BxGJoBFwcp8vvQzXx3xULMTr0I/jWPMlcJRXcEo5w2nvNIrsugPwu4OcFO/dI+gIpqOj6BSocbkx
YxDOxpW2AwfUMkVJMXk0fc4j9+i6YNR+n3qHrw1JcOhjhRfS/o7gJ2u+/pLZUmQexBWOkWpRwFyE
rlLKb8YjXbj8U4T0Ipz+9fOtddtEdeVOmpG2w6l3h0CpHudKEbIFFOM4pfROPoeDIhuW6whQYXOb
iinLOo2XJ1uQibHxio8f6cV7AIwfEveFkptLSL4ozhUz7whj6dJ4v7beJoo8wX/nMfmkGrF5AVhm
yE6zLLuTzlr9S9tLWbvyPA4SVF6pOqLoYXsrtP/EJy+/L+6CdKk9aZ4OOUC8dDWlq45AyehjeVrh
cdXXBGK7zPVFf3vrMi0WQH8HhH/OUzJNgTR7QJE5hPGjJeCG86uYFc+9GBspZ9CyFGl0D8Cqot87
e1IhgP2YZLiU66nWVVIypKMg/ms0fDDmVx1A71X7qdwX0OY08PKthGpDxNOimDRJMBtmo1b9NDeE
1lEj5l06Cp7PTE2L+Ba/lpMzn6iaR9+msU/NCHdC2REWUX+EAKho5n0xsALZygIR+3k/R5A1OJT/
f6vaPbfQVJ24Ch5uLeG5wAsbSWJwS5m32qzaByXqgm0qZxy6Mrq97NhWZEt7QYylgLSbG0SJ8A5J
Y/+3SJKErYOZ4gWmqwEcGuqukYQ7NYtaULou2VpFNKvSowi1H9gp+mOQOgqcrmmGDCvFhxppsmlN
5HtuyduLagRnEiKwzhLM26NEDviZn7IsrS579Wmcd1kSCKcoH6KX2dME3z5eNW82SofOD70rFgBN
8/vZt0DJI5KKSKK3/qob0y6L/p9P2lNbXHeHicmEgx92PQESIhYd5RTvt+dIlfzFfIUcrDlAa5yU
AnOgH3QYgXl4cc7TPZoKM55LZQkd9rdAzXXfsUYRl3VEe1WKULY1BsrIZS33KBY5zMqlpbSfBwYQ
li1EqIJ3KFoVKt88aQUIKe66Y5qoxscdD5mTQaoBtioebFoomcz79WzbOAf+TYwyThWNgQ1m1hKB
B5gBZlJ9IbxKz0Vtgku7lD/g8LtRjaD/J085UsdD8G/hA7IvPhqz8PvJKM3uFBbka+03PYatVhIk
GfbedOg6W6by53/XlH8DLJ2UeyYGPUeWkVABKUS2lJAUXUMy5fYHEZws+9+z9+g8NnqUNxHgwqCC
Ax/sXS5P/hcO+CsWLcDCwKd+nkLsBccYaVbH23slQzzP0o+BbP6zm3F+MzRsH3h/m3HPMKujCEwA
PdDNTk2dkqiNqoQxLixj4bRC0wNU08PknY31FpcZmV0Rh/UOfYg+6aLlwmr5DcSMsUvjgn6vuD1E
bz8SPL304SKHmxDEiKSkCkyfFqDrBEg7cZo/KwlzMK2faMcW9Ou3Ti+hZrSvg4kwElG1ZId5nJAT
kab3EVAxMh389sbMGs2OQi1E6CYe2fHoFy92PMHG5xz0RojKnyqihFl8w3du2kQyOThW7hcMNten
aa2hRb5eThU6AHgYxUX0MA6LXgMfDoW1bw1xH7DmY+fmYrFueQAOBUo5eZMA9f4WU4iYo04hFriY
4dOXQ6JK3qpoMg1t7XAwQgmT/hXz4I4HbtV0JpjhO5/Xr08J+aLkonDY8QUfF6AFdS/u31kFHbrB
tT5QeMafcXVKDsaNdYNQ9FB/OAKEoVNKhWX+oohe2+bvhoTrQbRTDAMTqagYQyplSxIR1Zsd0BLY
Qpi+o2/ySZdCtH7/vRV6W83wiHVgMnTXBHRR2f+ZKHCip0KHH3r3+r3xHDxRJhmLpgn7aVVxT+YR
iUlVofAHwrgbpiPHSYY2O7lAs62rvbkxyK5CBUowFJPbpwhKz+w75sYaBXpaFTJv21McxnEVHVpK
bfQPJVdvYf1vxY1L+qs7UqUB8CtfpbqXyPvlv94jTgdNsE5hTzu2SIo7H7b/tRHpUeOjNvL62QI2
ebJousE+I93ADZhH4RldQ6yzN5CIBD1rdwvqTyh2wRs3j8UkeL4ZtOwzeEWYb8gdJT0SOTsaVjoo
psnZj9SNC0IEWGZ8D+Ab4Cl+vVOScD0rPc6soF+VPfyb5GMM6ya9mfH6L/N1OFFLAgsvBFPEW+Uf
X7zEmfxh7NV9FCCccF5eGIVq92u5x7LSJgrbHzJ8TH1TjGhdcgRNsaCaCB6yLrcq6mxNdQuE8kD5
O1ykbPp3euei3TW1HV23eeNMRAM9DvQjo8+65Ukwft7U+TpeunD5Et9FgIuoNYoKSDCBrPzXOJqy
EyPjxbrNCsoA74kjM1A6F9kRmsxHitzCJt1avXtoaglLK8DrpkXFdoN8AKnAIxXesV+wle2IYrBI
5vQzWzZA3RHwoU0Pmk5JGDy8RN40Pjewne/sJ7EyJvUgfARx5KGsR/iAK5DSqoNn4Ug7Cy7/vITs
VmrtkHmOwDHGALlz3vO6SAKtkAv3C60zPXpfDTBYzVqLUUpNbX2VK/Z+ksjC4igMroa6Cu+V2YuB
TY7xDkZw/5NA6DLWXjyofQuS0mZ72W75h1jdT/Km8SHkEWXQO2Z7rihZoZrzVGP6cq4wYMoNVzXG
x93+u3Cuoh8ZGwR8MFeWTxqeh/XiPloGWdXfVD0WoLCv8xkbsElKv1Wo7S5x3YOj8hMrBjUg3LqN
5XS0e/6BduXIP8KRTtv7FISaAfU0sXxGjuKkOTXMsOEJ74CNUTr1JRUzc/ROyRbhZgftWQJ/c18d
d2sBFnRNOmAAv+H42QSHWwudEHglJKg/LSBdJRTX7iJ/4fVqSjJaNTELg0AG0cU2qLfoFDzlc5ps
I6gRM+1q1pLWSuLCX+7JhE2LbrN/N3/wdDSIhFhDafscVkI3Sq9NhlF8TE71pmchtlzfr/vTJsqU
icsZ92vnWD4KadVeLH2XBqZP8xMj+Lk7Os3R1CI5Q+tTlqDI8fHnHMdBJwotidTLs2JBE4yEdXsv
5TpdE2Zb+95tUJ2ECi1xfAXmm6V3IXGKwse9iKRuBbHqQ1GGOLclnFAr2nv2M5VxPveSInP0tTqT
GQIbDV0ruCoVxkZRcP2CQxdMdmlyKWnFsSRKWZOk1YF679cPa2tzuSWjBtTszNOanPYjxaHVpc8x
RVBsCranTM3RqGs147rKbyQKXeW+GBdj3+KYQUgcb3LXfCNqpw1qTswA4LIEYL9L3v26CY4c2HGX
Uj4c7uYw+9Gq/CB7M6Nb6OUsupy8NWYtujMIOZn7Iqvegh1neb5xc+FJxlEShjpnZeYaFfxqWJmP
249AwYmYJkL/ksAe2sFuqBfD/EXFnPeDIC2KadI02Y/+6m/QGtLaOMuXy+IkwLaw5MXJcVGsvbVg
lwBXDHWbe1KRIIh8DBIdt03JbXzi4YHSdtqRvNuWiz2RQKfBBeWIXhtVDxsOj4irb1hy6Q/Ubh5e
EWU5Ay1wJRbUdqcHcmqPBpJutWH1Z+ZRoWTdWMTGfVsjdxOVwPGONHNliCynxUKqTVOqPbLh8Ach
Z16kmD3lywDc7y0Mc0K7w9Om9Y5MT7rwC+pRHsxdwJrNgquaILbqmWjYp0CfCsk+QkUEGkp43PFX
7ctdblngMDFtA3+CGF7o6ktEeOrLv9JKIcmnEg9eFcIdT1ymG7HZDG5+Z+uPJcALX9ETEaQVwxj+
9KcVBzXDEXy9vU/wzFHQxiE0DamfWoQoQyf/RU2kWDYpU0OwmOJbdBQdYcRnG/OtBVdEKknYxg5g
5A2dLmH6aFeco2zXUQmWsoG9fLdFZT6C1w3kx0RLZ6uPkHoiZH+e7jsj0sO4DRWYURvY9VYUu1BD
7Pm8B5RBVC6T0JnOMreQ693wGMVRkluBi3cSr7/WHMquasOG4UM/BillbHhH8MdBDJiq+HcqbY+v
/Uo9cmKRLUgxIj/xP1C9UemQxWiHVmdjAJWgg7cvfj2aR4+1KQvX/g+JGG3opX6bsaPh/+yAHHAD
V8WuB/CxpbaZpLFb6nmlzYdQC+ehtr0O/shymAFsOJihupM0xsOP+VSimJ2dpO2EDaXcLBrNvxdK
hODszQFqr9Wl8nU6s+huXKMdkOtzIR0sqKDeqEBaZwunXWAfo7dVxZec4hJ8Mu0l2V94s9b6jbRj
ZmuVssnY9I9Y20aAmXbI2DTYPg6RuU7mvLdFyLQymrn/cqyiQrxEYrgRHM0r4adiZPtm7jxXY3YG
q3pYFdupKqUZ3ilOfU5xyIPuTYeeZTFXsq36rMIEiEEBziPXl3UKgF6YA239TWug3+YX7cwcJYkr
jzh0kZJM0wpQdI+k1KVjUSb3cZSkQ7PVntlv4sTcIaj9H3YVlr+Zi0fgMIlHGO3gClxCiIJxqfv0
IDQoHzNDb65GQ9c/vxUQC6eZDepA0VXA36a7VQBoZXP0Zw2db5dHP8Ls7CT0q2Grkiq7raXO+7jU
Xlz/FORkIENoBWU6S8yrxEq1jH3lMEjVABKXCBHB11eyOzlmsbnbc8e0xJe9hLA6jwA6Au+KzqIY
574lZ968AMukW1qeQTDzcmJsRYPXn5ba0+E1ErT9NozYX2+mX1hDJfq5VcX5g9QF+L4tNUZe/08Q
kyVj3RHCr/S2Nk+QmEcBsdJ8HssO+VNnfga+cvi8Bef5Qhl3BbrcgOXakl3Q03Y4sN1q9dZ8YMWk
+BJcQpIz26NWc0z+YaQJfPin9kknGHpT6GlC2AoM877b2caG+O5o0lbJ6vpuRRxQKRe2UHKfab1/
eBQP24lbLbxByHzD3Zatu0sfA6uua6xak3mViaKc7cRpIhKQXfDY2Kqv8EZP/QCLuAtOe+Ywg0z3
YEseu3N0jhc2SmN7XNtdnEjgbbLiNW9TUBxwPE5xKv6elltepvBV4dav5DcsnoHXFbbGrJYV6y4/
i0JxOVfesZkAL24PWIEaB33aM2XXgtHeG73D1cXBB3t5XTRsWvY0DlVX+kjEqlFEM+m5MfBf6yV3
XblsuknZStlioqoc7lDlE0q3ATw042VMAlK2iWGbYTToHT4A6i7hJHS9zcaKnbJ07gHutho/BqIV
4FcPBs63tXfYU2YaGqemVu9cPSxea4M956U8rG910RbS0Tjetoar/x8+CbamzR2v3bTpVEn5MBsM
/tdVBhkasJ4CfAFMwx+HkauQeDl+0wo6RRF2x6qgIvGOk0fsTbVi6tdAOXbCskBAI2D6QSUqkrDp
17nvb8ecj+KfbYKv2MfOOn5cdu7DM4P0rlUYR5mniGCR89/f/zh0zPvjPgh50W86C3e/I0iGiKpW
Cv/9+PRk84Rqt80tKv5lIfcRUEV+Mg+sNTFqaxtjBlpIlZxwAcpXKsBGtoRgRqI3+FKqupu2sgI+
dDz3BPuqGWb16xCniJLZxHE1e9a4ThNatcuA3eSkBT9DBLQtz9mHUoK0PEen1ZjocnDNr+YVKDU/
yjfBXnWbadv6tznH/dNxdNs9rvbs1QXV0f4maIYL9QQI2MB1CvT2EcHdYYlzOQYHbGyBsRjcjNn6
gL1w0XQalxR13fg1c+U5SFy/iU8aBE5ziKA6phZoWWHE7AC5cZJYO4pMgWYyoKIl4Ev6htmdpCTZ
6maz+tKInhAg3NsHxhU2m90bU2/u6Fa83YN+V+Exve7Q5lgxGibUgTHseLItAAUWgUTwI0N35+z3
z+tPvFXiJwPPq9s4xl69uwLr+2QGwFE9gc+KyhlNYlwNF7f+F9R+3ytc9UA8SDZ5fCw6VjoCXyJS
zO3ArvjGJlbkEeEMFuYeP99yD93idnh4VpWpQ9l+aaX/f1aYfgz+im9VBQ2C+rPBLP3SuYLt6KUc
U3LfIsXqu14ld3/t6eSY7tX/hcWRBAbsn5YIS4T/ic/kOoPxT2LxEFQA81BDWIetgNZRNFPouHRZ
hQoy+2zxVgGm0vq7H9LkzgFMhEplDyVz9r4GEMCSdpONEIv2l2DTxEYaOkgnssi8SePo0Upg81ME
G75o2z/RpmrNMaPqroyCyEcqyj7HJcqH+zHJJRX9+DhnFvBmNyEhkJhxKpUeMJAqrMDWdgZ+a4QY
hDeoNEYuIVBekiHcwjsjxTR7fJRLeYcHVTVnj2HaCXN+xOSA71ujXvn9FFMvw3jGnUKjBCdB+ovU
alGY+ZEb74BD8kDRTVZpOKfhRO8b3peKmCwmabKe0s/5vpXrfJVNh14MqxcXmOnjwsck7Ldgw3BR
A7gaENXOd4hKUI7XFzLsPxcsYIdM0rIub1g3Vhs/0UW9zZb1hc+DbyXIe6O85IKrqenVvZFNcqWG
iyLf7B3Kz5pSh8qM/TpWuajul1nQrWDu5dEhbARzOCeLTn9LFOk90RSzdJvlaoaxUv57rkr/FvXc
dZbzNJVUCxgbwIkrKLVFAiAzA6I8TUvgfkvnp6kofniYb2UyVYq8cYmm7Oxnj+jcya2AJI5FwE0y
5SNkMq8lj0PCrvm+mrxbptlAqun/iqgryiEid31jehfkbUWi4R7ukFId35vi5VqpZeu0QRSLRYDv
WksysSNE71yeTJkHeeivjfeJINTsnXA4YdJMQLywjqvqewTjmYVdRTyDqXTYYG4z52EGe2YBdEsQ
fIzXH4Yr6eupGL00emCJDM/myi6rtNhWBIWIWRvZt1+uzLqu4/wWdUO8Avrtus4PytXYv9zyt2wD
2BuMOYX5DYEr0U/wL5oUu1V5orY+zlrkbgFlbX5DWd1w0WU3WorLRKcJkU028OEUhGsc//sCLHWc
+igw/wSclVH/kKWzEUNu7w69k/WfZIp14PZ/WrhSJUdcF61FA5VjEPLOLh3k5ojJkQgoa217qK90
hrieB6LWtBJ8sSb0dkRmYK9pH3wzDg+sqIhHRrkOWf8b0EQo/0iC22cURlzC9lMTXpY7Iw6Q/3/F
j8meLAmTrdP1/c/pFfb9btGNziozSzO4m6f4Xfk08tMRkAzGO9v+1Y52GRuMIWNQIrr85BqLeNU4
rcBlq+fKRA7q/Etr38Syaiw4ba+MfUeDiag36v2CAJ26n5p4HmoR2+FplmqBgeuD5wct/l3tJ/yK
WFoWIq33tGHTD0hYxhdy3ZgWjfWCeB8RfB7HuDXeLTlPuGk379LOPxzHo8Ivro9OLaAE4UTgi8pY
H8VkbhzL1LSosu78Q2S8JgpJ7AzyD2SUsK9OEu+I+mkKHBwi3VItOr4XqX3Z5epcgIPA3J+Eqjij
NeLptT4ti59h8v4yJkM9jedU+tUpRvoamdHwI/IwJFcLi4TYGoFGpS63Vebsjcnh2lMxj8EbOzpe
UlzwmrAyC37HUiE3LNyDuQ0ArSMF0kIAA/hs5Hb2vH9sogi1f7wEXHk6am6J1/ioBrKZSYtiE8mN
77HrSQg/DYBcu5faKZjXgkH7aMpuJaE6OaOm4CU0JmWhpWVRSNEqdZ0M8bWhMV9W+VsIo1fD08j4
LGDE14tmhEDzy0XL6yeZeLp/YF/fFv6+L3d5ern3IoD1J+Q8htzOK5KR3guQGVv9RtcGOd9xeNma
YP5Ah+Uu37KIXujX0pDtposojtMU0gWM2lPMpnLRJ1YTHg9f178ZhdUFzGZW49DakpG5gLYeOrgg
NtYo1n582zKbQfmuUywlIqibdzvuahIPHBymAzDZ5hVPCJzivhc7ql1EISzetixN+hoGlrXAqR3L
4SfIL/USrO3ssjfqtevFl/22nw6e9/Mq7NxuSwo91z8PBZNI7gdFD6nTgSqF428NdoflWm1Q1qZU
IgENlbpumw78S7ok+hV2yos8yUxzS7n6tRBVhKEj200tOUvUEXGnqJ8CkZiHdAJV4YDsNaqcxY3U
Kk+PI4L568dLFfJg98dUS/lJHOQnVebbhXRgYIlqJuic1b65rBNMPo+Fgp3siOtRtrT9zN6M0t2V
V5CxIWQh6F0SUN/ZX3qwS3GBSm1BhPcgQ5oyaTMkqzs89Ezret1rGSf5eq/teMaZbA1wYnN29Jgl
4L7jW8A3sd19miPjwvVwBSeoWUr7/zAwJlxbMzKIX6mxzL3IBqGK9H5ILU5XQsIYMQir4i35yImr
wE7YGbsduEZkAFmCGH9HsjN8PP74+N1NthyNPaxYlsbUC8Cqq/tytED0UWMwEIsQwRDj5BkokB84
Q3FQhp3c0y/D3/JcpAe/Z50ciUNfe6p5gNCbyM1dtuJNjXOLiDYvcmBjsm3+YQ547S5rjjTESztD
ywjZVm8HzmSL7deyVOV8OTX28E83yWHObJbqOh5st427l1NR41fjh1wVBeKAf7RkJUXNkeb7eIe3
Lr11TX73SOYA20gUkxDXuI8p6KJiY+E6ntqMMKqL22IPJ2T/bR6xibKRL+veLLS1cm0N/pm01Nhn
rUPcuJi15hIcxno8mCBmcpLKajTODnLa3ZbrtaAWB4g2pWk1AvzTdM4aBkKTyS3cQnCIpgNE3dMf
Fc/ftjIsW/vY4H89SGT/U83JFPb0M8Rno/CWMEWmXxHgqI6WEshCO0WC3llEnmvvc1oMEU7PPfpq
6pNLcGDea1eHLN4SomenOK1VN0/Oa3xK8q+U/EiUg6QIh2Z15MuFzroUOWbsuFbG3aC/lfnGVL6d
m31h0xnfmx3GQn0LxtG7apdMbTZZ7LnlandC3HblrrCpGEuZowjB0UupT06fFhuE4Ogv9CtQRk6N
6UY1p392QqccVibyWLbG02dT1aVdlwxn1hWyUtyi6IOKXjIDMHGW+Ubyn4PP/aiWJ4UGlKc4eYHB
Yz8qcKm6bo9usev0wf6apT13cHUUq6nEG1XlIQSc4GjL/ZDG3fPVwE3/M/ntEuzVMf5YPNsIIeqN
WYG8WRyjYMJ/TOG85Pwxn7tTLxKEmqqfgmOGh3G3tt3PKU2TRg95WHBqm2yr/hTxfE5IO9xJzTHd
Jf3GvVU1dg/W91+mr11C1i37YXPVhuG+3M/386QRQEx41duRX9pfEthD6nWPPJ0eBFD4CgyE1VLE
vOxufZpq1MeGvKRa0YlFWph9HYqH1V4EgD/rjjNxvT+6bHZhHpjWuu0W8SIAGNFK3nVbV70YPJ06
TLfo6H9eYPdqN2j5TWFf3aPKxcrjEqvLyp3LUOw5NhGpGKdVZDA+ZMMs2rzHIZnTk0+J4fgD0m8D
eOhLML/2M4uFMxPHIv1FQdr0+MGhTAXIh9+SbqTRdsJA6doGhmYJTHPN0qPMNDnsvleus5WOUMts
RRqTP8fUhXyONxz69rPLki22q2P6bQ0BXzX4hit0kZQuUTvsVNMGeMo4+vEDXMR4+Ol4vxDjkFC0
9bcBN4roHJ/z/POyoIPDvyICGMv+uorULJDKmhTdofLQyxwYoHs0h1N4vLD6ChR/GXK5sBMX8WnT
d2rXzI8Q9IYZ0M3mAafW6kNb8XNJ+05oHucvcrmZUBMH947Af0ivm8dFvNsWZla2Kjp6m3YOQuSI
6yMemakRGOWdcgm7g9Tw56PqwOuePCeF3nHnqVyGspEoKIeXXnYFec6dE9CSoRe1RDLw6GHj+ij9
2hsGsxk4mppumQP/lMuY9471icf3KNFXlgR7dpAqryCBJhNfDKqT+zIj3Y+UqOsMH8VId/huPX6k
DouYPVHlJgy4Hr6Dy8t3LxRfz1+NqY8Wbw8ZgyxtzLN1UgqqY5j7OphDkTH4XGmdxsTZPIV0Dr2I
DQ9bLy00jnFNAJWmeoyIdncbS7fIC2n/mi18QTrzdJW3TlA00RinNBj3T/AKzB+bx4eIAenX2Roj
+Uxnhmd+XB4rTvqpTFpV26Wn2jZmQjLIuSjo7ZXeM5iszLdW07vCS507FFSx6qbSNNKoB22EWBt8
HNVvvLFcbnYJTAVYZfSuZ//tA3NWjSb5UoH66TDFpoXimKnxk8p7yDS+Qa4yAApRqoMmWPScLQ7I
bBEdcRKKfPYf/0aWrZJcwivOHLdC58Z4sYDTaxv+3NGqr6snijnAhMe9GwQP6DrA4R4JUb+WlWDz
JN1PRf1crwcyi2b8Z+/JSvdgKbGgiN8YSFGBY5FhNSj/fzDhPD2RlVQs0hF2/VKrN/69s2XLInVI
mAJW2/PIS/4nqOVCmbdiL8MQVxrtfLRrHaviYCgsM3y1bn+vUH5AUgePTdQb1ExomKIS1ksfGHwV
O4Lhd87mg3H9JKFpIps2haSzRDaY88V4NLM30cuv5mrrXAfzlphH8+MghrvejJUkK/AQrgj5I0q6
AvkbEPQI4V3mpCy2oAez2MJi8+jBEznpdKfn8jUXlwMivwqEFqt7UVRLX9RzAoYN2xCw+3GzVLIQ
xEw4ZFmDTdgcS6IwwNosibqcacH6qmhQCKs8DmvD3McbAik0P1J2RlsBxoWv5+3rX83kQIL7FM30
2ZFMwRr35q3rJGEk6fONjuOcpTDfF0biK0DwTGi5Bn63vwf7BBHCT3G70Ev9NPjwxzCUa/JDkw1g
YVee0zSR63LTmXGEgqD5NZKSM6gbB9VUNex86l9Uh+xVrnXYJIgH/CdQR4Q76FgS5Bw9xIz+fMc6
sNDyn3Xsv8mfw95aMtVmStlHTgRaMdQyqzjGDrmQ52mic87YxiqBh8yrXsNg/uy/rT5JhVd2vTN4
vk1hcn/iP1QveoZjVQWDhotyVlFLv8jfecKH0x36k0HUyJwdJ2aqBGaDbjpjAAAPnOXYI8im00Si
GDIPpr2EPn9m/H6wVRKArZHLZnU4FeHtM3FqiiFl53caYm8oZ52ZR9MQwmmAiA51V+06EoeNuV34
eTj3NLuEXEeQhotrHpLOExkh1xScA96z6ALOJD+6SPTRbVGAeTxO9qoHXw+SX6f+7mWBdzPl8GN8
Tqhzi+bFkD7fX6n8hqi6TZM0KkFDOxi39MGhJJYBjgbxDy4B9AKhFxMISixh2Rg6GKaJzA34xok6
mkNmUtZIQl9kEmgrBXpWoNRxTafjuHIxXls+OTcudKW57/b/lWee0ZWTMS9t9cgmjXANNNF537eV
PPP+IPlk7EwK0LM45Ajh0wfuSX7D3TWBVqy29uvjVAl0qsrXKn53IhLTyCIuVaBQeiHDIyvWGWg5
e++0UJyW4chgK4oEgavQbgMWPYfZugH0PJ/wg90Bz6x4QOugTpX5f3BWKRpeh6oePSxH5rZjIASQ
lakP3/tjOWIbfI7fEm/zhFlT2VfXJV7I5BLI6uPWtL3W0SDpoleIhseCwIyWMillpcyrz1HHgo0+
TNEz+oBmmJ/nqmLH2YJPmIQV3P3f20rFjA/udy60tCW1IJSY5DkZ9IAlNnUtHDNa5HafI4AFSXxa
4EPjOG9XYa8dLYjLGrhrfYQLOT2RcwSunva6fmcLUT6m4FitRBl8oDF3GYQo74REOH7fEKeIDP/P
XKpL8ByYV9cxtjPi96gWFi4YL7P2n6JKTJkWE1IkwkfhfaZMg6ALU71go5PLRcUdANYAetrQ8cXj
YEqFvgzdZh655K66GSa8Z11QWYLkhs/k2LaDyXpouMNWzvA31QBf5kvfqomF9QtI4avNxJHc0DFF
yXisk2Jb2+z3gghhLydtaT9RxcKDOlmP/DpE8gqZgeRbIEdw/7qH2bgD68jqbdN/Zj29YerXNNHT
2aY89aFJWpf2wgdoutm47QbrFdKCYNW/NiPpcl+GMZ8NfP/+hJM5j3iCtCbkRS4jrb1tismb6+FR
TRKHFfbmoXmXZMncs2o/rm94stTH1ccUOzLN/ApkT0kBvGMNJLiVQ3qEXVEWoF/ZbE+9jOasFuxs
JtRBzJviE4eunxE2YWnjOHx0yhmY8cbZU7gnetZa50CFn6VWWmzbayXyNLZUbF04MLVw7X5Rwrz4
quqT+2bu/3/SyKgZlMSK8NUukS9wwq3zfdLTyXrNZrb4CYn3Wwv52VMIXOoCBXtmWrvA3EkJ55s4
Ma1g4zNIh9paucnQd/6Dyh0uYphapLjCPcWIOowqHEEJHBe9LwuHaqVFc3bbCOEYPdeQphpJKhyu
vVtq4dB3sD1ppHx1YDe7oFWGQxmazYX5Ig7SPNEIrOWvmqv1v4I9HJQD0qDeHh8uq3Xsz2zjyB+N
PDiOm9Dsz7eHewpRQz9dumKljLwp/QSlkaf6+q+A9hIXdAZ2qgGmQmNKhDgYjdtSWfEtF9iBw/Gr
6jvJJvpCUCOMQDfLO6Fs3t588Wqlb6npQbnpFZnIAxqIKvN75FG5whau0M+NC/eQ3GAYQ7JwUjyo
OomwUI4em93zaiiKX9hx8w0rZQmyymp5xmrJ772QS2Ag5eGKe08z2FhNjFbDqrGxcMuE3kkCCMTw
bMLhNFegCuFGbkrAyU4+sT/YXlSy+DyY7eerXJl9rGWzva+IP/ThGOUnTgMKzXrg0mGvJ+9HNl5b
QqqwVo+PXkWoJzH8ycS4beVIhzs0EbpJG4uPrdxWVfr7KUE3hqIWmDwbzQrE/yFukbDLFSQWiWLw
4pd69PLaTil0Jzz7z3Ea6RafPYx22MOkDZhZNXp3QLeh3Vevd7HVQeCZZAhCv34DGfgPN3+84azc
QhlTBKGJboElKcmOkFcxSTvTjrkQpPQ5qhLLkoTiXmyncwoySm578PniO2jPueeKV8/ewfByutI/
7yfc+7Eqn64XwQW1HiHkca4I+9rli1LMnKBMzBNa43mhD5dsAsZQSyBCxJZi7B9xN2eoTwS8dtkm
mr+tX3BRXOPhsyL2SODTusmxS6P671erVA61th3WcJUZF2yhyopjgwGRajoEUE2TQ6XTMVdcM2vH
nguo4Z0xqS1yVpLuiXB4DV5NYneb55uEV/Sht3AxvFO/CN0e8cOtjlTyCGMTdECB5h1L8GLtIaSb
Z2C7xUn/1XTEINcBRM6cNvhTUfrC8bqioWlneL4swouBcuZrJ6bnkU63khj9/QwsXJh5uuhwbRJ2
Iv0CDy+hd2L98f06bR57uu6nDM63iXBCSUBjKPU9EotGEj82PJP+lgy0C6tm+K8enr48M6BaUJmB
xgABohVh0gDbS0a5I9msgeB2g8D81YCOMGehxPT7s1otyhTeZo0P6AerpCPi0YEUsE2HWjuPosmK
kc9Uv9lWd28WM4kE1pyndK1xu+xQEJxHOa2OF/VQRmy0bhwXdo9vxQAtQuKz07brWW4NQ9b6s411
9q6RZks2llxCitauYCElU++qFrBcvtU6jothvI8jTVs0Ruy1o7M0ii9Sif4jFL1X3c6fovTH+4Oi
XW6x0DXjEPyowOyTNtxNfOKtWB67jhKdcZ75GEy1CK3cp/WFtuQamW6QZ2uQsW6oZStZpPIrqf2C
gaA0qkpLeuOjf9B9GLgro2ufAoHll7BM7pQ1g8g2ktR6bLretzJyu52cLvqmHASrRdbsjcYFpGv8
fkkP2egqSaTd3ymvRIHtFsNPvshdvHtW/zkEmqhpiyfO9OWiohroSmGema2Ie2pGFHu3peYw81zb
5ncfQPA/7YZic3YE7I/fGiPlSvW6dqPgsj3FqocFC4TcaQR2U52k6f1nLfYHVN7sF/xXSe48GTqg
ilCc5aA7NneFYeUxYOouvQnVZdyMdD05B2iKYZd4vXGef7EwHmOh0OLngVwFj1ZVetn4CXrh+cN0
PctnqJU61QOy9WkDU07DrEG/iwdWzn9tBKO0VP2yD5PL9LRPDhqC7euJoOZudSvS9B1MHPoyZXy/
S00zXHatc/j1GhvXs+28ZWWwc28aRMREIEQ6l18dyEt3MsP6B7TepQ8VCMQCKp2E9xQROTPLlo9Q
Uq9V6aeZqlQSha6yLAJTEUFs2cU+Rt2QMSzM7Zg9b+jHN/AF7LQ0sy2hhWMi3XLhKIAaDYSHzyaw
PkHCEWYnv7zUAlfOHYSLbDBOQX4a3ZXauaSDD+dXJkxM3QrN/OtT780jiyEGIfyP+tNg4fkujmsc
4vmTEuksyVl2VnykVTyS/pHsHXE2+atg6N1mcSuOFJz1Sg1YywtaVHcmHk5e0qA7bxLm7A7LTuqS
01JwAE2lafOthmmACUGqa6NWBkrENCu7rN0O98Bs+PRa8Ra+vGXCi945DyKZBNbsWne/dJlceW2A
TVIb9uS6Bj6LjfrN7n50kw8yO1VZZ/grEZyzTASnG6Q3jZ8jRr3nmOil/50asE5EqC7Q3ZTOkejI
K5UfFVXJAVr3PyO3jtA5by3/MFFwuon3jGwv9K3/J1McjyfmNVfTYCNKp5KQkNOveQyliQ1PLIkT
7ZO4x1Pv/TpMVdZl3J8OuGX/pa4M93G098WMTRYzcqUiRzE22JKh4AWvWJvZBm5aLpuVbzUIDGhe
Se9df0ovDoLthMUiTEN1cPhHg1gQBIKp/pNA/D1ZHSmA4vWHW6yAyaD4ZiU0on877XQU851of3hP
m2p8zZvnKbazbeCoJmS834tbdTxmFxfoboXsjJvr7Gfz6/97LzycvJIjhRTudko1WGyVHE9vd29+
Kt3P5Gc5YEZagbZHfgMsSMAJYiaujRnNAjLU0am1KWkCRbkzJm3j8YpBPngAqqneA9Tomh+F1qva
5lKViMftFl8ZzWkmT0uYaJvrnMqqWbUWABcR3k2/pleqqayJXMzmefoCqGxUCg614tSgrh5zOFPa
H1trzEi7LsPF52AmZHcWDseVQ6lc9uiRgan89birNnDDpJ3Z/PTIiQ9Y7xmR7ytIvsBNu/BR0iCI
Tjmyhl1y5GSIuUY517eZoF9xH6Uu+kh0IZbe2BaMl3LfJ/chHWOhDi+KH0hoLlGlqmAJ2y+G9GyF
68G7h9dy++aQh450cKqo+N2hL1vMETHPa62tiMCEu5wrc3YZ1bb8mHfbPTBCzZjwHNftVG+K/CLR
dM4+u+R2bl+ZxPi3/KzcFsczW/2nhS75Wxako39LvUZKFCHLpeD3XVuxj4jb3OpgBrORB7WJ4abS
GvEKt00S18eKtds3BmxdQN5q2GUIsIYWihmptbp6dg8NqtWP+59//SVYIz8TkLfg8SpzO/6lycgp
FAiSLj59pxme4+tIhQ7JH9m0qac4jk8s6Cd0QEL2y6KyHc85BUdrK/+XKDwZiF4ljZVjAr7ruILw
9ead1TFg4mpBwPalNMZjcRVxXItTB7kAXDCJOmS/jIZqG3vqXgvFO0ENEMXUGsVPil4Py68HQqBn
gA3Ws6v2VXls5FDzUXAMHQoSVk0kd+GsD6F9tG3bEFzWggmd7hxZHOWZO0VyUUngZGtFqqDruDSs
M6RmC9whXmJ/h6Rjb+4TynnYT3ltG7Ex+IzPC95b9A1mcT4BafXJkC9jSmmntju+RQuqmS++yXlZ
y8eMYox69tqkpgfmqoo2/+LxrvIUpr0bLrkJGk3bYkLag/yJkEYd/pCkn5hu/mwAAvLIE1GiwreC
pYMYp3Q+lwlfBTfLzO2eZ6ZboH7CM9K39l+4auZr+Yd7wRRbvwEp/e1C9pUgBiqS5ppDjZaiGAiV
IiX7ZLVcL3P2RKJgSu/nukWhsVYBwenO3eS+LrL8YbAF6qjWHLKaFGknJTDaClungVJdDDiOJdFK
NHxpgZQ9+6IMQE+zUbtyNcavBw4XCj6fNnZg1KK+QIudKqsdVN6qvfrZviKuCyXdyQvCzWC38/x0
QY4dquRuPi6l0W4tIGc0kkY4afdA06ycwQNqeolpL+XvYFFiUlmI20B3RLUo3OtP5nP3LsfYsjzR
hUt1tgDQWdVCcz+gZszztmmfuIZUIlYVarc3lvcMahXSlfYStqIXQJrXRhRVI0XAT13uoundoUIu
X82na8gYUILJ2F0KJl2q6j6CAClJ8iLKHX4TMTe8rmitxlfkySWL4z/GtBfhYDVtcnxleoaZMBsc
m5ahWHpOpSoOxCAXcYkOAipHtZh1yuLvEIrH9RM9bDdlSBg3j83tRaoQmgxpHDGOsTr3oEqY0Zdc
GnvVZGXbOHVIUREbDhVaqxYvlpOAUW06y+fMSBmEWjpc2BV6WuUKBvfef/Tj3bJIeWr6DkcE/xEp
A2wfy9WZKsNu08QyfChsPVFk9Ol7cB323xkeLPkrcW/8ztWZheIbcVHX7DPwp6eCI5OX4ez5G66f
HIkQ+dt+6VU4/SKCnCgaG9uSkn6HAhL+0DjCfh1jck+ZRJeSYcPjOjsDmtscXBKMSqkACqHOZrZt
JSljFSwMQkzdIZHwmJDzNF9RubxVl8oKJCAHfawUYUnWK4XMZSkTa/dGnnv+mys5nYuIm+X5TTeN
MDhthaFYzoI6cvrJF1+jqtetDRjn46IuifKNV01RmxxCJ+IpbpRm/V8KTLFJY3hkp+tKtQH0gLPH
KzgMStDwdbde33727jI7KRtexITfLx8sMDVtB+lgAo45NtcId2ZhJ5//f7gl9kp5hDVS8kKlxTgB
dFtSSLE956AMJ97kfc6PZ3tP7NGJvm+jG0YaBQrmSYiLM0yqCSO37sk9aTbVjNYceyvgFH3xv4el
n2EScPCPHRBU2eebV8eq6thV0TZmp1s3Pm1Z5Uyqd0Tf3TguhJfCeOI37kbVahVPcoej33Ec6+rt
uNSy1N9+01ywicxUwvmVKycH1C9N2Cl19Jo1qjgCohsCJ6uOgD7u+wjsGPv0oHi+lB41dYNn+9Ci
Fm0/5UmK5y9w6ZYZDL0EB0kfdRCOcVrcNEpG8BKwMAxM2ki4Q6E8OMJ/lWq7QbcdOxTPuY8B407B
aqhOZjI5rOoPhJ5K/b04s4URP+8um+UIF5IuRjUXpI79Kv9GUrC5okQDHjcBFxaJLWktjzeeWM+U
YG2MbpVFrOBnoDnQYtYwdgnGxZjbwviJlySLuFiPOx8+BqVzcjacQmyUtn76dWODp9GcEcusUbAG
nJmHkH7qzDZlEcrqIIU8Wpg0YYanHiZdCUnyqQY1slAEjc1NcUdQIpkLcD+qIUUZbRN9GKKZXc+A
fE2dg72zHYh+qTnRvHqJi9hijrboHrRC+TzsHYy+8f59HAMi133eZIWQHJUjNtHJ9zKdaabKZ6wq
ROUXw6UL0/DionRGY3Ed/MCDWq1PwxXKGy5AFfJN9BCVdMHRvSGq2KcioBjrZJ6mqOFuaedvN/GK
pWQ0SlKER2MEFFjBT9TGD1V03bWjd2XHOpZb2feMDXMwVBIeVvMy7jB0lY76yTB3CTsdROaq4j0e
ItOFPPQNywngGF/aLz719NM5nyjDUq/IS1f1BfG2S90RTKfTlOKGAA1rRAwJ1hWfRoC/EA+jH1uc
ZpT4kFpT2xfE33U3MpMlwvQWqbUwQGK6kSQQaU3UCVO2KzieIBSMb5r1JXM4LQOyTp1uR6TECxqd
6EAwm95bfimuKC1XXkz/ZQxO+RqF88n87EDtSba+rnPK3KQB0MwqcWidNQkXGv7SHCQ1saxz9wvu
BWv5r/KzXTWnVGgXTFs+Jsop+wcUcxXxZ7L/nY34HWy+TD8EOk0T+3sJOhyArIvFeziT+U6/MIeD
46yuu9D5RyoRRSfwykIpS0IK79C+y3wDvO0HMRSEXQancu8E9DNRL+10CYSEOZ2heTR7tZwbzLAE
mbF4gxd1S392sGXlmn7TziUYBW7CDX8ivFRtW44+N04ylRI9DmfCaWukJ0ncb/9CUI4wyi7lsr8A
vYIx9qPoPp84C8L1mXl6stUMBQaBgZ+X5T+4XQ4z4oUgQdylfXRmQ3lNGzbAMM21criuAkXf69S1
tD0Ch1XHAXOH+b9kfXFfYwwxMqeLRCsSLQDDZlR8E9CQioPrFUWQm2KClTXge5PRS/debzCI04RD
IN8+pockpN5m029jIM9ALi74Z7+mET2GQEhciV7UOh5OC1OmZCHtJEsUvIKIJY4+LrHEZfDfcXu+
pe1OqfABbJ/JQILB2XLFntIHkvVpduaRE5r6HOgeziDWaZXL+LWvhvAFhoj7oe4Fw4QnR/5mM6aD
1CELmtAmFjcygeoUIznu0ZgWHGJQzRouCgcLScjH5hCwpGEfVecr6fNyj6cq8wC6Qs4GBTOFKgIT
leCQevCrs0+Pe0bAUzoIpss2A29uQl6t0MUB9ioKJwYXxpSDBcQ0I2zCQWBzNEX4m3cL/kRQNbXR
R4vphg5aOPNbPlrjSN16aAGpbBXa/aIAY3/d7+jeaV84NfEEjncucIDlQD9v82zLgw/QFFdY+5iu
f6dEiCmbgKmjVy0veN/D53yux9AU+oo+rz35UnYl4DCO3rOgMfj6LDpK9WO9XUcYxodhvP6MgbAE
cc7E9MYkG9nwLUCVaSjQRpyAGyp4/QQ0StvIti3oO1gbBRRqwAv4FfHnBVigmEJseSMtEs5UdUp6
Wd/HNv0UIzO4wjfOZhXDlO/FhAXk6x6+ljAEVFIb9aLsDnVlJknFXGFUvtpLu53eQGRYW/U0e7Py
1Pc8A8ucnoX5HaQJcWFmeE0/m72WezsL9mjwTYBv+22ph1ntDP6eomk/EvXQ1aiuwEU5Y9zVm3Kn
j3t5pLPLsJJHzKCnBCc5DuPmV0QmskeZDpqPFifBSLVrgIsB8PiN6Fd+iXInybHWdtcCrBya3VNc
vEVx1MwUNw0Ik9L00jsxPS8CbhAHyhoKk7FvgmJm4N/Af9ONO4rMbhksFlrPPWVW0eQy6bt07g3h
IzBuoG5TRIEeYJdOIawOI7Um5BxDfVVDlzm9fClgCqWt3iS0+JR2D2lRrs00crcV1dG/nNGbf3rW
CLbMpejBcjeduH4nCZgITWkJseoPKgTxgSQh+nFXtG9YVUWoFzcEiOuHP9zRuUM/oJzN3LuSqoW7
VKFHwt+aHW4GVHEvo1YE1IInwPfZB3CadehvzPsQVYm44Vdu737Ko/6TC2HHelRUPw+kPGKbxY8s
VLQDwUnkse9lbEw+ne6JLP7QOdBb7M1sw8AgY1xB1zHANU1PJFneVyN8/62eaMM3Ch1Wh8Tb9hwU
aiAGRrwsOaJQ7J9HWgb5+fwlNJATa/gfy+PWnxgJlVrRvCfcarrd0O6eGj7/DitC5jXky2o1ZxFK
KjTZyHP28B+HJUkKRGsqrnQ0+DjvPBh8Uz6ELfb+cBsXcbKmVFA67q1wDs2sjruavNB80ada7Zk4
9iARssrgqcB12GQSdQNFVV6cT5UY0Tm0NjFxFbrjWrYMoBm5Wm1xkoYBI0QLf4I0L65xfGdL0PlX
aePxnYA2FwUqREnzQ4a/YTaVJ1/fMe6gUoKWYBqJDAsfctTXqQs0k3mydsUm6WNiVi7Kgjl5gKF3
7WWUs8qB3MKPLw2+kNCGXT4jPBcXUA3KUk9rGgdr1uVQYVZdM3WSBocjLdhluaTblPEyKCDmRHoP
o/pEz2wREE4kkZlC7UtDB+Sbc7a67PnBL9RGtlf8Iw9Wx63OHPgm8WWQj/SuE7SWsFE5W0GezZ5P
LV57iBBy9AnHQXlFYascAW+XzGqEY09eIT1OjLpr8WzKqrRkFpmVM1F1diNHRycTj+JLiK9a3Qgq
S+jx5o6Y0hyFt7FWc5BZUG0Fo21jfcctsSxw2GqCVO/eFlob8YHW8Kp7esro0wsPZKgQsC2veGgA
VxjD/HfXOUOLUufp8KJoGKFbryVp7bUnjGBvSPTsyx/vxqTMTFrHfbMm9DFE8EJqN9RZQvRz3g9Y
3N0fOeNzENz8Fnlflfh8ZIc6yEHhk+bxTEQ33mu7zej97NhzDk0axzyC1zbhoxnpTrSGMWTgpFoR
DzD6fAwE0Tf3NcWUPJHrpkXIfKyvfj2RXBQNK7qTKAJxsDSYVnZdxb4SmgXEry2pObmBSBp3Ti0f
3BGVuTyBPU8aTt3wOYP4vK65O0Ipl5rb0/Am89WDdIjW1B6nbY31tVaXNuGtxm2/SErp1VCDATDe
7dPQ9Qod7+qCVu4Gl9sw7Plr8IUeKxGrmvxDwGX0rp7fbKNVXwyUZCf4qhtQcmMlTF/wIWHr2Tos
N0nkkJ+kgUkakwSuBAqEE3QUZjP/yUXOOklOgulW66PStzYe+a7rAUGjVNHXpEEGMiMFrhzqVzYO
TIISWixMpPnxFGbAyWj1M3JpnYPR/0TFjd3TRfoeBick0JPgl6KHZ+PIV0w0WOnccBzEuLnOoTRG
IOosWAtGwldFwYp+Gse5T7e6nDEf6CuSx1u/VHa0Z/iPjKD93kDroLbEf/y7RQnjcUivBgPwzpy/
AZWZoRkotTdFWy8ZRRSiVr2ZC4UHuZh/Dabes0v0bimedvOw6/S1gv3dJr0GBbvoh88hbcVVL9ej
PZofW0xyp+T0q0YJmbF3lZEv8UY1UtcJPWL+SZXBaSXLVhKYBTF9o+ibrubkOGPVN+E3tYLwWwXD
5LY/x9h/8IKUWx22l1FSGIDq+02yFna4BwsYt+xXSCnyeiOu0iFMv7LzsMzYPtz31b3F3iINBZEh
IxAGNa0pLsw1iPU8l8aUnz53TQFEXgbliQ0Zioj8evKW/xQfoWjvCrHN8/V5WCdbJaSomfX9Lv20
bmwCviIzQiJdHW64u14gl35gbQ/koYeFmadTNFH66pDBgu9IocFfOHGpBqaWSsF+oBOX3j8Fx+OG
pgPjQUEYYTA3fk1eMuQfK7XrySG2bB5mkj7Ls44keBNJomD13R1hSQnIl9FNMVKkOsmDU3CsOBNO
A7vaqk40dPEaiWrppR/PMHsEFZRHnGyflhu4bXhDM2GMVY9kpC1XJNS/UtO8x+2skFhvS0d83YsI
0xq3VIhnvJ1J5/0HAO2NhZ9Hb2fCJRnIZec57GmPQT88wYDkoiRyjd4p3cVL36WSrbrqdoEbkfl4
OPCzOYoF54jrOkZsz6lm3kxdjLQyKSnDUezF3qR6m3ZBlZRiQVJF0AHV8VBdIIDTyKtWxqsiYXZR
q7FgDyrmnHdUoZIr0MV37Xxqaw8Vzqv52ktyY2pMXVmuKGirTIL4kGV7+2dO5PlpnaW0eLn6tp9S
Ab6ADasfl/v0Z/bddDQfOj8m1ALijM8HJCcWjPuxbZULIKLpGZ3nlUVqMj+Vak9AMlNYPkAGCVkf
d9gYne4IH50ooIDQZjy09vScf/YP/epNrRq3+dLQRThUSQo2Rsp/44FcxSTwnCmXE3b1dohU+ncQ
Zan/gCv/Ix2zzTgqkiKkSRU8JLBLusjLxJ6j1PuQgndtMcYpFcn37y8lxCe/L3NSVnwxtlrcouda
M+wezwFMgBpM/XyczoEW/YwvKAK5iH3Z9+uiiYM/wEr86Z02J62xsBDr3/eCkvhkMzMK4bP8ADBn
MziAJ82qd9ULIsi7AybQL56x7rhYqy/MkTOBd0nMqXkRJNakPaTpG+a7CEhXoZzRxqFN3QW9ij+Y
5axLUs85tD5hFx1J/LmECPIeJtqFhcV1KLbKe4Tka1kVkxcWHkZXY4rAiwkL60Ya7Az8gdClZnCZ
6N2W9ImJR4TQuwUe/ebcVBJO1oUlPAhebq5MICH/9YWJHG6IYD5sx9ZZS38RYCrhAF3F+T7NilRk
jUMNuFhKEl47zcuJmMxCQxYeKQRSwUMyYAg5OmHghsRM9r0PbzkAq67ufmqVZmGSJDRiBJxDIlZT
bftuC70cxsT9GlsByWzL2iOzBfyg/VmDM7s+b4lJbISrm4lbwTYb2CaGZ++S+yEbVOI6j0fmdjKh
H+BPDrDnY0FwVlE/Yrl9Qu17KOkF9OeucE9X0r/K5/O4f8n6MJGSfKosdzLe6UpIrFRtOMh/JD5u
9awdE/Ely5snKxcE9IOeyMvLWcnxCVhnCTtUVxjFzVcnyW5DlUOWK+nOXkECC7+n8TcldrvPW3HK
WzssbCFcAFTjaQXkmXcIOE7VLvIjeuaRJ1R4IE51kfjgbOjjoYSaKnYu5CNWEowmuffUB52OkfpZ
QI46zAiSt5eDRjzjBJq0DD8NCk0PHz+gEZQP2Ifz7mf/wgj6ivA3tmRUFg8m43dvsyIxFfXDbS2N
h2BDhUqHYrIXK3D717tobmwNCs2HbuVyoaLZouzLQuIIthWqCO8XSgg7IgTzwbVKD1QvC2F9Ax3b
UH+pu2px3+HrU+p/ZB+PB/NJCK412i86SMet9NH6nXiCcHuSbx1r1tSoT07P6LwaOs5JqkLPPx8B
jBAgXuHJlRZ0RzTfQ3svl5SvUb9vHjaeQaIiVNF1skvSdyEdzsRTZ6G3baIBK/ucWH6Nt2ALG7aL
C0cjAUQ9ZFe4xcJ3GI2ipI/BRKVVHnoqcyjMGDpxlofKZNApxKp1M+mexNjq1qompXAwIfMFsSPp
yk15UBJPzXai+WFkL5VMvlTIu07ir+m+pKrlvj6W/nstfsNz/COAkEJgssr/aKZpSbwxTauCQ2Kz
/fJdnZiz4tRjDcgl3A5v4AxaXbAClIGJlghWRYYofAxWa0FFjJFAiVfZLEhdZdTznD51omXJI7+n
fER1yqcqvZiAQD12fBElMQUpsQa3TghZb47JzTdVHSz7Rs1AlrKmKycrq1J1RbGBbCvUG2S9thqO
zAyPv0GKivt3Tjcl4UU/lgD1aBGBrWxCW1CgBUFaF40wOgTRaByy4I2WZ+uN2fW23TwwgR1Dyum+
aEX1iEWtrO62zJergtVQQZUDFnlzvrXSdo24sQti/jFv6faij0aVmWXtlp+fYjd/RN0PlWhocVYk
blNevB1EluZj3ERI59b+97LXyxYMfjRedWQQbS72K6/5H6cwmhRg3DcCUxzoYAifKQFXaNXsNWZT
HetkZmstZomHzeLj9IQw1dQgbl3gjmCaeVn3GRllyoJE8ROxOgI8fzFXPsOdP/CViJrYwk4vm4Bz
ZI533bqscW0vO5vQ1OB/cAZx0lNMAQjC2KGis07cNbsYDCJLEF5NO5SaGgwL15i3eH9AorF4KaDL
JYXHJo9TJbvDiLIF48mFdbl0bAsyclDDdGgXYafqDOPC8HBx38DGW/LmfGhwNtg0+ck83WCJ0PGi
YNcjkWj3b0ozJmdGhRcdPxgT2YjKb1H4JVxuYlmyXzOOmYaE6xAOC7ajYtYMwnJ+I/ee7rmY4W/+
1rXEuj9DXvRKEgjBjBT7ewdaJZ74d1hMyoYyZ7KFfhefoRJaCYR+kB32PrC4NDPNLcCtLlmUd3rz
0ii5rRWZvu8YBTvSHcQZR7Kn+G2zpzVzv3bjdPbNKNCwFaWT1nivmUTcqpRachx45+ULUOB51bEh
PSzYo7WUHyXy4vP9j0sltNAAXsVkhq2a4wYXhhrcgTmeOTfmqkSXS7f+XpCVI7asdhi8MztjtfIk
cGwHBpQjq7jTZIlitovclVkMZ4lDl3nQzmTqCoVmtV/yBEKI7r/1rmhCA371l6NIQ9r+9aFV73y4
E5OL0t4pCm0hyhitbrHOMckJF6xzihMwQt6gwVrL/IJLzZRTTJPijwPGghs+shmlie3kfPvt/pik
U/9L+YnDv8ohG3UfgLv58aSvUIV9zcu80YjXlRuHtwvZrO/eaKZGnqrEwem5Um+MU6dm87nGIjL2
ByuiVxCcN0X+kOy6SejiZDBTRUYmn1uX2a3jq/2HYvQA0ObaXZ/MXSVivS/PHlNF2VCTB9qaishX
5eqPEn+2FH8TOB0ZxEE0A0RMQ3gy04QvGsIqA2HVwArjolUwwCGZsrJpgwh0Cd9V1N8KBhsj7Lli
7hZ7HIPFvmPaTcSXl6/kxdCImYYsweTlssFi6JgksTVFVJPfMQqXWOCi1CxKbVn6KqWJ2YUBvhQ/
yzCUPQsKGUsvbibi04Y9vIK+5W5QPTDWnyUQBPaL/CiyORhkomy+k23MkbeTlO9Bo42huIv62oGB
hc6Oy8bkKeUBbcJeCpmFlAQohrtRdx66W6psD3sIaaydPyTAe4iEQr8INjsWRZlI5cjt6NVYncEX
tRv4aN01IQ38I3RCCPmL5v9EmSjaOTcZzzk0fU/wrMiElZLS49fonWOr8CMt1vVzuReavOdvgINz
Eifz24smNeVblTYmwJXIuqrqekTgPo3YykeN+mGCyzCmfZoFjFOM6apdo67btlTkUUIp9a3y1H8g
wnxIn6TqxeTFd8xSWwg43AuG+nkfj4dFi11Uypg5vqdF97WFRvzhQLlNWmO3mfHOqTwhn14KVlji
FChVoZy5hLRAZre/KuyI1UV6lvg2JCZmctfWbAz56bT3t+PZy5ER4DzY7zxT1+PS55KKjBqLcz5k
iBrd3GatUBXPWBnP02UCqz3swLVjWkAQ+nmNVWEu0QB3p4EIOW0M5ansO2oHPFwe0Ua2EUEQV+pI
za0RSYLFSC0+Eh/AlMeVIGwEZqPc4u2vGaXAFBSi8hHn9pEA59E8PXk0MwLWCvhfoTZ0TDFXbyDx
cNagQCF5+iMcBb5QG83bXbzPYofproyGhykzxANyf/5Wiq1uyuhlfa2AtjUWuIUq4xVil2YDjBh1
nEl/EME5m4itcMhtx3OHKxoKF1MX0hr32PYEe83Xvwk4Iou3nyQP4Gh2rIJw7+bvywjM/ygpbcAs
XprRa3WFr7sQB7s0WlIa/xpHdsyjn2kxjNgw4wNgIn+Jw8/MXdidZE7oRs0mKUUWTwylTPVzjKT9
xC6a4nT8uRKVM6NRk4a/Jr2+yl30zxgWmomMlueYUrt0MpBcu1FVbGDOYWRKgeuBqV1vrRTfr8r4
/CUPHUVCHBxDwZu3NnhZOl922ekK7Zu+/R5EFIhT3BAkXiiu2pRXsnFY9J4ri1UwAI5xfjk6eb3R
RNPM14g/vBYvNQruFY+aSah7t0EMSWdz4ZxOnd2I66BtaSnhrIJY1ECJ4MLtc3cWSpXeFjkh4SDR
qlDXqgj6GQI8PMtRR9//Tfs6q0XLUaout3/0L9myIl9vwe3s7HBglExu68brk7OZDlbjgCQmgjdX
H2xgHzEm4B6FkUakP3As7uHAFc+GoIc/XcLEDRn0E0nq4ew2AAZASMiLBwzy+rR/CtcxAy6m6EWh
lml9n9yuVf3qUbR5T0vYYVSCyvtpz7VHAA3pncX7Jn5ML8SXh43rYeFOSJG8N0OXkRQtDZtAFaPx
Oq4VURgRQz1qB0CSZwzIjea5JGufQc56zVz9Q6tS4zxd4heZzTmPSHEV5EwCxXMMRedRxgsm7kW3
6nNnpu155m1be0EmB5GkhMvUxTyBRIzGHPC/YzMk3hy8oHk8PvBhQXQnPFCHnJPe05Pupmbl17EU
ezuPxncIJP4cwKyheeNh2vc8Q3G6tHatiV1p8nmnWMwMtajqdcPOj/NvdngQiZXFob1AWITUXizu
Zl1yAy1iw1fCyXVILOGM8ejQXN1pqMz9XDy2XknOSzmBOV+BKNTn9niLJQxrOoABvJQo0WRFpw+L
y2Ajzed0b32zybS1XO/xCcGJRMW3Vibm9w/0WWMn/oBRv7/y9fUiP0Mtpb8S/3obU3bqnxAmkqt1
7jNoY/IL6OtcxJR+JAp4IRbSvr7OSSfXaObzRXvBcuIPlfgE/p/CeK01lkooYZPNVeTYOPOkr7n4
/RcWObMfkZcWq0x1NBVNg35AI6b4ecJHxiwfFm0PiGTQS96bx5t6eI21WPRyULT6jTa+5DEYjhtu
STShvm6a/PGs+wGaT/ByC8yzOq9KUIphJwauvdj7IMtGZUvZUHMP1ukKEU7Xw7WxOw04dyds2FB5
2hJmu1+YEKOQ6fQUEVej2yYBo9HqHRBD/XjeN/tu3dV1KFk9CEvJGjPs85tFh2qYMQoROdBMdTii
tKIq9SFUsE3d4lQw4kemOEzYAK9Y9DMcy5V+gGxSIKx7HYiRrGGo8xTksMuMWEEgPDd9kThman9I
u/gQxeq81HhiiO7SGJ95bgyHoVguMtZHy4oU+YkiXW3oBspiGHD4MptGePczOV0u4zWOAcaDF6jI
2mp6CuLF5TPco74n5U4vGEkGxWdpcYfcbWCy5fmyKtFjk56hp+Ukva2lJ5fVtytkwfGhRgagKl20
Yrbi1dQftJEC8O6aejcLJJBESwUi1q36ELsI89KTILVRkjyjSNLCYeqHw5SHkUk67+rZ8RDOT9nd
Bw1zLrlQBpgvvDI70iLz9rAyjgcWx7s6Ufpf8tc1Br7oRqOvbdfI/iwAxn0mAtBtmIpodquYwEI4
bMnELmupbBAGv+amDNYc5FXJoxOBmXfUpnUAurbaP2EM6VJbdZewZuCpBL0vM1DV72yCOX6+DhCg
B2Ux1QHKygcwfMdHTU34BdJ08LwCmI7dtoqyeaGsIZy6xx4WiKEG4EBxZ/U/F17JB+4aiHlXuLh7
BK9eveaH8XzvEWrC6m+vntkKdmxXhOhsaQDmCdPDPOJGlEHMysRLubVcGVk0heW8EtWDBJEc9EQb
1/Hc4uxmcTsALTxcuoG/s89Pa5W3URQRlIz2/3g7m1Kca2hjloFTHcctdr0IeSP/D6Qwi+m1MB0e
dLWnDiz4BSF0XEsJfnkk+oD1QZsinGGNgeEatIR82hyowo6qsO38ME48CVVlK9Us7g9rozlfB31H
XLwVYLG6M6TgYD2Wz+inqC5ModJlEhSQpSgK0b97FRRrllg0bcozf/vMRcpAJyCq8UNYrJs5S/zg
IA+E7Fh7XLydB7cvmQzCBAR04m2Qq9oW4nms8queexBfKRoW+7qJ/KjYdj6brHlwREuKp2WvlYZy
l1biLsGFOO9vO8PwYcwMVDIYxJ5dkj7ifogPkEMBdy4rXOaWq9E770vpvi8iri1kYt9PQSqX0El0
g3jHOeuiVyd+anBOJqpXfIpWQ3DD+kMAN9aaeKTPIXW5lE1BLj/SLXmgia6mW8GD3y/7PLzcilps
pBSBylR9Tf6ns/3zDE94kYa0zcCa0ZaDS9Pe9OSTCYlmehDNUIIDfvGvCtHr4HR4XMFFwuDdr84q
+ROUG7ExI+7PpBO0IDnOvlwFBWukHrbd1CQ9QmgXzdcB/SJJFEOQyXrYQoTbAtDwMjeWDV4rm100
jIDXOEfcYTpcJ0GVkMxGVZOOrUABzBmaOWXJczPRh4bMjM09sZ6BY/6Sci9MWOlqrJsuchFBjSs2
sc+byOE9xSQXIo9WtUGWVyHnli8ZU8jBEigOK4rtyq5Td02qo4ct7fboxItu8ZC14cQOFp5YG9AM
IsxLS+Vb10mh0LzXrlU93nrNKUPMJkQRDzZFnHITkSSGuCJ3wBNRYonDw3ClezEk7rO8oxdK4QZS
U2aKSRpPyTUuNudQIDm8bzylhcmcfGeM9MSrgxzQlMYixL341QrkwXEUJodZtNh2M0lLoxD1CLe/
cr0D8HanN1H8sfpl3eOmfwmjwF7QKR8mdwwLX3F5rVkur7OOp9uMmGuHoII1TQhk1L6sfnNQeTsN
EcqGlt20qEC4R+ivPhOfXjFyDtE05NdtHSPHviNR7c7nQNrjZrP0GLNJK+l4X/JkdT/SOAOvUekA
ouAMZfCT65pTFwTw82xOBZPGpae2m+jQXUJ+9aAnurmFWKabkEIQrmP04K0RSRZwttRU8LSK+eRL
Ve9GXzh3nOYLojGq4pAe0IpLDa7o2rJk4s67lJxWJYw8BfUJ7fJv4Cu+pLMc7ZAnXOYEoYPU85NR
qYNNqHX9CsoG/58ukcBXbCwwEhp8xxskecgen4T00Nn1BO04c9nybQ4LD77ScO1nYCRHQxkknHq0
Txh47Y+0F0CkBBPHT8b9cUSpIgGWQZXsifnfhDmxaMAUf3lV928mNXpqrQD+A6CkPYZnMuh1U5ce
Njs/WNCc9PeOT0pcrUaZf+IUUaOQO/I2yFxB/PxiJn9XzINtOq3AobeJ9Tj5IzD5dae0dUetIV0+
/N/lRNqzDj8w9sCSKLKiFPrFmVxOHN7B2HZh2a1gpc2Sl6Pu1siXAplklnRBo1abcP9wbSCoyxgo
dV1Dh5Nyu/WpR0FTR0lUYcWaxuSQYJIeZINt8e36AeysfyGgRHmxWwu1uzNeqxu73IFbzFlkpjZc
s9KvjrbuIzeY/iHv8X/vXckjfLFLMihH+VmyouClZUbd2+sJm5EoVYrk3qh7pCE1Cy17ZfXIztlt
Yufq3zW7kK7DTxjJeZo0BhhORundiTmtwCjej0LntgUaVYOS5MsVkDBEXXRHjwlchowNavrszUnX
3W+K5AnqMmjT0NuJkAWePYNPJBdo+3kQZQfobJxq4PaYadSxYZt1f1sAHAkJ36JBBXFVrOAf0DK2
FtC4oei857X/N7rS9VYIviT2aw+O/r8oGSIJKId5AgrIjV/G/PpJTlU6CkF7pu151efNcsEvCyGV
Q3+1GQ50FdUf2bRBXJzbW2Wm4VIGEML+WPykMwnWURGGqz4vGTXZQAmaUrFBok0e4Wk8dBV7L0WE
BXpQcKgBPrPEOMOSVJBecWTyKxEZjAR9F68LjMtS5Tkn7ck1uj3mjh2HTgbhsn/w3FGojSuPKroQ
Gx8/tSGftXQfUp0J7gYAlIZRnMLT1aWJ8emSo7p3qcq0vgzdYARGdIVMHVU/xadNu/POTGlD8dJo
TUM4wS6bGIVfspngPGdIEM4mjaSRvTbCQ3WULRTzW1nrTN9tspH+NyWafmlnNJK1tozY/AsU2PRS
fyxWIiJOm9XHkmd3qMALtap8x9FDIxNh9bzL3pbTpJ5qzgIoqNimKIVgbHZrEyEerxOcX8F8HKEJ
Jo1eTU9PEhVB/B19qLUEIRgf4TylIrwkCv2m0JgZiUzvTB94UmP7lXDMA0ENjUCAJrKifYkTlCVg
cEd8AzfrXr9HEwD3URNj+9kx1Y1fpRUd9yraah3FgGdXm1B0MH7peuS3Skc0H/R+FRZBbA7pQrkp
S2Pg55A3+z+YkS1nDrUU82NJU+2qjN1BWZVZOfv4GABicpAQ0i7bjG7Qt+n10Q9TVccVsZf5KMN4
R89/TFvjg7Hn00IXTeeQ581W0A3TBNzxZ6sBgeKldvWCfoNo+8UETBNjktnmPfY3OKbTgzkfMK4d
FSGApAdDxTkV6hBbEWGK8DZwvLTYDnos7X78bew0z0QJeBAeSNkmzWqCTQmCtRoPmRu/uzXHTPQE
S0NxmuwDdh4uURni+I1I8EUfEuR0v5biIS0P29K+HYI6mUQA1gxavMNhXw+qLRD4qGwkf9EcksPW
SMJm3voqlaLH0bIH8MK53VIyO7rkFm3/fUZut/pVRq8rHMXT99m5behGoMNmoBLlK45E+66qthIr
KEjWsPiw1Pm/cewVIz9zQ+8yB2JPp/3I/Wg1RknA6NaYRGfDst2tNerZzvB/2bL6jAFSeOMIPyh7
I21PmG/WkA4IobHO24F4qeq/jzsr050/suMGOiYedeslHQsbk1TZg3T91tRv6CkzMYoF39QPpeei
g8OPyf3rwpuFhNvSjL/4L7TIhT9dGpAq+RHs/I7saegO3aCR1uAK0xZ/+MLYHvWQQqrttPeJxJRH
/+TL6IJQkrXEPePQ91xh2UGUOOgf3gEdygW5heBuiVsB6hpIScP04s+orl5ngLS9Q/xVW7jvoHYO
RHuy4QgTgjFu7RlVceEOqgvojoEJe5x8aOeusvGa9zn8Lrya1yNFnxbE1FDOM4tpkKLBVds6Qp07
lRtB/qaqpEbNPEEhAsqdCunBKV04a3BPsu7cy9YFYxuj+N+JoXBsa57EUY7oZWjpb6Th2l3FTMPF
3nUGPD6hEwHxvNug1Vz8hzKOxB6VWTXittXUzquOdLjrKMXpA5fjxUFsiKXizj52lVp+Y8MUeLw+
Obyai2TQcCKqYJ7VwhDgWd0G7aGpf7vBgX9kyWnnJN4gX+N7r3or9IX1bByRwF2onos+v1KpyfxT
2gVwwfNYOS5YE21Fwjg4i8HuEI4RcAssy2Jtv6Sc9plsC19pKp1C2wvVPB6FPQ62BrhEAlp1ixvu
Sgk4rti/2Ij8cXcS7i1J8mXBiCji6M8no7j4KgHLli93jdppLpwwiNpQ2nXyISgDdrpBVBIP3R8l
PuU4BcgnF7beBkeS7C9R6IrbNoFYfgkrBVhBW23opAe02VnAvXj4KUq5C3p0xwCwjf/Z1T36R4c6
FDyzWx5LHMPCN5tiwGpmAtyz9NaN4jlMJKRN1V2p0TlFJHFs1cYba6kxBWS4X5ZQ3s6wOYtTMSpX
JFUYNb6FqudZQOjnifJRvx68SqZl8x8puUB8uCSGaLWqAjbLmekjXpXq0dYDPTL4IeMvnlje+2BL
t3uxFiUWvfrtW/FXcAAXpxZJLWqox9HyRzqx7P7hikD+lD95OCblaOoHuaVNntlYmu2Nj8He9taT
e9mvG+KLeoC/1zViRLd+DCSRWy6tU1IZCmXo3tGPacXRq1Yq9RaDtfG0T1tb3DOSvXCcemmxn5Y2
Xp842aGeOkSFLl9033Ak4jLuOL4/nQjykrPKEHaWkWIGXnS8zKA/LbiQWDv+ENHaORxLb8Th2Ke9
hGbqq3xBgLdPbNEVrctcJsFeGx0D+1GG0ADMFYKSJJxewOXPYrz/8WyXRbu6yX6MyBx0EeSnkRrI
b+infLx/r2ksJ8bKqkZ4k+jAF3mWGLQA5aDvIRa3hM8bEQ/rZVchZiaAt/O9CXGzZyF7IFokWzO+
lw4M3uXmfPndBYB9TEncrXCIY+MmGh4grxcpIiPO0WRgQ4vFy7M1qP/2IlYND7tgdyEeX/mmZO7/
cKS1lM0F3nF8OziEawl88wQ6iZ9ly138wq5oBI41sYgul1xS5lcq/MLGzMYY4aghHyxtTi3EwW/e
g7EZfNIQzKTSzZOzYly6E7xCHnZl5Tc+sibtdGe9swLVlly9noLb9jhU9lMdS7sQupacfxq1ke6l
g4sYRkIVGyo6rN1ql9X+gUHf1LAzJ7aAsUMJgaVY0zXfIugGKNMp0xHkQKn0XrR/kmofqWfJwiSO
eclgqVXE5hJATiye/1Ba3XwsO5D+CFrxCOXJcI7ERLAam+eHMLUb0cZ0GgEX98SIGnzs/+haUn48
bxdyIGO+pXRdiVlQ8mqHO+FIrv7yCBUjAs2BmWbAfLdqM+7xGxuaQCOE/jD1HqaQCQeB4nK9JlZQ
FqGeSt+2eI3S/aqhPs91FCx1+YKIes5fprLunCKXLtPm/LfFlIItd7rmYA5fPogLEXXfzFAt45eb
fFhRN00aHz0+cY48aTURbdlh9jUvJfDpM9VWHiwZ4ZeWYG5PJQ+sNJmKHKHPGVj31zGycDOb/6pa
Em6hFYqeCZvKilX9iCbZYqoS2sZU48tW7XKwDkWWxabkykx/sIxc60egpkYeL0D1+gyEqCsvU0Z9
Rt05+fVWq3WAkELHqFQrIy5XTH3/qJ3AULLgn+ZEnfZ53INFsCnzP/h+2zLC4zQKFFa2uba7URGr
CDYL3vQm8KREFLE75VWrIroKJ+5uYC89ZdGZKhBGPhTVEWYM+9kad/llJZluLvnR/EJU+83U9+Lc
XVOzPgcIOSZOcQXV1oAM3TCbXwNHpLdoLslBHamNlLKkS6S1HC38M/sLTO2r6QBJQcsdyvtw54Mn
w/magtuGR1qQ715X92NcYJh2iQPen52Y9BO3tRhE3cszsnqrntUDxh40aVwQ58vEKz2qi4SIYwHF
jz+Cjog+FT0jCe+Geaui312VGccPvd1Y15y2YxVUuVpD4fAWrex/CWysVdypsGJK14MuOeyg4p1u
4LKwIxJMu00uKB3k6FlNLGDr8PC713p21xaiNzzqfKAxOwytM1KtTuABazegsE1JwWqJkQa8T8BG
i5KSxiPZHMrEHc/R/yndqDJFfezbNdkDuEp4+r+ZxE6MRIz1lruzRCjOP9iZT+MtWG48ZBCnB5aO
ZXKYfwQLAAZHcU/jBLBD4auxU3J62zeUSEFHQlXICnrauBBQz//uHD4e1dZUQfmHZXvN37/H05ow
jw4aq6u2RiNPHi0r1fN3nFUwZF3BmZvHyrsJU7K93buXK8281dmMiCZtdOfotBYp3m/O0/RwLt7A
cFp84RWm1sbONTnLPo7IIAv2c4ThuvOgwgL4bJpWeT8sM61TZ8jne+HZi0zUlOiZDXimyVUQbmvj
SmB2hygxtkJfaMeL5kyfK+ArdUa5lrSD0BloFNfZ23avdmFJ3ljaFVnEx+O2ZFRN/bySrGkgdR3j
3eELPeXy1R8J/9bK6hMP63jjtzJi20WtPvkwpA5vXL07bJvWyJLd1JKx3tT8ZmGjQ+T/LTaYSRyF
oKVt5uAyvrmIGYq6DbRreuo+6U8DajvlwrkCcG0pnQsjL7ORpLyz9UBce4yJ6ogIyevQZsRJj5hb
pfyOVBjbsgi8NYi3VpmUk4PL13sqFMRfOJ79nu4/PEp+IpPBkUtEOJ6wXRYE7ZO6y7C/NzB8CMx5
Zm17LFuw2JZvdXLfGM/gKaJPOI4IzWnPDjalbUD3YtbSxWX3c8fwoR/Qf7grxL50v4nseUTgkucM
8hUMvLxHUD+jZTfviWY44amyXFougy7tUf7pLvWf3QLh62TO3BJs+G26OEf+QjKQWI69gbOexxcL
O8Hj0nXOyjbHrOAD0ff4iOtT2t4FfhyrvCxjAAm9e5+2KvDxkpxcR1vF3T6+Lba/UCNgdPhkDoQS
qk1hWS1hGDKarN4Aj4U6FGv8p+3dfZRTogpZOVmr0vm+gg4MmjHa7/oDmxbycD+Zn3v2xO3PTfLQ
5/pC+mke3r64c0cCanixl3tnbFUz3dx3Hi9C+TUbQr3hULr4DpOV69wgctSNqViiDq5+CXWb4nlx
EEym48I7NZMIyqsmOX9xwDRU/pXmZ+hyRvSP5A8tKcNB0dP+qC8GZLIO6/09W4Ptx42g+lN8FBS+
fUczBTwfLzmcN3zJ4SwAEuKKm22mHMA2y5MtxrIDH43eKxD5hCdoWXfteS8Vks+EHwzyzbS77Alk
avYZIbutCM4dcAf4DqrC5WskT5NscSZbLD22g7KeDCdy5m2cCcPHKtpActjl8QdVVlx/Te3Q2FXg
XOKWKybFysQxgOHSByYqvNftMvVXGS3ntVabwLIxYBU9hLMa3CeZC/kyLLmmQwLAyQ1Gmicb2nCk
YIXE84RNgBBpp389jpPzmX7akEOjBf+2VmvV4TZhuAii6cwUiXMQa2rlBpfmX2M121G7TMvf8dZj
j8+twaKH39//FSc9MXDxo06H896Q/BQ1UtPq655xR7g+/LGwXoGrVtPEVeiKg6Z1nShWrvTGDES4
89Wjp+RGz6s+02je88O8RQMIP3DbfeLPpoKFgkLcPycZe4FDA1PFSV2V6Qe0CfljQ7dlzS7PToCo
QNr+WifIa9W6MQQB/HNEt3tcmo+ARjMAjK/0cFu0hXgPgFp5OlhgtEngENkkSN42taM4GA/8LAyz
nBJ2iWglf9T0KwxVudo3Uf7wZtth8rBNDJ6kG7ANXLWFFMrPCDxyMaKN/pVBqikTJ7gXQXWWMJTI
KwNGAJwJvtbGF0cqDTS+LOXvYnMoo+uOzDmxcMe5za/yWPjdyWeZaIdjS0YNSt8l1Xf7Kpkd7pSp
oMXBljku2njnnFDGzsKMKLWzbZrKGbAc+Usyx5QpCw75xZxWgjjAAmXoSWlBZUJOFD15qw02LT9o
Q9AhgXJBLNmVesaA0h+Tx0n9L7qLoEVGJ73/SM/xtqMR8ysJkLYQyvfgvskiry2Q15D/5/hxVypc
kI2KaMaBkwU3fyB5w7dBCIC9pQWugnqf3IOpZJaxJnVcAkTBDrmmeZ1aX6EJys+Bl3ifMIdmgwZD
kCMITMvh44JUOjkpCaIoKxMVQWNt5xLmVCwuXczPsftfF49P68CYFNy+uS6bI1W/ZzfE00JJRhRF
U/QFtTaj02IOzMSRRMcGXTTn2W6L14vo2Bl5YeKLEixqcO+EPloly6lultK6IRzWTvp3S7j2LI1S
PSWaoyTiDBensmYYK+ua9FB34No+Cos5i/S1zYicgPFtu1AtvrOWCFAaz79uSLwvYPBp6RCJYlQV
XjOzAHi1JbwzJDCqwWs7ZglHRCSVGp8dCEqhOkWcni61vhBrfLdgNtG/CVUFHXoKZgXrAuXwYhAp
trNlrP1NTdV10IxP8+B5uoxRAfAS4XuC2DPe6qs9Has4puBJdzss2XlXVRahrf1Z4p+Myb3hOfTU
GQrz6w4oy/mVsl2NKOu8RGm5dgoJ++UUuRxfNE713GocYaLMfumNIh3Wzm2dYFgAomwMfgs9qmnm
ZHJR/LaHAVg7s5H6IgV1l0nFyRovEN69gsPWs4n2G+3exuBT9JdT7Y/XbPric3tH0T11D3ow1+Jt
bPLpHl123R7uaz6Awe7qSvJoq8wf9Z1yLQ7Jdwsr9753I3z23ndlb1Bph/ylJ+tbN2dgN40lSr7+
ty4Cd8gTrQ/ajqjVTOS+MISBkUjOLRH4AmJ7dtr0+/sj5Mum+wUX9EK0jaI+6Gj8BSx9jfsioifC
geTiEAS77MF1Xk0LCM8nVlZUB/5zVMzKyoI9WpeGcRiNelSqSpM6ReQIMXReNtdm+i0av02GnWLG
cfXN/xprmmhSzDOk28IJkPsWxACo1vYxiEVmojmItjPy6Por7htcLNzvbltlYZvPu5RZpH9j0/XD
aE/oBfF1CQxcUZaUS9mddOri8J6fxHKcrnh9wefDp8XC5HLB5zir8JQ9o9HY9QUipLnY0WgOZzNF
l7cBtCFiovb8v+SJpEXLv+A5lWJq7owWpRuzsirnZcOqYCs6k0h3z9TExoWiE+b8zhB6v8zkOwHC
YAigLX+HgqmAOL/KBaDELaZSDGJUB5Dmwqah5ewjWTzea8NHpxRgtxuuahek9CNcRip+2lx7HW+c
+oNicaiuVVF34PiPYdzxi0fwCR5niQ8vgN/kDpsqC0AB1gDI/2VJLZI9OD+Fi+uMkbxBbHl2YAOV
3i4zzjSkecq1Ummmbnwg64MDwhPKzgPVlYBnRqwwHMccN8+P1VpqYzsTEBiOGyttUHGmsGmURdKn
kgGr4D9uHWjl7GmGV2s5XzRMof5UwvfH36HT4iWc35ZZKLU9KWF3LFxXE4JxAV5j7EUnjpQvC4fY
D+Y8Dbe1vv7Mnqbi1ZxRXgFb+2e+vQaec2ZAnDDKGwdn8v0F1iRGaGIqIy9RbEcabRvfhpepUhnt
0nhh/YI9J59W8Vgk2So2yqFtic2TgRtPipNJm8+2U2y6XXm47OPyz1hCbib7RRGuys7vf2uBdFXn
nsb00td05QAsaz4ZvYsS36PKUyweWLcIAsf/5rQMOTx8HEScugWW2hfYwozO1qlaCE9w3SzBEXUb
lcnPc8UdI2tDVI8M/wiCJxaCcJbfGWCFL8hPayERJfMgAwAk6ja1ZYwQnB2eoYh1hHo7cTktxroS
aoyWFXPYThkXjzVcujTbJlzb25N4Qx5O2DcKGWwhMdGBUQdrqL5Av/8s9aE9yySIJEt5AzYWvrQt
6ba+SiR8S7+Zwd8U8Johi8koUzl6ymFT75si8TGr65nfz44qg/eTeI/H66NRS3nbiLoCtHAiW+gm
dRkGnfBdWrfoRMtKkNZfhdFYqdDOCBmVQzb3Ivj7H3Y6bvogSCvj0e6pyt4dqWgTXCrV7zfnid2u
YhwgdUNHe7XVsE/R8IhmHLYvgvecZG8k2qAizd+Ppud54+sEfQTzv5W6hAwRfY3M2/VbzsU5ezZU
pkaoBVh0NmD5LvuVxnqkUuQjQIpi/iwjFIC/4vyn76ngxg8aroHcsjaYo97RxPZVdQ/3hhted27I
qL1cx/zUadTvx1K11upauxLlI0Oup5epSy+C8i8zpz4e38492Shl2Ue69JYbQFyg+dJuGx7eEIj4
calrzTY0yy6hVdQ0+detkMvAUEKktA0s/G0jXN+S+sMFq04TJs1pNObBSG4lrn0LrOOddomSqSb6
LTDwxqN/zJfFyK0kyag5P16Mkqw6yFrYDjjqTtkK4tJh3Ddo6z9V7wB3bRr4lF03WZ416nfzVT0J
U7/u1tg5aMeh0/9UE5jNY0n27X6ElOtKQ0wv7BnS1Xabjv9Al+tZtCzQ+z/c34udl8+4E1DeJYjW
2pMW37TKNsgyMasl67V6mSCfJD8P/NvqVtF91hewOfU0Eifj3KeSD0MtbUcJw6g1yfGU+R+EZAg0
4hl/bsYs1x7E1gmFLiIfz0pzZSKZJZN6mOMZgBOEjW7axxUD/Jwq708/w8Vc9ntc3RnLyv7HP9YB
1kp5gJsSwodEau8gXZKExgypUQKZWqVgS/ng1+KAJgsEEWxJgnVk2/AdG9kzy5UdtkIFMBi/Leqo
BHk8sWrFhlLlBB6YvXdJXUtGxHnITeyucqQPSrF4w961D3e1vQrhHPFzQggqMdoHKixUmrvgHGXy
46XRGpeXu1stJ8CDuWHM2nmjPwYzdtlHPaTQjoF//NX50dKydMdmN6xPtBYMlJm4jdwqjXkOU5dJ
mT3oYa9qjFFnMaVb8AuEpHJtAE9Xa6vVcmSfaoWLm0JnDnq/Tebl/DIp0ac7MLrK/eijVjlMNojA
BOmTbHrIWxsxiO35iaNcwtrVJTMEweI5XPCQqIwN5gTyqVaGpVjVPgzW81eof+1WfjMEAeon5O0a
QB3wt2JoSz3b+YL3PKsnoU+U07GuHJ2NA0+peZ3zl5YknMCsPiPHK62CGQF1rw7fgIM875yRnNIT
YUPG+0Z/HSxrRKrjfubflxNTAbwynUSEffAJ5i1m2cVtfXA8P2YJAiMVGnD3e8yift5HufBPn+bN
Q5UcJNLevqQKQ+UPmSzJ1NvxptPszEyMSR0ecT19BqijbDlqqE9u65MLAl1LODfCVSQSZypS/xft
w3ijexahPxwwuCHhhvdmgsYc4+Cow0tso+5bf/4bPBj+hcKpkCSY5e3aZjcA1hX62dqKY2cUjgpx
R2/2JulAk4almUXsTRgcwKOOLiKctAyt2trsyCxlPui4RGLhLgNe524dypAN7+JWSbPa9PGcqazn
RVaSgwP8B020p8KYZz/3/wDeqx+oqEV80GuCdDTiRye7V0XRtrO0KApjY+KVBd7yn9TUYPDtOFw9
rev5yGpSD5DAYDtQdq++kK47yYE65sziY1yTMH2BqXo35glw+VigQDhWOP5eLYqEmOQDbKdsyJOI
1gNbm5PMGS3vcPuwfcv8oNzXpk6osE+J/D/mKK8AZ2rCcl8aCR4xFvUCHFiZQ56GwhRxocK1EsDK
f4UszHmZssIv6BTmka/JrhfB6nFaMHLMbcYCe+t/Hw8mmQVAECVPaL5w6QJvFxIDCkFuhDsUvnsP
bMtT1nOUpf3rTuUkux2+SIF4yO1LivoyH2VSJXsiO91fpsqaBQ1CpKSwR2q+eiQaXdcfiatVao4t
/p9L8xdTIXxHQEmdaZb9xmujzQIndzcEbyVGeXIT3zZMizp1b/XmT+A87jK29+QnPqVdVARwzCF+
pHWP4XyW7y8evrm4UOAmf/iWc4lNR6dfkKOXn+cZkGCP/xJHftbcwwCatAyWRoqA4BoL9nzm3zTw
EgYf1iLR6NIrEBwTAytjeenCjuDTmD/UlG+37LEYzLjF0MiEoKMayX745MG6DZM0cbFdeCl6JX9Z
7VT8N1d1AI3TGoD5bV4ua9/BWZi98TItNp7o9XdBkm5KVbWVZIZfKMFbF1rcmP41P/ZhwrYVgXef
L8P0MDM4pD19Kch74JV4aANWJNZER7DMxjUJjUl5J+c9m6xljKDt/At3iz4Nux+db5a98eAvqcVf
eFEJygLP/QruvOyUzbgxi2vPXpY3zVPjTYxup/sxMF1PLhzN2QEQkUVJ655BkFtKqOZBv/hDgFDQ
NS0nvZP3dln6WP1xbtJejdk6dHfnnfTF1W088C3g3L3z0/yCQ6m+JmeFyAaDRalEfVp02MhfzbdP
kokdBiKxrimiT1olZStOVmTsFjvwV5zbM72VpmCk/UVXkHdrIytrFsU9ttxn202tpwcRjaeNh/rJ
5NsTxWGT9+UJFz8xYSlcgYjCbdbFUPgzOaQ6a4rwgXTJolY8CAgdspblf0NiJDGRJ78qD9qGoRgc
94eeZSk9zKDDbKzCy5DJJXqMVqwJDgMCSAeYzxu/tVvzJOsHicYtHz7IeHXHNf9Es8Rt1whyVygT
So531KIhm22V6ND6gHoze36brbPq4FeSTo1p7OcNwFPocdnJoCUXhieL2JGaOM6FBsWS48haesyZ
JPmSepMkdWvbLBJAkzCteof7lpo43SW4XFEzWB2zxbEYNlQzNhaOj3hkireTdybynMBB7asxrgpS
LIoRTPUMEuNcGhTmkO5V6X3mN7F9NTZ7tAvKKMxjalihfGacp5DyzQzYZt8DZwQMH6W7qmtgLmn8
d3G3QyDbMH1/01GUJl0ivN3tVrnDFfFHbs/iqjVdYTJpz+OjYqEKmncaUVo78xsaFmz4AXIZ3m2p
0znR5BKqk09/KI2L1n7ytOu4MEa0rmLbmabSev91pvvpDhDwJh8hQeVmilwYvEy3qTWAr3M70ocF
D27Oaih3FBwUd5HLirSwumrPmq+iaGBF1cC3CspZYmAeaKuW5Rih7IUbCnSjL4UlljesG62wylEQ
7+zpzAkvFPVgVSKhn3ZWF5zwL4Jyw1rOYLfoF4PyBatkQoWHMeslt+agFLMhbVkY/2mw6LDyO3HR
uHw/LEBWrTyp8Y5C4WyrVd/buzPGhqgphOjENANF+SoRJ7x+dXF4DJelmnCCaFKrhyjjBZix6WqL
fuejtrLKe0ClAAE6Ek+A9FQD6MDx4y6DHviqnTaPLxf57DU6/Sw9LjzldpLEcJUsbnRNqkpZt0aK
t/3NIDpdWJbPtGwOdheiRqEqYHaZx21xwe1AfiYvWNXzrlVZLrwCTlEkv1y/xx+roOguSbbs0ZGY
qJQgYeCI1BZpgN5w5Rof3i7nVRVlffLuX17v92AEzLf14SmOJo1TT11KSFi/nNUhrangWrfYyBG3
5MtlznB5ZAl25djkKKPkuo723CL4QyEKSd9tXZRjeKn/ZnLhlIJYFekC5p05jcDLNBpnSd86Fk2H
lE3dTCNywN5bnngfuWMBrXCNKyOo/hrZ+yxt6lY1FgSjKa9d2PL/bepVNvWtwM5POgxWPfTcE2b9
RY6ItoEjpcC97YWsTd5zv5xcRh8fyjsyRpGHDBVpM38yJIvWZerXb6vDXu82CXMeAcOBMs/TQR66
xmbXz3i+Ge7m34asReKHRVzCAoNLAlM2oBhi68sbeKtkTt64Hzkum99QuiP3Uhzvsb+on0tWaXFd
eCr3o9453azc6Gz6qPSebZnUkTjIxjlY+ECJHEQyt5lytkfBnJJZAlCJDROmitZMejU+gwGbKh/j
WpOPq4Re2QgFlygNUznpMXI8MyuCYmQQi1tEbfLXpr6wqY43AQstpMW1MxQlSkyHPWr8XwFDUm1O
h//3YRuWFwHXMnf3veStFuP+xS4A3iEdZQd8kuLE6FtE0ksr3TIWSuqvwmM8tIMjj+CBFSA+tTdd
IxY6LJCSizqIU7dAOUn1RJPnbeQ9KRP8md2ubxQqYcY7FMW/KqcgGE0kNg3eEIItoZnSBV+94e49
1ILUv3s2LZBdDpg5DJU8eP93vO+pyIwRWIVmTkqoMPghO8vlMZuJgGIkb1IE8E94rbFibry/u/y4
/v5UFNH/4obuuFrzpVVgDi78EmB4YZbhn1LthW394IitwMiDLdYTm/GFvRGg4rX+65oZfCZHGUbE
LNIiJHPB/X4c1EHBqPtgBJVUtAA7oXeND+LU9QVAV1oox42TxNaUJ516Uz2M+THB3eOERJEX31SO
DD7x/pXNcGgGHpy8QYvKHotOxzUe8zp1F77jrYRmn4+k1NpM8csUGLLFJtaBLsmvMxXLHVpvosgA
CE5mVvMtUPWuRfPvTsvQzbZPjwc8hWsFMlOi/xJI3D7YjfW9WzOKhPOfSf080MdH4v2CmVSiHj7Y
eBuvm6X/kIWTbCnzd+Djuf77iicixur3RPLFuED6oT8NsMfllbWF5/IdHOG9AqMknwKkzJmIYm+/
gTEKUVi5H3apB/ZxNKbkXbZiJElNBUzEd47MVSbMol13zj2HKtrqP3qR1vwbH1WDTtZGcb1GcS/m
kDgTKCOta/tp559/b38d8Kfa8poE/gfZCGWEbsrdM37yVaBrVnEfIdHA6bod1YUnTfnlHvLNtnR/
QhZApGjszHLtIqd/w7wiFze4hlXvtrBnKeWNoxEBKkBpuXgmfWq/9Fxwg9G4WnJAI14gBVSvFPeF
Yxm8aEfo7OAHQUVNwMflwLytVGIQeRPQI+93sJCo7HEEJBr9jJJnRtzil0pf93FovMoCUQ4ZvXsL
dVit/vGba4vniS9qu4PD34XHlcETyNAnbC0lQoy+oX1iGq0hWnxJFi7HaM9amlXWTE61SZ/0GC8X
FwQ/NRbszmJdL6lmqJSU4wGxzalTTWLC9JhtAtYEw7aaxdQ8EgX4aaOmnzgqUrIrNZxOYGtkOQW8
bF3iUbnW1YSjdCj88iw8EjWCLlShGTIbx4C0SW7m/WIuJWhVsyvsD9hEVrxbwUbU5tDJ/ZSkvpcD
quf84JutHHmN5eJDNrD1ANbR0bFNHEUk8W3RBviN3I7VGsEXVpj4PFsrone1VDj203oPf3xGSYBA
MPLDgGK04XcKchbHrF12wduJgVilMj6/oIrSzDjSRKee5ND9kAfOrlBT/6d/Pxf/hMJbQhlsAkf0
KNIMNHQ9IkrAOiEt6XBURcLpPcWUdaaqcEbuzL6r0d+MlxE7/jmHkYWV5QiA7EDxt1vJelSgirY4
29o8dtes4osOsVAxtetcioqvcbF4nAumLRrSISEF7tCZf9XjiTmtuJODWQskalmdf1He9hX+dt0E
0Dx8Kh4LQEvTz47u/r+b0HMphcrEgmYJmGv3QQpHPrL4/REZFha6Egk5dTxPnHcHzWP829HFy/2U
wmHs/CL6P/xK2fIhb3VMopfDaEEamRnvoiJA+uWWZAd8IDaWwjeGhGLojKTNZ3T51/mSSN5oLjOp
HZSjJ0KG1t/MvjYB7jV3SM116tFCGBhBsRojxuxx25I1iLINnd1ruLqiCnZTHXuvQ/b5Nf2Kl0GD
32CzwlYfGy316OWlUUybfmsYKBS0CQlA6wN+OYMetUs7T4YyLJ+7Xjbx1fRhXrX2DQRGHLzlwRj7
bb4LsHF5WJ4KaaDdilScX22nn90fc4+B95wIZGEa1WEmJhZHNvpkkiPgkEOhgPrBzoI5h0eCtyPM
+L4MOu9/Pi8f2wC5KDxZtNzEsNA8qK8xDcg+ezS3lW3Ou8Zr3L2dRMMlsdHM0uS0vcDbkCru6yH/
Dl8eaWwzET8HfxDIqnTUpSzvMMxpMayJ8LNXTyi40dq2ynbqsVbhAeTLtt71T/Ji9dsuCEyE3k75
y5EumCUpbcdFfZ1ly3LZg9AYbAYGRASH/Iygkt0DB9pDd9jRC4CXq1tAw0oUxx8uIDJflynKFJHA
oP+0UvsPsoaU87+kzQzCJP9DtOGe/e8Qx4GTTKCbK123UI5DM15i479xXfWITsenRQneYQo5Tx+B
+ayjxfAvVIM1KKQPkO6PXdM4ig6tImROsxTeFVcqA4Y2UpkpbvwWsRTYl7WWK61PkBoLDJrVBbB0
azR97mEDagNR5HbXiOVmsKTfYJP+d6yOlx1s7Y2ffLUrf66vCAQzrZFnBanh6iBFwK90oZXX5d7h
BfrUIJZMjAnO67kWpu34UfBguPxfD7coEvKoXz8crcregkjuZ7W9hL4Jypd44e9KchWY13YCQERr
gciLL/Ra+ZuGfNrL1m5hgHBHohy2e3RfSPD884POqhIDdc5VbsCGrq311XpXL2ciNBCZNXmtVupc
RHQfFp3zszZfn2u71zpOcSZmUIG/1FLl+Rz0Kp2uPnwploKbPN7z20M8MsfgknFzXAv9ckBwYQUq
6X2yJ2Jta7LzCeTLakJvXy6gI06VaxYBSF3aUitafSPOcRuda7wPPs8Ys8vrF7M/gnhNa8ngXlBp
5iAAi9F6KB9FgIhRJJVn8YhBkfz7VSQD6OaOVVF9nPZzDfkqMj+dWpfCuyDt+AREHvJudi9OrbRq
kM3MrORgotFr1zyB/dgHVnTEXCEB2nohBimzxqkDNfY3XGAU+HqhxZne7TiBrtBZCefCuc6MFUjN
uVLhiA2i+mko+KaWGTAJl5NDyZfD7ODQoU1lVKSY699Wrm9MdWOfG1Uz6JIPPrV56fb33g6Kigzd
lpNd0ZPswNrxopNffOxFy7FyLrmHursFV5I27dJeHPHqfUD7vAx8u2EUl+BE6AVcr0Y1o/OpUCXc
B4eL32Gni8nv2e3q1E3d2b/v7JBcRAxNyABBPKsj+qLAGeTAaNU+1HLa6Add78eEqzTgzH/WIjgv
Rt9xBctp5FVZ+MMQrpF3n78bcmIrvnZxCdEYsV7tRDU0X8j+UYoZIuM7S90hpGv6fbpl8Y/5r4Rr
4hAgDgFGLAyvLaA8uH7dcP8nIA1cTSncARCJI6lGP3OZn/4ZabhKeDK//UTXRTY1AuOIXepUhsQi
Fkkf43/Fxtqnn7OKnUwDjAWaMtE7SeYyPHT+5WMwFKk+J9e8ZyfBN5gkdouIMjuYt0QBn1YJEdTT
kfdNpEd+gmuuh0BHjSZPnLXj5r0ldfXL5NXkkmB84RZf4UZFYUNcRHB6zDBmVXH6n0nTUOJVPMnl
L3m9ncjZoG2WwZ83w0S/O4L3qrGcEGIYKyJaJG4dx7Ce5oE2jDt9Suz7x1LlIxmiDs4iTXOBjuIg
r/dFmImBxvAam+6XwjDPUz/NOXhGzvb1+zyZFlpcfEVY0gkNV+6AYD7dYUNY9lp0qtdKpnNXnd9l
5HHhreas0QSveabzyH3R74WXGbtAZR0U+GSzq7DogWjUbpkKuCEZ/bLL4C2xFSs//EpgZSKj9cT+
VBRIdM06xc3AZAD4H29wIhZTxVE1B70VZ9utTzOkLrk4DFlXj9uigcjDq6xMwRNyfvQB5ELWi7Fr
XS4mAdN+cPqwal1jhGyz5yD9EbuDKf/Yc9mvDtmZwBjBmqyBgSY6ZOGHUcQmjPiCSHsACEq4JkaW
ElvZFCtaWyVCGRasFGpCoTP0Uf7nT0DblgFbRTqqmVONC+hKc35uhlfv83FjepN2jzLthVEwO+Lr
iGAMaRTf7CnNqgM3jxcip2BvlemjSCxiOKdwCs/6opFVXI56FyPpmMa5OuTTClN6rlYkET4K3OXT
0c9VIUyHb4Y+gY6fzjgQgsP0GX03pLQMZpGLbc2M2/24t8xq84MO65r2WanRFuDI8hDXiY2eO324
O69GFXswacDCDyvRSVT6QMMvk4WYTQrdb9/mN0j+grHpp0Rd56zIs/t5Ve1mOQx2EqakChSTarQV
G+GSb1rVCrJ97a4hUTklffmN6CaZun2oPf5s0Vnz6P57qDgH4vZ6DdiOtC5ZRn+6ElNxGifhx1Sn
wlGv8T1II8+1lPqR7hwZGRrBDfBCyueTT+Jr3tgGyEezRCJN87JNjHgkP02nkHjX9FEsiL0hXPCg
XZcD/dHZx4JuBRXmRT457yLJS9Rx5rteOSlVfdaqqTsYi8LlT4zNsZN5MUndVtKf4eqWCqRscRP4
Fin1z4bcCD3UpVMuXzqBy3aEmoqpUvUSpkfa6mp94cilROGFsFgx9HHPRs/cIMr6zCJ+UJLZhdZm
Y80hOZKCAfmcGr5/lbyCTZ2AZUkelIEEuOyeqfOA6igkSIEMSUO9Hc6wDM0fhBj8aAA72dvcFU4C
8F8S22liB5WCfVpFDXaLIYis7rHdK/mMcplH1kLT+d50vawg9CCWz82jZhkUNZ+GM512ixpXwf88
NRfxkl9CrhT4trmyEA/PSvNCpGzareTgr1Ags151KdGzWJMKn2ds8fXYbh4tzkaMzfVCsAwdkkPW
dVyLNVk51W9dQqfySTUYlzGN35zz5bVtZD3jKgFf/V4NN4SE38CfyUYBaZAEPW+xy8UknWtCu/G1
3y7b023YuiQwHB+0ggfKghcolPudI3GDxawSeJ3a7YrAOsjSNcjR38peAAFyS0eYAcK375LAK+IB
2zIfx5MlgVFp5phpcKh8XEGjLTE6wx/trup3bvs2zcxuT3KknLi5jhJtaRo6+S7x/vU3Y/0TZ+s9
bF0Wzg8j0XZZh6ipFaWjwHz7a7vNsjoway9O4u3LBxOiSX61aDb18ZSObHdMUrTXCPh5iLYkwlWl
v+a+UbBgH+jdJ/kNH3dek6SKfyjbDyoWbNe8QPgwgPfOR3XU22sW5VcT0CkKwKmH/8Zwzcy65lo5
Mz24aF7j5Jjlvs1aQ5ZbmLkqAz5INDL3ao2rGw9tBZ3reJ83JsZsl1/j0Njj+HhqIpFTbioQedcu
kBDqHULF1/rQ6OpHlBqCX6vtYMDaLGxvn4u3egQ7gajTZEehy4zioSNXuiv2eE+Xq2bHuaEkSp9H
2aketYjOp76Klt3lIkr20Bw9BysbjMMNUvoVQoRaK7q3WeEMi8eM2VKvUDXQdIaKLl3etxUWl3Hr
L53QU4Clv8QPc5F+4kgcnBWhltySt5wcFolEAwHWr2mBQGNerWs1eTcGpafpz2xXNWVoKPcReBsn
XmZzm1LTp8RvkQwEVBOvzIjB8Vn1ywkad7VEJK1Jtpup+RY9eU7h61G0SC7o6UKkVI8KKUgX5Dfw
qNecC6ymQxyxJZXXjlKFSm+BAk/MKhw8FRgexYZZM+znCKmMQ+JezakuQbbI8tspNDnqnxadafrA
tOGA4XBmEI362RdOcV1/h8SaDqjF6ykjdIPrBUUYFsLv1GsYnicHhLeA/8X8rpUQwuq2NQUEnG5A
nrZvvaExWgFj+m18IiTWzoD55dVK9awHgE2ooNAdU0c2toQV1Vn1IhUhjFFDTQjCR4Nv1mWMcG3j
Be9O19/+CS15hsgEcyEjc/bL2PG71motP1BPidcdMubJEAJKeN8M+d0CxMe+h/04o+bnY+z1DKQO
o1ZtowfCmdkqPnnmuGUDipb7N6tIbjn85Bsh2nozB1tiEx+kIj7+YbocrNN/TPg/JS0lVoQdV5N3
Av1sOy2l6KAZmUkDQAyx3R7x0D3rFcDlkd9xNXAt3GTuvyOzhD7R/X58J6/kZrXXvGdrD7eST2xH
n8oBn0oQYwTqpQtHPu4Wk+0FdV/QzrJF3NhaIWEUVGXIrze7dUIwzKKHJLeAZAby7t2Y//UCfmTO
dTe7BPwAMrqhziM+GkzI1kILjh5LsT05VOK6qerZA528iMMf5PgK01nPCEoEgsRpfjCI0WDUO+y7
dAax3BKr54/ri31013REd8kNNaYL6wFivsaTQqffpVlh3DXAtcLY4INfJVhqVsu5R5rV6gXIhwFN
Y6m3wswv8tqTgS0q4I91o/8RJQbrsViVPSdrXBAa4JxeR+2JIyl5QdQYYqHSAOO33d+ME0cAw+Ln
PGyrHMF7wj2nv9lW0swmrTutnPLNbZ+vfrLAUDDQhzE7zvAF43j+QMRLhRy1xbTD131KtDaV1lSc
LsRgGK1jf9D1Bbc0L+CWIQyuI5oLuPY+RmgbN+SfC0HGkWImgplMfNSEG0A1wqJ2yxQB6ienv6pF
dxFhR5Qq9p5Muh90pL9PXTXic+s8qvEdRZGtZ8juvfV5wReywfyjDQ3wnqwqmvv3FPpZYv04JMiO
2owBWBW2iF83//+ecR/IuJ2BCLFBV/vtZUPrpqulEf8VcEvYjLQo7azr/IUBTwb0yrDy2Bd2D7vR
3aKfTDnIF6vqrK+qxalzRcihbUGeAeR4HbF1DCQyrb1D6nI1Wt+dIVpYUXARClPIWyJ6bSTUoi0b
1j6ITZqlLOhoqoRiAkl9Cws2eAw8mwXO62ELYIHtqJornasuKHARqDDRAZkmI92DhaD6gP5Om5dt
dRpMZCtD1+FQ7pWCG5dmpWDiY5yKpxFc15tzis7gC/DsZRKpNjccjNsnBaVk4PvPyiGggMfE1r+d
wxqWsARqDiyNvR/0roTzd0WM5LR7zrytprY3WeVgLkoyOrF+1hsGL8f6xZGa6KOA8R6E4GVgzeae
7+6bBOifoepfQ08TKh02WOaO8z1FgSVl0NCbe+QbYKquG5sB3jgovg1QEy0RQl/JwKTZRTNFttRF
gkstpF1awKfhG2//dPCGGkrV8FZc+6UBgulVD5KUru10xc+8ZIRxWls0qVhSHJNnQ4Wi4BZPSaaW
eDMttrSQKSj9xYFfsPJXnDzQKsPlx3PBpujrlzNA07oxOI1EJkd1t7dDFw+fsghJfcJ8NOhPOLrV
RMw1PCz64YskP/eIVgmEydxWSXFxxxnkOVo7+6nGQTPZLYfj5rK0ANYnhWHYIQTTYWFbzIeU6GPF
VCEVfKXiBuGjPQhYkdQWB2u99qP6RMffE3w0S2hxFsSibhdUuAICpMSrPq+tZ8Jzcwi+HbTgw3on
1XNrK+xJJQOMIFuo5DE3rKWARdqqphxRPaEjDrtOhHH1aq5p8nCWDeNj7WQd/uslU9APZRtqLrs/
svPRW++UowSYvBxfmQSfYR6SCw7R59VGg+QbQ2wBAAI4qFKRAu4Fb9A/nPq9DkpJbPrp4OUnBzi7
FUzdV3xiAzYxx7VN4NDEkOz2CN3H3sfwxlH3DZXqRk/LzkmJ8U8nyO440VO1tCn4ifjJEeTqc7KZ
wxpE3eHf5t6ukWaL41WO2n7J6Ow1Ryzc4n7R0Kz5dqJPXbJreVtK1n0jJqP6p2R5STs9+qSAjeR4
e7+p0xllnmR/TjiJi4Lm+F+0yHoufaE3qaKf0TA9O3nPPS7Bc/fmWV6uxYxME7CiAyp3nSP7eYQC
VDfKg7xopEoY7g3RCdOOVJg/vvx0Vwno4LY8/dze8RMTr5S0zATCN/uB+HK82MAU9hiOsNaeS2eg
Jcxbgq2FkvW2yA9efEiwBgRrH4m237vg3el3zhOMKix2VId4twgYHPveIhE2YQucf3OpxB9ZOtEL
cLvnR4+48w31mgKL3ufLP+zQtUVy4x82v51DBBKBJurac8mdKjH/9JAmQyi+5u8v9/gBd4QqFh1a
wtXBKQgCuJ+l6KyopP7wAjP2e4n2szQKnBzSU2ndy9XBnUjujz8U5WCVP064V2uUASuHwuVDzUNh
4oqE9bEH7PAtjj0KhMM11b1YsuIUUjCNYL3T6d2+nUFcnhX0ZDyuJjI12YNGlDq0lG9KP1pGRNcY
EckUqW1ew79IphBGtZ+l+D5TL76f0ECGnM6uvfAdkRyPEZd8Q2FAkvi5gV/33E9Dc5FgXu5eEAZD
yo3/itmRKn3erK2frzC1x968dL/GNylvdrNUQurZ4zUlsQXzLJ6mpZpaocJqu6x8weUdynFT/wLc
IEA3B6W7Cyt7PkksAuOeU6fGA04r7vTNqHeUrhsSgR/jKHL+mLY76pp8heNHWz5tdMtZyWP+2QuL
Xxj9TaXY3SPjVWnzwFbRYF3eBaymeW0WH0r2OCt9oO7icrc1EbE8WkQPBP9ACtmOOavAa4sR8x6t
5N5wHDEcxKdJTJrEYoppCfP0LDv91Mybd3iSzhLQfZd/sKiKsi13bRJVXQYs+8Tb52o721jI8FL3
hPORmWDnGvZ9JuYhHgOMOEy7nW/QQRYjZeYIzVQgA6D8zmkBZGDCksGfTThWxZc+21tUyo7N9fvD
f9M9UGTdRwmztAxswnOwHx8VcnkIWQUL2H/D+2K5FN+O6OAPu4fTC1aABHd+k22rOBRNAh6vdvsG
CYx9RaD6eS1LG3ENk37NLJV5deBvKteBV28rOIcTJ4zgxXujTbqSc1ECz0pYaQmYPR1a/hbouj6f
uVqQOVkpm8VQ1jHT+U68qKWJtRLDpw2FLi6bsgO0j8nyWZxoFMULWViiJ8K8mwk1Dh10ocied9r8
6qhWkmbBVs9pCxitSu9fCA18i70BVs2hze8A4W4MYaXRDbp6pysLkB/CXbtCE3R1wu2QfEWH1Tn6
2/RzNOVMXxCnLl7wUfMjHXu3SXT+uXbvDoLmHnn68Ujv7aDxegutrLtXoPts4mM7NlwGLOZ/dA6y
Y6mCBExEKGbvqdVGXsguirIVyhD8p3xYXFF9we6BMA+fa5K/lxTKsJIhNBXjmFSs9TDLGX1hh1ZS
//qk+PzofTG+u/S5zWsGO9F7r37kayXbev2yhUizoSKcA99BcRW8r0dNSPMxJkKDs0M69AJxOiL7
Y2he18t/+KTuRmyuLldyhuCl9sN+eCSfotk5qUBifuuBEcAzG0yMfgh3wTNI1mYH/hP9MeWkmIKm
WKefZ2S5ejH/NchsJowI1IRs0nJ7vUX+mUUXTn939yx07651z1VYf38QoPnzvWfwLQ/ffLH7Pv12
nLbwhq9J1DtZj2qD3knLkWsPc5QNY1aQbi1GypqN3qZAuY2FIw8Gs+BlFPqK178fiXhyzDHqx6d3
F+7RZEdC1aCIpnROwFR5U5wvbzI7buCidgWIi9N9vRTohqj2634BLLjAq47lXxiG7KMhjr6tsdbl
DLZokLIIi57D7d6fQG/Z/RWbsriy4nCxJbu0zDyt2iOXbXqF0gp5BK46x0zrfR2oZ/W1lr3Qlw/m
jQ5GlNZiCVbQHTOwmB/eH0OcD9uHbPZ/CesLqwwkmU5K2oFbfszOQ9+hMNPrK14rn5pV38RTfWFf
f0dQWtOJISmCpg1Zvp+66T/Fl0HizJhqxx4e7XF7bwRozpOJqWnooIuTi5fuJmDA2kKxzN/6EFfr
c7737vNYVORpAD7YkdyK2Dg5N96efd4uwLqDnoQHHoVMc3gKUB60vJ7++s5BqUqxNr9+dZObZRQO
CJmv1WUl7GJqruf22uRnbev8Zdo3ERPSFD0o2AqBJrGhcW+U3fryRorByJIDy6SanLAqZf3F+X5C
fE0XIMzk/JbKnsdMoJ5BuFhou+TkAOH95h9teoYd4zirqKVtOtDU8sEIUkgEb4uAy5b2/Ej4EnqN
mvOAqzl/jivESBLuJek3M5ZI+2R64C21cz0wVzBFHDByvOvRd2pZ57usYhFfmhTf3IobaGtR08aV
Fo29Ob/RbCED2ViMRitosm+GyOaDsOMyMkH4pP5Aad4Mn0MeIp1wLZVBFAj1fqotgRPvayW2dSrv
kTHIMR8LeMOYXymVIexVIqfw8wbAgRjbUKI77LlJQxLXz3b5NPQbIskerRo3VPLaRf1tbfFdsSQX
0KLLAoq5B1dJBxEosTMVA378ZUTvggm5SauTXr3WGbzQRrkqLEYKk2dwtDCYFSCx3qiMI3bTdVGV
jBIctkEmkFXeLDt8voa6KBz+c6ZJLQI1WB0F3GSqDkbNCIz63Z5RwQlGk0/xILzth8icAABXi6dD
ZC4C7H8f5qZukKinHe9CWXrYnlcxzLH/B21VfrWNLauHwW+lSuIG1x9/vfXlAvgzWDAQQ3hDyztL
v3jSNZS9bolGWbjweXAOcgA6NdyycBE8HNatK7TjGjp9VlDumwAgzPYmQCantPrORFfBUwvBvQaH
uC9V5auj1NSNSBZZRKQWC7P6JkFxDZLuf4FztlvEfc1208PCszXuLJf+LeY5m3JU/hxR/ZnmhLM+
4XSHLImPcWKWTfY7IQG4+ZKFkweORO/s3mPwEaEpbsPB8M45KHX3sS02e3vRcx6jR0YoEkc69fUD
v0MbSZU8S1xJsLhl/rV/ehW1VOGaCDxJLt10ArGu/hRRWTadmaDCePXulzK0xqN+i7fKcMtr5Gfq
QB8ue+yQ+dEiyP6qxO0YqMbya671eInBRRFotss8C8UfAj4MLoMYrM5TbRzMr4gVY9xH3K2owAHr
6+47KR13QwFbwjEc4JloQri0pKxdkALizYBQQYSCyOf6JgXjiQP85prAasmKPh+1IKvAsgDFIx8U
9jMtR0tLLPPKSJtNBc2P+ao6HyVDbUeVus67LoGId53udMJya1lPMgSfVEIX/1a5yBKPLRBGO+DH
D6XDACXLQr8k4ixv5Wxsmgao7BOjYrB/LL4rbTCRJR9i9XDw7Srs9tgBHG19E2WuuryhREpuLnpX
Xr/13LOvhUOlB69CqUb8KgXOaSgoZoUX85zeR4IJ+iWjKfIORGcn7/sNqUQ5bery4VPCTsbK0w8I
85UQj90vopwmo0RapFUT9ofrXH4tsnVz0nBmw9vW+iPHF+RwQiDvZhHgV9UiJJRyArof4KoY8Jlj
sQuzfiF7eqDlEY4UBieqIc7pk3mqmKny9NQVXKEh5+l9NODL187y82NFDbKSwa3xRJEu3DoYD9ZR
6tReqI0rcyPxv/QKUlasUsYBsklrjhDOr85ONOit3cuJWc3fXad5DwCEGuyYEJAQBGl7d0xJVDPg
BjiyHs7/JjIbit1Tdnl12/XzHTfYswK9mtBo+WYXZNLI3qUwyMRXO6s+bs1Tcvbh06Bhq6ygsn5W
NwgEnxU2sbsclccNIwifNhX9pkWTGKmd8/Qs2Jn0yFZfI5LCNOyV4aol43GACQcs+zDY4TdUDBi6
hUz3kJj/5EHM3NxBneDM7avisL2G0udcueXnbyOlE44yzCa+cbA8GGmsRc6PljiLlv9pgJzXUSzB
pRh+z4mNJNIV20J1RPMxiEFpR7PacGR12wkLerTFk6PPeKidpGp2O4xi/fOBkS2gAZk6FfTXy2rw
uiFMuK9Q6eKamRmBI2smBP1p+0JdyWkDAePUznFHLzJR+Z7QFvOWGKQBQ10E28R8B22Xsp2JBac/
WW7FfRj3DastLjXlocpXiSQLeCAPtMf/wAL1NYYSupAnxR81AItvY4PkuFa0iIv1tXrHj1mNftK1
XLg2M3ffTWplm04Vjsz6ZUGC6Ryv067yMSniTY/nAysZEzf8tvTqiY6z2azr35gybBDpE1HXIEhi
SP6GL1X+iBgRZJH34iGmLJysCKbtv8vGUsvnrMVYfTagAn66VzBx5BoB5obG2ieJTskNgVyqNLr4
Hb3oEjdfQUjRo1BX3HgGWgmqzYH8jWbtLoGB3V2Kg+CkWFhK8sMu3dqXQkRs1g6E2p16Jlr/4hGw
3npYni/0fPmkp7mqpb2TdENsODtOyMveKpuX+XEt3FV5t2+p8CbD6TN3yXMp5Wn7+fZG64Dav7rC
cZ0BK2b4i93CXcEK+3oELifY/hTOxq88nGIM3282Rc2JYpJQRuHLL8ZBZjKufcSJPymx1GlCUF3V
atHFpkKL000Hj6KegQGNIBtp4qGHdTIeV3xhUKW1lJQ6bVRzSIO7LvpU9JWeLmh9wjcI2XH8/aAV
C/WzBJTg41IeP8TKjmmQMvDiCwcFVSW+IgqpA1iGHaFZ2x3pudNUJcPjcTXB82PdWHluUVo0jx+y
Pj1OOMABcZLt3RBXdwPhqpg/ZAsyGA6NXp4qXh9yxrrdk0oEmV1ieg8G3YENoo6EB9/R9m/XH+oO
HWA8CmLvLWVzdjsNQmHGzIZh4E1maemUnxh1Yp4j8ocdOgLU42tePDXU+YKxpCa5R71V9lRz2m6v
SivMl72zI7Zgemg5lmloC8ONPTN1uM3GwIZtXI4n86wl28N97o35U0NJSptNgJabrL4Q8yFLYDPL
Ax7v+n/fe29jfWLMRrpvbZNySbOM5litNEnyWoMr29t/LelR3yRL1xCFcpmG0rYvLpYDUzrKrjBv
pbhtPR9jd5fTAQJxVtyegJ5BB8qFNlTap3rbrwmiwlFm9yaB7PdKewi4t50p9KEitXCErERKUzEk
pcxd1xGw0/poTc2IKbwn8jXzNEC8fPJICO6zdphiXy/fs9Dvw+/POsMvEtrEONdMMRQ+T5k6/XRa
oe+ZMNqSWlwFMFdqBQuHhK7a/+WPlHIy6wOQKXkiy9YybbLMQukHyITYd008Mcw0DK3cnlWBQG6I
kug9hbcgHwKdQ2E6+0BP7Bk+/QkhPP2pCe3BKZ0aGI1EYQFD6prfjg9+sZxJkOOz81guu2ehsQIG
MVeaZIW8UZ/itDSS3JsV3lz2O5ifYyOcMHGEYWN0StMMt5GkUxd0eWQA6LZ+4N+6LG+7d4S4idoq
ZZrVmX3umBnJH6299wLp6VrQ3kgvmZQ5We7Ok8WyR6CFUUIIhw9xk1XLWRYABWVRvl3MubjoUaQ3
UXGCcjnzZzz+ZlXqlVFiVWaJ1PY7ZxyTU9TMsUu8iGdjS59eLpMAkmCKHU3GmQ38HROM49iNs3SP
pL4u+hBSwnKuXpb7y+NSvsN8DxJ6zew9uX6L+cHIS3Q15l9UqXoPsvfw/T43fQkgW3J332TXeFEa
a7ocXQokgZYUgTqIJN+NeeHysTFk5f8XOJU7+Zzqbj3zLKz07BynLL0gvq1JrHzsxgjc9hP8r2Kc
jD/s6CZYhcC3ghot+xJds8zygGf4l00SEYqKtLTpN6DyJz1r+Mk29ILSVdqK90OGBKJbXuhTJyPp
vuH7cKnAdH/ipL2cfxEPnRYU2ixtLtvsl4HGXiMmbwrQDr7cuNKK8umWbnWTPW5BkZrHwbkq2KMW
9KmFo81tU0/omy9I2WOE1bTadT0TiXVGs526SKQrgLSIW1nJ1+bb8u9lm/dAabT5wbNwA1Jwe1kf
0KLi7c89y8i8DeRZnqQwjxvt44Z6tsTPc6OOxhCyngjAUukb+QqQD3eLv2D0ns/JjqvZxcKxLH0o
sDXRauoEciwXPa1+ronmwLSiGDGDTZisv7pddGVLsj+Ug45oI4/0j9LFVjNDtVp9Me/0WvkFvvhn
fwr0ANHf5U5ks1SdybcXeAVKlIDSk654jdTDh8udAEVHU322/48JttvfmukU6Fm4jMDnK+nS+k8w
+Qyokn7sLLZeSx8mzve6k0CZbRVEMa5ojYLRaQNN7D8SECjHimOhkeo1eGU+A3OW1WE9b9aGHdJ/
TsopCIebYD3BbNRvbaj+ANPhxgAABn3dV8UoeISxEwPdc7OuHn/rUYlYxMxaisABgApnnD/iKENc
wiwKjV31+mEaj1y+Sebbv86FIiTyaVp68/uJk92Nft/7St8CLnwzBfKW2DnyXjJ6FrAyELBpZ5V/
uGC5kGX+yzwFHbIz7nj9JX4lJNBij2K6Jt8tlFG8ghkZqnkuHfYWtV21OxeuT2ZMiKDKEn94LDW2
o2zI/S2UF0cSybnTKlENFh0duD5OeoN5n8xuK0/TRPkh6EK84zu3Y573dR9p04mDRsjYgjpmSseG
SNu3N9qR4uu/AZNEP25PCDKu3fyCwrd9Tk/nt7bWUeRo42EcTsLeYjk9NxiDcpHzaXv8idVs5mG6
uwvctDwEs+ra5yIi4xoxedgvetjXu6/XQBaOtq8XRpM+xZ0AWCnxgk8390bsZout+tpi7k+Loeru
nbRe8Y9ndSi6ercF0UNXgoVSdRNlKW4dKKMXpJyUQ7bc/kz8TWiCsPNjwoldc4ZlfCARooY2KSZJ
QxlGtCUE9N20fS8Fbss4klXpziJo2nXJPBpHVkheilQmefxZ2PVQJNqpqT/D5u0DtP593K2rc20h
XJpt+MtEbHUMxFDfAzEsr+liFdnE/U4nz0elSCTsghRVgtK0r1eoXkskBX11pqtD90k5aphOEPHJ
S399o+kWxJ8GoNMCiTInKqAaoauaqqatBrBy18+NS7dytLo2v2rs5XZINy1E5CWxv7LbtHfw5QYS
L4DMWZ42WStkxjAL1QmHmq11gyC9t+cUhO2llNP/Uc8CI3UI0XGmEBwXzfT77OJ5XaifpzIMzFT4
YsEiLWdA6L3mTlz4JGNwPGvKDBhsPTL+U0f8x66In58UWpXi5SQ2fP04uPDEiWN6AqSI6mk+XIOO
8luNWRhfY05ar1GlQL/x0eAA+tucfBUmgioGng6dUTF3yu648Q72vVsLFt8lqyurzYQFPWrYK3+T
cRxJc620g9VR9K4L2SFoSCh5DGQGK1UD/yPKxXjGKCpmVFfudR6hyvPZU9sLXz5+s76kRzPKep99
4vVYMRpbuPnIgM36FubXavWfFLaZNB97w45DF90wBa7r80bS92gIcLMN0SqKKaHN1ZF6gg9uOPLg
pieid54Wz+3zUIiXrLr9EpGiHpEo5bdH0wxE9LrSrMjPIzUgqnsxhKkWdKj+W/LosBAm+BTogvDd
ULiS+4Axeq6TpMLrd0W7WV01admdKKi3P/ateQQXCgCjk/gnMoBLVlz4IyahuX8zJNw06XZAofTZ
Xe7NUTWVrRiopVg2T4zedmRWDBWM9SFp0rnDNxsocP5SEI7xEMhhfkr/1NrCSH0eRpwq5Wrl4C70
PtwAwy84x927oLbCO+tQuDX8EfbyhIlIBH9GJZasDHxDYdWw38m3KpKemjnTHxU3ozkoP2O4cFyk
/LcKLSRPY6ybSu0e3iUFCNviNSMjNeWMfVPSmSKU4a6YeklHntEtNHqJFK3OyMwRKH8IeL96C5Kd
sUz7vn0D0VGSf/QKaGmYIQ9OebJGCzyQ+D7pzNpiKz25MnewNQrTe+BENzDxSmfWM2/UB0mGKJcE
SFyPmKNqjq/tHe0MIzfc2+6TdVVMwFqisBAa/N6X7Gnj5c6FnsgamzmLhnwEQdj8fUUCNVvSIVGv
l5zwWJrsL2TEkRMa8RgbFXK6hhlryPheG3SjgebLZaOzfJRjZB61Kk/Vqm/Qph/mg4Rqk8bPa8ei
Z8lmqMJ/V3yygyu6EsSa796IEbMaZRV2k3cSqidNxrQ/qy+1P9THv7pQNSIJECLLjJlm3N/Kjr1t
oZoVNl/ab7NaUDb7jEW8dlGT4Sefb7Mr58CMwVUwGtAddsyzadZvV3iUw6GDhcJl8KgrXIjVmaz4
73JE5ulI9jGlILtuJzNvMrhqvkFXSFrfYy1YBaA/sVah/iyBqOdtjXR8z11lsiVnzUeE3EhjWZqC
Yb9xj+nC7215JY6Qgxf5XstDIXFlCLI0lSswoJb+3apxWdQXDbFN9nDicf8OYmt0R/iVO5LWGk9m
E5a5KJ4gkMCfTu3ek0wpzlvv+4IqIggOjRnwCTdIT26/nFU1GUfy8iW1FLWsRj4deLVIz2EQp4Ke
OjkvsENw583BgyXc9P+rWc/eY/AtsCBu4c34mRyKTJy+2s8YgteckokWfmUVb6jFrfmm+2kBv11I
oKL/oxV9e9erdH5EPouvZEc9b3s/tOdPL209SQOunbA5e0x/lkaS0bvf7neuyUce13majMwP64yF
8CCq3gwtZFs1ZV6LrBo0ggawt0hjds8p8gtCTUtzX02Rt2w80hGy54WuGZ1TcttBc3TRLmOqa0ur
VVFzMsmlzJ2bV4jMQekU/QExI2abIA0IMzFsFas3flrSCFXd1rxCQviSLSOBGYXDmo2MxENJJgD9
9cKRkxDFA+3ttV0IbMQMG8hmopobj2+Cj+M50Vg1seKoPtE2CJkHQUIFcSG9r/zovC7xH4rVADOZ
Qg5rviFriMdhE2+E4DZy3nGu1BokZX8diIJ7ZtGjSU0WqayJsEVoK/tVGv8zq4NxBflPJ48cL8Cd
6Q34TjfIpkFgkAdkyWRl9AjjR4yzeMn5+Pmrn1OZWjPNwZ7Mny3+fOK5IV4wzusWVjRhHVhCWgoL
j8toNphg6BSdLSSupk5WjxLeCaBqUuGA2AZyt1EOJFWXrpRJBLiugLgnS24idOPPUTYZtiMdJ8bY
Zk3W/2Pbjjy27aLyJmcDWzNaf5ynm6mVWsYktX2f6TOLxi2htet+PcKGppruoFAZEagxH2ySOg6z
AQwsvg29/vEKcYljvi3QqsF86m4f80VB4WwFd5uf9kPBViYk9mUITOH5Nw0bKPVy2xgkjJmiA6qN
xMNiwdIWu+4DmLnEbyIP511pFe104v0Eyp1oUSjFfPcU720tNefZAPMbWwpAREXGEOLK7sAsP0YL
EyMzEwdRASG6VIH80gOOeHwRBkGe0xG/Zd4fRMJCWQt4yXnCsP3ExDBkChE9JZMdAoHFGY9K729u
/eFFSX6XmmLbXZKx5DrZPNsIRo0ISIF1OQCsBiDXVcomKpfqhRedD9dGkrdtZK8pJxIUBa+o8ZnH
cgO6MTsGsgtJ9q1Dc8W28wokCYuon0M1N3K73tBeOGUA4u3Y7waVvYSOFxz9z6NCVYsvqskbZO88
/LGUwL0vlnCyy+JNWa13qlW0DGUlneMUqEtIkCtrv9reZkgMC1mHdlHOjmXX6Eo7jghBNSEg5Nld
EGsNNDuO+Ob2wua1iFVy1WLa9LesEPlUXRrP2UV3XCCIo6UKsRsJrVs7lKk9jfO5cH1v5zBuj4xK
/4tEC9O8ykfH8dUY1jaFoEnI1kSzGt6D6vFSi9QcWl5797gAj0TnmFulZlzqAlxczlKUE9dyG3+F
k7ZPjwbhc2qKLU1TsMc5RTUGZJMKipRUvJN39QoTDqVY3CCREZFx/xSCXtYNmTkShh8SK/3CtXXj
6Bf7AUvta32RwIlMCZ+F5TBl14Rfiy6vybelgszFmAeNvCRtoKUGy/Fqyeuc5nhFWUezdHgUAwIO
OlJwo4OFqDsLSCQZqTychAN3sMNDv9pDJ4bZIkVYNnhbcQRwLyzWY+glTcj2WGrqp6gwae4yctkW
oDvAYmK03Zpygi4DCBzKlaQ19QpJRktfAhFQjm5VzXOHn/6W3V7wim0KwMxA8uhy0WbukwGqdF5u
Kzr3ZSh+BUlUWDKD9hA8iunTM9WXn4kGo+naAErS+FiDMw9uLBDsaEExPiPzchu3KfQgGR+BCyvF
ZIcuKDH+ZGTLJIU7Fcx0lD5Y1aecUfUJeGhhRzmI0bzCAP/sm070ts2yJGHRw5tzyHOAgTAAoeKS
dBjE3HXJuYGk2oTrGNTZrJkwQoe/dTPG8a3MIbGSp6JqN6omr5kDtzDq68UaMbOV8nzP8MhKOYf2
n3nDMoEisy8Y6d3Xn9pUG1vNzuJcRCpGNoMxPTmzYhYlt52vVKyK4/Auh+8A7IAhLiYEzJ5Hc0Rg
FYiDD37y3DpdRYpvL5lGyf157Q+TksFIhEhHTI/DYAmTqa7jceubrpbKD+jsYH7WDyB5abEi5KSb
EwyjCitldlfCPMoWemAXxUvNPnY19DrroKq7VQPxK/ylq/zHMusBEhRjFD+4zEZwbet+inqfLvMa
KTIB6ciOs3UBaxOHR3SPBI9ZtEQ1hJOqAs9mIigtHi8sDerqzHTNuOdC23wKz4IzGDysZNQunxyp
rqoXKaZ7AdH6L2KmNb7jkzCqGNU1LLzXNPfyO7n4sv0mC1faV5ZARNAhIADq0x5Q9/Gw/fJPHKHO
zqhv0R/4Hu1LdYTbjEKW73MaXBaoc4XY9yQK9ojyNiiuaPkjEw/3Wg624ZCXmbBowpoTUVPoqmeq
Ytlb1oSK986Gp+OFZjX1KCZmSWPMwUznBpRKvZIoHIwC5RyLE40R5zybDMIWS3u3CsWpJh8qX2u8
cDgNRiT0pEzASVoLpCnFeiSSjDGDqxXEUr5qqSJGFM6PueCHzqY2Bxqb2xwU4Giwsesf537J7tNM
ZOEpGg0sfPoG7Sp/zQI+GpNkhWCwrBgTi080Js9r8CG0iFJ0qRHAXQejakMqP6dCOKAMAFbtNe8p
NXDlUd/2osCs33QZRHmdXDb6/iZZxxjBVCLP4emzRp/iafM0l3hBoigTdIcdtuGExCBEGuLRGUsu
zbwMtWYGoOU6hZksj0gfOWqDgxp9Hc2oTiNzMl+Jy1wQF5G29BJSkSTrQ5MPvMDETOXkyYhX3gj/
EXzqLYUshEZ8sCXShKf5e3DMVR0TTB8KfdRg3hmvF8NqJ4JVMnBMPBVoAho9zEvMQ9Q9GpHJ+ISl
zdoCkxCSbqgvfeGubR9SD0KTTGLrVX90D6TBMYl4dhSNf2QxybXurf9uTAqko5+fC2yRYEuxbtcY
6B53gxaJHZr3fAehCqakbOIS+kpmZXno0rDhVX0Vb1cSYBny5Ianb+RROlvEyzkhChBuEIEw9U3w
2nox0ovT8m56SPRqcWlOqSfgNroSfApL8KOVYr5KyINfmPRYe+p5c1y1+i9HmCpStzV0xu/QDONy
l/WAw5TmkAIrFyJTcKXzVYY4g6bfYXTQG8qwBXbtlthwD37/j1EzREfXxf2mFHV3ikeDwoa4REgJ
r+335Q5QGM1M3+23MiXiOQ6tg31+Jj5IMjXZKh94oe//4gLARWCoiiKk/2yTgY0p6Y9gy7nbD+ly
faXRfhh8SeHGaJRxrmuGGZ3fUId0ozN9VEGT/hfR3Wk3Po8ss8GYP1Ebxx3HAW3foHWVIhMW/JRI
eVB67H4ymYo5l3Z04bjKvcd+ZHJdnFAUnwpb9fsCc1Y1xGmTCRZsZSIq8KvLFi6jdupSsyW0GPct
ul5+FZKf9ZbeRW070L8pNgYdfJypGxSTBQRo2VKUwHa//LwYG9PjHOTD+BTMGza5nuxghvPQB/aC
u810pE5m8sfb5WZu7dcFr0leR+bDElwWcKQUG+eXxEIRujp4hmbICVn6/H+B1KHCVWXzTFlY0vHd
YI0ps4p/hc15SGf7V0C1XyFxjvmr6a4KLHwZq/oyJuqzwKKmSV8k3cfdSVb7S/MQCwSISq1rek5a
Bedv07hlyFf9Hl3rr+yY6LElGWrXORNXbN9aaaOEXTqw/nOvMy1i3fh2ZAicxN/zOyrEdG9YSvK1
1Q9CLu1Gh0JRvlkPxmYHvXxG9BS9VmusUf6m9nHOC/JRS09GhAvE+Uu0T8NXrm8GaQQIXNUfLh5X
uYlNrQZz/ITXhqGi6tKLM3Y9lP1JuO4r+9vc6EfX4glVRmE9GE9DIGrFIsYGCmeP8Pel4hGlLjoz
yoekyGNHOQ/gcW4xjrCYhkphBXtGvcQTm9GscnhZ+3Sfs2W2sDU4Cnt8YVcYHsWzp6mNye/9jNqa
LLnnwaZ18LV7n93Z1ec+jeivkbtcx+E0MaQQpXVFfIRUriJfCIumMkEGRvlu6tj1S57QtYRtFLgx
z8dBFOOD95xChbhQtlQIPYPUT6u6m6sgomL1MOmTyRd8SWpzgZzXU4zehdu4SCbWBNvS7RC4nUGY
QzcHKybFoN9db78Z5nbQsTMxFBXfqnQw+0LOG+r2c9MsJ8nP8PyrTH7nxY/9LRvULBj2DtqU4kib
1mVWFwqnFAvt2jRymHqCCkJzBiJWzOiDsKCzLNBlC2rGfonsDYByI5x+83g4tQAZegxaHQLEv21c
3Blf0kKTUc7Cw70bqjf8fcvW9TVV+9GSTWvTSMCm3iPssryQFNqrhfAPgAAogXskgKnF8G3FsIJF
vA5DuLTWmOwAqxKfbu5i/ohyZXH1fOqdQmfFe5m9mCw1EO9aSdLFLc7fWzYC3lBfjCG9DO1L/E9W
lTF2OaI6BKozjqPrENk0WocTkHgRAVKS8xNm/xS/B+62o+rld0k9vx1YGrRI3k3qUmKQA/M8ku10
t+t+2uF5ninG0irVzg+lS7WycCj3oezsFQ3z5zOJR6+tI66r5Z6UWkc1bHRoGvPsdN98vN4I+3la
WB4HiT0AtnijysH4aotdZBldp1BKe0IOoFq0f+nb2TgXq8qcOMvRdiwzIfP7keAA8DBGAvpnrc/F
HmwUEKCGDQ4bFtAs1yGfpkJ6CpV8AOQuWijlIigwdCdTc7XuHQmpl7tjo50jdsXuRCjcxE/Y+Ug4
3Z940IaVUv/1UsE/kX9ShbBaqVXSM+G/V8+IJzIPWfZ6CYg7kPtODnBFbDqSB4P7Hgq4F6X9VIja
SGmXHcFmMXr8F5/m1xvKK4kmV60vaQP8YShxXL9WkN4yE/iMk2noQKZoQKvQBEHlX5HsuUadCDHs
nitqRmkCtzDITQBio4hziPNsrZb02kJA1ZdpnOXYnl56fOmQNyeBq/biTMvhMYXvISLTDJM2axqZ
LBG3mzbTGDui0rtp8BcWvh+hwBa9R/NpLJTfHyxzUuSi4+Vril0CGSjdSgIeN7mmkuobkUeQKLym
tiApiyJOJ6/UL/er5bzLAtFwOa+LCDNurXA+WpdplEzcFd9JvsovdNOfY4+IGVPg2G0twoLtYoxi
xz+douW5WX+Z8DaNoocWqLqs2/Nxb23oQvXwuH1uuRnBae6QteybHTU1PFXm1nb/Pp/fyf9LxLLI
0ajNRz2mYeYympx6306pFpGs9Dee9URRuETuY+bF2jftndRHnPULYt3TjpdoIr5iHwHpBGpcHWGH
PtAjO0JNECmPMyBP3gchO/nqghexdxtGl83pqWON/YuTC0p23B5CQizAVACfeWiMfmZ2GqIiABTJ
76GjS0S9UuQrEOBLJJ6FfjdenP3tk8AREKUGkHclYAEkFWGeta1v7N9uBgnbo6wSksuHkE04uoW7
aIO2M9MyBlafsVIunrs1mHrhrQpGzzTwklITfCQvhHeiCmSys/fjgC/XY8pa/9x4ypFFsLO4kptW
RZnutf0+EG/mYcyD59ErQHUBb2CJI8U6QXS175nX0vPKs1kzHp3Tto/RF4yrHjgJUQwp6php8o6X
l3b8xhVqnO26d1232/1mL8mAi9WDg6O/D4vYVvwxnMYcJ4tGE/jrVaTdGcUvet+cVL/YckPgXe5P
Zqpd1A4/0L9N5ZTeH0JPblDtVdGEiaeacLCY73QFX6/R7oi9fjTXhsYoN6KNwICVgGJ0cQCyQY1h
LE5ohTV1G791Ml2qBgfafQwWjluyuC/EGW2z84WwXgkaQ+GBATpTwrBiO3GuC/9keep7kxzwlMrX
7exSVsHepboht/mtnlfzEhPGJ99By9WG4fxVmYu1dRbfaiZvTdIIxmWrguz6BBhr+apjalIuy2Qk
8TfzJIe18Y5vQRm8E+see0gIJ2w9WR9Ew0OmptBUAc7re2gvhxTodPpfwExGa80dWiWcUQ3Joujv
ouuI0LomlW7HMukYK5hGGGougEWbz8Le4Prw5FmQKpvCgEcsdx+W5t2fMNyL5yyw0RQgMKP8/d0l
xNYxHdkp20Fn6gRilGshOjm2hcdIqJ4By7iJCiMVKiDlzTXQwV/JxJh5LW87nmGtZ21GU6xtfANK
k8rkR5iR4dhvB/nkcvvq6EltVU5298rReOqTef+DPYuD9Bj3M3Zw6+aNWgFt3LKgGy2Aw8Ce5gxk
qS47Sj/98xTVY8IQFXZ1uJ46E5UQlW1bB4pPBlAiyD11+KGPn2Oc1E4LIOkgNhDxO+XMJBnMfTgr
wnnU/nIguVI396x3OxO+Zy/W2WAWayBLrAJVE1AyPQbdOzrIRVXUfMJxZ5RUvw8t8smV8r67HRsZ
kRlzcfxlaUfGaI17j6QbGmQwRxrZsjU3riv+9grlCB+g3z6lgMgosi8ZsJvSjBDHvM06O0fZsuDS
KW2oWQ3TyOkxI7abzCY2TEQLaoHgkstqjieuiHC2wLSvW7Vzq6Fr4PDAJ8kYCQfEhjTBr0Wf3HVD
gnCp8DSTRCwZPPJ5k0IL9rMsqxBG0llCCtrXwUjmA228n293376TqODQWOmL5xrtlqVshiddzVUl
onUAi35GAVggkx7frQlVwUlR9ZJgs+vi5gN2YJtAXu2HwIdlrnlxJBh01/h4o4DyOYa4gS3wwekU
W42fVhEiQ9KrgGtj02TNxCRIrQ9HFgXlNhberP9wqHY7wEe5V7dFqrjedYymlZnIWfACl7AC/mA4
sowd5WL1fpFGYvmJBNeICnGXgLxyWBaRGKIGwchhD+a4iYf6bmJx3fNbbEgzleaGrSUXeitSqILE
C4u3MPV4J/tKcEF1so7NB+7+xwHkKyYo0ELFJLpwKVnnQN1GKTIobWM4cdrjmuZWyT7QVdgIIO9E
6d+ehnf5kcPVdRmLfQLSWVVEOFYlxlKRM/lBx1eIL1YkpVRj6G2fGG+ItPcS5dMH51j5UxiOx3co
+sLkW0S6UEeJia61b8+Tiv3r1JN+eE0s/071XG3JV7VUbRRE+vJ5Ror8b/fZAoGg7UGSWGzs1/+D
JRUbNJo/BBgrk6Och/bpxIUjVgeVhphYJmtAu6RJne1Y3VEu/0ukvLu7tdADKtmEMnUE95ZedcSm
8iibZrLxYT68K8GsI4lgjMPunHNnY5fp8QmbHw8D7micSEJA1l8MwM7m9ON2Cv9HeVAB8CRCDjcv
USOOqXWzAQKdpNyU+oapY4sC1DDgWVVhxW91Xu9YA8A+nD8mQ9btm22bUwRm3IQ57sIys+5ghAeS
bJ/LoY32mKoslJmDB3ZuuoylO0L7nWWB9AkaGKJb0/8xJE4tF9AyTpmWSAII3YJp381vyHdQHuT8
aBmOiNblr4TRuCemglNBHJv0B+qiZj5Gwu+nMATdG4P0Ct3ft6CreCCqXhVGlB3V9hZJB5lmUHJZ
Q7Sazq7Bf70VtKQW5trkVQ+et9qqDFzTjR3DSx0usqOMNox0K08TdRmve3uEr98EBzI5ZQnNKQyW
rWN99FZfEwkfob9afIxx0cX5AHuleZ0pd6f6OR1Vs+HxickzJR3/xAQ3fMh1zHYTi+SeMIRep7TW
kXvgVGIOBXpw4Exyo8kXVzGXKUNbR7P1OcBtxq3GI+Bxec6MO1YqiHMRh9cwXabDFtzA6uxZQsuh
RoiLoIaWgaMFVwz9eAUCEM4v1FfSN9pR6qefycVtKw46FZN7+9QHCnEWJdCin3FooAgJpIvUjOAB
7mvf4BWC8gtzXTWm5nQjtlR/1HJWVIR4xs/bouopoHlwhqVkRCrWR1MgmtSesk7IzUeOByn6jlRF
rNvnHsLd/admd5S06UCixhACWBqVoM1AmmVXr3D1kBwHC9cJu/NBtHgBB199jL9q9YAHfBry0/Uh
TsB9a+vvmYyHFZENvlPDeEfhLn7QEcIZPMWyVofbWOgZYKmpixGGrfmNaqcOENw9umy/6q7gmLjG
YsIEigJQWOUg1RTNpTpBLOowAb/MmTwdUFBHG2EVs650gcO8/eQB6cImdkeen0QCMTD2Ijk4atv6
ff5DUPDk8d9SeeCmk7FEZELRqjHnjcC8l7EZKGlxCu8OpkNlvPXgICXG5oPuWD8I0d2RE/5P43ZO
qY1f4joHslvkdEc3+HuW2SlfB9LV2MqGOWGf3XMwPkCAUJyMDRs1cZOmKWINUcQPFOm33LGzjD6g
uaVN7Ky/TqQRLUEXyxCK+w0zX9EYGClOLjlEKMmHeEF4wG4HvVzosWYnyE23awnimKlzkP1V5ZVe
HCpAXgxCesueswluLhjvZncoteJyR51/O5hDCbSuqJMAiByMOI0jYE1Vs7vylQxyus1suxSEh7Sq
pYac6wytND+OHCzzjpNz5uNa7d3k1O3rOpFlpasbO8iLkZytUJFFzqcP/U+bqBbftpAJALuOpcdX
1L4CD7NBYTaaU9HGqBzNtlMB+Pz97KU/KuS7Wx/6PnTdM3G7QJwxI4QG7khaNq/sjCaKQ1M9pj5G
23eEhhoR63x3UcZP5HmBF1F5MN/bV0PQObZoK/6jlPOr3er47MmqLqIMcqlLuvC1UXrPwokXRtIL
HsklwW7TsEZrYiMcHjzT6SxIiXeyXpZAGXmuJHtWwK6dX1DoaeG6C7rCHT2KyJXbbILVVkz47Map
3zAKeqHvC/OmPytHKfJhBuYc0sapbA3fychBlC2ByeS9hwxetqhI9AfOzU+S+7DFpptxETu39olk
qiwLjCpS1zSXUJ0TAMht+Mb+bh7Xqx+Ihxmxc2O7dxz5CffwYHV8W4SLog1VOdPr6mXipFagTbVr
olVziL+zNsrGoJkqjRlrIAHQ4otXneJClsEzkk5HRmFpkOlAFZpq5IxVLd/ZAnybnGmZY16Iq9EQ
ecOJj2jo7ZbxwjAN95sMPGvu1y5dX8lfVWDbOXnaxxuaa8ZxYyUKvw9HJEDpiVRUxeaDgEVq9TUV
xDvLpsu18bA6PoRiYiK3aQWMW8mIhX/Yu3+7okFxOD286RhFHj0DqDOxZc+Mo9JAhwcnTOSKuQWx
U0wVqL9F/c78U7GkpqB9ZOh5Iz/DKU9rRpE+9beRcHSC8Od4UNqUwUWySOUfEYACykACyg8/lS5d
BLz/lsPcHHHZvr6hZnUXzf0Sdfss64KAY4g4ywNimpB6BUeQE45bfENwyoDHPg/oViu4gosATuvA
qgWCLXltVY7kd6BjmKiCUtUkGMgUil7pz9407Cb9tjsLPXsQd8xlvZbdLZPPNsmeGjHLOShUoyYE
Po3VKN2eBU3fOBNodzsOVO2bUOd25ycWCmc/cdLH8qvfGeb7qQKGEF8kFjssX1DBU68MjXYSB18b
CPyl4rvcvkCY0gpNVhC5OiuoV8wyk3JiSJ6jIZJoJAGQHAsoYVwnoPtp5xDecERxUV4nFwwfx/J1
zWPTpXjLHqkj65ivkBMhnPme6BH3LPOfZ1Buywrzzt4t+6qPO0XIykZrKIrxwRQwVsvRmxl0lxvg
itF9/O2gALOHyhoBf/nVF9DN5KKKHhVzQ5XGg+AEpwB0B2P8m30tLfUa3DDy3F6342YMVNYNTXvT
prQH4K187ANdPVfx0O9YbVfwi8m5RGlN3BKihdoqRmkz0dCF3Lwtvg/d6BJmYRlA6GW51/f+Ha4o
T4EToYYM3WJGKPfXbiJG9TmI3JuRtGwOC28CssMJRfjNMDpeTRAsyv5tBwoPdZN0QMrlBsO5dFUy
9tGvCTAcWIJTeDwtgDpMhyZJQ5Zm93/orByCTJKS3AHJJT6nBDz3LgrPKAFUjUgYa8eze677w5tK
0TzAkkWO44Bp4Y0EXoRxhxJATMnPydnb/Zf6U3eOBF4MynKfz6f9d9lcmMJSEFTNwhdeuhIWcpIH
mKKTrCGKVN7VdClaAhNk8jlxwoIhm1jye4TQAypfDwKeZUAJ2QxlCdMbKIhdQG+AKssi1DEzGuyb
ekxE7vV36fSnzAkV4vxz21PjimzbYJLyN+o52I9zno2OmWxXGFuIR11R5qWCrI88yKzFTPGw68Zx
QROZ648CoVhJxRuvU61PXMHEabXVt/AW1PG+KWCGdM/GHzt/biBLF0x2TEq9G6ihx2sbSIsazSfP
k6UDxBnoTBPa+GH1q2qHk6rxsEHsXQHkdhB/kGz1elHWNqSpltjsTBalw6mUyb8w96nbvR/Ejz7a
pOWwW3UaNgcLXiFLdLOSC44Lo9PK61VYLFtIMUuAOqu9kAcxH5DCw2g6yBcdM8aA87SQ2KWcMwyz
ZFPdQ2znJ9gLNIDTwdwEMpsSRjr23+RDidYg5A5ES9uxJTRPiiYDXDZmQ1EStE7a0l3k2SaGo6Ot
6iSHawfwYu02Zi8+Nk/jq7CMEls83Lv/x1BL7EV6msU1Ns3SCaXdktNYJatp+ghnnNS0jfjjqjlc
MGUcQQH4MSMXpSL+lcpbLWIZwvwWsaHhY1N1T+qla1wz6qaGFeZ1SuwKK5x+tNPseijktxFRkshX
B33izhMulfIA+Q6h0ehMe3QkuZyOkNZo8h4GQeaPBHuiVeaFQBpjSaZ2SWDJZvA424mgXUWRA6fs
WOl29QFxj9cM5Aec56TVSg1IiYUIPLsqvIwSK/dYhXfGd9GwmlOsNLwR+6O057Vp/gH2nbljwmci
5f44JIhC0MCmAD5GsnNLA+lelRbUHJTZimoZMr5xxjGthcBwagZvVG9379oiSsSZ4SDNo3XjcP35
tKB/SofWCGHwOeeM8B2PZkDJv65NmQAkcgfmeTwyLx78gk6WloTgill0ta9yG5J9kpRiP7aPWZc6
u5T2eutUeTfSMLvdJoR5P5jBrTnxKtOsw4FQ+FxCxCscqGI1c95ITlTu/BDTEE5Wl7cWuCjBqHvr
k0z08iD2C5At/syLPtpgrasq83lpugdMPFkRZf2nMSgj451zeGqK9CGVTFpMSdrbkX9I2fZ9GNtd
Wt2v+qLLhvfAZx7SV9Keh0ieMAc1CStscSNKB9bDj7GfIVkP93TYzp2nsqSfn5nCqsgMNW0GEQU4
hw8cudr2L7RGjD1+49C9xflz3gJgbLm19mpHPKkXT2u+QUPRvgAzkb7zHoQhe9sOerZiPMzir3ON
fdQqnFpGRnHVd1sACtML8xai5j3mSO1x53/zMfVDSizEyw4JtQNNfWYQnlEeDB4eEH2Bkvhzj+dM
1FT+n7fdir+NdSe3MdGQvgGpFrGhATMQhp0Do7g5bEALphdjpB2yxfU8jcmSjbsbDcYCNltGm3Xi
HysltmItzAizXuc9h18omAES11hfY0WoYByaiRD0V+izqvwnqqc7T0roaD8QjIR6hkTsi7e8/NU0
eTXnMIegTl+WPrMOfAjJCgIuYiDyx6u5NmrILnWtgINT+8aqWptTt3SG5AnynthZHHZsX7gkB6VY
SQGRoX/dEXKVkyhbNjFWynJRYqphnJaSS/d2mmTd9If4czPGn27/bEGh/jzzeuK6D5yERMK/PBP+
PDApL+gFJVcN7Bw8akinttZoyQD4GJ4qeUJsjEyBYbhxFdfrvXRhCugY3YXdIxxBqhoYmy/xPAxw
XbmHcTaAqTbsBF26Q72d/unqfRpCd6x4VREagcAmXd1vDarz28XtKkvaQICKU6yFmYk36s5gatrX
sCMTMftmW3YJB/GIm+kFWAWN2Zvb1Ay6fCRU2NKm8bvg6vVqp+35EUxIRnKfw8dNUf7oXNDF4fZG
MFrHHHibQbSjDCyPmeD9FR/3hTg+6N8cg2qwY2yQyaU+GXgXbTgt6P1ENKKB077xTfnNP3PWNGcY
gzXlKaz4fxAVZWsmeXiZRV5pU1fwTexsWUM2X65zg676Hy/7AHuby6D6gUE3w3lOxbNhY0NCo98V
CJUS2GFXkFk4F9VNHUbVvsSk0au6ie5wXS8+l24C++wMMkCgAaKHQ/PojCfNeWSmphk7aZH2AtFl
Ow8MOhGSCALmTap3/X3/KBqAjVrRqwz6rlPOkqWTfErEY0/K5MKyrvCEcsi2gUgvFNz+MfEOf7FN
aVKvTArxbKGnrWJwrJA6t5iZYhJs7pSRr7JAiyKQ7i/GcLU/lZCjVRSkDCxf0MQdMNDlmxKrRg4J
q8uQjWqGBW3NBLFVhsdt0CwPnb+u+t5eJSMTmCl6YDBygDEFSmG89o+oUl6V6Z28ORJbNou7c7YN
/JMqV+LuDVTeZtV6WMq+uUWE1qiALDg1dN13w2ZssqcrKOhIzrslACfHIViWJsN4/1No0cEuaSnZ
POatPWCUnOqi6f4woHmcZRt76FBS8Z97QIzCauzZVmijmNE/hz7GePA9KHEIdmBAn8fnc4aAqTu7
LM+uqibjIXNBExK82TmZpveRA0MRAd/tOqpKE8vKdG0FT92JLl2NZ5b1gatpg2GL8tJ1u/XCDbCl
1AtbD6e9jwUPqkYtjUDGu0SAi9EtzXHlVDhtqSSRI0+RGGEE2wJSe08JpDryj8MbHhM8FEwN+P0V
ABgNtz5iLFWRhB2Ix5l8eVNuuzj4XKODHiSsAtP7OUkCQYt/LBt3uTm0NbcDGASMK/S1yupekfTM
XIoC+1O3s77kEuO+xawIDcYjgUAByJ/fLQm9T0r9Jw0zwHxxzQdvhhHTUuDk89dX21THJoaIMA+R
WTi5/CflodXjGSo+gq1gQVzIeDJnlN3iIA3E5RuPXP2i0QAd3Q9muhKK6HXqRNJ7wC3RzNy/Z4x3
hHk3uDiHfGFLuISo8qoBD53Qz6my3Yzb8DCSNS/1aXtOXGHkoHLQS05LQ1BnjAfGtfkViwrYA1j/
D37HWy2PP5Iougq71gIEDv3/V++mZkZRnMmQ+nRvMgniVZqW8v3pUt3p7nUC6GoesbTvLx0J14R8
vMTZn7G/yAMl+EDlHF6Rcxqo0++5+x+ixyXJjU+U6upof9HOf6e+iC9+Oyz1ZpTzNHAgY/Z+ke2J
sv3ojvtGnI56G4e246LMN3Qn8l0mbsfqvIp2JSd8ocEDDgWYvNl/dWtN27S5blThSOCuZAhFVSqb
Sk0wn/aN/6V5/Qt+xcTwYbJIVhsm2ebUmw6K2sDlici9GTQSsIv1M/eXd/kyWiN3viT1g/F2PjOU
wngSdHr0WWapGSkkzrUKfeQkmEyWUYeZMstEyAl9Yzp/AQGmPP8b9rNFv1EGnaxa10CcK5uZr4iC
I51cTZilqZTvrDaGHgj2jV+d8b/RNAmt2Pzfn3s9yDxSUd42u9wgXNFlSsxY1fdaVis+31r08bTO
URN0RyUtPBAiSvEN5W1joF5+zyEjuxQMmwz7KmM1UoGQ4fxtagq6b5vJ+Bq0co/Y9ycleGasu/v1
wvFLchFnMNSMIv7dFOvWrpm8HzljOV2HS7lGC5tUvAkJW+m0yV1Uw9arrVwjszssH14cHK76LITf
L5rEbnZXjlMPvS/N5DO8gOhIpbg3r8cDI2YaqW3wnmiS3FUW9JvVN2rI4vieJGd5oo3w/zDp7IOV
+DMMxzNhQY/2C6lzkAv9oewVgFXWv8HLEHQrKLSb9fc3pm8GwTN4b9V6UACpW7J4JSYJUOWU42/3
HA6r3otes1q8CjbpaQSbyOTLxPXD3OUIeNqRrxcMx6bEtU4paGioILy/1Bme2hygrir4w91pkGj9
7LWkIpcrpurKEdOAiiaPThsXTb1FA8T0oxpm5OkV5Z6ZvYLC35FR24CWkq2IyUbgIMTJ5Q6Vvjd4
S6F6HHfR52eoMsRd5RKTTdkXd+kKVkdQQQ6UzqJDlY3wrtIFhGnTlmVwbRTK9NpJTJExIZKdNfqY
lRHwFqdoV35O8pwyyhy3PXH8/v6w92x5nr9StT0YZAVNIbzsJcbCi/zeDfFWwi9seULJr8+LIHmy
l2CWPToTvpUf2m87Xogeo3ivAlLmKtt390mdbNwB5Sf4MnxetDvDPXbILkET1sooJVS0e/nVihkY
rWY3WNyz21NKViB/gSVJVDAizlrMxKfPRsMs7iJYVHr74bxHXL+H41RJHLGqs0f6ZgbXhpLTqYhB
5w4OY/L9JyV2UudgDcBT6nbGri5Mg7+N1HwzOwcACAQ/ua81oFqvn0+FhlLj9rmfiN1onEmrwRb4
C+1TQsOfcPlQiSbvGBLZEFWW7ySAKhm9wh2VnuTH02A41Wf+Hv3z78s5R8ot1UmEXUnzrul73i/0
fkn1kamiHNx7eJxGzw1sBhzyDtjT4HbOR5EMB7VvyTKVqsX0hVJ01pjNaYRGh0iNRJ6bBCCjgteT
BUxHlCQBIk1hI7D+hn/exMh6BcbDlVuFLnMolNzizOwPuX1vGBrVGHxIow62ZZks6Rqmi5R94Yl7
A1zoGjzNBx1lLJOwoBNwXlfenh3wfBuBOzC+YbFk3yU6yftIiLB55BqBpkKdgkVp0rknKpxjkqLl
DsJSRaRRVwn2XZNyKBHVEqEKI6D/2kJKn5aTCKN5/PGhtWv6qBcJpgGYl5fhTVyyuD9uXwLWOk4m
Ib3M1mhGLPZUb88mDNpIXlZOVQFYC7zLmXePyG7S/3ZtcZV52jYf89EH6qUxlzlsuDEHWmF5Hiym
/ktZwE0TrKgiTjTRf8bqSu2MJ8bC+5fCnQoU2EHKq3G/imvEPKpYmOrUXPvGZPQ7YkTQfW23Ttt1
kxuwIyHd9uSJNlZorTsROrEjfS8pZlrytCAIzpuYCUECIgCPZgjVrhRcN1JFa/0rHXYbVz9EFz/i
tug2Me7b1WZXFrC9mSOR6ti4xjohuGqX3RE9OqFcWVLMDkUZnKxe5+eGcp6fqIqFvwfcnoP4iMTD
EyPIi+98CxLdBohFLHz4s65aLDMxMtP+iriOxB1tJv/ibMS3VGAPPt0rRh2Ql4DqkBLhdPBov8Jn
Qu9CNRgwG04/KRK0pK1iDZKB5AUG1sO2kot4p11hSVFJn5OhHAi324AJURy4ETiVT9UgKBy+GjlX
lmaTmizHh2ih76QE42am2si0+oCkxA+WFoNgZ1fveC1aaSRMkH4a+PUD/yeXQA5whlsnhIr/QqCP
Uih8Pw83HOe9RnC7N+hAcF2f3dxYWRHdLYQi3YIJGVP05bM8k/4+tyGwerHUEFJNGymaS031iomw
nSEsXkxTxwRu1QkCCUY6ch3Bkvbd8uTkK0rqe3AywMb5zVQ6MllFvhAV2WfxnYIKJqQJWkhW0XuZ
y9cwFHWLMAZ+Kmt7hfs2N8qoapiS+nVQFnfHMJF+WUTgw4RhYkZDoI6NGG1tITlFgTAhCc1Mcprk
SxeZH0Dxy26lia9QN0WC8WP/vCAf8XRK5iHPQvACmQeUqmsNfA4DJ7spERX7jaXrgeOVf9mLDuJc
buHQkCg7ZkNxCLCK1ql9qvPeeN1/jISOWq53/tmnj3T30K6TQHfL+vysc95CacCvqwSl2DlEj3O1
ZHAE5BYfSGxPkOfkjfgd/9bhINrZNKilseGCCuOR+yvyeaS15xLhJ//utvQgQFvnlTt/GS1HThur
Io31WUR/R8xm1OsWZKCGcufU/XCgOvfIlGC7ySbZHc5O47t5xNs/OLOYQBMIkblT4v8l2XfGCUJn
CjmP3GX7E5QXhrwJQ84KIoggyTOQ1sQn1AtTU/JXfYvXF6x8rqhAhmt5NVzf9crtnTRlH8twuzCh
JJUtbsadxRtJaFbJB5TOmHLwMvZorhJbODQ9yOCsNn6FGh2kc0/d5bhl4SlQRCMOt2jsfw9z0wj8
8UZhqAPYg69s9WddL2oGpwpGOr8eWmTgRfOfxiuRDLbGVwiIYNF06XR8Z0hh9jO8xo3UjaXkB+z/
2w7meAKGkNvJ6jZu50y76IpcNqKClIcs5g7FgdTprKVCfX+YizmPtjRkAQ1hpTcPVnnzaUnLimk/
3pzm6jM230QtQQ6ElPHA74JpSm7uLifC3B/fc6XwI+8aXqxPA31nE3sEA8/lvXM2PuykTLwlFqaG
ZdNLvPunP21mviSoyHpNs8EOLMc1YtiowcZp2pc6UqESIPjZLFrQKfR/NkDXDlqlvRoADsfK4aJk
i1g3Q0L9rpQXqQReqzjjmG7mECNRohkfJmu2iyYgOIZ0/3dU71rA4tlVD22IIuiwiRtEEO+dyDRD
2co+i8q4lwSIBXbxtX5RoN7O+6akMSDNP8nnj156mlGHM9FAOp9xwCd54cfnnX7TZIU853Fs72nT
kQTDu2H2rBaJbyZ/64hzZH6x67p0QzICUkAyEJHJDk/RkbPe06uSAdcD8287vYxDqwckJuh6l6Nu
PPa/3U0XPnNSexc4f6QcdmqkAIGCz18QHezoI3fazCLRddlPR+7rAhqKk8YikduMS5OX58lAHdcQ
ktJln8ASPXoOVfu9MTHZz4WhTZtJyXyfmoQaldVCtiA1QyEYz0QPAWfL8t/G0+y+ySsx+zet5PHG
juusXDNDOljBOa6xebWpvGsMCT8XCCl/AbyLnleOJ5p6Vr/onge+1ENOq3Hng8ziRWNV+MLL5S8Y
PQVJuEXyytd+fw5eEMXgVDv1v6B4t42yYVcUc7anH5wGrUwEXVOL+v4VvYR0nPV2zM23jiLtCKKL
dThWtIcV2TXWJSgYd+SeUD4ciPmJdMKCfPZjr5hDCnZajuVLRyaKJR1gwp97pGlb0ew38+hhOOZ0
YaMNCRGwPNMbeSiTzfRkOX3AiFU5hbpA4Z4NLYtjqT6tK6M/w+UVDPzyaBoypyE3pef6/WMALsTX
at4j87/iijV5fSnETPpHOk9+FhIKZhhfcpN5q/22IoMAeMil/VDFGfoseOi5JzJcAYQbTIKBzoqI
DwhgEgqDPfHsi6XMv4i8PGzCeRiesSdxo2uAdK8KHc/4CqzIvWG+xlDwzJCLypptTZYwGhV7uM8l
OlTYtqsdL6rdq1n0lAQ1T/f7b8aohVcjxST+KAhCwiXyA1JUy+WG9p2bMfZyWhqr4BiB6LRMLYpO
8RWv1nkdDNxpC1kJSRvDyfQFqunBOMv0dAPCPywxY7UTkAbsyK2wVIsd7LF8BXLofGuscZhYUxBq
jWAWmuAp4/7uMc60KsUaCh9Rg3pnEZIoJPgiW/7N+f9WE+SOOgKbyCMzK+ABMEoOkQEvRqAanaNd
ImMqm1HKktRy0BhMtoC6kmB4RLhR/D8qynShIpoiZzOso4Rc85Bpn+bYTt3e6O3XIGZaBXkri2HZ
Y2/fWwAwEh7y0G5KCVXpCwWMZQCj84RMzSV16MdKROkQMpAZszvikfS/04R2B0ANQIvxG6UcNwLd
OhXF7dsil4rgp/3Wu1NdqdFNC8ZLS9mY7+b0ESVYDuozpSwrPQE5NiFSNL9riGnbQgDpSrd/ZA05
6Bnnt1vyIaOf0l4u1WfeioJStWiJS45P/vWOkC04nXomt14iU02/LS9G95tD6yi8+dSwryjEU6Gh
cIPb05r9VPyBKBq/iUefqoPxtEk+l8y8T2PkkxEsFi2O0Ne7MwkRKpOLAaGRhtfRKSH0fSwzKcnD
ZFCJKkT9+VwQGVchEKLzbix++KAnoStx7ZyCsV0Ih8q0KBun6XCmr5zEdLp2QO9Y1AK8LhtN3EZp
69oOpy4WLDavmOCK0w0G706I1CDrfa1nj3bdm1s+eBZymiU3tCtQ4/rk3daMk4ncZJL+ayz8TFVC
cPYw6RXoYnlqV06E/F9luyN49CjMwLa6s3WeaXDpiBq1EUhIbAPn3zf1fnrvfzNYPKW+Kwt1KP4d
Jc+pde4t+TbrPDHQDHZSffR9TlglDGwoU17+nEZNm8ZQLVc57FDVOGnizPE6KlAjITV9fxJqkhpx
OhMgnWu9o0otEkSnczqE0uYIjW291M9G6sRlV+DJERWQRqNy1kSU+oZkky/b55JKAuz1gIA2496l
4bggztKF90BkYDM462CzcXYtTeuNtkwCQ80qxIU/y2IT0PGmpze2XoAGh2EwRs2BvOFqF4vrFV70
EDsdF4hn3yq/QQLBDx2S2GyKC2FJKCfFN6zo4QrG3QannrIMZDZOZRiQ/Rdt3bsEnEzSE3cUWAPb
+aljzn40Lg/9gClSC8K6P+8NdIlUD4JuGu0btrqI03wzArdb8PLwjY6FO2+0SXyHI31rtKwXouvO
eY+Ep/2RzbSd73gksz8oL4o9aAhe0LSL8YQdP5GsmK7hZFZY+vBPB7X2GxPpT7wZJijB9tdTq1IC
bSsHjmFEeqzh2VxEd/Rc3KeGEDbLO78v3bNoZVn58oJRvng5VNJYdmd9GRiU5FVJV9ZNPsoU2WAO
TQGXtm0wek0eozRPyEJbJt4dObm7s9KrKKqBH1SLa+Rbm6qyNxv/fVDAnFw0/rTgVLykD6q8Fup/
LMM5fFDI/lzmRcr5cUMSr3/Mvk5DpZQ7lSI3KKtZB2ZZ/mGLbjOfUAOhxlK0XARuLQqfYot4cb3O
ONweqgnrObpO+TH2tAzDo1lFgR5SoLwTgJ/bLSRG2TRvFoUafXZ9F2vySEf7OyNgnkJt+SgRKGpk
EqbDnQ8OEtJua01I3Hl08o+zxdFPmfEumUCZFmxohNpFm1FBgx4AMs3a8s7lHnpbwDumLEtM4MXu
WwZAD7GqqQ4WoRkXo2RwjeQEdBv8Alow414svBqWOIPMVPdq/AbN7kDfgA4ZlZskcCe5deH6ivs0
G86F2+6rV3/+AvdQ26MInl9FvXGK58+V8isau72Cb4XlM12lMTFmlbSm9L1FNnqTW5O6mx6WnGWI
VnVVjHU8LOIioe02ix36LxEGNEdHWLwjNj054TGww7l/MbL5KHnGhDzLVGu82wqn2tQc+a0PPKc3
rbXPwYjtHy0uqcn10AjzviopQIHd1JYeEOA22GNaBFUvqRfU13m37h9QJIECb5DX6jsO8rJFB8iv
RB9lND+OYwkg4OJIN6pdAXvfJ24Mu6nPtFWSHghb/By1SSkIIYnjw/ioxl48kzeCw+mlv7M9eERJ
36zIRCmnT73Cp6dNw/46GPrzY/Hxd7umoNlBw4mGcIGv5a5N3wmix3lDsQROYCiTcbAZuR5UrMLU
pYm1h2HEHxImvmNYRT/jWx2pEP7y79K/1GUdF7DUfYLCXxAM7eNAGF4x3A5tUcOT0pORTbyJjYfV
oSHqG01PiVTqxZuTne/ryN5wHrqUAzZ5TXJqDb3Yv4KaLyfsIsQPdRTlTKeO2Wfh0skrN7NYebwk
DUVFAYiAH4Jo9Jt2Wd4RdYl+MCDY4WlIMKsSSr9ren/G8k2vwklOyAG7bZVN5tb7Ib7DAf9wJaBh
ak6kTS3jzycaPN1hCqTNbU/fNq9dmNQq52REpL/KmXvpdmmHo9Im1GNoRxXTgdSBgXKvQynckK0w
eCVkru+aVj6+5V/6hktQ6vJO2YcPSkpBaMgvH+rZzntBOYleyJhToJ/TrfsNoKs7uS2MvNU5bNUb
qQEftwtrFGFMtffU6GKF7Oh3C1dVinrGw9q/6HhCjxJ2FVtOTeNalZTiNadbVvh+yMWzziq8fz7Z
AqxHoYqVHNMdkE/unVg3qv50XJ07PNAsDhSmT0/bN2RAs4ggft6XJVD5A9dv0eP2InPuWiQYWp0l
bTc7kyT4KHL7qZq6d7WM68yFl5AGpBEMrzBA8lcx+aAQ1b/UbnSPqH6ilMC0R8EJ9xZangiolKuQ
XpFjPKHT6RvOgpBDhHW/636Pg4X3y+qlXYr5Do84GteglT2GnVTyrfQcr1GUMpYzyG4xCoXnvitA
vjEunQvfaJ/i3rDOz3kN07etvvUFhgr39K8bPo8vuBmy7bzyxUG1spqDuxEeUiymXEo/wfkBtbMa
ERwfAi78/KyTgf8IhlV8QFnN2cLQ1nrsnaGOZxKItS7rhK1HMEbyl8G2KG3g23BG/xWqxhoo+pbl
Im4Kc5brPn0aV0+Cd2jGhAlV/kL3W4byekT3SmDYmL4asURp9z5gEnLMrfQg+N2cLF41ddngX2bl
mrd36MEmb/D1TbuI7SSdfDHF/kWM4pCGAz0LqsFzlejiIvc9yadnu89byWFckmlWcrHk1ElxlbEm
6LnnKkfDKSFCh/FaLkdgzwOoiYzSX/hIzzn6VHruYaPudB/65gUYP+WlxviYmXrAEPMBxfYTxYgn
Rt8Tr8AV6qPoMYnKvJP0hoHkfQS26bKO2gJlb9Zf6P5JFbHDynbX4k65eccAWrSxZ2dX7lMlvcBU
fxN/pD33iV8rxuAg95hEcnhJJDv4iuxeNa49o1rxThM0khbhrdPTQcSs9d4GbUMZX0skRanecjBE
DNZ/lAmw/sfkGAH2sHvwbfmFPN6m/xBtD5oUgxpjNfrJKlKNYAlm1QncKIqPl9FETDV4GEXPc5WG
n3L+KsNE0ZPLuLXvKdhcRi7XvAoWCctty7AvzAb3VORlOQbcU8UNetZ9yEgYIZVXNcrSBrFT5gIL
+Nwuq7uJPqY/wQzcMPzj7b0468RkIxwH5WcbTPsa4STWY7gd3cLg/yfR3CKFR581yiW20hgDwAgq
ZQ4TuhgS1UMQ5UwIrK4dAltiKo3GImVUzicauWJEUX9ucxSY4Slq5GUQ7KqMlMLl2wGTYN+xY3SQ
cxNrHe/P/AXgPvaAnWogXvF8rfnYv0N10FxpYYpwwtoVDlYw70q+fZPEzdl3E6okGNidlof29csT
1zrjBvkhhe7BAMIBMpKgh5yRROig7Mv/Jh1raUWi0bvUU7BLD/vKSwKEMeK7eBj9396kUs8ItI9M
rdcuQOc1tcz++Aw8x0yDlLPQrxlULYJeHUy2hn+VBqlhqlzRl9TC5VKTE6tKHFjqXx/SPeRLcbV6
02hDf61HY2O9T1KQNNb9DkXbQlrvyIFZFPknSVQC1uMkYGUtI+/68r7tBoogQVdHA3vmYmSEeNGo
aLSn5bZ+ZIQM+Rwxc1XvLSQegs75D9zNTgWxRoxJX7VCaEF5yFazx3kLNP06auhDmued8u0Mmlu7
b9qv3AnbdbyenlxJvgeXCoyo4tPedmb1qSCHqrMygiK8kXTlGXMx5JR2KsnZp1Ob7SKzRDEtI2yk
vIwXHB+Sv2DB1YbAsrz7beOoOmICxpo9r2I51Ii9kvJ3pb2pddotjjsw6qAw4UkKz6qtMgfaSNBM
NfLGbELY1myiRm9exm8080fstVqidMqYkJjbIHEhp82h4KXAjCxpOdSsTidHrz3F8RQUI/IoJQgu
4M86PiQgK3YWMcJNZ/1O4K8EOopqfYEg+8FyD6mS0V4qq2pXxg8l4nB9aqC2Wy1zPNhB2RUTF51o
40Ns+yAh2sHUcwOqyTIvO3OppfjqvrWwRx5OJoJWtCf1Sn2F5TndmlzYb9cyfmswE9r7slvJNf0G
2azs7KKcumd8p4SfPHfeTVN6Oe5tR+CYFE5AFXAJ+pBiZrvZZRb7e6N4IR7KYqkcehhwaBocTO8P
LPe/ZfK2VGqpGR28PYvlht7TUCKPFIdhBcSTC7Hx6+0U2Erp2tcyGCO4hXPeeWka9DChZWzr3rxs
el56xjQCPJNmpVj2HaBnCfTeOGrngbAajrHtIOnGB7ZKctumFTjzG3rcxg9oCRLs3PRsanSOIAR5
UuARYP/nnNRblXskMQIwD0o+iPWnK0FyODIuj44LnArz/8Nu8IBBS+uRQoR/q3we1XOsnUe90ot6
Zx2Vk1aJgjJWfVi82ZrVSR9ba00OPKndepDODDVqxRUh6d0+RT5BMNFt1qAp+gN+l3rLNF6seJeb
8RbubduFH26rK0r44+CQ1MtHx3samp/K8lJrajUqiayUatS+Ce/AWuDojZ36WR4kzEcA+D8qKoqH
TFL4fQVWc7rVcOjRpMW0pMlvEVaz5iIyrv+zs2qPcnXsVZkLe2ezGzQYGxxyi0DUQ8zZ/pwD0c3k
wXKAnQ2bK0lDXJ+sT1V+viUhAg2j6iYsqIrVK7Is1LtBelS+BBVO2pgR5kYeQGNsAQQZ97zSOYRe
/jJ71RfNjzOwiS87hwQsYlvu0S+yBPMGsUrfACJpOfeYi1M7ys312CWQtwrd3ryb+P+rHeGLFO94
WC7+XeFXnS4nfNgYXhAcQ9UvMPilUxeF85djIGfsnX1Q5qUMjz+RxFl+QHFYD5v/PtpE0jI/4pyS
8s1LyaETE49HhtbyQls0q4OXb4Gd/3sJxRlkurJW+k3BQAJMBnA1MUuZlNvNn6FCp32juvkdqY4X
XvLyIekJdK+9vPzsGx8kWzuKuqrjILgWnM++AKv11AD16WnFNFwzCTfdSCBcVB0dYLZHTKlxppkB
rT8ZeFRe2cpjzYsIyHRxSEW/+LHDcDKWWGLC8Bna9seUPOdXVlJBOyGXSgXd2+Rlzt33dy4giEcD
jXU5ElAOhGYedCLtftpGvkFvr+bt6+Q2MR+AoPTbqiCHwoH8+cmfXf56VtnOam0b16C8G3yB38NI
6R4vVwx4e3GnkqSjJ3wHudyA3NTt58YcK+zEr0aSA5sCqTBqJ/PsHLmc18o3DLdVRxQ9vCf+Zgym
4IzjwdOs2QUct2dWJ4pi25lBP3Vzyg+kjMP/Cum1OPdooEC0w483VRJfxN36fBG8cW/QSfVFSUYh
2yenLtsAFisitEuxz+aD8QOuxhRew6WNriD2Hhu8JOFtmsnYS/BOnhEkftgg0LqsZhS4xlbXNU3P
Uvl2MUcwtBzyHgerVmU1CorSOQxwSmYGWMWbOA8ZLoCtwg2B+E9oEpXdk2wHgxK6Cfpe6hQhyjmQ
TffaRaPyIp198gwGl/+Ap7aA9FBRnpxxdaokBrDiq100kaoZJVW+THhjkeXqawHe7Ob7Oci9RNh6
21OebctCHwCtII63l0hHBRCNzKYE0htepX5uL/vn7hNag1lnMhsPVDls6FmRhEZbe/O2//DCGHVw
7SlkzU5U0hbdZ9T9ju/NIEvcDdV70h3UpsyB+6hpWhXdS1FvgS3bt3reKeTZ3LO81PA7NCvkbaSv
fh46wZP69kJ+ufjhm/RnjD7o5ctcQrx5Al06zJ/GsQDBhGIym6fs8SJL5vOuI2lG1l6kB7XCB/Df
CvAxNKsiuUFCz9389hCbSuFllNqXWUSYEN/xPZdzxZTPhU1iN9+FKdruF1a9UgzWNfk99YBnrpCT
coV/rvlFxP0qq7yas0S+56pBLLL/yFfMeTVoq3ftjUV03kCZsl7GdX+LKrU9Cnvhq1dEE8lnWBY8
nIozi/krrykgpj185dZPjuQV5wLfM0s6mGpVEeMqHW1Zb+35ZJRWAargq2U7uKfnWZ7m6W8PSDwy
dj9CcpvfLKVePvA6qf4UUu0WKPjNVdi1voeRhANneshRl/mpwbWyKFDUq/TBEfIZMvHOQkg/J/Kn
zVIV7B8PXuW0Lh2McsPPKEwnVRObuIM35kxf+IOwq+2uinfekd0qJpuxcA+lgQtRuf6+K06hj1xM
7wobO7Xiu6/OxMityDaZQPSW9NfEm/iPj6Mi7ZxQqwCFWQuGaOP1W8EP/nNxdNY48YiIy1oRVc8r
NT1aq+4Ta2x4nErH23dKXY3fzgXhgGU5T+YtxfU+uAQpNYIOakXwehSPAoSEsZoJvdLfe7YH76m2
QLvO7pY4OJtfwaWKU8Q8AfcbxZNJouNx/AtMuBXI/ZW36CkdJR2McJV/UCPFMSTCQBVxtgy2Qb/i
jiLh7BzFVWNZtTXEcMNIcEeOaOE8gwzkQrvBTJwB3ExxIQ8LZ5r0EznFe3xTAAv6FMyi7W60ZV5H
mHAUNV/+Lf8vTYo8QUap1frluLDvLp5t51/DeOumYhkfBIdAbiD8+w3gm4/aF5O0RjPnJIkkleZ8
pZv3ESVgC3kmRkHipldXdn9exsAVBEIg3UvXpF9oEa7cvwuwIam5T23xEx3h3xav49BZm+dsd8hK
DAp8+PJd8m8Tl3dSZH5JSppr3GGrpC/Rs4WJsmW4Qr1opbjuBIoI8KaBPIvXQKKE5y8SdFuSuWuE
uNXBiL3UnHlpTnRPhCNXiXASObRGg6duxyoU1k9VYQL38aOmsC7D62m6qqwjH3wNCNQerFZWfqCy
9tLzSaG9cYcxff/jTmYgCbCbr0+2f1FhMwkSK8kKmYkis7i79odC1Xv0AaccGxaMsJvYdIS3XFCO
VzgX3f3HgMRcpJuKAUa0sY6bIxGxG6R5so7KYfCjGEOyfOEDVy71oi5EJudt1x1T98Xh/4+r6yX5
G7vO5Fm/1CwhNzr+/aBUyEGcot4gRdgWjiLQZ7FpUquSnoti2UtfTBBVNYVrdBHNvvgCjyY1lmnS
5nGLqOr7/jU73obaoskSDsRV2IZ2DK4qqNZKR0f8nO9d+fWyc8NeEYd3hEnrOgbmgCkcVhfEtpPh
CPh7pLnoN7zHKfpmkAXCXZ35fo6FlKXyNVvLeMGaTC1gniXW4DiVGOizihXJDcKzTkoPff7a3Tjr
+ug9rpyVPCN+aml7LDHihZxmhS4SuPyz040NSypexXwaGGZDJlj8DdFwuJ2GJ2qzyndkWNUC2TcR
d/k0h4Eq9NZLz6DZK4vaRjsVZ83RmV4AEZhBPBECd2l0ADRunQWJ+told+ZZYoGAcLZhKOSf9t0m
PVUORtnlEyjXKu+zlJgq0nNNk/KP9AO/LBO/DCVkvaURtkOQaR0TlrrQw+Ra6bIEJF2r8rCmO0hw
8PsUe4ZTIXmgZeAWvGOffa4ZGL4vLZlZGK5zlXfuce385oZB4h09msYUYBYgTh2I0HdbABZMafET
nwGHq79JrJvGdnMz1DdFElJIRvVxlWxOPD/W3aEIEX3T4z7JjEUTMcEDZWovHYupmdWw27GpdtSu
zmsOlEmJrn9qWAtbpjI6vTQsUgZPV3cv6lJUUaY/ZPUkyaGFdoNIGOfXNeW0CAdK1omOMnDbrbAE
Ktso9DRq32JCFUyIqql8xfBO4yPy3EYdC3ovXIH3nRMPN+xW3krmBAjzTshB6PwizfXV61DzHA8Y
bivVWYMVYirKkc4p+Rw4SAQPkH5gadXVuPv8ZOcZnguIRiy3CSz3SRvMJiaM/tj2NJfaq53Ilqov
W6El1BTNSm9tLjU21ZcHbOXoiPfhhf86yuQkjMefnklvHl4inuIzXSWgAEMNaEeuAltmDS32xD03
jTYGWRov2OMQA1XM7QRiT6KnWqW6v+1x/y08uEegGCrkvQmKJuP4mYydbl/CUldlGyDpZk3xQO1W
P/gI3x5TXd45PRwbBoIxN/mTIP+YgB9VaRBXZK6vBnpMI8cBe/n8Xo+WVd0sicSTmeWTTIEdEd1p
xAmkKxhoaXKEV6A+lgwXLYmUvpN0VDhARcxp9HX3IPwpJBHuU3CdfLhQ85uTFV6ECpjIAe75WowH
0/5sNDzAIZSBkTT90kHd06jq7p9tjr2JykF8cntLj5WhjIPsQK+6QAV/pwDy1kPiJjcm2cffmUds
99XirjmcmaJ4V4Q65gmraFrDhsVfKTcwtQpTqYPWw+LGCknvPFeD/IO/aLbn2tqjzQ9fpE7RyWsq
IB5H6NPquKqeOhG+wfJCrweIpooRKlJcUhWLmP3ncY6KmesUC9j+pGxF4XsIcHyGz0j246DQhyqS
Z3dL2EOQGNPELZqHMkcl8phdU/1j7COa+g+pr4Ch1cJ5zbGgzv8Gp9epijd8JjXcfLtAqXfHqu+J
a5DeX2IT+KlEF0PO97XaYSy6G9DC067mKQ+SCc+LYe5ZzLdCD6ta4+o8lWAdRmHfhdUhkUnSBvNQ
7BFzgvYcI4YIVcjDP4r2LDIyG2VbbgW/j84ICET+5JYrwqSXfCmQgefIS/CrIBSb7ms8XuQSE6h2
wZre1ZV0mSLV+V5kAiT4GNUICGgaPTAfdZVpzZl7vPtP8fXtqghk4EeX+lOYOrazHwKwx0JafQ2X
OJIOSncM8b+M5YKqKj0h4JBNmYNp3BR7pL4h/CPlGwQZ47/4iOLte/2IvTeUn98Blm8UvoaVvvrh
MYBHq6yuNk2U3hH9YE//bnMVtoE3TKDODFonGw+hIqnZeb8auzvZOLn4N8sNF+xmCBhQw9gIUt4D
jnyWtWx63ob5C/CRtKrjC0TAv8Iu/u0ey6dxQoIyKhsXzuwK1eVdzC73bMCucZPKjgROSa1U0sj0
royiTSYVQv6DKCIayUF4WTNPZGz2lFHuF6r4wksJLa4oz/oRg1Y+eYQW7WdgBecXqWzL86RiCvpl
hNQs3wE7ZDU6zWWHisS8FJoJwxWzlaofGk5j+V5CUhUTqSyg3Xf9qSA1wbIbygNUkqLsH255WiZI
WpAGEQ2BI2oPN+Uw3It7cQVGXzXrp3gXbrvtxdGHLauNGa6PBJo50v6/dG6Z0hvmMRXnug5Moy+Z
1CEqB9VcEHU3ot4j2HBC08r3M3G0PyGAUHj7pIODQoptfVnIOZ6nvMkJ2E+erfzSi05IX8rXVF0n
e+0j14/uhbZXf4SKDSoUzMtzMgRRXlOHhmeDy6G/uzQSoCOYBHxVSg3HsdRzykkGTuf9zsqCGU3n
qpgh+aF/moxgzlYz4TfZbZkrCQMbYAE11nQKARr0bXXgEif+3zFzMep16TtwYuRPGpql3Xz4CXNh
iM1NIQFnSEBcK/l1NsSjzohAAX+H1Sgd0IoA625dAiOnlsWg8mni8sXfiSxGT1EURgzFbrL1puej
2UK0NeSsJgUEKPTP09vxeRQ3TEp/qC4CT7i/V8DnL84JnHAjUXLGnfjm7AaffgY7O6HuAlSU5N9x
1w2apgYzwtL+k5JmnLVxZ7b7Pl5BrR2JYSEymmeO3uCtd8j8EYCjJSG1ioHPU67A8uQtvibqKi6r
bt6sI7kn5Or1bqXhUg0heIZmJGEW7zTZtLhRTQbnSz71DiRl9033tbhvkMFBVCTgnmQnDin166dx
M/Z1zltYG+OaovI1mnqkaU7u9f0JVAhgyGZXli0/not224+ViZepwzxGEyYwKYXVuz05tUZHsTKV
qB03PcxDGh0kbedNOciHbJdZdvyNiiw22oNIHXvfN7+t4pTEb+VSTGapgHMrjkaBbb+X4vA8+Mlh
8fBE91G2yERsMoQ+iDsaByuBYU+G89QAVCFLJEtOzrIQ/OVQispVoJCpnkhWS6z6ZFLGxjRJ/RZq
NP2jUb/o2Vh5AS9kOgDOLGW6lYDtpdLxoyx9hd6ecxVLeBREWP8mNhoRpzNMqIfrkDwUeJ2PGCwr
QatmyqRE7J3Rf+F1ehKEM6Ll7LxwAjyj/R4rxR9Tf0cjE1B6N7el3sWBM/QSddVCRrRGgXJK5mD8
e2cFVwJyKUVHZi8/oTdu99rv6cZqep7rQzb4izhN2X7x4jxzF+CmsWTl3bLtn4SK6+zebsO+qMtx
hPwVc2I0tuFCSRvtscS68w9V9FM1oNm/lO4A4uQz119HYUxu7jnZp1l0nufAZB6aOrp9uEXlsqjQ
nd4G6zP1a+Ek24N84VWv6GV89wIiicKE9Qg4HXQT4lhuRPHEBkDE8Tvc8Ti435466YuHESDG+vu8
CK4WZxFP/7Hvn6j7zlqGf2ExXBLbs5keif35FwC/1tMS8xFcnryRRBfFLPGVPoym4Yqe+51qj5u0
9bhMcg8TcSuGqnA5IKEjDf5lXNO8rwxKVdhkhGNYJaPWLihmOVupvSIQK1p0nH7H5ELHDBaLb+KD
Id+Havx35Y5IZB2++jGBc4urJqvR2oqS5Kip3FSQchnY6tzqmDNYh9f/Nx8AgAUv1q9vUY/Q8Cp7
LReqeXKRX1JKASnxrn/ulsqrAHj5d2w6l+NIGtM+DpcL8LZHDFw6Xxlpsr6emgBwZoxrkZ4gV94w
PvMmBDybsEmdA31uLe/xY48YuDtJCIt4U/OdKmpX17I5doaf/LVPtsA6zXEwF4FuM+2atVpddfg7
eBqiVbgJ49pJx3Cus00U5KcraD3RwYzyCBnQgLh9kmT03J2O8QKiYHk7R/2SYzVddok8vJaGlPsC
ce54Vc5JhP2knQd08mnyji423sNnTtH0L5jynTUeYsG+fNAJ+q5peAOvPEsLSEBdmtePZHAAmjYq
vk8STFPaIe4R23XLwTXsUwLspIB7IX4haqSAuC+hf8jeJFYRxIcB15Ym36F8rPEo9t03kbMfiW74
+a8QGPQkOOgp/obT9IUMaQoCKxURksjBv0n5kkLgJFthMLUnZ823NiyfNenvdjWdsLK6/UGJE+3f
628ExJggXvpF2W28TLsjYr406pmR5v4lanLIX71/ZJWZk2iaT7Uq4/FERzZrp+sfMGbEsHYBXN5R
LREl/+N39M+ahcrsbJxFJzTApkfv+1lQG+++oqAHBvtkl+YGe+XDGEBnd4HAIWCLwNDZP0HlMMfc
9H9CFdYAoRK6AremLXAiAX6UNy3UbXSpaI5LOu5rRj8oyYgR9h/es4QJHR/0JWBUq0894lvcq0Dg
T56mU8XAV9qQzPC5U7s1aYFVJKwbrVN7uDJG2q+wzWWMnImlyRNsSXIeFpBCkwJ6OjUp5bgspu3C
qYHSe73BL+6xSV+v+EI7qbIyk5fMgks0Is7eIA9yFZsPHTPen5ECoRiGSL329hPIHsAHDKpbAZIS
1Zvq0HNQLa07M7gX2YtORC0o8etMTg+PVTYQF3BYja3sY7OqKey/T9en2KPIkEIxiQEQkAQPz0kj
nuLjt68MaPlo0gt1ROGVeg8+80v8s6iQtkbgtTEwUmRCJ8R5Ycz5B8edBmYDSA2jjqPBgizM29K9
8dT1FiKQUSB7RNwuR93L3bxxS6UOeY+ZFj/dJl1BjGsabBHaRi44n1/9fU0sQ4oxweXRUVk7fMUi
NWNh0Qu2CP/cYhAwMtAjd4srD2HhNgCSU+HDZcbBedD4Eu2gmfl4KNRvfIkcNuagE8EvhgEdLTkO
wrIEzNYCm6xxy9sko7DcIF3E1L2GULfhuGgO4csVCn1rFG2YXNAaaEhWZeWvamnyh9RnkrqGD+Ut
OpwuiNn6ocHNa/AhycNZnbC7vHKPG2dBfU5v4+ZkcvIqk/si2hZEXsyUvW1uxKCRccJiNem+zAWE
HFP8duOT2iAV4X36/KxB1SF8MmIrRnrPX0T2AnXUfmZ0ut929N7NLCBlKPIAbRoieVAVVYHMcgvc
t7pQFGshMl5fYp1NTUTdcw81t+u5DElMNvhwgaXHU+KapX/FmvEKd+xvJx835EmNCIeS8Pk3dkL3
6Ru6tR+8OYgPyZupnobmDMYkpRJxi3d9u5/q9nDSNybiTtHgmukhFgmEtTeD4oOD6VH/RAu3aLJY
bctWc1XXpZTVts01tjy0HXvCWKX9mA4ikpBEVQGAuKIaY9LvQNJEBm8b5yhljP66zZhfigcVUVBw
Z+7B3ZiZfNLzS0r9/30pg0Pm3apro4TkKsrMPPymjMe/ewaXINxcaG+ZsoubhkpLy6JX0AM2EIUJ
tXl3btI/1RrwKrrTpUOin0TnVvrCm9mkZsbAVptj/NpOACBfbluVRo4fQsNFNi2uu2F6EiXT0US+
GLVojKxnBedtPDHl1izkScwC5vewBe7JyA708j8fOP2TtbdL/r/SdZKpq/36m3I/Wac1V35GWOW5
lwqESEJHEAvj1h0mE+7OH8S8GTR8bBqh6Srj3sUMkwg+Ir2hmdQzLAOj8MpyWMTOCtLyeCpKbJRz
KuDwRvAdvxLcVcwzvU3SZ9sTn30Egdoz6HsfsDDl5ye5wqMCh+99h8n9K8kSY6ryXDZqt5zJr3R8
+zN1KvjubU1kk+zeF+byq8WbWAL0fOCL73o8c+6V3Ux+2PR3/1LqfCEbDCKVKHqU18NyfCe71Z9c
RMMvfpmkc0ufRbhXmjwEXrj/ePM+SwEDH4RtQxbXSREeUz35Apq4i0MiUSdZf00SpcUITd4ADgL7
oXw1YnU/Bax0zKgGkCAGMOy94RtTpSO7adfI5vk320SE++QXoayz9i7tAM8tUC4q8Wc0zh+i4qFw
pcK5Zb10HcG5nwXYf5LRc3b3SVit0uyImL/uxsz/4y2vVDIzqRPA+FOwvSFB3N455SpJiImD9oxw
r+w6bDpfVC+XnEvD8+CGtBd1/gFBM4NhfHtJ38hEjNNpBYt/ehqS4jWE/BRNf8MHJKzhNx8Dvsk3
gofaQJ5djMEizPXhRswYPlbxMd3jGGoMRu1AD+eLwtTset8E2SPXIlLd5MnA1luqFctTkPxOyOkS
K4x5CQlV+I4k97IcP9asPPTkcNBapotYCLdPWeHyAbc2EcLpYp5HYSCgdRgN+OnI5pO2YkWehVZq
UvalQijjNn23DBTs80AtZR0/VyAra4FxFsBMr+OTZrGu1pgdXcoPj7KxfVWvQDl5A2JJnU+Q7cwA
dhrwXhqfjcNtbDrM+r/nV/16kZQxex27XkCfqKAw/d6EcUGXkR/0ctEAT4x2aTRcd8ewjKs05chr
6M53f+LBIDoDriZpEyUQkr+/Qrz4LxPtg5XYHoyaFKGMZ2VipOS6JhKdhIq38Dsd2WqovpQc0XaI
V38gg1qQMLzYcJpRR7QeK6zcnXjX2LaVAjgChgLV1zPc1WglSK0+K4C3inUfEkdDc44R18hqQDZy
jKBbMF5EnxNTk6LvSiUkEUng1+yHJ/oMkbQWd+KWHBxMeu9O/1mNFVeHDEdYpnwfVj3++so0akME
dZ6vzi86nryIVniMnSm2j/73432ze193qm6E3fcA6RzGScFao8LOqu6ieu21V8SKdrKytlR0/K4v
RN1f2Jkk93GMblO6UZ0FUqpgjdLDc1uc6KiUT86h/KR81PvHGB5dKbkOLOkJqI13rUzGO6ScVL21
96FpHbDlqSjNAu9jNVomfzRzDFs32XJWFFoAca1oIFYILTxXzUL91zhvb5MHYR17gX6erj9Zm2uE
1tXy+OndwuxF0zqtGsBYZxywPbODU3QhIl36lD1YMcD5kSwYQdS/fHMxCC29sVKncb71moUiSQhv
OsN2GjWEc+VLj0JJYT3hBjXTQNPSqqaWHShFyZwoQo0ltLrmmOsMNnXI5k/DdOW/hEEka1VZYo7D
/gFgIBBA9RtQoSgPzFz4KaCQBuhiKxI7oSQ8HCqnUc6u/gd9ZUlYs5eNh3Wv3cEmPvupNhvLRQEG
aMYIlIZRlI56KqebhJadUyfo3OYqf1tbWpKDJAqGNuHKVnpYutaoSiI4ozpThb+Pf7FF9Su38MkG
eajtUWXgGkLpmkyl73FZUx9xS4bvpUgZmOaGMYNPR/IRtBDMD8Owqr+VLD7J4l0iC6282ASauWjl
cGN99IOpkTd9afkVRcaMglF3RNnLearoLb3EsWpscgZ4jqrLcuUYtK2k7tEp33M5ZPiBrdl/q21I
goAG9mIS9Keg97XlgFITnCD0Whr+1ph33B0GhGXGSXXeKLb/aSz8BJrvgYylGbgqSIMnfye+XmyC
e6bzHSO+bxpINHsxGUU4IrJL1Hobgumw4PMJ3F5RuA2S6sccoJoH61iELEjyJHqitPmSrnF9NhwI
6kbuymxyzLqORrFoG2D8M7tUvmIWEHApXPAzC/U/MM4qplM0Wtqyv3jKHczjPUnRNk8GNDa13tfr
xhb1PqndHPzpv018yIg+KF6YPBWB
`protect end_protected

